`include "formal/assumptions/frv_core_di_asm.sv"
`include "formal/assumptions/frv_core_ti_asm.sv"
