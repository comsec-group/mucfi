// kceesay@ee-tik-cn105:/data/kceesay/workspace/cellift-designs/cellift-picorv32/cellift/generated$ git log -1
// commit eb41d95179d5064eb1a8f435df46879702022c92 (HEAD -> master, origin/master, origin/HEAD)
// Author: Flavien Solt <flsolt@ethz.ch>
// Date:   Thu Nov 16 10:41:00 2023 +0100

//     Accelerate mem bandwidth by using the lookahead interface
// kceesay@ee-tik-cn105:/data/kceesay/workspace/cellift-designs/cellift-picorv32/cellift/generated$ git branch
// * master

// update condition Yosys

/* Generated by Yosys 0.29+11 (git sha1 eb3eaeb79, gcc 11.4.0-1ubuntu1~22.04 -Og -fPIC) */



/* cellift =  1  */
/* dynports =  1  */
/* hdlname = "\\picorv32" */
/* src = "generated/out/vanilla.sv:1.1-1811.10" */
module cellift_picorv32 (clk, resetn, trap, mem_valid, mem_instr, mem_ready, mem_addr, mem_wdata, mem_wstrb, mem_rdata, mem_la_read, mem_la_write, mem_la_addr, mem_la_wdata, mem_la_wstrb, pcpi_valid, pcpi_insn, pcpi_rs1, pcpi_rs2, pcpi_wr, pcpi_rd
, pcpi_wait, pcpi_ready, irq, eoi, rvfi_valid, rvfi_order, rvfi_insn, rvfi_trap, rvfi_halt, rvfi_intr, rvfi_mode, rvfi_ixl, rvfi_rs1_addr, rvfi_rs2_addr, rvfi_rs1_rdata, rvfi_rs2_rdata, rvfi_rd_addr, rvfi_rd_wdata, rvfi_pc_rdata, rvfi_pc_wdata, rvfi_mem_addr
, rvfi_mem_rmask, rvfi_mem_wmask, rvfi_mem_rdata, rvfi_mem_wdata, rvfi_csr_mcycle_rmask, rvfi_csr_mcycle_wmask, rvfi_csr_mcycle_rdata, rvfi_csr_mcycle_wdata, rvfi_csr_minstret_rmask, rvfi_csr_minstret_wmask, rvfi_csr_minstret_rdata, rvfi_csr_minstret_wdata, trace_valid, trace_data, trap_t0, trace_valid_t0, trace_data_t0, rvfi_valid_t0, rvfi_trap_t0, rvfi_rs2_rdata_t0, rvfi_rs2_addr_t0
, rvfi_rs1_rdata_t0, rvfi_rs1_addr_t0, pcpi_insn_t0, rvfi_rd_wdata_t0, pcpi_rd_t0, pcpi_ready_t0, pcpi_rs1_t0, pcpi_rs2_t0, pcpi_valid_t0, pcpi_wait_t0, pcpi_wr_t0, rvfi_rd_addr_t0, rvfi_pc_wdata_t0, rvfi_pc_rdata_t0, rvfi_order_t0, rvfi_mode_t0, rvfi_mem_wmask_t0, rvfi_mem_wdata_t0, rvfi_mem_rmask_t0, rvfi_mem_rdata_t0, rvfi_mem_addr_t0
, rvfi_ixl_t0, rvfi_intr_t0, rvfi_insn_t0, rvfi_halt_t0, rvfi_csr_minstret_wmask_t0, rvfi_csr_minstret_wdata_t0, rvfi_csr_minstret_rmask_t0, rvfi_csr_minstret_rdata_t0, rvfi_csr_mcycle_wmask_t0, rvfi_csr_mcycle_wdata_t0, rvfi_csr_mcycle_rmask_t0, rvfi_csr_mcycle_rdata_t0, mem_wstrb_t0, mem_wdata_t0, mem_valid_t0, mem_ready_t0, mem_rdata_t0, mem_la_wstrb_t0, mem_la_write_t0, mem_la_wdata_t0, mem_la_read_t0
, mem_la_addr_t0, mem_instr_t0, mem_addr_t0, irq_t0, eoi_t0);
  /* src = "generated/out/vanilla.sv:1180.2-1182.42" */
  wire [4:0] _00000_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1180.2-1182.42" */
  wire [4:0] _00001_;
  /* src = "generated/out/vanilla.sv:1180.2-1182.42" */
  wire [31:0] _00002_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1180.2-1182.42" */
  wire [31:0] _00003_;
  /* src = "generated/out/vanilla.sv:1180.2-1182.42" */
  wire [31:0] _00004_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1180.2-1182.42" */
  wire [31:0] _00005_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [31:0] _00006_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [31:0] _00007_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _00008_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [31:0] _00009_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [31:0] _00010_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _00011_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _00012_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _00013_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
  wire _00014_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
  wire _00015_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
  wire _00016_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
  wire _00017_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
  wire _00018_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
  wire _00019_;
  /* src = "generated/out/vanilla.sv:339.2-446.5" */
  /* unused_bits = "0 1 2 3 4 5 6" */
  wire [31:0] _00020_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:339.2-446.5" */
  /* unused_bits = "0 1 2 3 4 5 6" */
  wire [31:0] _00021_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
  wire [1:0] _00022_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
  wire [1:0] _00023_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
  wire _00024_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
  wire _00025_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [31:0] _00026_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [31:0] _00027_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [4:0] _00028_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [4:0] _00029_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
  wire _00030_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
  wire _00031_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _00032_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _00033_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _00034_;
  /* src = "generated/out/vanilla.sv:1144.2-1150.5" */
  wire _00035_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1144.2-1150.5" */
  wire _00036_;
  /* src = "generated/out/vanilla.sv:1156.2-1179.5" */
  wire [31:0] _00037_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1156.2-1179.5" */
  wire [31:0] _00038_;
  /* src = "generated/out/vanilla.sv:1156.2-1179.5" */
  wire _00039_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1156.2-1179.5" */
  wire _00040_;
  /* src = "generated/out/vanilla.sv:761.2-788.5" */
  wire [31:0] _00041_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:761.2-788.5" */
  wire [31:0] _00042_;
  /* src = "generated/out/vanilla.sv:761.2-788.5" */
  wire [4:0] _00043_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:761.2-788.5" */
  wire [4:0] _00044_;
  /* src = "generated/out/vanilla.sv:761.2-788.5" */
  wire [4:0] _00045_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:761.2-788.5" */
  wire [4:0] _00046_;
  /* src = "generated/out/vanilla.sv:312.2-338.10" */
  wire [31:0] _00047_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:312.2-338.10" */
  wire [31:0] _00048_;
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _00049_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _00050_;
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _00051_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _00052_;
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _00053_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _00054_;
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _00055_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _00056_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _00057_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _00058_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _00059_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [31:0] _00060_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [31:0] _00061_;
  /* src = "generated/out/vanilla.sv:761.2-788.5" */
  wire [31:0] _00062_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:761.2-788.5" */
  wire [31:0] _00063_;
  /* src = "generated/out/vanilla.sv:312.2-338.10" */
  wire [31:0] _00064_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:312.2-338.10" */
  wire [31:0] _00065_;
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _00066_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _00067_;
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _00068_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _00069_;
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _00070_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _00071_;
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _00072_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _00073_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _00074_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _00075_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _00076_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _00077_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _00078_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _00079_;
  reg [4:0] _00080_;
  /* cellift = 32'd1 */
  reg [4:0] _00081_;
  reg [4:0] _00082_;
  /* cellift = 32'd1 */
  reg [4:0] _00083_;
  /* src = "generated/out/vanilla.sv:1110.52-1110.69" */
  wire [31:0] _00084_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1110.52-1110.69" */
  wire [31:0] _00085_;
  /* src = "generated/out/vanilla.sv:1163.23-1163.55" */
  wire [31:0] _00086_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1163.23-1163.55" */
  wire [31:0] _00087_;
  /* src = "generated/out/vanilla.sv:1223.29-1223.44" */
  wire [63:0] _00088_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1223.29-1223.44" */
  wire [63:0] _00089_;
  /* src = "generated/out/vanilla.sv:1323.23-1323.62" */
  wire [31:0] _00090_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1323.23-1323.62" */
  wire [31:0] _00091_;
  /* src = "generated/out/vanilla.sv:1335.23-1335.38" */
  wire [63:0] _00092_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1335.23-1335.38" */
  wire [63:0] _00093_;
  /* src = "generated/out/vanilla.sv:1341.23-1341.49" */
  wire [31:0] _00094_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1341.23-1341.49" */
  wire [31:0] _00095_;
  /* src = "generated/out/vanilla.sv:1554.17-1554.37" */
  wire [31:0] _00096_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1554.17-1554.37" */
  wire [31:0] _00097_;
  /* src = "generated/out/vanilla.sv:1618.19-1618.40" */
  wire [31:0] _00098_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1618.19-1618.40" */
  wire [31:0] _00099_;
  /* src = "generated/out/vanilla.sv:1716.27-1716.50" */
  wire [63:0] _00100_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1716.27-1716.50" */
  wire [63:0] _00101_;
  /* src = "generated/out/vanilla.sv:299.59-299.96" */
  wire [29:0] _00102_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:299.59-299.96" */
  wire [29:0] _00103_;
  /* src = "generated/out/vanilla.sv:829.23-829.49" */
  /* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _00104_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:829.23-829.49" */
  /* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _00105_;
  /* src = "generated/out/vanilla.sv:833.24-833.50" */
  /* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _00106_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:833.24-833.50" */
  /* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _00107_;
  /* src = "generated/out/vanilla.sv:1137.39-1137.56" */
  wire [31:0] _00108_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1137.39-1137.56" */
  wire [31:0] _00109_;
  /* src = "generated/out/vanilla.sv:1280.53-1280.95" */
  wire [31:0] _00110_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1280.53-1280.95" */
  wire [31:0] _00111_;
  /* src = "generated/out/vanilla.sv:472.18-472.51" */
  wire [3:0] _00112_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:472.18-472.51" */
  wire [3:0] _00113_;
  wire [31:0] _00114_;
  wire [31:0] _00115_;
  wire [63:0] _00116_;
  wire [31:0] _00117_;
  wire [63:0] _00118_;
  wire [63:0] _00119_;
  wire [29:0] _00120_;
  wire [31:0] _00121_;
  wire [31:0] _00122_;
  wire [31:0] _00123_;
  wire [31:0] _00124_;
  wire [31:0] _00125_;
  wire [63:0] _00126_;
  wire [29:0] _00127_;
  wire [31:0] _00128_;
  wire [31:0] _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire [1:0] _00226_;
  wire [1:0] _00227_;
  wire [1:0] _00228_;
  wire [2:0] _00229_;
  wire [3:0] _00230_;
  wire [2:0] _00231_;
  wire [2:0] _00232_;
  wire [3:0] _00233_;
  wire [1:0] _00234_;
  wire [1:0] _00235_;
  wire [2:0] _00236_;
  wire [1:0] _00237_;
  wire [2:0] _00238_;
  wire [1:0] _00239_;
  wire [7:0] _00240_;
  wire [3:0] _00241_;
  wire [3:0] _00242_;
  wire [3:0] _00243_;
  wire [5:0] _00244_;
  wire [2:0] _00245_;
  wire [5:0] _00246_;
  wire [3:0] _00247_;
  wire [1:0] _00248_;
  wire [1:0] _00249_;
  wire [5:0] _00250_;
  wire [5:0] _00251_;
  wire [1:0] _00252_;
  wire [31:0] _00253_;
  wire [6:0] _00254_;
  wire [1:0] _00255_;
  wire [11:0] _00256_;
  wire [1:0] _00257_;
  wire [1:0] _00258_;
  wire [6:0] _00259_;
  wire [4:0] _00260_;
  wire [2:0] _00261_;
  wire [11:0] _00262_;
  wire [6:0] _00263_;
  wire [15:0] _00264_;
  wire [2:0] _00265_;
  wire [6:0] _00266_;
  wire [1:0] _00267_;
  wire [7:0] _00268_;
  wire [2:0] _00269_;
  wire [1:0] _00270_;
  wire [1:0] _00271_;
  wire [1:0] _00272_;
  wire [30:0] _00273_;
  wire _00274_;
  wire [4:0] _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire [2:0] _00335_;
  wire [4:0] _00336_;
  wire [1:0] _00337_;
  wire [3:0] _00338_;
  wire [1:0] _00339_;
  wire [1:0] _00340_;
  wire [1:0] _00341_;
  wire [1:0] _00342_;
  wire [4:0] _00343_;
  wire [1:0] _00344_;
  wire [3:0] _00345_;
  wire [2:0] _00346_;
  wire [1:0] _00347_;
  wire [1:0] _00348_;
  wire [1:0] _00349_;
  wire [6:0] _00350_;
  wire [1:0] _00351_;
  wire [1:0] _00352_;
  wire [1:0] _00353_;
  wire [4:0] _00354_;
  wire [4:0] _00355_;
  wire [1:0] _00356_;
  wire [5:0] _00357_;
  wire [1:0] _00358_;
  wire [1:0] _00359_;
  wire [7:0] _00360_;
  wire [4:0] _00361_;
  wire [1:0] _00362_;
  wire [1:0] _00363_;
  wire [2:0] _00364_;
  wire [1:0] _00365_;
  wire [3:0] _00366_;
  wire [3:0] _00367_;
  wire [2:0] _00368_;
  wire [4:0] _00369_;
  wire [4:0] _00370_;
  wire [2:0] _00371_;
  wire [4:0] _00372_;
  wire [3:0] _00373_;
  wire [47:0] _00374_;
  wire [10:0] _00375_;
  wire [12:0] _00376_;
  wire [3:0] _00377_;
  wire [1:0] _00378_;
  wire [4:0] _00379_;
  wire [4:0] _00380_;
  wire [3:0] _00381_;
  wire [1:0] _00382_;
  wire [3:0] _00383_;
  wire [2:0] _00384_;
  wire [2:0] _00385_;
  wire [2:0] _00386_;
  wire [4:0] _00387_;
  wire [7:0] _00388_;
  wire [5:0] _00389_;
  wire [2:0] _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire [30:0] _00511_;
  wire _00512_;
  wire [30:0] _00513_;
  wire _00514_;
  wire [4:0] _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire [31:0] _00519_;
  wire [31:0] _00520_;
  wire [31:0] _00521_;
  wire [31:0] _00522_;
  wire [31:0] _00523_;
  wire [31:0] _00524_;
  wire [31:0] _00525_;
  wire [31:0] _00526_;
  wire [31:0] _00527_;
  wire [31:0] _00528_;
  wire [4:0] _00529_;
  wire [4:0] _00530_;
  wire [4:0] _00531_;
  wire [4:0] _00532_;
  wire [4:0] _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire [7:0] _00539_;
  wire [7:0] _00540_;
  wire [7:0] _00541_;
  wire [7:0] _00542_;
  wire [7:0] _00543_;
  wire [7:0] _00544_;
  wire [7:0] _00545_;
  wire [7:0] _00546_;
  wire [7:0] _00547_;
  wire [7:0] _00548_;
  wire [7:0] _00549_;
  wire [7:0] _00550_;
  wire [31:0] _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire [1:0] _00561_;
  wire [1:0] _00562_;
  wire [1:0] _00563_;
  wire [31:0] _00564_;
  wire [31:0] _00565_;
  wire [31:0] _00566_;
  wire [31:0] _00567_;
  wire [31:0] _00568_;
  wire [31:0] _00569_;
  wire [31:0] _00570_;
  wire [31:0] _00571_;
  wire [31:0] _00572_;
  wire [31:0] _00573_;
  wire [31:0] _00574_;
  wire [31:0] _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire [3:0] _00589_;
  wire [3:0] _00590_;
  wire [3:0] _00591_;
  wire [3:0] _00592_;
  wire [3:0] _00593_;
  wire [3:0] _00594_;
  wire [3:0] _00595_;
  wire [3:0] _00596_;
  wire [3:0] _00597_;
  wire [3:0] _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire [31:0] _00602_;
  wire [31:0] _00603_;
  wire [31:0] _00604_;
  wire [31:0] _00605_;
  wire [31:0] _00606_;
  wire [4:0] _00607_;
  wire [4:0] _00608_;
  wire [4:0] _00609_;
  wire [4:0] _00610_;
  wire [4:0] _00611_;
  wire [4:0] _00612_;
  wire [4:0] _00613_;
  wire [4:0] _00614_;
  wire [4:0] _00615_;
  wire [4:0] _00616_;
  wire [1:0] _00617_;
  wire [1:0] _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire [4:0] _00624_;
  wire [2:0] _00625_;
  wire [2:0] _00626_;
  wire [2:0] _00627_;
  wire [2:0] _00628_;
  wire [2:0] _00629_;
  wire [2:0] _00630_;
  wire [2:0] _00631_;
  wire [2:0] _00632_;
  wire [2:0] _00633_;
  wire [5:0] _00634_;
  wire [5:0] _00635_;
  wire [5:0] _00636_;
  wire [5:0] _00637_;
  wire [5:0] _00638_;
  wire [5:0] _00639_;
  wire [5:0] _00640_;
  wire [5:0] _00641_;
  wire [5:0] _00642_;
  wire [5:0] _00643_;
  wire [5:0] _00644_;
  wire [5:0] _00645_;
  wire [31:0] _00646_;
  wire [31:0] _00647_;
  wire [31:0] _00648_;
  wire [31:0] _00649_;
  wire [31:0] _00650_;
  wire [31:0] _00651_;
  wire [3:0] _00652_;
  wire [31:0] _00653_;
  wire _00654_;
  wire [31:0] _00655_;
  wire [31:0] _00656_;
  wire [31:0] _00657_;
  wire [31:0] _00658_;
  wire [31:0] _00659_;
  wire [31:0] _00660_;
  wire [31:0] _00661_;
  wire [31:0] _00662_;
  wire [31:0] _00663_;
  wire [31:0] _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire [31:0] _00668_;
  wire [31:0] _00669_;
  wire _00670_;
  wire _00671_;
  wire [31:0] _00672_;
  wire [4:0] _00673_;
  wire [4:0] _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire [7:0] _00678_;
  wire [7:0] _00679_;
  wire [7:0] _00680_;
  wire [7:0] _00681_;
  wire [7:0] _00682_;
  wire [7:0] _00683_;
  wire [7:0] _00684_;
  wire [7:0] _00685_;
  wire [7:0] _00686_;
  wire [7:0] _00687_;
  wire [31:0] _00688_;
  wire [31:0] _00689_;
  wire [31:0] _00690_;
  wire _00691_;
  wire [1:0] _00692_;
  wire [1:0] _00693_;
  wire [31:0] _00694_;
  wire [31:0] _00695_;
  wire [31:0] _00696_;
  wire [31:0] _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire [2:0] _00712_;
  wire [1:0] _00713_;
  wire [11:0] _00714_;
  wire [3:0] _00715_;
  wire [3:0] _00716_;
  wire [3:0] _00717_;
  wire [3:0] _00718_;
  wire [3:0] _00719_;
  wire [3:0] _00720_;
  wire [3:0] _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire [4:0] _00725_;
  wire [4:0] _00726_;
  wire [4:0] _00727_;
  wire [4:0] _00728_;
  wire [7:0] _00729_;
  wire [4:0] _00730_;
  wire [4:0] _00731_;
  wire _00732_;
  wire [4:0] _00733_;
  wire [31:0] _00734_;
  wire [4:0] _00735_;
  wire [31:0] _00736_;
  wire [31:0] _00737_;
  wire [15:0] _00738_;
  wire [15:0] _00739_;
  wire [15:0] _00740_;
  wire [1:0] _00741_;
  wire [1:0] _00742_;
  wire [3:0] _00743_;
  wire [3:0] _00744_;
  wire [3:0] _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire [4:0] _00750_;
  wire [4:0] _00751_;
  wire [4:0] _00752_;
  wire [4:0] _00753_;
  wire [4:0] _00754_;
  wire [4:0] _00755_;
  wire [2:0] _00756_;
  wire [2:0] _00757_;
  wire [2:0] _00758_;
  wire [2:0] _00759_;
  wire [2:0] _00760_;
  wire [2:0] _00761_;
  wire [2:0] _00762_;
  wire [2:0] _00763_;
  wire [2:0] _00764_;
  wire [2:0] _00765_;
  wire [2:0] _00766_;
  wire [2:0] _00767_;
  wire [2:0] _00768_;
  wire [2:0] _00769_;
  wire [2:0] _00770_;
  wire [3:0] _00771_;
  wire [3:0] _00772_;
  wire [5:0] _00773_;
  wire [5:0] _00774_;
  wire [5:0] _00775_;
  wire [5:0] _00776_;
  wire [5:0] _00777_;
  wire [5:0] _00778_;
  wire [5:0] _00779_;
  wire [5:0] _00780_;
  wire [5:0] _00781_;
  wire [5:0] _00782_;
  wire [5:0] _00783_;
  wire _00784_;
  wire [63:0] _00785_;
  wire [63:0] _00786_;
  wire [31:0] _00787_;
  wire [31:0] _00788_;
  wire [31:0] _00789_;
  wire [31:0] _00790_;
  wire [31:0] _00791_;
  wire [31:0] _00792_;
  wire [31:0] _00793_;
  wire [31:0] _00794_;
  wire [31:0] _00795_;
  wire [31:0] _00796_;
  /* cellift = 32'd1 */
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire [3:0] _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire [1:0] _00831_;
  wire [1:0] _00832_;
  wire [2:0] _00833_;
  wire _00834_;
  wire [1:0] _00835_;
  wire [2:0] _00836_;
  wire _00837_;
  wire _00838_;
  wire [31:0] _00839_;
  wire [31:0] _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire [31:0] _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire [31:0] _00854_;
  wire _00855_;
  /* cellift = 32'd1 */
  wire _00856_;
  wire _00857_;
  /* cellift = 32'd1 */
  wire _00858_;
  wire _00859_;
  /* cellift = 32'd1 */
  wire _00860_;
  wire _00861_;
  /* cellift = 32'd1 */
  wire _00862_;
  wire _00863_;
  /* cellift = 32'd1 */
  wire _00864_;
  wire _00865_;
  /* cellift = 32'd1 */
  wire _00866_;
  wire _00867_;
  /* cellift = 32'd1 */
  wire _00868_;
  wire _00869_;
  /* cellift = 32'd1 */
  wire _00870_;
  wire _00871_;
  /* cellift = 32'd1 */
  wire _00872_;
  wire _00873_;
  /* cellift = 32'd1 */
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire [31:0] _00935_;
  wire [31:0] _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  /* cellift = 32'd1 */
  wire _00944_;
  wire _00945_;
  /* cellift = 32'd1 */
  wire _00946_;
  wire _00947_;
  /* cellift = 32'd1 */
  wire _00948_;
  wire _00949_;
  /* cellift = 32'd1 */
  wire _00950_;
  wire _00951_;
  /* cellift = 32'd1 */
  wire _00952_;
  wire _00953_;
  /* cellift = 32'd1 */
  wire _00954_;
  wire _00955_;
  /* cellift = 32'd1 */
  wire _00956_;
  wire _00957_;
  /* cellift = 32'd1 */
  wire _00958_;
  wire _00959_;
  /* cellift = 32'd1 */
  wire _00960_;
  wire _00961_;
  /* cellift = 32'd1 */
  wire _00962_;
  wire _00963_;
  /* cellift = 32'd1 */
  wire _00964_;
  wire _00965_;
  /* cellift = 32'd1 */
  wire _00966_;
  wire _00967_;
  /* cellift = 32'd1 */
  wire _00968_;
  wire _00969_;
  /* cellift = 32'd1 */
  wire _00970_;
  wire _00971_;
  /* cellift = 32'd1 */
  wire _00972_;
  wire _00973_;
  /* cellift = 32'd1 */
  wire _00974_;
  wire _00975_;
  /* cellift = 32'd1 */
  wire _00976_;
  wire _00977_;
  /* cellift = 32'd1 */
  wire _00978_;
  wire _00979_;
  /* cellift = 32'd1 */
  wire _00980_;
  wire _00981_;
  /* cellift = 32'd1 */
  wire _00982_;
  wire _00983_;
  /* cellift = 32'd1 */
  wire _00984_;
  wire _00985_;
  /* cellift = 32'd1 */
  wire _00986_;
  wire _00987_;
  /* cellift = 32'd1 */
  wire _00988_;
  wire _00989_;
  /* cellift = 32'd1 */
  wire _00990_;
  wire _00991_;
  /* cellift = 32'd1 */
  wire _00992_;
  wire _00993_;
  /* cellift = 32'd1 */
  wire _00994_;
  wire _00995_;
  /* cellift = 32'd1 */
  wire _00996_;
  wire _00997_;
  /* cellift = 32'd1 */
  wire _00998_;
  wire _00999_;
  /* cellift = 32'd1 */
  wire _01000_;
  wire _01001_;
  /* cellift = 32'd1 */
  wire _01002_;
  wire _01003_;
  /* cellift = 32'd1 */
  wire _01004_;
  wire _01005_;
  /* cellift = 32'd1 */
  wire _01006_;
  wire _01007_;
  /* cellift = 32'd1 */
  wire _01008_;
  wire _01009_;
  /* cellift = 32'd1 */
  wire _01010_;
  wire _01011_;
  /* cellift = 32'd1 */
  wire _01012_;
  wire _01013_;
  /* cellift = 32'd1 */
  wire _01014_;
  wire _01015_;
  /* cellift = 32'd1 */
  wire _01016_;
  wire _01017_;
  /* cellift = 32'd1 */
  wire _01018_;
  wire _01019_;
  /* cellift = 32'd1 */
  wire _01020_;
  wire _01021_;
  /* cellift = 32'd1 */
  wire _01022_;
  wire _01023_;
  /* cellift = 32'd1 */
  wire _01024_;
  wire _01025_;
  /* cellift = 32'd1 */
  wire _01026_;
  wire _01027_;
  /* cellift = 32'd1 */
  wire _01028_;
  wire _01029_;
  /* cellift = 32'd1 */
  wire _01030_;
  wire _01031_;
  /* cellift = 32'd1 */
  wire _01032_;
  wire _01033_;
  /* cellift = 32'd1 */
  wire _01034_;
  wire _01035_;
  /* cellift = 32'd1 */
  wire _01036_;
  wire _01037_;
  /* cellift = 32'd1 */
  wire _01038_;
  wire _01039_;
  /* cellift = 32'd1 */
  wire _01040_;
  wire _01041_;
  /* cellift = 32'd1 */
  wire _01042_;
  wire _01043_;
  /* cellift = 32'd1 */
  wire _01044_;
  wire _01045_;
  /* cellift = 32'd1 */
  wire _01046_;
  wire _01047_;
  /* cellift = 32'd1 */
  wire _01048_;
  wire _01049_;
  /* cellift = 32'd1 */
  wire _01050_;
  wire _01051_;
  /* cellift = 32'd1 */
  wire _01052_;
  wire _01053_;
  /* cellift = 32'd1 */
  wire _01054_;
  wire _01055_;
  /* cellift = 32'd1 */
  wire _01056_;
  wire _01057_;
  /* cellift = 32'd1 */
  wire _01058_;
  wire _01059_;
  /* cellift = 32'd1 */
  wire _01060_;
  wire _01061_;
  /* cellift = 32'd1 */
  wire _01062_;
  wire _01063_;
  /* cellift = 32'd1 */
  wire _01064_;
  wire _01065_;
  /* cellift = 32'd1 */
  wire _01066_;
  wire _01067_;
  /* cellift = 32'd1 */
  wire _01068_;
  wire _01069_;
  /* cellift = 32'd1 */
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  /* cellift = 32'd1 */
  wire _01077_;
  wire _01078_;
  /* cellift = 32'd1 */
  wire _01079_;
  wire _01080_;
  /* cellift = 32'd1 */
  wire _01081_;
  wire _01082_;
  /* cellift = 32'd1 */
  wire _01083_;
  wire _01084_;
  /* cellift = 32'd1 */
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  /* cellift = 32'd1 */
  wire _01089_;
  wire _01090_;
  /* cellift = 32'd1 */
  wire _01091_;
  wire _01092_;
  /* cellift = 32'd1 */
  wire _01093_;
  wire _01094_;
  wire _01095_;
  /* cellift = 32'd1 */
  wire _01096_;
  wire _01097_;
  /* cellift = 32'd1 */
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire [31:0] _01140_;
  wire [31:0] _01141_;
  wire [31:0] _01142_;
  wire [3:0] _01143_;
  wire [3:0] _01144_;
  wire [3:0] _01145_;
  wire [4:0] _01146_;
  wire [4:0] _01147_;
  wire [4:0] _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire [31:0] _01167_;
  wire [31:0] _01168_;
  wire [31:0] _01169_;
  wire [31:0] _01170_;
  wire [31:0] _01171_;
  wire [31:0] _01172_;
  wire [3:0] _01173_;
  wire [3:0] _01174_;
  wire [3:0] _01175_;
  wire [3:0] _01176_;
  wire [3:0] _01177_;
  wire [3:0] _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire [31:0] _01186_;
  wire [31:0] _01187_;
  wire [31:0] _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire [30:0] _01192_;
  wire [30:0] _01193_;
  wire [30:0] _01194_;
  wire [31:0] _01195_;
  wire [31:0] _01196_;
  wire [31:0] _01197_;
  wire [1:0] _01198_;
  wire [1:0] _01199_;
  wire [1:0] _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire [31:0] _01204_;
  wire [31:0] _01205_;
  wire [31:0] _01206_;
  wire [31:0] _01207_;
  wire [31:0] _01208_;
  wire [31:0] _01209_;
  wire [4:0] _01210_;
  wire [4:0] _01211_;
  wire [4:0] _01212_;
  wire [7:0] _01213_;
  wire [7:0] _01214_;
  wire [7:0] _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire [63:0] _01219_;
  wire [63:0] _01220_;
  wire [63:0] _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire [30:0] _01228_;
  wire [30:0] _01229_;
  wire [30:0] _01230_;
  wire [31:0] _01231_;
  wire [31:0] _01232_;
  wire [31:0] _01233_;
  wire [31:0] _01234_;
  wire [31:0] _01235_;
  wire [31:0] _01236_;
  wire [31:0] _01237_;
  wire [31:0] _01238_;
  wire [31:0] _01239_;
  wire [31:0] _01240_;
  wire [31:0] _01241_;
  wire [31:0] _01242_;
  wire [31:0] _01243_;
  wire [31:0] _01244_;
  wire [31:0] _01245_;
  wire [31:0] _01246_;
  wire [31:0] _01247_;
  wire [31:0] _01248_;
  wire [31:0] _01249_;
  wire [31:0] _01250_;
  wire [31:0] _01251_;
  wire [31:0] _01252_;
  wire [31:0] _01253_;
  wire [31:0] _01254_;
  wire [31:0] _01255_;
  wire [31:0] _01256_;
  wire [31:0] _01257_;
  wire [31:0] _01258_;
  wire [31:0] _01259_;
  wire [31:0] _01260_;
  wire [31:0] _01261_;
  wire [31:0] _01262_;
  wire [31:0] _01263_;
  wire [31:0] _01264_;
  wire [31:0] _01265_;
  wire [31:0] _01266_;
  wire [31:0] _01267_;
  wire [31:0] _01268_;
  wire [31:0] _01269_;
  wire [31:0] _01270_;
  wire [31:0] _01271_;
  wire [31:0] _01272_;
  wire [31:0] _01273_;
  wire [31:0] _01274_;
  wire [31:0] _01275_;
  wire [31:0] _01276_;
  wire [31:0] _01277_;
  wire [31:0] _01278_;
  wire [31:0] _01279_;
  wire [31:0] _01280_;
  wire [31:0] _01281_;
  wire [31:0] _01282_;
  wire [31:0] _01283_;
  wire [31:0] _01284_;
  wire [31:0] _01285_;
  wire [31:0] _01286_;
  wire [31:0] _01287_;
  wire [31:0] _01288_;
  wire [31:0] _01289_;
  wire [31:0] _01290_;
  wire [31:0] _01291_;
  wire [31:0] _01292_;
  wire [31:0] _01293_;
  wire [31:0] _01294_;
  wire [31:0] _01295_;
  wire [31:0] _01296_;
  wire [31:0] _01297_;
  wire [31:0] _01298_;
  wire [31:0] _01299_;
  wire [31:0] _01300_;
  wire [31:0] _01301_;
  wire [31:0] _01302_;
  wire [31:0] _01303_;
  wire [31:0] _01304_;
  wire [31:0] _01305_;
  wire [31:0] _01306_;
  wire [31:0] _01307_;
  wire [31:0] _01308_;
  wire [31:0] _01309_;
  wire [31:0] _01310_;
  wire [31:0] _01311_;
  wire [31:0] _01312_;
  wire [31:0] _01313_;
  wire [31:0] _01314_;
  wire [31:0] _01315_;
  wire [31:0] _01316_;
  wire [31:0] _01317_;
  wire [31:0] _01318_;
  wire [31:0] _01319_;
  wire [31:0] _01320_;
  wire [31:0] _01321_;
  wire [31:0] _01322_;
  wire [31:0] _01323_;
  wire [31:0] _01324_;
  wire [31:0] _01325_;
  wire [31:0] _01326_;
  wire [4:0] _01327_;
  wire [4:0] _01328_;
  wire [4:0] _01329_;
  wire [4:0] _01330_;
  wire [4:0] _01331_;
  wire [4:0] _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire [2:0] _01455_;
  wire [1:0] _01456_;
  wire [1:0] _01457_;
  wire [1:0] _01458_;
  wire [2:0] _01459_;
  wire [3:0] _01460_;
  wire [2:0] _01461_;
  wire [2:0] _01462_;
  wire [3:0] _01463_;
  wire [4:0] _01464_;
  wire [1:0] _01465_;
  wire [1:0] _01466_;
  wire [3:0] _01467_;
  wire [1:0] _01468_;
  wire [1:0] _01469_;
  wire [1:0] _01470_;
  wire [1:0] _01471_;
  wire [2:0] _01472_;
  wire [1:0] _01473_;
  wire [1:0] _01474_;
  wire [2:0] _01475_;
  wire [1:0] _01476_;
  wire [4:0] _01477_;
  wire [1:0] _01478_;
  wire [7:0] _01479_;
  wire [3:0] _01480_;
  wire [3:0] _01481_;
  wire [3:0] _01482_;
  wire [5:0] _01483_;
  wire [2:0] _01484_;
  wire [5:0] _01485_;
  wire [3:0] _01486_;
  wire [1:0] _01487_;
  wire [1:0] _01488_;
  wire [3:0] _01489_;
  wire [5:0] _01490_;
  wire [5:0] _01491_;
  wire [2:0] _01492_;
  wire [1:0] _01493_;
  wire [1:0] _01494_;
  wire [1:0] _01495_;
  wire [1:0] _01496_;
  wire [6:0] _01497_;
  wire [1:0] _01498_;
  wire [1:0] _01499_;
  wire [1:0] _01500_;
  wire [4:0] _01501_;
  wire [4:0] _01502_;
  wire [1:0] _01503_;
  wire [5:0] _01504_;
  wire [1:0] _01505_;
  wire [1:0] _01506_;
  wire [7:0] _01507_;
  wire [4:0] _01508_;
  wire [1:0] _01509_;
  wire [1:0] _01510_;
  wire [2:0] _01511_;
  wire [1:0] _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire [3:0] _01567_;
  wire [3:0] _01568_;
  wire [2:0] _01569_;
  wire [4:0] _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire [31:0] _01577_;
  wire [31:0] _01578_;
  wire [31:0] _01579_;
  wire [31:0] _01580_;
  wire [31:0] _01581_;
  wire [31:0] _01582_;
  wire [31:0] _01583_;
  wire [31:0] _01584_;
  wire [31:0] _01585_;
  wire [31:0] _01586_;
  wire [31:0] _01587_;
  wire [31:0] _01588_;
  wire [31:0] _01589_;
  wire [31:0] _01590_;
  wire [31:0] _01591_;
  wire [31:0] _01592_;
  wire [31:0] _01593_;
  wire [31:0] _01594_;
  wire [31:0] _01595_;
  wire [31:0] _01596_;
  wire [31:0] _01597_;
  wire [31:0] _01598_;
  wire [31:0] _01599_;
  wire [31:0] _01600_;
  wire [31:0] _01601_;
  wire [31:0] _01602_;
  wire [31:0] _01603_;
  wire [31:0] _01604_;
  wire [31:0] _01605_;
  wire [31:0] _01606_;
  wire [4:0] _01607_;
  wire [4:0] _01608_;
  wire [4:0] _01609_;
  wire [4:0] _01610_;
  wire [4:0] _01611_;
  wire [4:0] _01612_;
  wire [4:0] _01613_;
  wire [4:0] _01614_;
  wire [4:0] _01615_;
  wire [4:0] _01616_;
  wire [4:0] _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire [7:0] _01637_;
  wire [7:0] _01638_;
  wire [7:0] _01639_;
  wire [7:0] _01640_;
  wire [7:0] _01641_;
  wire [7:0] _01642_;
  wire [7:0] _01643_;
  wire [7:0] _01644_;
  wire [7:0] _01645_;
  wire [7:0] _01646_;
  wire [7:0] _01647_;
  wire [7:0] _01648_;
  wire [7:0] _01649_;
  wire [7:0] _01650_;
  wire [7:0] _01651_;
  wire [7:0] _01652_;
  wire [7:0] _01653_;
  wire [7:0] _01654_;
  wire [7:0] _01655_;
  wire [7:0] _01656_;
  wire [7:0] _01657_;
  wire [7:0] _01658_;
  wire [7:0] _01659_;
  wire [7:0] _01660_;
  wire [7:0] _01661_;
  wire [7:0] _01662_;
  wire [7:0] _01663_;
  wire [7:0] _01664_;
  wire [7:0] _01665_;
  wire [7:0] _01666_;
  wire [7:0] _01667_;
  wire [7:0] _01668_;
  wire [7:0] _01669_;
  wire [7:0] _01670_;
  wire [31:0] _01671_;
  wire [31:0] _01672_;
  wire [31:0] _01673_;
  wire [31:0] _01674_;
  wire [31:0] _01675_;
  wire [31:0] _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire [1:0] _01700_;
  wire [1:0] _01701_;
  wire [1:0] _01702_;
  wire [1:0] _01703_;
  wire [1:0] _01704_;
  wire [1:0] _01705_;
  wire [1:0] _01706_;
  wire [1:0] _01707_;
  wire [1:0] _01708_;
  wire [31:0] _01709_;
  wire [31:0] _01710_;
  wire [31:0] _01711_;
  wire [31:0] _01712_;
  wire [31:0] _01713_;
  wire [31:0] _01714_;
  wire [31:0] _01715_;
  wire [31:0] _01716_;
  wire [31:0] _01717_;
  wire [31:0] _01718_;
  wire [31:0] _01719_;
  wire [31:0] _01720_;
  wire [31:0] _01721_;
  wire [31:0] _01722_;
  wire [31:0] _01723_;
  wire [31:0] _01724_;
  wire [31:0] _01725_;
  wire [31:0] _01726_;
  wire [31:0] _01727_;
  wire [31:0] _01728_;
  wire [31:0] _01729_;
  wire [31:0] _01730_;
  wire [31:0] _01731_;
  wire [31:0] _01732_;
  wire [31:0] _01733_;
  wire [31:0] _01734_;
  wire [31:0] _01735_;
  wire [31:0] _01736_;
  wire [31:0] _01737_;
  wire [31:0] _01738_;
  wire [31:0] _01739_;
  wire [31:0] _01740_;
  wire [31:0] _01741_;
  wire [31:0] _01742_;
  wire [31:0] _01743_;
  wire [31:0] _01744_;
  wire [31:0] _01745_;
  wire [31:0] _01746_;
  wire [31:0] _01747_;
  wire [31:0] _01748_;
  wire [31:0] _01749_;
  wire [31:0] _01750_;
  wire [31:0] _01751_;
  wire [31:0] _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire [3:0] _01792_;
  wire [3:0] _01793_;
  wire [3:0] _01794_;
  wire [3:0] _01795_;
  wire [3:0] _01796_;
  wire [3:0] _01797_;
  wire [3:0] _01798_;
  wire [3:0] _01799_;
  wire [3:0] _01800_;
  wire [3:0] _01801_;
  wire [3:0] _01802_;
  wire [3:0] _01803_;
  wire [3:0] _01804_;
  wire [3:0] _01805_;
  wire [3:0] _01806_;
  wire [3:0] _01807_;
  wire [3:0] _01808_;
  wire [3:0] _01809_;
  wire [3:0] _01810_;
  wire [3:0] _01811_;
  wire [3:0] _01812_;
  wire [3:0] _01813_;
  wire [3:0] _01814_;
  wire [3:0] _01815_;
  wire [3:0] _01816_;
  wire [3:0] _01817_;
  wire [3:0] _01818_;
  wire [3:0] _01819_;
  wire [3:0] _01820_;
  wire [3:0] _01821_;
  wire [3:0] _01822_;
  wire [3:0] _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire [31:0] _01853_;
  wire [31:0] _01854_;
  wire [31:0] _01855_;
  wire [31:0] _01856_;
  wire [31:0] _01857_;
  wire [31:0] _01858_;
  wire [31:0] _01859_;
  wire [31:0] _01860_;
  wire [31:0] _01861_;
  wire [31:0] _01862_;
  wire [31:0] _01863_;
  wire [31:0] _01864_;
  wire [31:0] _01865_;
  wire [31:0] _01866_;
  wire [4:0] _01867_;
  wire [4:0] _01868_;
  wire [4:0] _01869_;
  wire [4:0] _01870_;
  wire [4:0] _01871_;
  wire [4:0] _01872_;
  wire [4:0] _01873_;
  wire [4:0] _01874_;
  wire [4:0] _01875_;
  wire [4:0] _01876_;
  wire [4:0] _01877_;
  wire [4:0] _01878_;
  wire [4:0] _01879_;
  wire [4:0] _01880_;
  wire [4:0] _01881_;
  wire [4:0] _01882_;
  wire [4:0] _01883_;
  wire [4:0] _01884_;
  wire [4:0] _01885_;
  wire [4:0] _01886_;
  wire [4:0] _01887_;
  wire [4:0] _01888_;
  wire [4:0] _01889_;
  wire [4:0] _01890_;
  wire [4:0] _01891_;
  wire [4:0] _01892_;
  wire [4:0] _01893_;
  wire [4:0] _01894_;
  wire [4:0] _01895_;
  wire [4:0] _01896_;
  wire [4:0] _01897_;
  wire [4:0] _01898_;
  wire [4:0] _01899_;
  wire [4:0] _01900_;
  wire [4:0] _01901_;
  wire [4:0] _01902_;
  wire [4:0] _01903_;
  wire [4:0] _01904_;
  wire [4:0] _01905_;
  wire [4:0] _01906_;
  wire [4:0] _01907_;
  wire [1:0] _01908_;
  wire [1:0] _01909_;
  wire [1:0] _01910_;
  wire [1:0] _01911_;
  wire [1:0] _01912_;
  wire [1:0] _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire [4:0] _01944_;
  wire [4:0] _01945_;
  wire [4:0] _01946_;
  wire [4:0] _01947_;
  wire [4:0] _01948_;
  wire [4:0] _01949_;
  wire [4:0] _01950_;
  wire [4:0] _01951_;
  wire [4:0] _01952_;
  wire [4:0] _01953_;
  wire [4:0] _01954_;
  wire [4:0] _01955_;
  wire [4:0] _01956_;
  wire [4:0] _01957_;
  wire [4:0] _01958_;
  wire [4:0] _01959_;
  wire [4:0] _01960_;
  wire [4:0] _01961_;
  wire [4:0] _01962_;
  wire [4:0] _01963_;
  wire [4:0] _01964_;
  wire [4:0] _01965_;
  wire [4:0] _01966_;
  wire [4:0] _01967_;
  wire [4:0] _01968_;
  wire [4:0] _01969_;
  wire [4:0] _01970_;
  wire [4:0] _01971_;
  wire [4:0] _01972_;
  wire [4:0] _01973_;
  wire [2:0] _01974_;
  wire [2:0] _01975_;
  wire [2:0] _01976_;
  wire [2:0] _01977_;
  wire [2:0] _01978_;
  wire [2:0] _01979_;
  wire [2:0] _01980_;
  wire [2:0] _01981_;
  wire [2:0] _01982_;
  wire [2:0] _01983_;
  wire [2:0] _01984_;
  wire [2:0] _01985_;
  wire [2:0] _01986_;
  wire [2:0] _01987_;
  wire [2:0] _01988_;
  wire [2:0] _01989_;
  wire [2:0] _01990_;
  wire [2:0] _01991_;
  wire [2:0] _01992_;
  wire [2:0] _01993_;
  wire [2:0] _01994_;
  wire [2:0] _01995_;
  wire [2:0] _01996_;
  wire [2:0] _01997_;
  wire [2:0] _01998_;
  wire [2:0] _01999_;
  wire [2:0] _02000_;
  wire [2:0] _02001_;
  wire [3:0] _02002_;
  wire [3:0] _02003_;
  wire [3:0] _02004_;
  wire [3:0] _02005_;
  wire [3:0] _02006_;
  wire [3:0] _02007_;
  wire [3:0] _02008_;
  wire [3:0] _02009_;
  wire [3:0] _02010_;
  wire [5:0] _02011_;
  wire [5:0] _02012_;
  wire [5:0] _02013_;
  wire [5:0] _02014_;
  wire [5:0] _02015_;
  wire [5:0] _02016_;
  wire [5:0] _02017_;
  wire [5:0] _02018_;
  wire [5:0] _02019_;
  wire [5:0] _02020_;
  wire [5:0] _02021_;
  wire [5:0] _02022_;
  wire [5:0] _02023_;
  wire [5:0] _02024_;
  wire [5:0] _02025_;
  wire [5:0] _02026_;
  wire [5:0] _02027_;
  wire [5:0] _02028_;
  wire [5:0] _02029_;
  wire [5:0] _02030_;
  wire [5:0] _02031_;
  wire [5:0] _02032_;
  wire [5:0] _02033_;
  wire [5:0] _02034_;
  wire [5:0] _02035_;
  wire [5:0] _02036_;
  wire [5:0] _02037_;
  wire [5:0] _02038_;
  wire [5:0] _02039_;
  wire [5:0] _02040_;
  wire [5:0] _02041_;
  wire [5:0] _02042_;
  wire [5:0] _02043_;
  wire [5:0] _02044_;
  wire [5:0] _02045_;
  wire [5:0] _02046_;
  wire [5:0] _02047_;
  wire [31:0] _02048_;
  wire [31:0] _02049_;
  wire [31:0] _02050_;
  wire [31:0] _02051_;
  wire [31:0] _02052_;
  wire [31:0] _02053_;
  wire [31:0] _02054_;
  wire [31:0] _02055_;
  wire [31:0] _02056_;
  wire [31:0] _02057_;
  wire [31:0] _02058_;
  wire [31:0] _02059_;
  wire [31:0] _02060_;
  wire [31:0] _02061_;
  wire [31:0] _02062_;
  wire [31:0] _02063_;
  wire [31:0] _02064_;
  wire [31:0] _02065_;
  wire [3:0] _02066_;
  wire [3:0] _02067_;
  wire [3:0] _02068_;
  wire [3:0] _02069_;
  wire [3:0] _02070_;
  wire [31:0] _02071_;
  wire [31:0] _02072_;
  wire [31:0] _02073_;
  wire [31:0] _02074_;
  wire [31:0] _02075_;
  wire [31:0] _02076_;
  wire [31:0] _02077_;
  wire [31:0] _02078_;
  wire [31:0] _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire [31:0] _02085_;
  wire [31:0] _02086_;
  wire [4:0] _02087_;
  wire [6:0] _02088_;
  wire [1:0] _02089_;
  wire [11:0] _02090_;
  wire [1:0] _02091_;
  wire [1:0] _02092_;
  wire [6:0] _02093_;
  wire [2:0] _02094_;
  wire [4:0] _02095_;
  wire [2:0] _02096_;
  wire [4:0] _02097_;
  wire [11:0] _02098_;
  wire [6:0] _02099_;
  wire [15:0] _02100_;
  wire [2:0] _02101_;
  wire [6:0] _02102_;
  wire [30:0] _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire [4:0] _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire [3:0] _02409_;
  wire [47:0] _02410_;
  wire [10:0] _02411_;
  wire [12:0] _02412_;
  wire [3:0] _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire [30:0] _02493_;
  wire [30:0] _02494_;
  wire [31:0] _02495_;
  wire [31:0] _02496_;
  wire [31:0] _02497_;
  wire [31:0] _02498_;
  wire [31:0] _02499_;
  wire [31:0] _02500_;
  wire [31:0] _02501_;
  wire [31:0] _02502_;
  wire [31:0] _02503_;
  wire [31:0] _02504_;
  wire [31:0] _02505_;
  wire [31:0] _02506_;
  wire [31:0] _02507_;
  wire [31:0] _02508_;
  wire [31:0] _02509_;
  wire [31:0] _02510_;
  wire [31:0] _02511_;
  wire [31:0] _02512_;
  wire [31:0] _02513_;
  wire [31:0] _02514_;
  wire [31:0] _02515_;
  wire [31:0] _02516_;
  wire [31:0] _02517_;
  wire [31:0] _02518_;
  wire [31:0] _02519_;
  wire [31:0] _02520_;
  wire [31:0] _02521_;
  wire [31:0] _02522_;
  wire [31:0] _02523_;
  wire [31:0] _02524_;
  wire [31:0] _02525_;
  wire [31:0] _02526_;
  wire [31:0] _02527_;
  wire [31:0] _02528_;
  wire [31:0] _02529_;
  wire [31:0] _02530_;
  wire [31:0] _02531_;
  wire [31:0] _02532_;
  wire [31:0] _02533_;
  wire [31:0] _02534_;
  wire [31:0] _02535_;
  wire [31:0] _02536_;
  wire [31:0] _02537_;
  wire [31:0] _02538_;
  wire [31:0] _02539_;
  wire [31:0] _02540_;
  wire [31:0] _02541_;
  wire [31:0] _02542_;
  wire [31:0] _02543_;
  wire [31:0] _02544_;
  wire [31:0] _02545_;
  wire [31:0] _02546_;
  wire [31:0] _02547_;
  wire [31:0] _02548_;
  wire [31:0] _02549_;
  wire [31:0] _02550_;
  wire [31:0] _02551_;
  wire [31:0] _02552_;
  wire [31:0] _02553_;
  wire [31:0] _02554_;
  wire [31:0] _02555_;
  wire [31:0] _02556_;
  wire [31:0] _02557_;
  wire [31:0] _02558_;
  wire [31:0] _02559_;
  wire [31:0] _02560_;
  wire [31:0] _02561_;
  wire [31:0] _02562_;
  wire [31:0] _02563_;
  wire [31:0] _02564_;
  wire [31:0] _02565_;
  wire [31:0] _02566_;
  wire [31:0] _02567_;
  wire [31:0] _02568_;
  wire [31:0] _02569_;
  wire [31:0] _02570_;
  wire [31:0] _02571_;
  wire [31:0] _02572_;
  wire [31:0] _02573_;
  wire [31:0] _02574_;
  wire [31:0] _02575_;
  wire [31:0] _02576_;
  wire [31:0] _02577_;
  wire [31:0] _02578_;
  wire [31:0] _02579_;
  wire [31:0] _02580_;
  wire [31:0] _02581_;
  wire [31:0] _02582_;
  wire [31:0] _02583_;
  wire [31:0] _02584_;
  wire [31:0] _02585_;
  wire [31:0] _02586_;
  wire [31:0] _02587_;
  wire [31:0] _02588_;
  wire [31:0] _02589_;
  wire [31:0] _02590_;
  wire [31:0] _02591_;
  wire [31:0] _02592_;
  wire [31:0] _02593_;
  wire [31:0] _02594_;
  wire [31:0] _02595_;
  wire [31:0] _02596_;
  wire [31:0] _02597_;
  wire [31:0] _02598_;
  wire [31:0] _02599_;
  wire [31:0] _02600_;
  wire [31:0] _02601_;
  wire [31:0] _02602_;
  wire [31:0] _02603_;
  wire [31:0] _02604_;
  wire [31:0] _02605_;
  wire [31:0] _02606_;
  wire [31:0] _02607_;
  wire [31:0] _02608_;
  wire [31:0] _02609_;
  wire [31:0] _02610_;
  wire [31:0] _02611_;
  wire [31:0] _02612_;
  wire [31:0] _02613_;
  wire [31:0] _02614_;
  wire [31:0] _02615_;
  wire [31:0] _02616_;
  wire [31:0] _02617_;
  wire [31:0] _02618_;
  wire [31:0] _02619_;
  wire [31:0] _02620_;
  wire [31:0] _02621_;
  wire [31:0] _02622_;
  wire [31:0] _02623_;
  wire [31:0] _02624_;
  wire [31:0] _02625_;
  wire [31:0] _02626_;
  wire [31:0] _02627_;
  wire [31:0] _02628_;
  wire [31:0] _02629_;
  wire [31:0] _02630_;
  wire [31:0] _02631_;
  wire [31:0] _02632_;
  wire [31:0] _02633_;
  wire [31:0] _02634_;
  wire [31:0] _02635_;
  wire [31:0] _02636_;
  wire [31:0] _02637_;
  wire [31:0] _02638_;
  wire [31:0] _02639_;
  wire [31:0] _02640_;
  wire [31:0] _02641_;
  wire [31:0] _02642_;
  wire [31:0] _02643_;
  wire [31:0] _02644_;
  wire [31:0] _02645_;
  wire [31:0] _02646_;
  wire [31:0] _02647_;
  wire [31:0] _02648_;
  wire [31:0] _02649_;
  wire [31:0] _02650_;
  wire [31:0] _02651_;
  wire [31:0] _02652_;
  wire [31:0] _02653_;
  wire [31:0] _02654_;
  wire [31:0] _02655_;
  wire [31:0] _02656_;
  wire [31:0] _02657_;
  wire [31:0] _02658_;
  wire [31:0] _02659_;
  wire [31:0] _02660_;
  wire [31:0] _02661_;
  wire [31:0] _02662_;
  wire [31:0] _02663_;
  wire [31:0] _02664_;
  wire [31:0] _02665_;
  wire [31:0] _02666_;
  wire [31:0] _02667_;
  wire [31:0] _02668_;
  wire [31:0] _02669_;
  wire [31:0] _02670_;
  wire [31:0] _02671_;
  wire [31:0] _02672_;
  wire [31:0] _02673_;
  wire [31:0] _02674_;
  wire [31:0] _02675_;
  wire [31:0] _02676_;
  wire [31:0] _02677_;
  wire [31:0] _02678_;
  wire [31:0] _02679_;
  wire [31:0] _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire [1:0] _02777_;
  wire [1:0] _02778_;
  wire [1:0] _02779_;
  wire [31:0] _02780_;
  wire [31:0] _02781_;
  wire [31:0] _02782_;
  wire [63:0] _02783_;
  wire [63:0] _02784_;
  wire [63:0] _02785_;
  wire [63:0] _02786_;
  wire [63:0] _02787_;
  wire [63:0] _02788_;
  wire [63:0] _02789_;
  wire [63:0] _02790_;
  wire [31:0] _02791_;
  wire [31:0] _02792_;
  wire [4:0] _02793_;
  wire [4:0] _02794_;
  wire _02795_;
  wire [31:0] _02796_;
  wire [31:0] _02797_;
  wire [31:0] _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire [4:0] _02811_;
  wire [4:0] _02812_;
  wire [4:0] _02813_;
  wire [7:0] _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire [7:0] _02823_;
  wire [7:0] _02824_;
  wire [7:0] _02825_;
  wire [7:0] _02826_;
  wire [7:0] _02827_;
  wire [7:0] _02828_;
  wire [7:0] _02829_;
  wire [7:0] _02830_;
  wire [7:0] _02831_;
  wire [7:0] _02832_;
  wire [7:0] _02833_;
  wire [7:0] _02834_;
  wire [7:0] _02835_;
  wire [7:0] _02836_;
  wire [7:0] _02837_;
  wire [7:0] _02838_;
  wire [7:0] _02839_;
  wire [7:0] _02840_;
  wire [7:0] _02841_;
  wire [7:0] _02842_;
  wire [7:0] _02843_;
  wire [7:0] _02844_;
  wire [7:0] _02845_;
  wire [7:0] _02846_;
  wire [7:0] _02847_;
  wire [7:0] _02848_;
  wire [7:0] _02849_;
  wire [31:0] _02850_;
  wire [31:0] _02851_;
  wire [31:0] _02852_;
  wire [31:0] _02853_;
  wire [31:0] _02854_;
  wire [31:0] _02855_;
  wire [31:0] _02856_;
  wire [31:0] _02857_;
  wire [31:0] _02858_;
  wire [31:0] _02859_;
  wire [31:0] _02860_;
  wire [31:0] _02861_;
  wire [31:0] _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire [31:0] _02869_;
  wire [31:0] _02870_;
  wire [31:0] _02871_;
  wire [31:0] _02872_;
  wire [31:0] _02873_;
  wire [31:0] _02874_;
  wire [31:0] _02875_;
  wire [31:0] _02876_;
  wire [31:0] _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire [2:0] _02924_;
  wire [2:0] _02925_;
  wire [2:0] _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire [1:0] _02930_;
  wire [1:0] _02931_;
  wire [1:0] _02932_;
  wire [11:0] _02933_;
  wire [11:0] _02934_;
  wire [11:0] _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire [3:0] _02942_;
  wire [3:0] _02943_;
  wire [3:0] _02944_;
  wire [3:0] _02945_;
  wire [3:0] _02946_;
  wire [3:0] _02947_;
  wire [3:0] _02948_;
  wire [3:0] _02949_;
  wire [3:0] _02950_;
  wire [3:0] _02951_;
  wire [3:0] _02952_;
  wire [3:0] _02953_;
  wire [3:0] _02954_;
  wire [3:0] _02955_;
  wire [3:0] _02956_;
  wire [3:0] _02957_;
  wire [3:0] _02958_;
  wire [3:0] _02959_;
  wire [3:0] _02960_;
  wire [3:0] _02961_;
  wire [3:0] _02962_;
  wire [3:0] _02963_;
  wire [3:0] _02964_;
  wire [3:0] _02965_;
  wire [3:0] _02966_;
  wire [3:0] _02967_;
  wire [3:0] _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire [4:0] _03027_;
  wire [4:0] _03028_;
  wire [4:0] _03029_;
  wire [4:0] _03030_;
  wire [4:0] _03031_;
  wire [4:0] _03032_;
  wire [4:0] _03033_;
  wire [4:0] _03034_;
  wire [4:0] _03035_;
  wire [4:0] _03036_;
  wire [4:0] _03037_;
  wire [4:0] _03038_;
  wire [4:0] _03039_;
  wire [4:0] _03040_;
  wire [4:0] _03041_;
  wire [4:0] _03042_;
  wire [2:0] _03043_;
  wire [4:0] _03044_;
  wire [4:0] _03045_;
  wire [4:0] _03046_;
  wire [7:0] _03047_;
  wire [7:0] _03048_;
  wire [7:0] _03049_;
  wire [4:0] _03050_;
  wire [4:0] _03051_;
  wire [4:0] _03052_;
  wire [4:0] _03053_;
  wire [4:0] _03054_;
  wire [4:0] _03055_;
  wire [4:0] _03056_;
  wire [4:0] _03057_;
  wire [4:0] _03058_;
  wire [4:0] _03059_;
  wire [4:0] _03060_;
  wire [4:0] _03061_;
  wire [4:0] _03062_;
  wire [4:0] _03063_;
  wire [4:0] _03064_;
  wire [4:0] _03065_;
  wire [4:0] _03066_;
  wire [4:0] _03067_;
  wire [4:0] _03068_;
  wire [4:0] _03069_;
  wire [4:0] _03070_;
  wire [4:0] _03071_;
  wire [4:0] _03072_;
  wire [4:0] _03073_;
  wire [4:0] _03074_;
  wire [4:0] _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire [4:0] _03111_;
  wire [4:0] _03112_;
  wire [4:0] _03113_;
  wire [4:0] _03114_;
  wire [4:0] _03115_;
  wire [4:0] _03116_;
  wire [31:0] _03117_;
  wire [31:0] _03118_;
  wire [31:0] _03119_;
  wire [4:0] _03120_;
  wire [4:0] _03121_;
  wire [4:0] _03122_;
  wire [4:0] _03123_;
  wire [4:0] _03124_;
  wire [4:0] _03125_;
  wire [31:0] _03126_;
  wire [31:0] _03127_;
  wire [31:0] _03128_;
  wire [31:0] _03129_;
  wire [31:0] _03130_;
  wire [31:0] _03131_;
  wire [15:0] _03132_;
  wire [15:0] _03133_;
  wire [15:0] _03134_;
  wire [1:0] _03135_;
  wire [1:0] _03136_;
  wire [1:0] _03137_;
  wire [3:0] _03138_;
  wire [3:0] _03139_;
  wire [3:0] _03140_;
  wire [3:0] _03141_;
  wire [3:0] _03142_;
  wire [3:0] _03143_;
  wire [3:0] _03144_;
  wire [3:0] _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire [4:0] _03186_;
  wire [4:0] _03187_;
  wire [4:0] _03188_;
  wire [4:0] _03189_;
  wire [4:0] _03190_;
  wire [4:0] _03191_;
  wire [4:0] _03192_;
  wire [4:0] _03193_;
  wire [4:0] _03194_;
  wire [4:0] _03195_;
  wire [4:0] _03196_;
  wire [4:0] _03197_;
  wire [4:0] _03198_;
  wire [4:0] _03199_;
  wire [4:0] _03200_;
  wire [4:0] _03201_;
  wire [4:0] _03202_;
  wire [4:0] _03203_;
  wire [4:0] _03204_;
  wire [4:0] _03205_;
  wire [4:0] _03206_;
  wire [4:0] _03207_;
  wire [4:0] _03208_;
  wire [4:0] _03209_;
  wire [4:0] _03210_;
  wire [4:0] _03211_;
  wire [4:0] _03212_;
  wire [4:0] _03213_;
  wire [4:0] _03214_;
  wire [4:0] _03215_;
  wire [4:0] _03216_;
  wire [2:0] _03217_;
  wire [2:0] _03218_;
  wire [2:0] _03219_;
  wire [2:0] _03220_;
  wire [2:0] _03221_;
  wire [2:0] _03222_;
  wire [2:0] _03223_;
  wire [2:0] _03224_;
  wire [2:0] _03225_;
  wire [2:0] _03226_;
  wire [2:0] _03227_;
  wire [2:0] _03228_;
  wire [2:0] _03229_;
  wire [2:0] _03230_;
  wire [2:0] _03231_;
  wire [2:0] _03232_;
  wire [2:0] _03233_;
  wire [2:0] _03234_;
  wire [2:0] _03235_;
  wire [2:0] _03236_;
  wire [2:0] _03237_;
  wire [2:0] _03238_;
  wire [2:0] _03239_;
  wire [2:0] _03240_;
  wire [2:0] _03241_;
  wire [2:0] _03242_;
  wire [2:0] _03243_;
  wire [2:0] _03244_;
  wire [2:0] _03245_;
  wire [2:0] _03246_;
  wire [2:0] _03247_;
  wire [2:0] _03248_;
  wire [2:0] _03249_;
  wire [3:0] _03250_;
  wire [3:0] _03251_;
  wire [3:0] _03252_;
  wire [3:0] _03253_;
  wire [3:0] _03254_;
  wire [3:0] _03255_;
  wire [3:0] _03256_;
  wire [3:0] _03257_;
  wire [3:0] _03258_;
  wire [3:0] _03259_;
  wire [3:0] _03260_;
  wire [3:0] _03261_;
  wire [3:0] _03262_;
  wire [3:0] _03263_;
  wire [5:0] _03264_;
  wire [5:0] _03265_;
  wire [5:0] _03266_;
  wire [5:0] _03267_;
  wire [5:0] _03268_;
  wire [5:0] _03269_;
  wire [5:0] _03270_;
  wire [5:0] _03271_;
  wire [5:0] _03272_;
  wire [5:0] _03273_;
  wire [5:0] _03274_;
  wire [5:0] _03275_;
  wire [5:0] _03276_;
  wire [5:0] _03277_;
  wire [5:0] _03278_;
  wire [5:0] _03279_;
  wire [5:0] _03280_;
  wire [5:0] _03281_;
  wire [5:0] _03282_;
  wire [5:0] _03283_;
  wire [5:0] _03284_;
  wire [5:0] _03285_;
  wire [5:0] _03286_;
  wire [5:0] _03287_;
  wire [5:0] _03288_;
  wire [5:0] _03289_;
  wire [5:0] _03290_;
  wire [1:0] _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire [63:0] _03295_;
  wire [63:0] _03296_;
  wire [63:0] _03297_;
  wire [63:0] _03298_;
  wire [63:0] _03299_;
  wire [63:0] _03300_;
  wire [63:0] _03301_;
  wire [63:0] _03302_;
  wire [63:0] _03303_;
  wire [63:0] _03304_;
  wire [63:0] _03305_;
  wire [63:0] _03306_;
  wire [63:0] _03307_;
  wire [63:0] _03308_;
  wire [4:0] _03309_;
  wire [4:0] _03310_;
  wire [3:0] _03311_;
  wire [1:0] _03312_;
  wire [3:0] _03313_;
  wire [2:0] _03314_;
  wire [2:0] _03315_;
  wire [2:0] _03316_;
  wire [4:0] _03317_;
  wire [7:0] _03318_;
  wire [5:0] _03319_;
  wire [2:0] _03320_;
  wire [31:0] _03321_;
  wire [31:0] _03322_;
  wire [31:0] _03323_;
  wire [31:0] _03324_;
  wire [31:0] _03325_;
  wire [31:0] _03326_;
  wire [31:0] _03327_;
  wire [31:0] _03328_;
  wire [31:0] _03329_;
  wire [31:0] _03330_;
  wire [31:0] _03331_;
  wire [31:0] _03332_;
  wire [31:0] _03333_;
  wire [31:0] _03334_;
  wire [31:0] _03335_;
  wire [31:0] _03336_;
  wire [31:0] _03337_;
  wire [31:0] _03338_;
  wire [31:0] _03339_;
  wire [31:0] _03340_;
  wire [31:0] _03341_;
  wire [31:0] _03342_;
  wire [31:0] _03343_;
  wire [31:0] _03344_;
  wire [31:0] _03345_;
  wire [31:0] _03346_;
  wire [31:0] _03347_;
  wire [31:0] _03348_;
  wire [31:0] _03349_;
  wire [31:0] _03350_;
  wire [31:0] _03351_;
  wire [31:0] _03352_;
  wire [31:0] _03353_;
  wire [31:0] _03354_;
  wire [31:0] _03355_;
  wire [31:0] _03356_;
  wire [31:0] _03357_;
  wire [31:0] _03358_;
  wire [31:0] _03359_;
  wire _03360_;
  /* cellift = 32'd1 */
  wire _03361_;
  wire _03362_;
  /* cellift = 32'd1 */
  wire _03363_;
  wire _03364_;
  /* cellift = 32'd1 */
  wire _03365_;
  wire _03366_;
  /* cellift = 32'd1 */
  wire _03367_;
  wire _03368_;
  /* cellift = 32'd1 */
  wire _03369_;
  wire _03370_;
  /* cellift = 32'd1 */
  wire _03371_;
  wire _03372_;
  /* cellift = 32'd1 */
  wire _03373_;
  wire _03374_;
  /* cellift = 32'd1 */
  wire _03375_;
  wire _03376_;
  /* cellift = 32'd1 */
  wire _03377_;
  wire _03378_;
  /* cellift = 32'd1 */
  wire _03379_;
  wire _03380_;
  /* cellift = 32'd1 */
  wire _03381_;
  wire _03382_;
  /* cellift = 32'd1 */
  wire _03383_;
  wire _03384_;
  /* cellift = 32'd1 */
  wire _03385_;
  wire _03386_;
  /* cellift = 32'd1 */
  wire _03387_;
  wire _03388_;
  /* cellift = 32'd1 */
  wire _03389_;
  wire _03390_;
  /* cellift = 32'd1 */
  wire _03391_;
  wire _03392_;
  /* cellift = 32'd1 */
  wire _03393_;
  wire _03394_;
  /* cellift = 32'd1 */
  wire _03395_;
  wire _03396_;
  /* cellift = 32'd1 */
  wire _03397_;
  wire _03398_;
  /* cellift = 32'd1 */
  wire _03399_;
  wire _03400_;
  /* cellift = 32'd1 */
  wire _03401_;
  wire _03402_;
  /* cellift = 32'd1 */
  wire _03403_;
  wire _03404_;
  /* cellift = 32'd1 */
  wire _03405_;
  wire _03406_;
  /* cellift = 32'd1 */
  wire _03407_;
  wire _03408_;
  /* cellift = 32'd1 */
  wire _03409_;
  wire _03410_;
  /* cellift = 32'd1 */
  wire _03411_;
  wire _03412_;
  /* cellift = 32'd1 */
  wire _03413_;
  wire _03414_;
  /* cellift = 32'd1 */
  wire _03415_;
  wire _03416_;
  /* cellift = 32'd1 */
  wire _03417_;
  wire _03418_;
  /* cellift = 32'd1 */
  wire _03419_;
  wire _03420_;
  /* cellift = 32'd1 */
  wire _03421_;
  wire _03422_;
  /* cellift = 32'd1 */
  wire _03423_;
  wire _03424_;
  /* cellift = 32'd1 */
  wire _03425_;
  wire _03426_;
  /* cellift = 32'd1 */
  wire _03427_;
  wire _03428_;
  /* cellift = 32'd1 */
  wire _03429_;
  wire _03430_;
  /* cellift = 32'd1 */
  wire _03431_;
  wire _03432_;
  /* cellift = 32'd1 */
  wire _03433_;
  wire _03434_;
  /* cellift = 32'd1 */
  wire _03435_;
  wire _03436_;
  /* cellift = 32'd1 */
  wire _03437_;
  wire _03438_;
  /* cellift = 32'd1 */
  wire _03439_;
  wire _03440_;
  /* cellift = 32'd1 */
  wire _03441_;
  wire _03442_;
  /* cellift = 32'd1 */
  wire _03443_;
  wire _03444_;
  /* cellift = 32'd1 */
  wire _03445_;
  wire _03446_;
  /* cellift = 32'd1 */
  wire _03447_;
  wire _03448_;
  /* cellift = 32'd1 */
  wire _03449_;
  wire _03450_;
  /* cellift = 32'd1 */
  wire _03451_;
  wire _03452_;
  /* cellift = 32'd1 */
  wire _03453_;
  wire _03454_;
  /* cellift = 32'd1 */
  wire _03455_;
  wire [31:0] _03456_;
  wire [31:0] _03457_;
  wire [63:0] _03458_;
  wire [31:0] _03459_;
  wire [31:0] _03460_;
  wire [63:0] _03461_;
  wire [31:0] _03462_;
  wire [31:0] _03463_;
  wire [63:0] _03464_;
  wire [63:0] _03465_;
  wire [29:0] _03466_;
  wire [29:0] _03467_;
  wire [31:0] _03468_;
  wire [31:0] _03469_;
  wire [31:0] _03470_;
  wire [31:0] _03471_;
  wire [3:0] _03472_;
  wire [3:0] _03473_;
  wire [3:0] _03474_;
  wire [6:0] _03475_;
  wire [6:0] _03476_;
  wire [6:0] _03477_;
  wire [31:0] _03478_;
  wire [31:0] _03479_;
  wire [31:0] _03480_;
  wire [15:0] _03481_;
  wire [15:0] _03482_;
  wire [15:0] _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire [1:0] _03490_;
  wire [1:0] _03491_;
  wire [1:0] _03492_;
  wire [3:0] _03493_;
  wire [3:0] _03494_;
  wire [3:0] _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire [31:0] _03499_;
  wire [31:0] _03500_;
  wire [31:0] _03501_;
  wire [31:0] _03502_;
  wire [31:0] _03503_;
  wire [31:0] _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire [4:0] _03508_;
  wire [4:0] _03509_;
  wire [4:0] _03510_;
  wire [4:0] _03511_;
  wire [4:0] _03512_;
  wire [4:0] _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire [2:0] _03558_;
  wire [2:0] _03559_;
  wire [2:0] _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire [1:0] _03564_;
  wire [1:0] _03565_;
  wire [1:0] _03566_;
  wire [11:0] _03567_;
  wire [11:0] _03568_;
  wire [11:0] _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire [7:0] _03576_;
  wire [7:0] _03577_;
  wire [7:0] _03578_;
  wire [31:0] _03579_;
  wire [31:0] _03580_;
  wire [31:0] _03581_;
  wire [4:0] _03582_;
  wire [4:0] _03583_;
  wire [4:0] _03584_;
  wire [31:0] _03585_;
  wire [31:0] _03586_;
  wire [31:0] _03587_;
  wire [31:0] _03588_;
  wire [31:0] _03589_;
  wire [31:0] _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire [3:0] _03594_;
  wire [3:0] _03595_;
  wire [3:0] _03596_;
  wire [4:0] _03597_;
  wire [4:0] _03598_;
  wire [4:0] _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire [31:0] _03733_;
  wire [31:0] _03734_;
  wire [31:0] _03735_;
  wire [31:0] _03736_;
  wire [3:0] _03737_;
  wire [3:0] _03738_;
  wire [3:0] _03739_;
  wire [3:0] _03740_;
  wire [4:0] _03741_;
  wire [4:0] _03742_;
  wire [4:0] _03743_;
  wire [4:0] _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire [31:0] _03769_;
  wire [31:0] _03770_;
  wire [31:0] _03771_;
  wire [31:0] _03772_;
  wire [31:0] _03773_;
  wire [31:0] _03774_;
  wire [31:0] _03775_;
  wire [31:0] _03776_;
  wire [3:0] _03777_;
  wire [3:0] _03778_;
  wire [3:0] _03779_;
  wire [3:0] _03780_;
  wire [3:0] _03781_;
  wire [3:0] _03782_;
  wire [3:0] _03783_;
  wire [3:0] _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire [31:0] _03793_;
  wire [31:0] _03794_;
  wire [31:0] _03795_;
  wire [31:0] _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire [30:0] _03801_;
  wire [30:0] _03802_;
  wire [30:0] _03803_;
  wire [30:0] _03804_;
  wire [31:0] _03805_;
  wire [31:0] _03806_;
  wire [31:0] _03807_;
  wire [31:0] _03808_;
  wire [1:0] _03809_;
  wire [1:0] _03810_;
  wire [1:0] _03811_;
  wire [1:0] _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire [31:0] _03817_;
  wire [31:0] _03818_;
  wire [31:0] _03819_;
  wire [31:0] _03820_;
  wire [31:0] _03821_;
  wire [31:0] _03822_;
  wire [31:0] _03823_;
  wire [31:0] _03824_;
  wire [4:0] _03825_;
  wire [4:0] _03826_;
  wire [4:0] _03827_;
  wire [4:0] _03828_;
  wire [7:0] _03829_;
  wire [7:0] _03830_;
  wire [7:0] _03831_;
  wire [7:0] _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire [63:0] _03837_;
  wire [63:0] _03838_;
  wire [63:0] _03839_;
  wire [63:0] _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire [30:0] _03849_;
  wire [30:0] _03850_;
  wire [30:0] _03851_;
  wire [30:0] _03852_;
  wire [31:0] _03853_;
  wire [31:0] _03854_;
  wire [31:0] _03855_;
  wire [31:0] _03856_;
  wire [31:0] _03857_;
  wire [31:0] _03858_;
  wire [31:0] _03859_;
  wire [31:0] _03860_;
  wire [31:0] _03861_;
  wire [31:0] _03862_;
  wire [31:0] _03863_;
  wire [31:0] _03864_;
  wire [31:0] _03865_;
  wire [31:0] _03866_;
  wire [31:0] _03867_;
  wire [31:0] _03868_;
  wire [31:0] _03869_;
  wire [31:0] _03870_;
  wire [31:0] _03871_;
  wire [31:0] _03872_;
  wire [31:0] _03873_;
  wire [31:0] _03874_;
  wire [31:0] _03875_;
  wire [31:0] _03876_;
  wire [31:0] _03877_;
  wire [31:0] _03878_;
  wire [31:0] _03879_;
  wire [31:0] _03880_;
  wire [31:0] _03881_;
  wire [31:0] _03882_;
  wire [31:0] _03883_;
  wire [31:0] _03884_;
  wire [31:0] _03885_;
  wire [31:0] _03886_;
  wire [31:0] _03887_;
  wire [31:0] _03888_;
  wire [31:0] _03889_;
  wire [31:0] _03890_;
  wire [31:0] _03891_;
  wire [31:0] _03892_;
  wire [31:0] _03893_;
  wire [31:0] _03894_;
  wire [31:0] _03895_;
  wire [31:0] _03896_;
  wire [31:0] _03897_;
  wire [31:0] _03898_;
  wire [31:0] _03899_;
  wire [31:0] _03900_;
  wire [31:0] _03901_;
  wire [31:0] _03902_;
  wire [31:0] _03903_;
  wire [31:0] _03904_;
  wire [31:0] _03905_;
  wire [31:0] _03906_;
  wire [31:0] _03907_;
  wire [31:0] _03908_;
  wire [31:0] _03909_;
  wire [31:0] _03910_;
  wire [31:0] _03911_;
  wire [31:0] _03912_;
  wire [31:0] _03913_;
  wire [31:0] _03914_;
  wire [31:0] _03915_;
  wire [31:0] _03916_;
  wire [31:0] _03917_;
  wire [31:0] _03918_;
  wire [31:0] _03919_;
  wire [31:0] _03920_;
  wire [31:0] _03921_;
  wire [31:0] _03922_;
  wire [31:0] _03923_;
  wire [31:0] _03924_;
  wire [31:0] _03925_;
  wire [31:0] _03926_;
  wire [31:0] _03927_;
  wire [31:0] _03928_;
  wire [31:0] _03929_;
  wire [31:0] _03930_;
  wire [31:0] _03931_;
  wire [31:0] _03932_;
  wire [31:0] _03933_;
  wire [31:0] _03934_;
  wire [31:0] _03935_;
  wire [31:0] _03936_;
  wire [31:0] _03937_;
  wire [31:0] _03938_;
  wire [31:0] _03939_;
  wire [31:0] _03940_;
  wire [31:0] _03941_;
  wire [31:0] _03942_;
  wire [31:0] _03943_;
  wire [31:0] _03944_;
  wire [31:0] _03945_;
  wire [31:0] _03946_;
  wire [31:0] _03947_;
  wire [31:0] _03948_;
  wire [31:0] _03949_;
  wire [31:0] _03950_;
  wire [31:0] _03951_;
  wire [31:0] _03952_;
  wire [31:0] _03953_;
  wire [31:0] _03954_;
  wire [31:0] _03955_;
  wire [31:0] _03956_;
  wire [31:0] _03957_;
  wire [31:0] _03958_;
  wire [31:0] _03959_;
  wire [31:0] _03960_;
  wire [31:0] _03961_;
  wire [31:0] _03962_;
  wire [31:0] _03963_;
  wire [31:0] _03964_;
  wire [31:0] _03965_;
  wire [31:0] _03966_;
  wire [31:0] _03967_;
  wire [31:0] _03968_;
  wire [31:0] _03969_;
  wire [31:0] _03970_;
  wire [31:0] _03971_;
  wire [31:0] _03972_;
  wire [31:0] _03973_;
  wire [31:0] _03974_;
  wire [31:0] _03975_;
  wire [31:0] _03976_;
  wire [31:0] _03977_;
  wire [31:0] _03978_;
  wire [31:0] _03979_;
  wire [31:0] _03980_;
  wire [4:0] _03981_;
  wire [4:0] _03982_;
  wire [4:0] _03983_;
  wire [4:0] _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire [5:0] _04033_;
  wire [3:0] _04034_;
  wire [1:0] _04035_;
  wire [6:0] _04036_;
  wire [2:0] _04037_;
  wire [1:0] _04038_;
  wire [4:0] _04039_;
  wire [1:0] _04040_;
  wire [2:0] _04041_;
  wire [2:0] _04042_;
  wire [1:0] _04043_;
  wire [1:0] _04044_;
  wire [2:0] _04045_;
  wire [5:0] _04046_;
  wire [1:0] _04047_;
  wire [10:0] _04048_;
  wire [8:0] _04049_;
  wire [7:0] _04050_;
  wire [3:0] _04051_;
  wire [1:0] _04052_;
  wire [1:0] _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire [31:0] _04079_;
  wire [31:0] _04080_;
  wire [31:0] _04081_;
  wire [31:0] _04082_;
  wire [31:0] _04083_;
  wire [31:0] _04084_;
  wire [31:0] _04085_;
  wire [31:0] _04086_;
  wire [31:0] _04087_;
  wire [31:0] _04088_;
  wire [31:0] _04089_;
  wire [31:0] _04090_;
  wire [31:0] _04091_;
  wire [31:0] _04092_;
  wire [31:0] _04093_;
  wire [31:0] _04094_;
  wire [31:0] _04095_;
  wire [31:0] _04096_;
  wire [31:0] _04097_;
  wire [31:0] _04098_;
  wire [31:0] _04099_;
  wire [31:0] _04100_;
  wire [31:0] _04101_;
  wire [31:0] _04102_;
  wire [31:0] _04103_;
  wire [31:0] _04104_;
  wire [31:0] _04105_;
  wire [31:0] _04106_;
  wire [31:0] _04107_;
  wire [31:0] _04108_;
  wire [4:0] _04109_;
  wire [4:0] _04110_;
  wire [4:0] _04111_;
  wire [4:0] _04112_;
  wire [4:0] _04113_;
  wire [4:0] _04114_;
  wire [4:0] _04115_;
  wire [4:0] _04116_;
  wire [4:0] _04117_;
  wire [4:0] _04118_;
  wire [4:0] _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire [7:0] _04131_;
  wire [7:0] _04132_;
  wire [7:0] _04133_;
  wire [7:0] _04134_;
  wire [7:0] _04135_;
  wire [7:0] _04136_;
  wire [7:0] _04137_;
  wire [7:0] _04138_;
  wire [7:0] _04139_;
  wire [7:0] _04140_;
  wire [7:0] _04141_;
  wire [7:0] _04142_;
  wire [7:0] _04143_;
  wire [7:0] _04144_;
  wire [7:0] _04145_;
  wire [7:0] _04146_;
  wire [7:0] _04147_;
  wire [7:0] _04148_;
  wire [7:0] _04149_;
  wire [7:0] _04150_;
  wire [7:0] _04151_;
  wire [7:0] _04152_;
  wire [7:0] _04153_;
  wire [7:0] _04154_;
  wire [7:0] _04155_;
  wire [7:0] _04156_;
  wire [7:0] _04157_;
  wire [7:0] _04158_;
  wire [7:0] _04159_;
  wire [7:0] _04160_;
  wire [31:0] _04161_;
  wire [31:0] _04162_;
  wire [31:0] _04163_;
  wire [31:0] _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire [1:0] _04184_;
  wire [1:0] _04185_;
  wire [1:0] _04186_;
  wire [1:0] _04187_;
  wire [1:0] _04188_;
  wire [1:0] _04189_;
  wire [31:0] _04190_;
  wire [31:0] _04191_;
  wire [31:0] _04192_;
  wire [31:0] _04193_;
  wire [31:0] _04194_;
  wire [31:0] _04195_;
  wire [31:0] _04196_;
  wire [31:0] _04197_;
  wire [31:0] _04198_;
  wire [31:0] _04199_;
  wire [31:0] _04200_;
  wire [31:0] _04201_;
  wire [31:0] _04202_;
  wire [31:0] _04203_;
  wire [31:0] _04204_;
  wire [31:0] _04205_;
  wire [31:0] _04206_;
  wire [31:0] _04207_;
  wire [31:0] _04208_;
  wire [31:0] _04209_;
  wire [31:0] _04210_;
  wire [31:0] _04211_;
  wire [31:0] _04212_;
  wire [31:0] _04213_;
  wire [31:0] _04214_;
  wire [31:0] _04215_;
  wire [31:0] _04216_;
  wire [31:0] _04217_;
  wire [31:0] _04218_;
  wire [31:0] _04219_;
  wire [31:0] _04220_;
  wire [31:0] _04221_;
  wire [31:0] _04222_;
  wire [31:0] _04223_;
  wire [31:0] _04224_;
  wire [31:0] _04225_;
  wire [31:0] _04226_;
  wire [31:0] _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire [3:0] _04265_;
  wire [3:0] _04266_;
  wire [3:0] _04267_;
  wire [3:0] _04268_;
  wire [3:0] _04269_;
  wire [3:0] _04270_;
  wire [3:0] _04271_;
  wire [3:0] _04272_;
  wire [3:0] _04273_;
  wire [3:0] _04274_;
  wire [3:0] _04275_;
  wire [3:0] _04276_;
  wire [3:0] _04277_;
  wire [3:0] _04278_;
  wire [3:0] _04279_;
  wire [3:0] _04280_;
  wire [3:0] _04281_;
  wire [3:0] _04282_;
  wire [3:0] _04283_;
  wire [3:0] _04284_;
  wire [3:0] _04285_;
  wire [3:0] _04286_;
  wire [3:0] _04287_;
  wire [3:0] _04288_;
  wire [3:0] _04289_;
  wire [3:0] _04290_;
  wire [3:0] _04291_;
  wire [3:0] _04292_;
  wire [3:0] _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire [31:0] _04308_;
  wire [31:0] _04309_;
  wire [31:0] _04310_;
  wire [31:0] _04311_;
  wire [31:0] _04312_;
  wire [31:0] _04313_;
  wire [31:0] _04314_;
  wire [31:0] _04315_;
  wire [31:0] _04316_;
  wire [31:0] _04317_;
  wire [31:0] _04318_;
  wire [31:0] _04319_;
  wire [31:0] _04320_;
  wire [31:0] _04321_;
  wire [4:0] _04322_;
  wire [4:0] _04323_;
  wire [4:0] _04324_;
  wire [4:0] _04325_;
  wire [4:0] _04326_;
  wire [4:0] _04327_;
  wire [4:0] _04328_;
  wire [4:0] _04329_;
  wire [4:0] _04330_;
  wire [4:0] _04331_;
  wire [4:0] _04332_;
  wire [4:0] _04333_;
  wire [4:0] _04334_;
  wire [4:0] _04335_;
  wire [4:0] _04336_;
  wire [4:0] _04337_;
  wire [4:0] _04338_;
  wire [4:0] _04339_;
  wire [4:0] _04340_;
  wire [4:0] _04341_;
  wire [4:0] _04342_;
  wire [4:0] _04343_;
  wire [4:0] _04344_;
  wire [4:0] _04345_;
  wire [4:0] _04346_;
  wire [4:0] _04347_;
  wire [4:0] _04348_;
  wire [4:0] _04349_;
  wire [4:0] _04350_;
  wire [4:0] _04351_;
  wire [4:0] _04352_;
  wire [1:0] _04353_;
  wire [1:0] _04354_;
  wire [1:0] _04355_;
  wire [1:0] _04356_;
  wire [1:0] _04357_;
  wire [1:0] _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire [4:0] _04376_;
  wire [4:0] _04377_;
  wire [4:0] _04378_;
  wire [4:0] _04379_;
  wire [4:0] _04380_;
  wire [4:0] _04381_;
  wire [4:0] _04382_;
  wire [4:0] _04383_;
  wire [4:0] _04384_;
  wire [4:0] _04385_;
  wire [4:0] _04386_;
  wire [4:0] _04387_;
  wire [2:0] _04388_;
  wire [2:0] _04389_;
  wire [2:0] _04390_;
  wire [2:0] _04391_;
  wire [2:0] _04392_;
  wire [2:0] _04393_;
  wire [2:0] _04394_;
  wire [2:0] _04395_;
  wire [2:0] _04396_;
  wire [2:0] _04397_;
  wire [2:0] _04398_;
  wire [2:0] _04399_;
  wire [2:0] _04400_;
  wire [2:0] _04401_;
  wire [2:0] _04402_;
  wire [2:0] _04403_;
  wire [2:0] _04404_;
  wire [2:0] _04405_;
  wire [2:0] _04406_;
  wire [2:0] _04407_;
  wire [2:0] _04408_;
  wire [2:0] _04409_;
  wire [2:0] _04410_;
  wire [3:0] _04411_;
  wire [3:0] _04412_;
  wire [3:0] _04413_;
  wire [5:0] _04414_;
  wire [5:0] _04415_;
  wire [5:0] _04416_;
  wire [5:0] _04417_;
  wire [5:0] _04418_;
  wire [5:0] _04419_;
  wire [5:0] _04420_;
  wire [5:0] _04421_;
  wire [5:0] _04422_;
  wire [5:0] _04423_;
  wire [5:0] _04424_;
  wire [5:0] _04425_;
  wire [5:0] _04426_;
  wire [5:0] _04427_;
  wire [5:0] _04428_;
  wire [5:0] _04429_;
  wire [5:0] _04430_;
  wire [5:0] _04431_;
  wire [5:0] _04432_;
  wire [5:0] _04433_;
  wire [5:0] _04434_;
  wire [5:0] _04435_;
  wire [5:0] _04436_;
  wire [5:0] _04437_;
  wire [5:0] _04438_;
  wire [5:0] _04439_;
  wire [5:0] _04440_;
  wire [5:0] _04441_;
  wire [5:0] _04442_;
  wire [5:0] _04443_;
  wire [5:0] _04444_;
  wire [5:0] _04445_;
  wire [5:0] _04446_;
  wire [5:0] _04447_;
  wire [5:0] _04448_;
  wire [5:0] _04449_;
  wire [31:0] _04450_;
  wire [31:0] _04451_;
  wire [31:0] _04452_;
  wire [31:0] _04453_;
  wire [31:0] _04454_;
  wire [31:0] _04455_;
  wire [31:0] _04456_;
  wire [31:0] _04457_;
  wire [31:0] _04458_;
  wire [31:0] _04459_;
  wire [31:0] _04460_;
  wire [31:0] _04461_;
  wire [31:0] _04462_;
  wire [31:0] _04463_;
  wire [31:0] _04464_;
  wire [31:0] _04465_;
  wire [31:0] _04466_;
  wire [31:0] _04467_;
  wire [3:0] _04468_;
  wire [3:0] _04469_;
  wire [3:0] _04470_;
  wire [3:0] _04471_;
  wire [31:0] _04472_;
  wire [31:0] _04473_;
  wire [31:0] _04474_;
  wire [31:0] _04475_;
  wire [31:0] _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire [30:0] _04481_;
  wire _04482_;
  wire [4:0] _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire [4:0] _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire [30:0] _04618_;
  wire [30:0] _04619_;
  wire [31:0] _04620_;
  wire [31:0] _04621_;
  wire [31:0] _04622_;
  wire [31:0] _04623_;
  wire [31:0] _04624_;
  wire [31:0] _04625_;
  wire [31:0] _04626_;
  wire [31:0] _04627_;
  wire [31:0] _04628_;
  wire [31:0] _04629_;
  wire [31:0] _04630_;
  wire [31:0] _04631_;
  wire [31:0] _04632_;
  wire [31:0] _04633_;
  wire [31:0] _04634_;
  wire [31:0] _04635_;
  wire [31:0] _04636_;
  wire [31:0] _04637_;
  wire [31:0] _04638_;
  wire [31:0] _04639_;
  wire [31:0] _04640_;
  wire [31:0] _04641_;
  wire [31:0] _04642_;
  wire [31:0] _04643_;
  wire [31:0] _04644_;
  wire [31:0] _04645_;
  wire [31:0] _04646_;
  wire [31:0] _04647_;
  wire [31:0] _04648_;
  wire [31:0] _04649_;
  wire [31:0] _04650_;
  wire [31:0] _04651_;
  wire [31:0] _04652_;
  wire [31:0] _04653_;
  wire [31:0] _04654_;
  wire [31:0] _04655_;
  wire [31:0] _04656_;
  wire [31:0] _04657_;
  wire [31:0] _04658_;
  wire [31:0] _04659_;
  wire [31:0] _04660_;
  wire [31:0] _04661_;
  wire [31:0] _04662_;
  wire [31:0] _04663_;
  wire [31:0] _04664_;
  wire [31:0] _04665_;
  wire [31:0] _04666_;
  wire [31:0] _04667_;
  wire [31:0] _04668_;
  wire [31:0] _04669_;
  wire [31:0] _04670_;
  wire [31:0] _04671_;
  wire [31:0] _04672_;
  wire [31:0] _04673_;
  wire [31:0] _04674_;
  wire [31:0] _04675_;
  wire [31:0] _04676_;
  wire [31:0] _04677_;
  wire [31:0] _04678_;
  wire [31:0] _04679_;
  wire [31:0] _04680_;
  wire [31:0] _04681_;
  wire [31:0] _04682_;
  wire [31:0] _04683_;
  wire [31:0] _04684_;
  wire [31:0] _04685_;
  wire [31:0] _04686_;
  wire [31:0] _04687_;
  wire [31:0] _04688_;
  wire [31:0] _04689_;
  wire [31:0] _04690_;
  wire [31:0] _04691_;
  wire [31:0] _04692_;
  wire [31:0] _04693_;
  wire [31:0] _04694_;
  wire [31:0] _04695_;
  wire [31:0] _04696_;
  wire [31:0] _04697_;
  wire [31:0] _04698_;
  wire [31:0] _04699_;
  wire [31:0] _04700_;
  wire [31:0] _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire [31:0] _04734_;
  wire [63:0] _04735_;
  wire [63:0] _04736_;
  wire [31:0] _04737_;
  wire [3:0] _04738_;
  wire [31:0] _04739_;
  wire [4:0] _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire [31:0] _04748_;
  wire [31:0] _04749_;
  wire [31:0] _04750_;
  wire [31:0] _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire [31:0] _04755_;
  wire [31:0] _04756_;
  wire [31:0] _04757_;
  wire [31:0] _04758_;
  wire [31:0] _04759_;
  wire [31:0] _04760_;
  wire [4:0] _04761_;
  wire [4:0] _04762_;
  wire [4:0] _04763_;
  wire [4:0] _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire [7:0] _04771_;
  wire [7:0] _04772_;
  wire [7:0] _04773_;
  wire [7:0] _04774_;
  wire [7:0] _04775_;
  wire [7:0] _04776_;
  wire [7:0] _04777_;
  wire [7:0] _04778_;
  wire [7:0] _04779_;
  wire [7:0] _04780_;
  wire [7:0] _04781_;
  wire [7:0] _04782_;
  wire [7:0] _04783_;
  wire [7:0] _04784_;
  wire [7:0] _04785_;
  wire [7:0] _04786_;
  wire [7:0] _04787_;
  wire [7:0] _04788_;
  wire [31:0] _04789_;
  wire [31:0] _04790_;
  wire [31:0] _04791_;
  wire [31:0] _04792_;
  wire [31:0] _04793_;
  wire [31:0] _04794_;
  wire [31:0] _04795_;
  wire [31:0] _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire [1:0] _04800_;
  wire [1:0] _04801_;
  wire [1:0] _04802_;
  wire [31:0] _04803_;
  wire [31:0] _04804_;
  wire [31:0] _04805_;
  wire [31:0] _04806_;
  wire [31:0] _04807_;
  wire [31:0] _04808_;
  wire [31:0] _04809_;
  wire [31:0] _04810_;
  wire [31:0] _04811_;
  wire _04812_;
  wire [31:0] _04813_;
  wire [4:0] _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire [2:0] _04847_;
  wire [2:0] _04848_;
  wire [2:0] _04849_;
  wire _04850_;
  wire [1:0] _04851_;
  wire [1:0] _04852_;
  wire [1:0] _04853_;
  wire [11:0] _04854_;
  wire [11:0] _04855_;
  wire [11:0] _04856_;
  wire _04857_;
  wire _04858_;
  wire [3:0] _04859_;
  wire [3:0] _04860_;
  wire [3:0] _04861_;
  wire [3:0] _04862_;
  wire [3:0] _04863_;
  wire [3:0] _04864_;
  wire [3:0] _04865_;
  wire [3:0] _04866_;
  wire [3:0] _04867_;
  wire [3:0] _04868_;
  wire [3:0] _04869_;
  wire [3:0] _04870_;
  wire [3:0] _04871_;
  wire [3:0] _04872_;
  wire [3:0] _04873_;
  wire [3:0] _04874_;
  wire [3:0] _04875_;
  wire [3:0] _04876_;
  wire [3:0] _04877_;
  wire [3:0] _04878_;
  wire [3:0] _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire [4:0] _04897_;
  wire [4:0] _04898_;
  wire [4:0] _04899_;
  wire [4:0] _04900_;
  wire [4:0] _04901_;
  wire [4:0] _04902_;
  wire [4:0] _04903_;
  wire [4:0] _04904_;
  wire [4:0] _04905_;
  wire [4:0] _04906_;
  wire [4:0] _04907_;
  wire [4:0] _04908_;
  wire [7:0] _04909_;
  wire [7:0] _04910_;
  wire [7:0] _04911_;
  wire [4:0] _04912_;
  wire [4:0] _04913_;
  wire [4:0] _04914_;
  wire [4:0] _04915_;
  wire [4:0] _04916_;
  wire [4:0] _04917_;
  wire [4:0] _04918_;
  wire [4:0] _04919_;
  wire [4:0] _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire [4:0] _04931_;
  wire [4:0] _04932_;
  wire [4:0] _04933_;
  wire [4:0] _04934_;
  wire [31:0] _04935_;
  wire [31:0] _04936_;
  wire [31:0] _04937_;
  wire [4:0] _04938_;
  wire [4:0] _04939_;
  wire [4:0] _04940_;
  wire [4:0] _04941_;
  wire [31:0] _04942_;
  wire [31:0] _04943_;
  wire [31:0] _04944_;
  wire [31:0] _04945_;
  wire [31:0] _04946_;
  wire [31:0] _04947_;
  wire [15:0] _04948_;
  wire [15:0] _04949_;
  wire [15:0] _04950_;
  wire [15:0] _04951_;
  wire [15:0] _04952_;
  wire [15:0] _04953_;
  wire [1:0] _04954_;
  wire [1:0] _04955_;
  wire [1:0] _04956_;
  wire [3:0] _04957_;
  wire [3:0] _04958_;
  wire [3:0] _04959_;
  wire [3:0] _04960_;
  wire [3:0] _04961_;
  wire [3:0] _04962_;
  wire [3:0] _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire [4:0] _04979_;
  wire [4:0] _04980_;
  wire [4:0] _04981_;
  wire [4:0] _04982_;
  wire [4:0] _04983_;
  wire [4:0] _04984_;
  wire [4:0] _04985_;
  wire [4:0] _04986_;
  wire [4:0] _04987_;
  wire [4:0] _04988_;
  wire [4:0] _04989_;
  wire [4:0] _04990_;
  wire [4:0] _04991_;
  wire [4:0] _04992_;
  wire [4:0] _04993_;
  wire [4:0] _04994_;
  wire [4:0] _04995_;
  wire [4:0] _04996_;
  wire [4:0] _04997_;
  wire [4:0] _04998_;
  wire [2:0] _04999_;
  wire [2:0] _05000_;
  wire [2:0] _05001_;
  wire [2:0] _05002_;
  wire [2:0] _05003_;
  wire [2:0] _05004_;
  wire [2:0] _05005_;
  wire [2:0] _05006_;
  wire [2:0] _05007_;
  wire [2:0] _05008_;
  wire [2:0] _05009_;
  wire [2:0] _05010_;
  wire [2:0] _05011_;
  wire [2:0] _05012_;
  wire [2:0] _05013_;
  wire [2:0] _05014_;
  wire [2:0] _05015_;
  wire [2:0] _05016_;
  wire [2:0] _05017_;
  wire [2:0] _05018_;
  wire [2:0] _05019_;
  wire [3:0] _05020_;
  wire [3:0] _05021_;
  wire [3:0] _05022_;
  wire [3:0] _05023_;
  wire [3:0] _05024_;
  wire [3:0] _05025_;
  wire [3:0] _05026_;
  wire [3:0] _05027_;
  wire [3:0] _05028_;
  wire [5:0] _05029_;
  wire [5:0] _05030_;
  wire [5:0] _05031_;
  wire [5:0] _05032_;
  wire [5:0] _05033_;
  wire [5:0] _05034_;
  wire [5:0] _05035_;
  wire [5:0] _05036_;
  wire [5:0] _05037_;
  wire [5:0] _05038_;
  wire [5:0] _05039_;
  wire [5:0] _05040_;
  wire [5:0] _05041_;
  wire [5:0] _05042_;
  wire [5:0] _05043_;
  wire [5:0] _05044_;
  wire [5:0] _05045_;
  wire [5:0] _05046_;
  wire [5:0] _05047_;
  wire [5:0] _05048_;
  wire [5:0] _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire [63:0] _05053_;
  wire [63:0] _05054_;
  wire [63:0] _05055_;
  wire [63:0] _05056_;
  wire [63:0] _05057_;
  wire [63:0] _05058_;
  wire [63:0] _05059_;
  wire [1:0] _05060_;
  wire [1:0] _05061_;
  wire [1:0] _05062_;
  wire [1:0] _05063_;
  wire [31:0] _05064_;
  wire [31:0] _05065_;
  wire [31:0] _05066_;
  wire [31:0] _05067_;
  wire [31:0] _05068_;
  wire [31:0] _05069_;
  wire [31:0] _05070_;
  wire [31:0] _05071_;
  wire [31:0] _05072_;
  wire [31:0] _05073_;
  wire [31:0] _05074_;
  wire [31:0] _05075_;
  wire [31:0] _05076_;
  wire [31:0] _05077_;
  wire [31:0] _05078_;
  wire [31:0] _05079_;
  wire [31:0] _05080_;
  wire [31:0] _05081_;
  wire [31:0] _05082_;
  wire [31:0] _05083_;
  wire [31:0] _05084_;
  wire [31:0] _05085_;
  wire [31:0] _05086_;
  wire [31:0] _05087_;
  wire [31:0] _05088_;
  wire [31:0] _05089_;
  wire [31:0] _05090_;
  wire [31:0] _05091_;
  wire [31:0] _05092_;
  wire [31:0] _05093_;
  wire [31:0] _05094_;
  wire [31:0] _05095_;
  wire [31:0] _05096_;
  wire [31:0] _05097_;
  wire [31:0] _05098_;
  wire [31:0] _05099_;
  wire _05100_;
  /* cellift = 32'd1 */
  wire _05101_;
  wire _05102_;
  /* cellift = 32'd1 */
  wire _05103_;
  wire _05104_;
  /* cellift = 32'd1 */
  wire _05105_;
  wire _05106_;
  /* cellift = 32'd1 */
  wire _05107_;
  wire _05108_;
  /* cellift = 32'd1 */
  wire _05109_;
  wire _05110_;
  /* cellift = 32'd1 */
  wire _05111_;
  wire _05112_;
  /* cellift = 32'd1 */
  wire _05113_;
  wire _05114_;
  /* cellift = 32'd1 */
  wire _05115_;
  wire _05116_;
  /* cellift = 32'd1 */
  wire _05117_;
  wire _05118_;
  /* cellift = 32'd1 */
  wire _05119_;
  wire _05120_;
  /* cellift = 32'd1 */
  wire _05121_;
  wire _05122_;
  /* cellift = 32'd1 */
  wire _05123_;
  wire _05124_;
  /* cellift = 32'd1 */
  wire _05125_;
  wire _05126_;
  /* cellift = 32'd1 */
  wire _05127_;
  wire _05128_;
  /* cellift = 32'd1 */
  wire _05129_;
  wire _05130_;
  /* cellift = 32'd1 */
  wire _05131_;
  wire _05132_;
  /* cellift = 32'd1 */
  wire _05133_;
  wire _05134_;
  /* cellift = 32'd1 */
  wire _05135_;
  wire [31:0] _05136_;
  wire [31:0] _05137_;
  wire [31:0] _05138_;
  wire [31:0] _05139_;
  wire [63:0] _05140_;
  wire [31:0] _05141_;
  wire [31:0] _05142_;
  wire [31:0] _05143_;
  wire [63:0] _05144_;
  wire [31:0] _05145_;
  wire [31:0] _05146_;
  wire [31:0] _05147_;
  wire [31:0] _05148_;
  wire [31:0] _05149_;
  wire [63:0] _05150_;
  wire [63:0] _05151_;
  wire [63:0] _05152_;
  wire [29:0] _05153_;
  wire [29:0] _05154_;
  wire [29:0] _05155_;
  wire [31:0] _05156_;
  wire [31:0] _05157_;
  wire [31:0] _05158_;
  wire [31:0] _05159_;
  wire [31:0] _05160_;
  wire [3:0] _05161_;
  wire [6:0] _05162_;
  wire [6:0] _05163_;
  wire [6:0] _05164_;
  wire [6:0] _05165_;
  wire [31:0] _05166_;
  wire [31:0] _05167_;
  wire [31:0] _05168_;
  wire [31:0] _05169_;
  wire [15:0] _05170_;
  wire [15:0] _05171_;
  wire [15:0] _05172_;
  wire [15:0] _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire [1:0] _05182_;
  wire [1:0] _05183_;
  wire [1:0] _05184_;
  wire [1:0] _05185_;
  wire [3:0] _05186_;
  wire [3:0] _05187_;
  wire [3:0] _05188_;
  wire [3:0] _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire [31:0] _05194_;
  wire [31:0] _05195_;
  wire [31:0] _05196_;
  wire [31:0] _05197_;
  wire [31:0] _05198_;
  wire [31:0] _05199_;
  wire [31:0] _05200_;
  wire [31:0] _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire [4:0] _05206_;
  wire [4:0] _05207_;
  wire [4:0] _05208_;
  wire [4:0] _05209_;
  wire [4:0] _05210_;
  wire [4:0] _05211_;
  wire [4:0] _05212_;
  wire [4:0] _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire [2:0] _05272_;
  wire [2:0] _05273_;
  wire [2:0] _05274_;
  wire [2:0] _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire [1:0] _05280_;
  wire [1:0] _05281_;
  wire [1:0] _05282_;
  wire [1:0] _05283_;
  wire [11:0] _05284_;
  wire [11:0] _05285_;
  wire [11:0] _05286_;
  wire [11:0] _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire [7:0] _05296_;
  wire [7:0] _05297_;
  wire [7:0] _05298_;
  wire [7:0] _05299_;
  wire [31:0] _05300_;
  wire [31:0] _05301_;
  wire [31:0] _05302_;
  wire [31:0] _05303_;
  wire [4:0] _05304_;
  wire [4:0] _05305_;
  wire [4:0] _05306_;
  wire [4:0] _05307_;
  wire [31:0] _05308_;
  wire [31:0] _05309_;
  wire [31:0] _05310_;
  wire [31:0] _05311_;
  wire [31:0] _05312_;
  wire [31:0] _05313_;
  wire [31:0] _05314_;
  wire [31:0] _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire [3:0] _05320_;
  wire [3:0] _05321_;
  wire [3:0] _05322_;
  wire [3:0] _05323_;
  wire [4:0] _05324_;
  wire [4:0] _05325_;
  wire [4:0] _05326_;
  wire [4:0] _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire [31:0] _05447_;
  wire [3:0] _05448_;
  wire [4:0] _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire [31:0] _05456_;
  wire [31:0] _05457_;
  wire [3:0] _05458_;
  wire [3:0] _05459_;
  wire _05460_;
  wire [31:0] _05461_;
  wire _05462_;
  wire [30:0] _05463_;
  wire [31:0] _05464_;
  wire [1:0] _05465_;
  wire _05466_;
  wire [31:0] _05467_;
  wire [31:0] _05468_;
  wire [4:0] _05469_;
  wire [7:0] _05470_;
  wire _05471_;
  wire [63:0] _05472_;
  wire _05473_;
  wire _05474_;
  wire [30:0] _05475_;
  wire [31:0] _05476_;
  wire [31:0] _05477_;
  wire [31:0] _05478_;
  wire [31:0] _05479_;
  wire [31:0] _05480_;
  wire [31:0] _05481_;
  wire [31:0] _05482_;
  wire [31:0] _05483_;
  wire [31:0] _05484_;
  wire [31:0] _05485_;
  wire [31:0] _05486_;
  wire [31:0] _05487_;
  wire [31:0] _05488_;
  wire [31:0] _05489_;
  wire [31:0] _05490_;
  wire [31:0] _05491_;
  wire [31:0] _05492_;
  wire [31:0] _05493_;
  wire [31:0] _05494_;
  wire [31:0] _05495_;
  wire [31:0] _05496_;
  wire [31:0] _05497_;
  wire [31:0] _05498_;
  wire [31:0] _05499_;
  wire [31:0] _05500_;
  wire [31:0] _05501_;
  wire [31:0] _05502_;
  wire [31:0] _05503_;
  wire [31:0] _05504_;
  wire [31:0] _05505_;
  wire [31:0] _05506_;
  wire [31:0] _05507_;
  wire [4:0] _05508_;
  wire [4:0] _05509_;
  wire _05510_;
  wire _05511_;
  wire [31:0] _05512_;
  wire [31:0] _05513_;
  wire [31:0] _05514_;
  wire [31:0] _05515_;
  wire [31:0] _05516_;
  wire [31:0] _05517_;
  wire [31:0] _05518_;
  wire [31:0] _05519_;
  wire [31:0] _05520_;
  wire [31:0] _05521_;
  wire [4:0] _05522_;
  wire [4:0] _05523_;
  wire [4:0] _05524_;
  wire [4:0] _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire [7:0] _05533_;
  wire [7:0] _05534_;
  wire [7:0] _05535_;
  wire [7:0] _05536_;
  wire [7:0] _05537_;
  wire [7:0] _05538_;
  wire [7:0] _05539_;
  wire [7:0] _05540_;
  wire [7:0] _05541_;
  wire [7:0] _05542_;
  wire [7:0] _05543_;
  wire [7:0] _05544_;
  wire [7:0] _05545_;
  wire [31:0] _05546_;
  wire [31:0] _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire [1:0] _05555_;
  wire [1:0] _05556_;
  wire [1:0] _05557_;
  wire [1:0] _05558_;
  wire [31:0] _05559_;
  wire [31:0] _05560_;
  wire [31:0] _05561_;
  wire [31:0] _05562_;
  wire [31:0] _05563_;
  wire [31:0] _05564_;
  wire [31:0] _05565_;
  wire [31:0] _05566_;
  wire [31:0] _05567_;
  wire [31:0] _05568_;
  wire [31:0] _05569_;
  wire [31:0] _05570_;
  wire [31:0] _05571_;
  wire [31:0] _05572_;
  wire [31:0] _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire [3:0] _05587_;
  wire [3:0] _05588_;
  wire [3:0] _05589_;
  wire [3:0] _05590_;
  wire [3:0] _05591_;
  wire [3:0] _05592_;
  wire [3:0] _05593_;
  wire [3:0] _05594_;
  wire [3:0] _05595_;
  wire [3:0] _05596_;
  wire [3:0] _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire [31:0] _05607_;
  wire [31:0] _05608_;
  wire [31:0] _05609_;
  wire [31:0] _05610_;
  wire [4:0] _05611_;
  wire [4:0] _05612_;
  wire [4:0] _05613_;
  wire [4:0] _05614_;
  wire [4:0] _05615_;
  wire [4:0] _05616_;
  wire [4:0] _05617_;
  wire [4:0] _05618_;
  wire [4:0] _05619_;
  wire [4:0] _05620_;
  wire [4:0] _05621_;
  wire [4:0] _05622_;
  wire [4:0] _05623_;
  wire [4:0] _05624_;
  wire [4:0] _05625_;
  wire [1:0] _05626_;
  wire [1:0] _05627_;
  wire [1:0] _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire [4:0] _05640_;
  wire [4:0] _05641_;
  wire [4:0] _05642_;
  wire [4:0] _05643_;
  wire [4:0] _05644_;
  wire [4:0] _05645_;
  wire [4:0] _05646_;
  wire [4:0] _05647_;
  wire [4:0] _05648_;
  wire [4:0] _05649_;
  wire [2:0] _05650_;
  wire [2:0] _05651_;
  wire [2:0] _05652_;
  wire [2:0] _05653_;
  wire [2:0] _05654_;
  wire [2:0] _05655_;
  wire [2:0] _05656_;
  wire [2:0] _05657_;
  wire [2:0] _05658_;
  wire [2:0] _05659_;
  wire [2:0] _05660_;
  wire [3:0] _05661_;
  wire [3:0] _05662_;
  wire [3:0] _05663_;
  wire [5:0] _05664_;
  wire [5:0] _05665_;
  wire [5:0] _05666_;
  wire [5:0] _05667_;
  wire [5:0] _05668_;
  wire [5:0] _05669_;
  wire [5:0] _05670_;
  wire [5:0] _05671_;
  wire [5:0] _05672_;
  wire [5:0] _05673_;
  wire [5:0] _05674_;
  wire [5:0] _05675_;
  wire [5:0] _05676_;
  wire [31:0] _05677_;
  wire [31:0] _05678_;
  wire [31:0] _05679_;
  wire [31:0] _05680_;
  wire [31:0] _05681_;
  wire [31:0] _05682_;
  wire [3:0] _05683_;
  wire [31:0] _05684_;
  wire [31:0] _05685_;
  wire [31:0] _05686_;
  wire _05687_;
  wire [31:0] _05688_;
  wire [31:0] _05689_;
  wire [31:0] _05690_;
  wire [31:0] _05691_;
  wire [31:0] _05692_;
  wire [31:0] _05693_;
  wire [31:0] _05694_;
  wire [31:0] _05695_;
  wire [31:0] _05696_;
  wire [31:0] _05697_;
  wire [31:0] _05698_;
  wire [31:0] _05699_;
  wire [31:0] _05700_;
  wire [31:0] _05701_;
  wire [31:0] _05702_;
  wire [31:0] _05703_;
  wire [31:0] _05704_;
  wire [31:0] _05705_;
  wire [31:0] _05706_;
  wire [31:0] _05707_;
  wire [31:0] _05708_;
  wire [31:0] _05709_;
  wire [31:0] _05710_;
  wire [31:0] _05711_;
  wire [31:0] _05712_;
  wire [31:0] _05713_;
  wire [31:0] _05714_;
  wire [31:0] _05715_;
  wire [31:0] _05716_;
  wire [31:0] _05717_;
  wire [31:0] _05718_;
  wire [31:0] _05719_;
  wire [31:0] _05720_;
  wire [31:0] _05721_;
  wire [31:0] _05722_;
  wire [31:0] _05723_;
  wire [31:0] _05724_;
  wire [31:0] _05725_;
  wire [31:0] _05726_;
  wire [31:0] _05727_;
  wire [31:0] _05728_;
  wire [31:0] _05729_;
  wire [31:0] _05730_;
  wire [31:0] _05731_;
  wire [31:0] _05732_;
  wire [31:0] _05733_;
  wire [31:0] _05734_;
  wire [4:0] _05735_;
  wire [31:0] _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire [4:0] _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire [7:0] _05744_;
  wire [7:0] _05745_;
  wire [7:0] _05746_;
  wire [7:0] _05747_;
  /* unused_bits = "6" */
  wire [7:0] _05748_;
  wire [7:0] _05749_;
  wire [7:0] _05750_;
  wire [7:0] _05751_;
  wire [31:0] _05752_;
  wire [31:0] _05753_;
  wire [31:0] _05754_;
  wire _05755_;
  wire _05756_;
  wire [31:0] _05757_;
  wire [31:0] _05758_;
  wire [31:0] _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire [2:0] _05771_;
  wire _05772_;
  wire [1:0] _05773_;
  wire [11:0] _05774_;
  wire _05775_;
  wire _05776_;
  wire [3:0] _05777_;
  wire [3:0] _05778_;
  wire [3:0] _05779_;
  wire [3:0] _05780_;
  wire [3:0] _05781_;
  wire [3:0] _05782_;
  wire [3:0] _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire [4:0] _05797_;
  wire [4:0] _05798_;
  wire [4:0] _05799_;
  wire [4:0] _05800_;
  wire [7:0] _05801_;
  wire [4:0] _05802_;
  wire [4:0] _05803_;
  wire [4:0] _05804_;
  wire [4:0] _05805_;
  wire [4:0] _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire [4:0] _05816_;
  wire [4:0] _05817_;
  wire [31:0] _05818_;
  wire [4:0] _05819_;
  wire [4:0] _05820_;
  wire [31:0] _05821_;
  wire [31:0] _05822_;
  wire [15:0] _05823_;
  wire [1:0] _05824_;
  wire [1:0] _05825_;
  wire [3:0] _05826_;
  wire [3:0] _05827_;
  wire [3:0] _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire [4:0] _05843_;
  wire [4:0] _05844_;
  wire [4:0] _05845_;
  wire [4:0] _05846_;
  wire [4:0] _05847_;
  wire [4:0] _05848_;
  wire [4:0] _05849_;
  wire [4:0] _05850_;
  wire [4:0] _05851_;
  wire [4:0] _05852_;
  wire [2:0] _05853_;
  wire [2:0] _05854_;
  wire [2:0] _05855_;
  wire [2:0] _05856_;
  wire [2:0] _05857_;
  wire [2:0] _05858_;
  wire [2:0] _05859_;
  wire [2:0] _05860_;
  wire [2:0] _05861_;
  wire [2:0] _05862_;
  wire [3:0] _05863_;
  wire [3:0] _05864_;
  wire [3:0] _05865_;
  wire [3:0] _05866_;
  wire [3:0] _05867_;
  wire [5:0] _05868_;
  wire [5:0] _05869_;
  wire [5:0] _05870_;
  wire [5:0] _05871_;
  wire [5:0] _05872_;
  wire [5:0] _05873_;
  wire [5:0] _05874_;
  wire [5:0] _05875_;
  wire [5:0] _05876_;
  wire _05877_;
  wire [63:0] _05878_;
  wire [63:0] _05879_;
  wire [31:0] _05880_;
  wire [31:0] _05881_;
  wire [31:0] _05882_;
  wire [31:0] _05883_;
  wire [31:0] _05884_;
  wire [31:0] _05885_;
  wire [31:0] _05886_;
  wire [31:0] _05887_;
  wire [31:0] _05888_;
  wire [31:0] _05889_;
  wire [31:0] _05890_;
  wire [31:0] _05891_;
  wire [31:0] _05892_;
  wire [31:0] _05893_;
  wire [31:0] _05894_;
  wire [31:0] _05895_;
  wire [31:0] _05896_;
  wire [63:0] _05897_;
  wire [31:0] _05898_;
  wire [63:0] _05899_;
  wire [31:0] _05900_;
  wire [31:0] _05901_;
  wire [31:0] _05902_;
  wire [63:0] _05903_;
  wire [29:0] _05904_;
  wire [6:0] _05905_;
  wire [31:0] _05906_;
  wire [15:0] _05907_;
  wire _05908_;
  wire _05909_;
  wire [1:0] _05910_;
  wire [3:0] _05911_;
  wire _05912_;
  wire [31:0] _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire [2:0] _05929_;
  wire _05930_;
  wire [1:0] _05931_;
  wire [11:0] _05932_;
  wire _05933_;
  wire _05934_;
  wire [7:0] _05935_;
  wire [31:0] _05936_;
  wire [31:0] _05937_;
  wire [31:0] _05938_;
  wire _05939_;
  wire [3:0] _05940_;
  wire [4:0] _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire [31:0] _06070_;
  wire [31:0] _06071_;
  wire [31:0] _06072_;
  wire [31:0] _06073_;
  wire [63:0] _06074_;
  wire [63:0] _06075_;
  wire [31:0] _06076_;
  wire [31:0] _06077_;
  wire [63:0] _06078_;
  wire [63:0] _06079_;
  wire [31:0] _06080_;
  wire [31:0] _06081_;
  wire [31:0] _06082_;
  wire [31:0] _06083_;
  wire [31:0] _06084_;
  wire [31:0] _06085_;
  wire [63:0] _06086_;
  wire [63:0] _06087_;
  wire [29:0] _06088_;
  wire [29:0] _06089_;
  wire [31:0] _06090_;
  wire [31:0] _06091_;
  wire [31:0] _06092_;
  wire [31:0] _06093_;
  wire [31:0] _06094_;
  wire [31:0] _06095_;
  wire [31:0] _06096_;
  wire [31:0] _06097_;
  wire [31:0] _06098_;
  wire [31:0] _06099_;
  wire [31:0] _06100_;
  wire [31:0] _06101_;
  wire [4:0] _06102_;
  /* cellift = 32'd1 */
  wire [4:0] _06103_;
  wire [4:0] _06104_;
  /* cellift = 32'd1 */
  wire [4:0] _06105_;
  wire _06106_;
  /* cellift = 32'd1 */
  wire _06107_;
  wire _06108_;
  /* cellift = 32'd1 */
  wire _06109_;
  wire [31:0] _06110_;
  /* cellift = 32'd1 */
  wire [31:0] _06111_;
  wire [31:0] _06112_;
  /* cellift = 32'd1 */
  wire [31:0] _06113_;
  wire [31:0] _06114_;
  /* cellift = 32'd1 */
  wire [31:0] _06115_;
  wire [31:0] _06116_;
  /* cellift = 32'd1 */
  wire [31:0] _06117_;
  wire [31:0] _06118_;
  /* cellift = 32'd1 */
  wire [31:0] _06119_;
  wire [31:0] _06120_;
  /* cellift = 32'd1 */
  wire [31:0] _06121_;
  wire [31:0] _06122_;
  /* cellift = 32'd1 */
  wire [31:0] _06123_;
  wire [31:0] _06124_;
  /* cellift = 32'd1 */
  wire [31:0] _06125_;
  wire [31:0] _06126_;
  /* cellift = 32'd1 */
  wire [31:0] _06127_;
  wire [31:0] _06128_;
  /* cellift = 32'd1 */
  wire [31:0] _06129_;
  wire [4:0] _06130_;
  /* cellift = 32'd1 */
  wire [4:0] _06131_;
  wire [4:0] _06132_;
  /* cellift = 32'd1 */
  wire [4:0] _06133_;
  wire [4:0] _06134_;
  /* cellift = 32'd1 */
  wire [4:0] _06135_;
  wire [4:0] _06136_;
  /* cellift = 32'd1 */
  wire [4:0] _06137_;
  wire [4:0] _06138_;
  /* cellift = 32'd1 */
  wire [4:0] _06139_;
  wire _06140_;
  /* cellift = 32'd1 */
  wire _06141_;
  wire _06142_;
  /* cellift = 32'd1 */
  wire _06143_;
  wire _06144_;
  /* cellift = 32'd1 */
  wire _06145_;
  wire _06146_;
  /* cellift = 32'd1 */
  wire _06147_;
  wire _06148_;
  /* cellift = 32'd1 */
  wire _06149_;
  wire _06150_;
  /* cellift = 32'd1 */
  wire _06151_;
  wire _06152_;
  /* cellift = 32'd1 */
  wire _06153_;
  wire _06154_;
  /* cellift = 32'd1 */
  wire _06155_;
  /* cellift = 32'd1 */
  wire _06156_;
  wire [7:0] _06157_;
  /* cellift = 32'd1 */
  wire [7:0] _06158_;
  wire [7:0] _06159_;
  /* cellift = 32'd1 */
  wire [7:0] _06160_;
  wire [7:0] _06161_;
  /* cellift = 32'd1 */
  wire [7:0] _06162_;
  wire [7:0] _06163_;
  /* cellift = 32'd1 */
  wire [7:0] _06164_;
  wire [7:0] _06165_;
  /* cellift = 32'd1 */
  wire [7:0] _06166_;
  wire [7:0] _06167_;
  /* cellift = 32'd1 */
  wire [7:0] _06168_;
  wire [7:0] _06169_;
  wire [7:0] _06170_;
  /* cellift = 32'd1 */
  wire [7:0] _06171_;
  wire [7:0] _06172_;
  /* cellift = 32'd1 */
  wire [7:0] _06173_;
  wire [7:0] _06174_;
  wire [7:0] _06175_;
  /* cellift = 32'd1 */
  wire [7:0] _06176_;
  wire [7:0] _06177_;
  wire [7:0] _06178_;
  /* cellift = 32'd1 */
  wire [7:0] _06179_;
  wire [7:0] _06180_;
  /* cellift = 32'd1 */
  wire [7:0] _06181_;
  wire [7:0] _06182_;
  /* cellift = 32'd1 */
  wire [7:0] _06183_;
  wire [7:0] _06184_;
  /* cellift = 32'd1 */
  wire [7:0] _06185_;
  wire _06186_;
  wire _06187_;
  wire [31:0] _06188_;
  /* cellift = 32'd1 */
  wire [31:0] _06189_;
  wire [31:0] _06190_;
  /* cellift = 32'd1 */
  wire [31:0] _06191_;
  wire _06192_;
  /* cellift = 32'd1 */
  wire _06193_;
  wire _06194_;
  /* cellift = 32'd1 */
  wire _06195_;
  wire _06196_;
  /* cellift = 32'd1 */
  wire _06197_;
  wire _06198_;
  wire _06199_;
  /* cellift = 32'd1 */
  wire _06200_;
  wire _06201_;
  /* cellift = 32'd1 */
  wire _06202_;
  wire _06203_;
  /* cellift = 32'd1 */
  wire _06204_;
  wire _06205_;
  /* cellift = 32'd1 */
  wire _06206_;
  wire _06207_;
  /* cellift = 32'd1 */
  wire _06208_;
  wire _06209_;
  /* cellift = 32'd1 */
  wire _06210_;
  wire _06211_;
  /* cellift = 32'd1 */
  wire _06212_;
  wire _06213_;
  /* cellift = 32'd1 */
  wire _06214_;
  /* cellift = 32'd1 */
  wire [1:0] _06215_;
  wire [1:0] _06216_;
  /* cellift = 32'd1 */
  wire [1:0] _06217_;
  wire [1:0] _06218_;
  /* cellift = 32'd1 */
  wire [1:0] _06219_;
  wire [1:0] _06220_;
  /* cellift = 32'd1 */
  wire [1:0] _06221_;
  wire [1:0] _06222_;
  /* cellift = 32'd1 */
  wire [1:0] _06223_;
  wire [31:0] _06224_;
  /* cellift = 32'd1 */
  wire [31:0] _06225_;
  wire [31:0] _06226_;
  /* cellift = 32'd1 */
  wire [31:0] _06227_;
  wire [31:0] _06228_;
  /* cellift = 32'd1 */
  wire [31:0] _06229_;
  wire [31:0] _06230_;
  /* cellift = 32'd1 */
  wire [31:0] _06231_;
  wire [31:0] _06232_;
  /* cellift = 32'd1 */
  wire [31:0] _06233_;
  wire [31:0] _06234_;
  /* cellift = 32'd1 */
  wire [31:0] _06235_;
  wire [31:0] _06236_;
  /* cellift = 32'd1 */
  wire [31:0] _06237_;
  wire [31:0] _06238_;
  /* cellift = 32'd1 */
  wire [31:0] _06239_;
  wire [31:0] _06240_;
  /* cellift = 32'd1 */
  wire [31:0] _06241_;
  wire [31:0] _06242_;
  /* cellift = 32'd1 */
  wire [31:0] _06243_;
  wire [31:0] _06244_;
  /* cellift = 32'd1 */
  wire [31:0] _06245_;
  wire [31:0] _06246_;
  /* cellift = 32'd1 */
  wire [31:0] _06247_;
  wire [31:0] _06248_;
  /* cellift = 32'd1 */
  wire [31:0] _06249_;
  wire [31:0] _06250_;
  /* cellift = 32'd1 */
  wire [31:0] _06251_;
  wire [31:0] _06252_;
  /* cellift = 32'd1 */
  wire [31:0] _06253_;
  wire _06254_;
  /* cellift = 32'd1 */
  wire _06255_;
  wire _06256_;
  /* cellift = 32'd1 */
  wire _06257_;
  wire _06258_;
  /* cellift = 32'd1 */
  wire _06259_;
  wire _06260_;
  /* cellift = 32'd1 */
  wire _06261_;
  wire _06262_;
  /* cellift = 32'd1 */
  wire _06263_;
  wire _06264_;
  /* cellift = 32'd1 */
  wire _06265_;
  wire _06266_;
  /* cellift = 32'd1 */
  wire _06267_;
  wire _06268_;
  /* cellift = 32'd1 */
  wire _06269_;
  wire _06270_;
  /* cellift = 32'd1 */
  wire _06271_;
  wire _06272_;
  /* cellift = 32'd1 */
  wire _06273_;
  wire _06274_;
  /* cellift = 32'd1 */
  wire _06275_;
  wire _06276_;
  /* cellift = 32'd1 */
  wire _06277_;
  wire _06278_;
  /* cellift = 32'd1 */
  wire _06279_;
  wire [3:0] _06280_;
  /* cellift = 32'd1 */
  wire [3:0] _06281_;
  wire [3:0] _06282_;
  /* cellift = 32'd1 */
  wire [3:0] _06283_;
  wire [3:0] _06284_;
  /* cellift = 32'd1 */
  wire [3:0] _06285_;
  wire [3:0] _06286_;
  /* cellift = 32'd1 */
  wire [3:0] _06287_;
  wire [3:0] _06288_;
  /* cellift = 32'd1 */
  wire [3:0] _06289_;
  wire [3:0] _06290_;
  /* cellift = 32'd1 */
  wire [3:0] _06291_;
  wire [3:0] _06292_;
  /* cellift = 32'd1 */
  wire [3:0] _06293_;
  wire [3:0] _06294_;
  /* cellift = 32'd1 */
  wire [3:0] _06295_;
  wire [3:0] _06296_;
  /* cellift = 32'd1 */
  wire [3:0] _06297_;
  wire [3:0] _06298_;
  /* cellift = 32'd1 */
  wire [3:0] _06299_;
  wire [3:0] _06300_;
  /* cellift = 32'd1 */
  wire [3:0] _06301_;
  wire [3:0] _06302_;
  /* cellift = 32'd1 */
  wire [3:0] _06303_;
  /* cellift = 32'd1 */
  wire [3:0] _06304_;
  wire _06305_;
  /* cellift = 32'd1 */
  wire _06306_;
  wire _06307_;
  /* cellift = 32'd1 */
  wire _06308_;
  wire _06309_;
  /* cellift = 32'd1 */
  wire _06310_;
  wire _06311_;
  /* cellift = 32'd1 */
  wire _06312_;
  wire _06313_;
  /* cellift = 32'd1 */
  wire _06314_;
  wire _06315_;
  /* cellift = 32'd1 */
  wire _06316_;
  wire _06317_;
  /* cellift = 32'd1 */
  wire _06318_;
  wire _06319_;
  /* cellift = 32'd1 */
  wire _06320_;
  wire _06321_;
  /* cellift = 32'd1 */
  wire _06322_;
  wire _06323_;
  /* cellift = 32'd1 */
  wire _06324_;
  wire [31:0] _06325_;
  /* cellift = 32'd1 */
  wire [31:0] _06326_;
  wire [31:0] _06327_;
  /* cellift = 32'd1 */
  wire [31:0] _06328_;
  wire [31:0] _06329_;
  /* cellift = 32'd1 */
  wire [31:0] _06330_;
  wire [31:0] _06331_;
  /* cellift = 32'd1 */
  wire [31:0] _06332_;
  wire [31:0] _06333_;
  /* cellift = 32'd1 */
  wire [31:0] _06334_;
  wire [4:0] _06335_;
  /* cellift = 32'd1 */
  wire [4:0] _06336_;
  wire [4:0] _06337_;
  /* cellift = 32'd1 */
  wire [4:0] _06338_;
  wire [4:0] _06339_;
  /* cellift = 32'd1 */
  wire [4:0] _06340_;
  wire [4:0] _06341_;
  /* cellift = 32'd1 */
  wire [4:0] _06342_;
  wire [4:0] _06343_;
  /* cellift = 32'd1 */
  wire [4:0] _06344_;
  wire [4:0] _06345_;
  /* cellift = 32'd1 */
  wire [4:0] _06346_;
  wire [4:0] _06347_;
  /* cellift = 32'd1 */
  wire [4:0] _06348_;
  wire [4:0] _06349_;
  /* cellift = 32'd1 */
  wire [4:0] _06350_;
  wire [4:0] _06351_;
  /* cellift = 32'd1 */
  wire [4:0] _06352_;
  wire [4:0] _06353_;
  /* cellift = 32'd1 */
  wire [4:0] _06354_;
  wire [4:0] _06355_;
  /* cellift = 32'd1 */
  wire [4:0] _06356_;
  wire [4:0] _06357_;
  /* cellift = 32'd1 */
  wire [4:0] _06358_;
  wire [4:0] _06359_;
  /* cellift = 32'd1 */
  wire [4:0] _06360_;
  wire [4:0] _06361_;
  /* cellift = 32'd1 */
  wire [4:0] _06362_;
  wire [4:0] _06363_;
  /* cellift = 32'd1 */
  wire [4:0] _06364_;
  wire [4:0] _06365_;
  /* cellift = 32'd1 */
  wire [4:0] _06366_;
  wire [1:0] _06367_;
  /* cellift = 32'd1 */
  wire [1:0] _06368_;
  wire [1:0] _06369_;
  /* cellift = 32'd1 */
  wire [1:0] _06370_;
  wire [1:0] _06371_;
  /* cellift = 32'd1 */
  wire [1:0] _06372_;
  wire _06373_;
  /* cellift = 32'd1 */
  wire _06374_;
  wire _06375_;
  /* cellift = 32'd1 */
  wire _06376_;
  /* cellift = 32'd1 */
  wire _06377_;
  wire _06378_;
  /* cellift = 32'd1 */
  wire _06379_;
  wire _06380_;
  /* cellift = 32'd1 */
  wire _06381_;
  wire _06382_;
  /* cellift = 32'd1 */
  wire _06383_;
  wire _06384_;
  /* cellift = 32'd1 */
  wire _06385_;
  wire _06386_;
  /* cellift = 32'd1 */
  wire _06387_;
  wire _06388_;
  /* cellift = 32'd1 */
  wire _06389_;
  wire _06390_;
  /* cellift = 32'd1 */
  wire _06391_;
  wire _06392_;
  /* cellift = 32'd1 */
  wire _06393_;
  wire [4:0] _06394_;
  /* cellift = 32'd1 */
  wire [4:0] _06395_;
  wire [4:0] _06396_;
  /* cellift = 32'd1 */
  wire [4:0] _06397_;
  wire [4:0] _06398_;
  /* cellift = 32'd1 */
  wire [4:0] _06399_;
  wire [4:0] _06400_;
  /* cellift = 32'd1 */
  wire [4:0] _06401_;
  wire [4:0] _06402_;
  /* cellift = 32'd1 */
  wire [4:0] _06403_;
  wire [4:0] _06404_;
  /* cellift = 32'd1 */
  wire [4:0] _06405_;
  wire [4:0] _06406_;
  /* cellift = 32'd1 */
  wire [4:0] _06407_;
  wire [4:0] _06408_;
  /* cellift = 32'd1 */
  wire [4:0] _06409_;
  wire [4:0] _06410_;
  /* cellift = 32'd1 */
  wire [4:0] _06411_;
  wire [4:0] _06412_;
  /* cellift = 32'd1 */
  wire [4:0] _06413_;
  wire [2:0] _06414_;
  /* cellift = 32'd1 */
  wire [2:0] _06415_;
  wire [2:0] _06416_;
  /* cellift = 32'd1 */
  wire [2:0] _06417_;
  wire [2:0] _06418_;
  /* cellift = 32'd1 */
  wire [2:0] _06419_;
  wire [2:0] _06420_;
  /* cellift = 32'd1 */
  wire [2:0] _06421_;
  wire [2:0] _06422_;
  /* cellift = 32'd1 */
  wire [2:0] _06423_;
  wire [2:0] _06424_;
  /* cellift = 32'd1 */
  wire [2:0] _06425_;
  wire [2:0] _06426_;
  /* cellift = 32'd1 */
  wire [2:0] _06427_;
  wire [2:0] _06428_;
  /* cellift = 32'd1 */
  wire [2:0] _06429_;
  wire [2:0] _06430_;
  /* cellift = 32'd1 */
  wire [2:0] _06431_;
  wire [2:0] _06432_;
  /* cellift = 32'd1 */
  wire [2:0] _06433_;
  wire [2:0] _06434_;
  /* cellift = 32'd1 */
  wire [2:0] _06435_;
  wire [2:0] _06436_;
  /* cellift = 32'd1 */
  wire [2:0] _06437_;
  wire [3:0] _06438_;
  /* cellift = 32'd1 */
  wire [3:0] _06439_;
  wire [3:0] _06440_;
  /* cellift = 32'd1 */
  wire [3:0] _06441_;
  wire [3:0] _06442_;
  /* cellift = 32'd1 */
  wire [3:0] _06443_;
  wire [5:0] _06444_;
  /* cellift = 32'd1 */
  wire [5:0] _06445_;
  wire [5:0] _06446_;
  /* cellift = 32'd1 */
  wire [5:0] _06447_;
  wire [5:0] _06448_;
  /* cellift = 32'd1 */
  wire [5:0] _06449_;
  wire [5:0] _06450_;
  /* cellift = 32'd1 */
  wire [5:0] _06451_;
  wire [5:0] _06452_;
  /* cellift = 32'd1 */
  wire [5:0] _06453_;
  wire [5:0] _06454_;
  /* cellift = 32'd1 */
  wire [5:0] _06455_;
  wire [5:0] _06456_;
  /* cellift = 32'd1 */
  wire [5:0] _06457_;
  wire [5:0] _06458_;
  /* cellift = 32'd1 */
  wire [5:0] _06459_;
  wire [5:0] _06460_;
  /* cellift = 32'd1 */
  wire [5:0] _06461_;
  wire [5:0] _06462_;
  /* cellift = 32'd1 */
  wire [5:0] _06463_;
  wire [5:0] _06464_;
  /* cellift = 32'd1 */
  wire [5:0] _06465_;
  wire [5:0] _06466_;
  /* cellift = 32'd1 */
  wire [5:0] _06467_;
  wire [5:0] _06468_;
  /* cellift = 32'd1 */
  wire [5:0] _06469_;
  wire [31:0] _06470_;
  /* cellift = 32'd1 */
  wire [31:0] _06471_;
  wire [31:0] _06472_;
  /* cellift = 32'd1 */
  wire [31:0] _06473_;
  wire [31:0] _06474_;
  /* cellift = 32'd1 */
  wire [31:0] _06475_;
  wire [3:0] _06476_;
  /* cellift = 32'd1 */
  wire [3:0] _06477_;
  wire [31:0] _06478_;
  /* cellift = 32'd1 */
  wire [31:0] _06479_;
  wire _06480_;
  /* cellift = 32'd1 */
  wire _06481_;
  wire [3:0] _06482_;
  /* src = "generated/out/vanilla.sv:1050.7-1050.34" */
  wire _06483_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1050.7-1050.34" */
  wire _06484_;
  /* src = "generated/out/vanilla.sv:1052.7-1052.35" */
  wire _06485_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1052.7-1052.35" */
  wire _06486_;
  /* src = "generated/out/vanilla.sv:1054.7-1054.36" */
  wire _06487_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1054.7-1054.36" */
  wire _06488_;
  /* src = "generated/out/vanilla.sv:1056.7-1056.36" */
  wire _06489_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1056.7-1056.36" */
  wire _06490_;
  /* src = "generated/out/vanilla.sv:1058.7-1058.34" */
  wire _06491_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1058.7-1058.34" */
  wire _06492_;
  /* src = "generated/out/vanilla.sv:1060.7-1060.35" */
  wire _06493_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1060.7-1060.35" */
  wire _06494_;
  /* src = "generated/out/vanilla.sv:1062.7-1062.35" */
  wire _06495_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1062.7-1062.35" */
  wire _06496_;
  /* src = "generated/out/vanilla.sv:1064.7-1064.35" */
  wire _06497_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1064.7-1064.35" */
  wire _06498_;
  /* src = "generated/out/vanilla.sv:1579.10-1579.21" */
  wire _06499_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1579.10-1579.21" */
  wire _06500_;
  /* src = "generated/out/vanilla.sv:1669.9-1669.26" */
  wire _06501_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1669.9-1669.26" */
  wire _06502_;
  /* src = "generated/out/vanilla.sv:1674.9-1674.26" */
  wire _06503_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1674.9-1674.26" */
  wire _06504_;
  /* src = "generated/out/vanilla.sv:1792.23-1792.51" */
  wire _06505_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1792.23-1792.51" */
  wire _06506_;
  /* src = "generated/out/vanilla.sv:1792.58-1792.84" */
  wire _06507_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1792.58-1792.84" */
  wire _06508_;
  /* src = "generated/out/vanilla.sv:1793.8-1793.35" */
  wire _06509_;
  /* src = "generated/out/vanilla.sv:1797.8-1797.35" */
  wire _06510_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1797.8-1797.35" */
  wire _06511_;
  /* src = "generated/out/vanilla.sv:1801.8-1801.35" */
  wire _06512_;
  /* src = "generated/out/vanilla.sv:1805.8-1805.35" */
  wire _06513_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1805.8-1805.35" */
  wire _06514_;
  /* src = "generated/out/vanilla.sv:372.12-372.40" */
  wire _06515_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:372.12-372.40" */
  wire _06516_;
  /* src = "generated/out/vanilla.sv:379.12-379.45" */
  wire _06517_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:379.12-379.45" */
  wire _06518_;
  /* src = "generated/out/vanilla.sv:383.12-383.45" */
  wire _06519_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:383.12-383.45" */
  wire _06520_;
  /* src = "generated/out/vanilla.sv:387.12-387.45" */
  wire _06521_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:387.12-387.45" */
  wire _06522_;
  /* src = "generated/out/vanilla.sv:391.12-391.46" */
  wire _06523_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:391.12-391.46" */
  wire _06524_;
  /* src = "generated/out/vanilla.sv:392.13-392.44" */
  wire _06525_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:392.13-392.44" */
  wire _06526_;
  /* src = "generated/out/vanilla.sv:394.13-394.44" */
  wire _06527_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:394.13-394.44" */
  wire _06528_;
  /* src = "generated/out/vanilla.sv:396.13-396.44" */
  wire _06529_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:396.13-396.44" */
  wire _06530_;
  /* src = "generated/out/vanilla.sv:398.13-398.44" */
  wire _06531_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:398.13-398.44" */
  wire _06532_;
  /* src = "generated/out/vanilla.sv:423.45-423.72" */
  wire _06533_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:423.45-423.72" */
  wire _06534_;
  /* src = "generated/out/vanilla.sv:457.9-457.23" */
  wire _06535_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:457.9-457.23" */
  wire _06536_;
  /* src = "generated/out/vanilla.sv:457.29-457.43" */
  wire _06537_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:457.29-457.43" */
  wire _06538_;
  /* src = "generated/out/vanilla.sv:797.17-797.53" */
  wire _06539_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:797.17-797.53" */
  wire _06540_;
  /* src = "generated/out/vanilla.sv:798.19-798.55" */
  wire _06541_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:798.19-798.55" */
  wire _06542_;
  /* src = "generated/out/vanilla.sv:799.17-799.53" */
  wire _06543_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:799.17-799.53" */
  wire _06544_;
  /* src = "generated/out/vanilla.sv:800.19-800.55" */
  wire _06545_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:800.19-800.55" */
  wire _06546_;
  /* src = "generated/out/vanilla.sv:800.61-800.95" */
  wire _06547_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:800.61-800.95" */
  wire _06548_;
  /* src = "generated/out/vanilla.sv:803.36-803.72" */
  wire _06549_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:803.36-803.72" */
  wire _06550_;
  /* src = "generated/out/vanilla.sv:804.27-804.63" */
  wire _06551_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:804.27-804.63" */
  wire _06552_;
  /* src = "generated/out/vanilla.sv:805.19-805.55" */
  wire _06553_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:805.19-805.55" */
  wire _06554_;
  /* src = "generated/out/vanilla.sv:806.22-806.58" */
  wire _06555_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:806.22-806.58" */
  wire _06556_;
  /* src = "generated/out/vanilla.sv:807.22-807.58" */
  wire _06557_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:807.22-807.58" */
  wire _06558_;
  /* src = "generated/out/vanilla.sv:951.50-951.78" */
  wire _06559_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:951.50-951.78" */
  wire _06560_;
  /* src = "generated/out/vanilla.sv:952.50-952.78" */
  wire _06561_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:952.50-952.78" */
  wire _06562_;
  /* src = "generated/out/vanilla.sv:953.50-953.78" */
  wire _06563_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:953.50-953.78" */
  wire _06564_;
  /* src = "generated/out/vanilla.sv:954.50-954.78" */
  wire _06565_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:954.50-954.78" */
  wire _06566_;
  /* src = "generated/out/vanilla.sv:955.51-955.79" */
  wire _06567_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:955.51-955.79" */
  wire _06568_;
  /* src = "generated/out/vanilla.sv:956.51-956.79" */
  wire _06569_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:956.51-956.79" */
  wire _06570_;
  /* src = "generated/out/vanilla.sv:959.40-959.68" */
  wire _06571_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:959.40-959.68" */
  wire _06572_;
  /* src = "generated/out/vanilla.sv:967.38-967.66" */
  wire _06573_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:967.38-967.66" */
  wire _06574_;
  /* src = "generated/out/vanilla.sv:971.73-971.105" */
  wire _06575_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:971.73-971.105" */
  wire _06576_;
  /* src = "generated/out/vanilla.sv:973.73-973.105" */
  wire _06577_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:973.73-973.105" */
  wire _06578_;
  /* src = "generated/out/vanilla.sv:984.25-984.55" */
  wire _06579_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:984.25-984.55" */
  wire _06580_;
  /* src = "generated/out/vanilla.sv:984.61-984.97" */
  wire _06581_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:984.61-984.97" */
  wire _06582_;
  /* src = "generated/out/vanilla.sv:984.174-984.210" */
  wire _06583_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:984.174-984.210" */
  wire _06584_;
  /* src = "generated/out/vanilla.sv:985.63-985.99" */
  wire _06585_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:985.63-985.99" */
  wire _06586_;
  /* src = "generated/out/vanilla.sv:985.176-985.212" */
  wire _06587_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:985.176-985.212" */
  wire _06588_;
  /* src = "generated/out/vanilla.sv:986.60-986.96" */
  wire _06589_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:986.60-986.96" */
  wire _06590_;
  /* src = "generated/out/vanilla.sv:987.62-987.98" */
  wire _06591_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:987.62-987.98" */
  wire _06592_;
  /* src = "generated/out/vanilla.sv:988.131-988.160" */
  wire _06593_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:988.131-988.160" */
  wire _06594_;
  /* src = "generated/out/vanilla.sv:989.20-989.50" */
  wire _06595_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:989.20-989.50" */
  wire _06596_;
  /* src = "generated/out/vanilla.sv:1584.35-1584.46" */
  wire _06597_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1584.35-1584.46" */
  wire _06598_;
  /* src = "generated/out/vanilla.sv:1080.20-1080.51" */
  wire _06599_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1080.20-1080.51" */
  wire _06600_;
  /* src = "generated/out/vanilla.sv:1166.5-1166.37" */
  wire _06601_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1166.5-1166.37" */
  wire _06602_;
  /* src = "generated/out/vanilla.sv:1181.8-1181.31" */
  wire _06603_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1181.8-1181.31" */
  wire _06604_;
  /* src = "generated/out/vanilla.sv:1181.7-1181.46" */
  wire _06605_;
  /* src = "generated/out/vanilla.sv:1214.9-1214.29" */
  wire _06606_;
  /* src = "generated/out/vanilla.sv:1214.8-1214.48" */
  wire _06607_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1234.22-1234.46" */
  wire _06608_;
  /* src = "generated/out/vanilla.sv:1275.22-1275.53" */
  wire _06609_;
  /* src = "generated/out/vanilla.sv:1346.27-1346.55" */
  wire _06610_;
  /* src = "generated/out/vanilla.sv:1374.19-1374.72" */
  wire _06611_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1374.19-1374.72" */
  wire _06612_;
  /* src = "generated/out/vanilla.sv:1454.7-1454.41" */
  wire _06613_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1454.7-1454.41" */
  wire _06614_;
  /* src = "generated/out/vanilla.sv:1621.11-1621.39" */
  wire _06615_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1621.11-1621.39" */
  wire _06616_;
  /* src = "generated/out/vanilla.sv:1668.7-1668.67" */
  wire _06617_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1668.7-1668.67" */
  wire _06618_;
  /* src = "generated/out/vanilla.sv:1669.8-1669.50" */
  wire _06619_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1669.8-1669.50" */
  wire _06620_;
  /* src = "generated/out/vanilla.sv:1674.8-1674.48" */
  wire _06621_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1674.8-1674.48" */
  wire _06622_;
  /* src = "generated/out/vanilla.sv:1680.8-1680.50" */
  wire _06623_;
  /* src = "generated/out/vanilla.sv:1680.7-1680.98" */
  wire _06624_;
  /* src = "generated/out/vanilla.sv:1715.18-1715.54" */
  wire _06625_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1715.18-1715.54" */
  wire _06626_;
  /* src = "generated/out/vanilla.sv:1774.13-1774.43" */
  wire _06627_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1774.13-1774.43" */
  wire _06628_;
  /* src = "generated/out/vanilla.sv:1792.8-1792.52" */
  wire _06629_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1792.8-1792.52" */
  wire _06630_;
  /* src = "generated/out/vanilla.sv:1792.7-1792.85" */
  wire _06631_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1792.7-1792.85" */
  wire _06632_;
  /* src = "generated/out/vanilla.sv:286.28-286.79" */
  wire _06633_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:286.28-286.79" */
  wire _06634_;
  /* src = "generated/out/vanilla.sv:286.27-286.94" */
  wire _06635_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:286.27-286.94" */
  wire _06636_;
  /* src = "generated/out/vanilla.sv:293.42-293.102" */
  wire _06637_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:293.42-293.102" */
  wire _06638_;
  /* src = "generated/out/vanilla.sv:294.49-294.96" */
  wire _06639_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:294.49-294.96" */
  wire _06640_;
  /* src = "generated/out/vanilla.sv:296.32-296.54" */
  wire _06641_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:296.32-296.54" */
  wire _06642_;
  /* src = "generated/out/vanilla.sv:296.31-296.107" */
  wire _06643_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:296.31-296.107" */
  wire _06644_;
  /* src = "generated/out/vanilla.sv:296.113-296.139" */
  wire _06645_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:296.113-296.139" */
  wire _06646_;
  /* src = "generated/out/vanilla.sv:296.19-296.141" */
  wire _06647_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:296.19-296.141" */
  wire _06648_;
  /* src = "generated/out/vanilla.sv:296.169-296.205" */
  wire _06649_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:296.169-296.205" */
  wire _06650_;
  /* src = "generated/out/vanilla.sv:297.25-297.45" */
  wire _06651_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:297.25-297.45" */
  wire _06652_;
  /* src = "generated/out/vanilla.sv:298.36-298.82" */
  wire _06653_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:298.36-298.82" */
  wire _06654_;
  /* src = "generated/out/vanilla.sv:298.35-298.138" */
  wire _06655_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:298.35-298.138" */
  wire _06656_;
  /* src = "generated/out/vanilla.sv:298.145-298.260" */
  wire _06657_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:298.145-298.260" */
  wire _06658_;
  /* src = "generated/out/vanilla.sv:298.144-298.288" */
  wire _06659_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:298.144-298.288" */
  wire _06660_;
  /* src = "generated/out/vanilla.sv:310.22-310.45" */
  wire _06661_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:310.22-310.45" */
  wire _06662_;
  /* src = "generated/out/vanilla.sv:344.7-344.72" */
  wire _06663_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:344.7-344.72" */
  wire _06664_;
  /* src = "generated/out/vanilla.sv:423.12-423.73" */
  wire _06665_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:423.12-423.73" */
  wire _06666_;
  /* src = "generated/out/vanilla.sv:427.12-427.73" */
  wire _06667_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:427.12-427.73" */
  wire _06668_;
  /* src = "generated/out/vanilla.sv:431.13-431.75" */
  wire _06669_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:431.13-431.75" */
  wire _06670_;
  /* src = "generated/out/vanilla.sv:431.12-431.109" */
  wire _06671_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:431.12-431.109" */
  wire _06672_;
  /* src = "generated/out/vanilla.sv:435.12-435.73" */
  wire _06673_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:435.12-435.73" */
  wire _06674_;
  /* src = "generated/out/vanilla.sv:800.18-800.96" */
  wire _06675_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:800.18-800.96" */
  wire _06676_;
  /* src = "generated/out/vanilla.sv:817.8-817.59" */
  wire _06677_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:817.8-817.59" */
  wire _06678_;
  /* src = "generated/out/vanilla.sv:871.13-871.61" */
  wire _06679_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:871.13-871.61" */
  wire _06680_;
  /* src = "generated/out/vanilla.sv:917.14-917.76" */
  wire _06681_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:917.14-917.76" */
  wire _06682_;
  /* src = "generated/out/vanilla.sv:917.13-917.110" */
  wire _06683_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:917.13-917.110" */
  wire _06684_;
  /* src = "generated/out/vanilla.sv:949.7-949.49" */
  wire _06685_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:949.7-949.49" */
  wire _06686_;
  /* src = "generated/out/vanilla.sv:951.17-951.79" */
  wire _06687_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:951.17-951.79" */
  wire _06688_;
  /* src = "generated/out/vanilla.sv:952.17-952.79" */
  wire _06689_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:952.17-952.79" */
  wire _06690_;
  /* src = "generated/out/vanilla.sv:953.17-953.79" */
  wire _06691_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:953.17-953.79" */
  wire _06692_;
  /* src = "generated/out/vanilla.sv:954.17-954.79" */
  wire _06693_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:954.17-954.79" */
  wire _06694_;
  /* src = "generated/out/vanilla.sv:955.18-955.80" */
  wire _06695_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:955.18-955.80" */
  wire _06696_;
  /* src = "generated/out/vanilla.sv:956.18-956.80" */
  wire _06697_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:956.18-956.80" */
  wire _06698_;
  /* src = "generated/out/vanilla.sv:957.16-957.69" */
  wire _06699_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:957.16-957.69" */
  wire _06700_;
  /* src = "generated/out/vanilla.sv:958.16-958.69" */
  wire _06701_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:958.16-958.69" */
  wire _06702_;
  /* src = "generated/out/vanilla.sv:959.16-959.69" */
  wire _06703_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:959.16-959.69" */
  wire _06704_;
  /* src = "generated/out/vanilla.sv:960.17-960.70" */
  wire _06705_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:960.17-960.70" */
  wire _06706_;
  /* src = "generated/out/vanilla.sv:961.17-961.70" */
  wire _06707_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:961.17-961.70" */
  wire _06708_;
  /* src = "generated/out/vanilla.sv:962.16-962.61" */
  wire _06709_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:962.16-962.61" */
  wire _06710_;
  /* src = "generated/out/vanilla.sv:963.16-963.61" */
  wire _06711_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:963.16-963.61" */
  wire _06712_;
  /* src = "generated/out/vanilla.sv:964.16-964.61" */
  wire _06713_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:964.16-964.61" */
  wire _06714_;
  /* src = "generated/out/vanilla.sv:965.18-965.66" */
  wire _06715_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:965.18-965.66" */
  wire _06716_;
  /* src = "generated/out/vanilla.sv:966.18-966.66" */
  wire _06717_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:966.18-966.66" */
  wire _06718_;
  /* src = "generated/out/vanilla.sv:967.19-967.67" */
  wire _06719_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:967.19-967.67" */
  wire _06720_;
  /* src = "generated/out/vanilla.sv:968.18-968.66" */
  wire _06721_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:968.18-968.66" */
  wire _06722_;
  /* src = "generated/out/vanilla.sv:969.17-969.65" */
  wire _06723_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:969.17-969.65" */
  wire _06724_;
  /* src = "generated/out/vanilla.sv:970.18-970.66" */
  wire _06725_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:970.18-970.66" */
  wire _06726_;
  /* src = "generated/out/vanilla.sv:971.19-971.67" */
  wire _06727_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:971.19-971.67" */
  wire _06728_;
  /* src = "generated/out/vanilla.sv:971.18-971.106" */
  wire _06729_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:971.18-971.106" */
  wire _06730_;
  /* src = "generated/out/vanilla.sv:972.19-972.67" */
  wire _06731_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:972.19-972.67" */
  wire _06732_;
  /* src = "generated/out/vanilla.sv:972.18-972.106" */
  wire _06733_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:972.18-972.106" */
  wire _06734_;
  /* src = "generated/out/vanilla.sv:973.18-973.106" */
  wire _06735_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:973.18-973.106" */
  wire _06736_;
  /* src = "generated/out/vanilla.sv:974.18-974.66" */
  wire _06737_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:974.18-974.66" */
  wire _06738_;
  /* src = "generated/out/vanilla.sv:974.17-974.105" */
  wire _06739_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:974.17-974.105" */
  wire _06740_;
  /* src = "generated/out/vanilla.sv:975.17-975.105" */
  wire _06741_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:975.17-975.105" */
  wire _06742_;
  /* src = "generated/out/vanilla.sv:976.18-976.66" */
  wire _06743_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:976.18-976.66" */
  wire _06744_;
  /* src = "generated/out/vanilla.sv:976.17-976.105" */
  wire _06745_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:976.17-976.105" */
  wire _06746_;
  /* src = "generated/out/vanilla.sv:977.18-977.66" */
  wire _06747_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:977.18-977.66" */
  wire _06748_;
  /* src = "generated/out/vanilla.sv:977.17-977.105" */
  wire _06749_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:977.17-977.105" */
  wire _06750_;
  /* src = "generated/out/vanilla.sv:978.19-978.67" */
  wire _06751_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:978.19-978.67" */
  wire _06752_;
  /* src = "generated/out/vanilla.sv:978.18-978.106" */
  wire _06753_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:978.18-978.106" */
  wire _06754_;
  /* src = "generated/out/vanilla.sv:979.18-979.66" */
  wire _06755_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:979.18-979.66" */
  wire _06756_;
  /* src = "generated/out/vanilla.sv:979.17-979.105" */
  wire _06757_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:979.17-979.105" */
  wire _06758_;
  /* src = "generated/out/vanilla.sv:980.18-980.66" */
  wire _06759_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:980.18-980.66" */
  wire _06760_;
  /* src = "generated/out/vanilla.sv:980.17-980.105" */
  wire _06761_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:980.17-980.105" */
  wire _06762_;
  /* src = "generated/out/vanilla.sv:981.17-981.105" */
  wire _06763_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:981.17-981.105" */
  wire _06764_;
  /* src = "generated/out/vanilla.sv:982.17-982.65" */
  wire _06765_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:982.17-982.65" */
  wire _06766_;
  /* src = "generated/out/vanilla.sv:982.16-982.104" */
  wire _06767_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:982.16-982.104" */
  wire _06768_;
  /* src = "generated/out/vanilla.sv:983.18-983.66" */
  wire _06769_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:983.18-983.66" */
  wire _06770_;
  /* src = "generated/out/vanilla.sv:983.17-983.105" */
  wire _06771_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:983.17-983.105" */
  wire _06772_;
  /* src = "generated/out/vanilla.sv:984.24-984.98" */
  wire _06773_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:984.24-984.98" */
  wire _06774_;
  /* src = "generated/out/vanilla.sv:984.23-984.130" */
  wire _06775_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:984.23-984.130" */
  wire _06776_;
  /* src = "generated/out/vanilla.sv:984.137-984.211" */
  wire _06777_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:984.137-984.211" */
  wire _06778_;
  /* src = "generated/out/vanilla.sv:984.136-984.243" */
  wire _06779_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:984.136-984.243" */
  wire _06780_;
  /* src = "generated/out/vanilla.sv:984.21-984.264" */
  wire _06781_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:984.21-984.264" */
  wire _06782_;
  /* src = "generated/out/vanilla.sv:985.26-985.100" */
  wire _06783_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:985.26-985.100" */
  wire _06784_;
  /* src = "generated/out/vanilla.sv:985.25-985.132" */
  wire _06785_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:985.25-985.132" */
  wire _06786_;
  /* src = "generated/out/vanilla.sv:985.139-985.213" */
  wire _06787_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:985.139-985.213" */
  wire _06788_;
  /* src = "generated/out/vanilla.sv:985.138-985.245" */
  wire _06789_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:985.138-985.245" */
  wire _06790_;
  /* src = "generated/out/vanilla.sv:985.23-985.266" */
  wire _06791_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:985.23-985.266" */
  wire _06792_;
  /* src = "generated/out/vanilla.sv:986.23-986.97" */
  wire _06793_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:986.23-986.97" */
  wire _06794_;
  /* src = "generated/out/vanilla.sv:986.22-986.129" */
  wire _06795_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:986.22-986.129" */
  wire _06796_;
  /* src = "generated/out/vanilla.sv:987.25-987.99" */
  wire _06797_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:987.25-987.99" */
  wire _06798_;
  /* src = "generated/out/vanilla.sv:987.24-987.131" */
  wire _06799_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:987.24-987.131" */
  wire _06800_;
  /* src = "generated/out/vanilla.sv:988.28-988.83" */
  wire _06801_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:988.28-988.83" */
  wire _06802_;
  /* src = "generated/out/vanilla.sv:988.27-988.106" */
  wire _06803_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:988.27-988.106" */
  wire _06804_;
  /* src = "generated/out/vanilla.sv:989.19-989.74" */
  wire _06805_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:989.19-989.74" */
  wire _06806_;
  /* src = "generated/out/vanilla.sv:994.185-994.253" */
  wire _06807_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:994.185-994.253" */
  wire _06808_;
  /* src = "generated/out/vanilla.sv:994.115-994.183" */
  wire _06809_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:994.115-994.183" */
  wire _06810_;
  /* src = "generated/out/vanilla.sv:994.45-994.113" */
  wire _06811_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:994.45-994.113" */
  wire _06812_;
  /* src = "generated/out/vanilla.sv:994.25-994.254" */
  wire _06813_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:994.25-994.254" */
  wire _06814_;
  /* src = "generated/out/vanilla.sv:995.60-995.259" */
  wire _06815_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:995.60-995.259" */
  wire _06816_;
  /* src = "generated/out/vanilla.sv:996.22-996.251" */
  wire _06817_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:996.22-996.251" */
  wire _06818_;
  /* src = "generated/out/vanilla.sv:0.0-0.0" */
  wire _06819_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:0.0-0.0" */
  wire _06820_;
  /* src = "generated/out/vanilla.sv:0.0-0.0" */
  wire _06821_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:0.0-0.0" */
  wire _06822_;
  /* src = "generated/out/vanilla.sv:1009.7-1009.14" */
  wire _06823_;
  /* src = "generated/out/vanilla.sv:1124.27-1124.34" */
  wire _06824_;
  /* src = "generated/out/vanilla.sv:1125.27-1125.35" */
  wire _06825_;
  /* src = "generated/out/vanilla.sv:1126.28-1126.36" */
  wire _06826_;
  /* src = "generated/out/vanilla.sv:1166.22-1166.37" */
  wire _06827_;
  /* src = "generated/out/vanilla.sv:1214.34-1214.48" */
  wire _06828_;
  /* src = "generated/out/vanilla.sv:1220.20-1220.41" */
  wire _06829_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1220.20-1220.41" */
  wire _06830_;
  /* src = "generated/out/vanilla.sv:1454.30-1454.41" */
  wire _06831_;
  /* src = "generated/out/vanilla.sv:1606.10-1606.26" */
  wire _06832_;
  /* src = "generated/out/vanilla.sv:286.99-286.117" */
  wire _06833_;
  /* src = "generated/out/vanilla.sv:293.107-293.134" */
  wire _06834_;
  /* src = "generated/out/vanilla.sv:296.147-296.164" */
  wire _06835_;
  /* src = "generated/out/vanilla.sv:297.35-297.45" */
  wire _06836_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:297.35-297.45" */
  wire _06837_;
  /* src = "generated/out/vanilla.sv:298.36-298.68" */
  wire _06838_;
  /* src = "generated/out/vanilla.sv:310.35-310.45" */
  wire _06839_;
  /* src = "generated/out/vanilla.sv:871.13-871.35" */
  wire _06840_;
  /* src = "generated/out/vanilla.sv:871.39-871.61" */
  wire _06841_;
  /* src = "generated/out/vanilla.sv:949.26-949.49" */
  wire _06842_;
  /* src = "generated/out/vanilla.sv:988.64-988.83" */
  wire _06843_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:988.64-988.83" */
  wire _06844_;
  /* src = "generated/out/vanilla.sv:988.88-988.106" */
  wire _06845_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:988.88-988.106" */
  wire _06846_;
  /* src = "generated/out/vanilla.sv:989.55-989.74" */
  wire _06847_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:989.55-989.74" */
  wire _06848_;
  /* src = "generated/out/vanilla.sv:1115.25-1115.48" */
  wire _06849_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1115.25-1115.48" */
  wire _06850_;
  /* src = "generated/out/vanilla.sv:1135.4-1135.27" */
  wire _06851_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1135.4-1135.27" */
  wire _06852_;
  /* src = "generated/out/vanilla.sv:1136.4-1136.25" */
  wire _06853_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1136.4-1136.25" */
  wire _06854_;
  /* src = "generated/out/vanilla.sv:1137.4-1137.27" */
  wire _06855_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1137.4-1137.27" */
  wire _06856_;
  /* src = "generated/out/vanilla.sv:1138.23-1138.46" */
  wire _06857_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1138.23-1138.46" */
  wire _06858_;
  /* src = "generated/out/vanilla.sv:1139.25-1139.48" */
  wire _06859_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1139.25-1139.48" */
  wire _06860_;
  /* src = "generated/out/vanilla.sv:1148.8-1148.35" */
  wire _06861_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1148.8-1148.35" */
  wire _06862_;
  /* src = "generated/out/vanilla.sv:1148.7-1148.47" */
  wire _06863_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1148.7-1148.47" */
  wire _06864_;
  /* src = "generated/out/vanilla.sv:1606.10-1606.38" */
  wire _06865_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1606.10-1606.38" */
  wire _06866_;
  /* src = "generated/out/vanilla.sv:1634.9-1634.30" */
  wire _06867_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1634.9-1634.30" */
  wire _06868_;
  /* src = "generated/out/vanilla.sv:1635.9-1635.30" */
  wire _06869_;
  /* src = "generated/out/vanilla.sv:1668.38-1668.66" */
  wire _06870_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1668.38-1668.66" */
  wire _06871_;
  /* src = "generated/out/vanilla.sv:1687.7-1687.26" */
  wire _06872_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1687.7-1687.26" */
  wire _06873_;
  /* src = "generated/out/vanilla.sv:1715.29-1715.53" */
  wire _06874_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1715.29-1715.53" */
  wire _06875_;
  /* src = "generated/out/vanilla.sv:296.61-296.89" */
  wire _06876_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:296.61-296.89" */
  wire _06877_;
  /* src = "generated/out/vanilla.sv:296.60-296.106" */
  wire _06878_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:296.60-296.106" */
  wire _06879_;
  /* src = "generated/out/vanilla.sv:296.30-296.140" */
  wire _06880_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:296.30-296.140" */
  wire _06881_;
  /* src = "generated/out/vanilla.sv:296.147-296.206" */
  wire _06882_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:296.147-296.206" */
  wire _06883_;
  /* src = "generated/out/vanilla.sv:298.88-298.137" */
  wire _06884_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:298.88-298.137" */
  wire _06885_;
  /* src = "generated/out/vanilla.sv:298.34-298.289" */
  wire _06886_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:298.34-298.289" */
  wire _06887_;
  /* src = "generated/out/vanilla.sv:461.7-461.22" */
  wire _06888_;
  /* src = "generated/out/vanilla.sv:464.8-464.28" */
  wire _06889_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:464.8-464.28" */
  wire _06890_;
  /* src = "generated/out/vanilla.sv:470.8-470.35" */
  wire _06891_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:470.8-470.35" */
  wire _06892_;
  /* src = "generated/out/vanilla.sv:506.13-506.50" */
  wire _06893_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:506.13-506.50" */
  wire _06894_;
  /* src = "generated/out/vanilla.sv:859.13-859.60" */
  wire _06895_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:859.13-859.60" */
  wire _06896_;
  /* src = "generated/out/vanilla.sv:988.26-988.162" */
  wire _06897_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:988.26-988.162" */
  wire _06898_;
  /* src = "generated/out/vanilla.sv:995.45-995.260" */
  wire _06899_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:995.45-995.260" */
  wire _06900_;
  wire [31:0] _06901_;
  /* cellift = 32'd1 */
  wire [31:0] _06902_;
  wire [31:0] _06903_;
  /* cellift = 32'd1 */
  wire [31:0] _06904_;
  wire [31:0] _06905_;
  /* cellift = 32'd1 */
  wire [31:0] _06906_;
  wire [31:0] _06907_;
  /* cellift = 32'd1 */
  wire [31:0] _06908_;
  wire [31:0] _06909_;
  /* cellift = 32'd1 */
  wire [31:0] _06910_;
  wire [31:0] _06911_;
  /* cellift = 32'd1 */
  wire [31:0] _06912_;
  wire [31:0] _06913_;
  /* cellift = 32'd1 */
  wire [31:0] _06914_;
  wire [31:0] _06915_;
  /* cellift = 32'd1 */
  wire [31:0] _06916_;
  wire [31:0] _06917_;
  /* cellift = 32'd1 */
  wire [31:0] _06918_;
  wire [31:0] _06919_;
  /* cellift = 32'd1 */
  wire [31:0] _06920_;
  wire [31:0] _06921_;
  /* cellift = 32'd1 */
  wire [31:0] _06922_;
  wire [31:0] _06923_;
  /* cellift = 32'd1 */
  wire [31:0] _06924_;
  wire [31:0] _06925_;
  /* cellift = 32'd1 */
  wire [31:0] _06926_;
  wire [31:0] _06927_;
  /* cellift = 32'd1 */
  wire [31:0] _06928_;
  wire [31:0] _06929_;
  /* cellift = 32'd1 */
  wire [31:0] _06930_;
  wire [31:0] _06931_;
  /* cellift = 32'd1 */
  wire [31:0] _06932_;
  wire [31:0] _06933_;
  /* cellift = 32'd1 */
  wire [31:0] _06934_;
  wire [31:0] _06935_;
  /* cellift = 32'd1 */
  wire [31:0] _06936_;
  wire [31:0] _06937_;
  /* cellift = 32'd1 */
  wire [31:0] _06938_;
  wire [31:0] _06939_;
  /* cellift = 32'd1 */
  wire [31:0] _06940_;
  wire [31:0] _06941_;
  /* cellift = 32'd1 */
  wire [31:0] _06942_;
  wire [31:0] _06943_;
  /* cellift = 32'd1 */
  wire [31:0] _06944_;
  wire [31:0] _06945_;
  /* cellift = 32'd1 */
  wire [31:0] _06946_;
  wire [31:0] _06947_;
  /* cellift = 32'd1 */
  wire [31:0] _06948_;
  wire [31:0] _06949_;
  /* cellift = 32'd1 */
  wire [31:0] _06950_;
  wire [31:0] _06951_;
  /* cellift = 32'd1 */
  wire [31:0] _06952_;
  wire [31:0] _06953_;
  /* cellift = 32'd1 */
  wire [31:0] _06954_;
  wire [31:0] _06955_;
  /* cellift = 32'd1 */
  wire [31:0] _06956_;
  wire [31:0] _06957_;
  /* cellift = 32'd1 */
  wire [31:0] _06958_;
  wire [31:0] _06959_;
  /* cellift = 32'd1 */
  wire [31:0] _06960_;
  wire [31:0] _06961_;
  /* cellift = 32'd1 */
  wire [31:0] _06962_;
  wire [31:0] _06963_;
  /* cellift = 32'd1 */
  wire [31:0] _06964_;
  wire [31:0] _06965_;
  /* cellift = 32'd1 */
  wire [31:0] _06966_;
  wire [31:0] _06967_;
  /* cellift = 32'd1 */
  wire [31:0] _06968_;
  wire [31:0] _06969_;
  /* cellift = 32'd1 */
  wire [31:0] _06970_;
  wire [31:0] _06971_;
  /* cellift = 32'd1 */
  wire [31:0] _06972_;
  wire [31:0] _06973_;
  /* cellift = 32'd1 */
  wire [31:0] _06974_;
  wire [31:0] _06975_;
  /* cellift = 32'd1 */
  wire [31:0] _06976_;
  wire [31:0] _06977_;
  /* cellift = 32'd1 */
  wire [31:0] _06978_;
  wire [31:0] _06979_;
  /* cellift = 32'd1 */
  wire [31:0] _06980_;
  wire [31:0] _06981_;
  /* cellift = 32'd1 */
  wire [31:0] _06982_;
  wire [31:0] _06983_;
  /* cellift = 32'd1 */
  wire [31:0] _06984_;
  wire [31:0] _06985_;
  /* cellift = 32'd1 */
  wire [31:0] _06986_;
  wire [31:0] _06987_;
  /* cellift = 32'd1 */
  wire [31:0] _06988_;
  wire [31:0] _06989_;
  /* cellift = 32'd1 */
  wire [31:0] _06990_;
  wire [31:0] _06991_;
  /* cellift = 32'd1 */
  wire [31:0] _06992_;
  wire [31:0] _06993_;
  /* cellift = 32'd1 */
  wire [31:0] _06994_;
  wire [31:0] _06995_;
  /* cellift = 32'd1 */
  wire [31:0] _06996_;
  wire [31:0] _06997_;
  /* cellift = 32'd1 */
  wire [31:0] _06998_;
  wire [31:0] _06999_;
  /* cellift = 32'd1 */
  wire [31:0] _07000_;
  wire [31:0] _07001_;
  /* cellift = 32'd1 */
  wire [31:0] _07002_;
  wire [31:0] _07003_;
  /* cellift = 32'd1 */
  wire [31:0] _07004_;
  wire [31:0] _07005_;
  /* cellift = 32'd1 */
  wire [31:0] _07006_;
  wire [31:0] _07007_;
  /* cellift = 32'd1 */
  wire [31:0] _07008_;
  wire [31:0] _07009_;
  /* cellift = 32'd1 */
  wire [31:0] _07010_;
  wire [31:0] _07011_;
  /* cellift = 32'd1 */
  wire [31:0] _07012_;
  wire [31:0] _07013_;
  /* cellift = 32'd1 */
  wire [31:0] _07014_;
  wire [31:0] _07015_;
  /* cellift = 32'd1 */
  wire [31:0] _07016_;
  wire [31:0] _07017_;
  /* cellift = 32'd1 */
  wire [31:0] _07018_;
  wire [31:0] _07019_;
  /* cellift = 32'd1 */
  wire [31:0] _07020_;
  wire _07021_;
  /* cellift = 32'd1 */
  wire _07022_;
  wire _07023_;
  /* cellift = 32'd1 */
  wire _07024_;
  wire _07025_;
  /* cellift = 32'd1 */
  wire _07026_;
  wire _07027_;
  /* cellift = 32'd1 */
  wire _07028_;
  wire _07029_;
  /* cellift = 32'd1 */
  wire _07030_;
  wire _07031_;
  /* cellift = 32'd1 */
  wire _07032_;
  wire _07033_;
  /* cellift = 32'd1 */
  wire _07034_;
  wire _07035_;
  /* cellift = 32'd1 */
  wire _07036_;
  wire _07037_;
  /* cellift = 32'd1 */
  wire _07038_;
  wire _07039_;
  /* cellift = 32'd1 */
  wire _07040_;
  wire _07041_;
  /* cellift = 32'd1 */
  wire _07042_;
  wire _07043_;
  /* cellift = 32'd1 */
  wire _07044_;
  wire _07045_;
  /* cellift = 32'd1 */
  wire _07046_;
  wire _07047_;
  /* cellift = 32'd1 */
  wire _07048_;
  wire _07049_;
  /* cellift = 32'd1 */
  wire _07050_;
  wire _07051_;
  /* cellift = 32'd1 */
  wire _07052_;
  wire _07053_;
  /* cellift = 32'd1 */
  wire _07054_;
  wire _07055_;
  /* cellift = 32'd1 */
  wire _07056_;
  wire _07057_;
  /* cellift = 32'd1 */
  wire _07058_;
  wire _07059_;
  /* cellift = 32'd1 */
  wire _07060_;
  wire _07061_;
  /* cellift = 32'd1 */
  wire _07062_;
  wire _07063_;
  /* cellift = 32'd1 */
  wire _07064_;
  wire _07065_;
  /* cellift = 32'd1 */
  wire _07066_;
  wire _07067_;
  /* cellift = 32'd1 */
  wire _07068_;
  wire _07069_;
  /* cellift = 32'd1 */
  wire _07070_;
  wire _07071_;
  /* cellift = 32'd1 */
  wire _07072_;
  wire _07073_;
  /* cellift = 32'd1 */
  wire _07074_;
  wire _07075_;
  /* cellift = 32'd1 */
  wire _07076_;
  wire _07077_;
  /* cellift = 32'd1 */
  wire _07078_;
  wire _07079_;
  /* cellift = 32'd1 */
  wire _07080_;
  wire _07081_;
  /* cellift = 32'd1 */
  wire _07082_;
  wire _07083_;
  /* cellift = 32'd1 */
  wire _07084_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1186.33-1186.40" */
  wire [31:0] _07085_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1187.33-1187.40" */
  wire [31:0] _07086_;
  /* src = "generated/out/vanilla.sv:1669.32-1669.49" */
  wire _07087_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1669.32-1669.49" */
  wire _07088_;
  /* src = "generated/out/vanilla.sv:427.45-427.72" */
  wire _07089_;
  /* src = "generated/out/vanilla.sv:431.46-431.74" */
  wire _07090_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:431.46-431.74" */
  wire _07091_;
  /* src = "generated/out/vanilla.sv:984.104-984.129" */
  wire _07092_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:984.104-984.129" */
  wire _07093_;
  /* src = "generated/out/vanilla.sv:1136.37-1136.54" */
  wire [31:0] _07094_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1136.37-1136.54" */
  wire [31:0] _07095_;
  wire _07096_;
  wire _07097_;
  wire [31:0] _07098_;
  /* cellift = 32'd1 */
  wire [31:0] _07099_;
  wire [31:0] _07100_;
  /* cellift = 32'd1 */
  wire [31:0] _07101_;
  wire [3:0] _07102_;
  /* cellift = 32'd1 */
  wire [3:0] _07103_;
  wire [3:0] _07104_;
  /* cellift = 32'd1 */
  wire [3:0] _07105_;
  wire [31:0] _07106_;
  /* cellift = 32'd1 */
  wire [31:0] _07107_;
  wire [31:0] _07108_;
  wire [31:0] _07109_;
  /* cellift = 32'd1 */
  wire [31:0] _07110_;
  wire _07111_;
  wire [4:0] _07112_;
  wire [4:0] _07113_;
  /* cellift = 32'd1 */
  wire [4:0] _07114_;
  wire [31:0] _07115_;
  /* cellift = 32'd1 */
  wire [31:0] _07116_;
  wire [31:0] _07117_;
  /* cellift = 32'd1 */
  wire [31:0] _07118_;
  wire _07119_;
  wire _07120_;
  /* cellift = 32'd1 */
  wire _07121_;
  wire _07122_;
  /* cellift = 32'd1 */
  wire _07123_;
  wire _07124_;
  /* cellift = 32'd1 */
  wire _07125_;
  wire _07126_;
  /* cellift = 32'd1 */
  wire _07127_;
  wire [31:0] _07128_;
  /* cellift = 32'd1 */
  wire [31:0] _07129_;
  wire [31:0] _07130_;
  /* cellift = 32'd1 */
  wire [31:0] _07131_;
  wire [31:0] _07132_;
  /* cellift = 32'd1 */
  wire [31:0] _07133_;
  wire [31:0] _07134_;
  /* cellift = 32'd1 */
  wire [31:0] _07135_;
  wire [31:0] _07136_;
  /* cellift = 32'd1 */
  wire [31:0] _07137_;
  wire [4:0] _07138_;
  /* cellift = 32'd1 */
  wire [4:0] _07139_;
  wire [4:0] _07140_;
  /* cellift = 32'd1 */
  wire [4:0] _07141_;
  wire _07142_;
  wire _07143_;
  wire [4:0] _07144_;
  wire _07145_;
  /* cellift = 32'd1 */
  wire _07146_;
  /* cellift = 32'd1 */
  wire _07147_;
  wire _07148_;
  /* cellift = 32'd1 */
  wire _07149_;
  /* cellift = 32'd1 */
  wire _07150_;
  wire _07151_;
  /* cellift = 32'd1 */
  wire _07152_;
  wire _07153_;
  /* cellift = 32'd1 */
  wire _07154_;
  wire _07155_;
  /* cellift = 32'd1 */
  wire _07156_;
  wire _07157_;
  /* cellift = 32'd1 */
  wire _07158_;
  wire _07159_;
  /* cellift = 32'd1 */
  wire _07160_;
  wire [7:0] _07161_;
  /* cellift = 32'd1 */
  wire [7:0] _07162_;
  wire [7:0] _07163_;
  /* cellift = 32'd1 */
  wire [7:0] _07164_;
  wire [7:0] _07165_;
  /* cellift = 32'd1 */
  wire [7:0] _07166_;
  wire [7:0] _07167_;
  /* cellift = 32'd1 */
  wire [7:0] _07168_;
  wire [7:0] _07169_;
  /* cellift = 32'd1 */
  wire [7:0] _07170_;
  wire [7:0] _07171_;
  /* cellift = 32'd1 */
  wire [7:0] _07172_;
  wire [7:0] _07173_;
  /* cellift = 32'd1 */
  wire [7:0] _07174_;
  wire [7:0] _07175_;
  /* cellift = 32'd1 */
  wire [7:0] _07176_;
  wire [7:0] _07177_;
  /* cellift = 32'd1 */
  wire [7:0] _07178_;
  wire [7:0] _07179_;
  /* cellift = 32'd1 */
  wire [7:0] _07180_;
  wire [7:0] _07181_;
  /* cellift = 32'd1 */
  wire [7:0] _07182_;
  wire [7:0] _07183_;
  /* cellift = 32'd1 */
  wire [7:0] _07184_;
  wire [7:0] _07185_;
  /* cellift = 32'd1 */
  wire [7:0] _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire [31:0] _07192_;
  /* cellift = 32'd1 */
  wire [31:0] _07193_;
  wire [31:0] _07194_;
  /* cellift = 32'd1 */
  wire [31:0] _07195_;
  wire [31:0] _07196_;
  /* cellift = 32'd1 */
  wire [31:0] _07197_;
  wire [31:0] _07198_;
  /* cellift = 32'd1 */
  wire [31:0] _07199_;
  wire [31:0] _07200_;
  /* cellift = 32'd1 */
  wire [31:0] _07201_;
  wire _07202_;
  /* cellift = 32'd1 */
  wire _07203_;
  wire _07204_;
  /* cellift = 32'd1 */
  wire _07205_;
  wire _07206_;
  /* cellift = 32'd1 */
  wire _07207_;
  /* cellift = 32'd1 */
  wire _07208_;
  wire _07209_;
  /* cellift = 32'd1 */
  wire _07210_;
  wire [1:0] _07211_;
  /* cellift = 32'd1 */
  wire [1:0] _07212_;
  wire [1:0] _07213_;
  /* cellift = 32'd1 */
  wire [1:0] _07214_;
  wire [1:0] _07215_;
  /* cellift = 32'd1 */
  wire [1:0] _07216_;
  /* cellift = 32'd1 */
  wire [1:0] _07217_;
  wire [31:0] _07218_;
  /* cellift = 32'd1 */
  wire [31:0] _07219_;
  wire [31:0] _07220_;
  /* cellift = 32'd1 */
  wire [31:0] _07221_;
  wire [31:0] _07222_;
  /* cellift = 32'd1 */
  wire [31:0] _07223_;
  wire [31:0] _07224_;
  /* cellift = 32'd1 */
  wire [31:0] _07225_;
  wire [31:0] _07226_;
  /* cellift = 32'd1 */
  wire [31:0] _07227_;
  wire [31:0] _07228_;
  /* cellift = 32'd1 */
  wire [31:0] _07229_;
  wire [31:0] _07230_;
  /* cellift = 32'd1 */
  wire [31:0] _07231_;
  wire [31:0] _07232_;
  /* cellift = 32'd1 */
  wire [31:0] _07233_;
  wire _07234_;
  /* cellift = 32'd1 */
  wire _07235_;
  wire _07236_;
  /* cellift = 32'd1 */
  wire _07237_;
  wire _07238_;
  /* cellift = 32'd1 */
  wire _07239_;
  /* cellift = 32'd1 */
  wire _07240_;
  wire _07241_;
  /* cellift = 32'd1 */
  wire _07242_;
  wire _07243_;
  /* cellift = 32'd1 */
  wire _07244_;
  wire _07245_;
  /* cellift = 32'd1 */
  wire _07246_;
  wire _07247_;
  /* cellift = 32'd1 */
  wire _07248_;
  /* cellift = 32'd1 */
  wire _07249_;
  wire _07250_;
  wire _07251_;
  /* cellift = 32'd1 */
  wire _07252_;
  wire _07253_;
  wire _07254_;
  /* cellift = 32'd1 */
  wire _07255_;
  wire _07256_;
  /* cellift = 32'd1 */
  wire _07257_;
  wire _07258_;
  /* cellift = 32'd1 */
  wire _07259_;
  wire _07260_;
  /* cellift = 32'd1 */
  wire _07261_;
  /* cellift = 32'd1 */
  wire _07262_;
  wire _07263_;
  /* cellift = 32'd1 */
  wire _07264_;
  wire _07265_;
  /* cellift = 32'd1 */
  wire _07266_;
  wire _07267_;
  /* cellift = 32'd1 */
  wire _07268_;
  /* cellift = 32'd1 */
  wire _07269_;
  wire _07270_;
  /* cellift = 32'd1 */
  wire _07271_;
  wire _07272_;
  /* cellift = 32'd1 */
  wire _07273_;
  wire _07274_;
  /* cellift = 32'd1 */
  wire _07275_;
  wire _07276_;
  /* cellift = 32'd1 */
  wire _07277_;
  wire _07278_;
  /* cellift = 32'd1 */
  wire _07279_;
  wire _07280_;
  /* cellift = 32'd1 */
  wire _07281_;
  wire [2:0] _07282_;
  /* cellift = 32'd1 */
  wire [2:0] _07283_;
  wire _07284_;
  /* cellift = 32'd1 */
  wire _07285_;
  wire [1:0] _07286_;
  /* cellift = 32'd1 */
  wire [1:0] _07287_;
  wire [11:0] _07288_;
  /* cellift = 32'd1 */
  wire [11:0] _07289_;
  wire _07290_;
  /* cellift = 32'd1 */
  wire _07291_;
  wire _07292_;
  /* cellift = 32'd1 */
  wire _07293_;
  /* cellift = 32'd1 */
  wire [3:0] _07294_;
  wire [3:0] _07295_;
  /* cellift = 32'd1 */
  wire [3:0] _07296_;
  wire [3:0] _07297_;
  /* cellift = 32'd1 */
  wire [3:0] _07298_;
  wire [3:0] _07299_;
  /* cellift = 32'd1 */
  wire [3:0] _07300_;
  wire [3:0] _07301_;
  /* cellift = 32'd1 */
  wire [3:0] _07302_;
  wire [3:0] _07303_;
  /* cellift = 32'd1 */
  wire [3:0] _07304_;
  wire [3:0] _07305_;
  /* cellift = 32'd1 */
  wire [3:0] _07306_;
  wire [3:0] _07307_;
  /* cellift = 32'd1 */
  wire [3:0] _07308_;
  /* cellift = 32'd1 */
  wire [3:0] _07309_;
  wire [3:0] _07310_;
  /* cellift = 32'd1 */
  wire [3:0] _07311_;
  wire [3:0] _07312_;
  /* cellift = 32'd1 */
  wire [3:0] _07313_;
  wire _07314_;
  /* cellift = 32'd1 */
  wire _07315_;
  wire _07316_;
  /* cellift = 32'd1 */
  wire _07317_;
  wire _07318_;
  /* cellift = 32'd1 */
  wire _07319_;
  wire _07320_;
  /* cellift = 32'd1 */
  wire _07321_;
  wire _07322_;
  /* cellift = 32'd1 */
  wire _07323_;
  wire _07324_;
  /* cellift = 32'd1 */
  wire _07325_;
  wire _07326_;
  /* cellift = 32'd1 */
  wire _07327_;
  wire _07328_;
  /* cellift = 32'd1 */
  wire _07329_;
  wire _07330_;
  /* cellift = 32'd1 */
  wire _07331_;
  wire _07332_;
  /* cellift = 32'd1 */
  wire _07333_;
  wire _07334_;
  /* cellift = 32'd1 */
  wire _07335_;
  wire _07336_;
  /* cellift = 32'd1 */
  wire _07337_;
  wire _07338_;
  /* cellift = 32'd1 */
  wire _07339_;
  wire _07340_;
  /* cellift = 32'd1 */
  wire _07341_;
  wire _07342_;
  /* cellift = 32'd1 */
  wire _07343_;
  wire _07344_;
  /* cellift = 32'd1 */
  wire _07345_;
  wire _07346_;
  /* cellift = 32'd1 */
  wire _07347_;
  wire _07348_;
  /* cellift = 32'd1 */
  wire _07349_;
  wire _07350_;
  /* cellift = 32'd1 */
  wire _07351_;
  wire _07352_;
  /* cellift = 32'd1 */
  wire _07353_;
  wire _07354_;
  /* cellift = 32'd1 */
  wire _07355_;
  wire _07356_;
  /* cellift = 32'd1 */
  wire _07357_;
  wire _07358_;
  /* cellift = 32'd1 */
  wire _07359_;
  wire _07360_;
  /* cellift = 32'd1 */
  wire _07361_;
  wire _07362_;
  wire _07363_;
  /* cellift = 32'd1 */
  wire _07364_;
  wire [4:0] _07365_;
  /* cellift = 32'd1 */
  wire [4:0] _07366_;
  wire [4:0] _07367_;
  /* cellift = 32'd1 */
  wire [4:0] _07368_;
  /* cellift = 32'd1 */
  wire [4:0] _07369_;
  wire [4:0] _07370_;
  /* cellift = 32'd1 */
  wire [4:0] _07371_;
  /* cellift = 32'd1 */
  wire [4:0] _07372_;
  wire [4:0] _07373_;
  /* cellift = 32'd1 */
  wire [4:0] _07374_;
  /* cellift = 32'd1 */
  wire [4:0] _07375_;
  wire [4:0] _07376_;
  /* cellift = 32'd1 */
  wire [4:0] _07377_;
  wire [7:0] _07378_;
  /* cellift = 32'd1 */
  wire [7:0] _07379_;
  wire [4:0] _07380_;
  /* cellift = 32'd1 */
  wire [4:0] _07381_;
  wire [4:0] _07382_;
  /* cellift = 32'd1 */
  wire [4:0] _07383_;
  wire [4:0] _07384_;
  /* cellift = 32'd1 */
  wire [4:0] _07385_;
  wire [4:0] _07386_;
  /* cellift = 32'd1 */
  wire [4:0] _07387_;
  /* cellift = 32'd1 */
  wire [4:0] _07388_;
  wire [4:0] _07389_;
  /* cellift = 32'd1 */
  wire [4:0] _07390_;
  wire [4:0] _07391_;
  /* cellift = 32'd1 */
  wire [4:0] _07392_;
  wire [4:0] _07393_;
  /* cellift = 32'd1 */
  wire [4:0] _07394_;
  wire [4:0] _07395_;
  /* cellift = 32'd1 */
  wire [4:0] _07396_;
  wire _07397_;
  /* cellift = 32'd1 */
  wire [4:0] _07398_;
  wire [4:0] _07399_;
  /* cellift = 32'd1 */
  wire [4:0] _07400_;
  wire _07401_;
  /* cellift = 32'd1 */
  wire _07402_;
  wire _07403_;
  /* cellift = 32'd1 */
  wire _07404_;
  wire _07405_;
  /* cellift = 32'd1 */
  wire _07406_;
  wire _07407_;
  /* cellift = 32'd1 */
  wire _07408_;
  wire _07409_;
  /* cellift = 32'd1 */
  wire _07410_;
  wire _07411_;
  /* cellift = 32'd1 */
  wire _07412_;
  wire _07413_;
  /* cellift = 32'd1 */
  wire _07414_;
  wire _07415_;
  /* cellift = 32'd1 */
  wire _07416_;
  wire _07417_;
  /* cellift = 32'd1 */
  wire _07418_;
  wire _07419_;
  /* cellift = 32'd1 */
  wire _07420_;
  wire _07421_;
  /* cellift = 32'd1 */
  wire _07422_;
  wire _07423_;
  /* cellift = 32'd1 */
  wire _07424_;
  wire _07425_;
  /* cellift = 32'd1 */
  wire _07426_;
  wire _07427_;
  /* cellift = 32'd1 */
  wire _07428_;
  wire _07429_;
  /* cellift = 32'd1 */
  wire _07430_;
  wire [15:0] _07431_;
  /* cellift = 32'd1 */
  wire [15:0] _07432_;
  wire [15:0] _07433_;
  /* cellift = 32'd1 */
  wire [15:0] _07434_;
  wire [15:0] _07435_;
  /* cellift = 32'd1 */
  wire [15:0] _07436_;
  wire [15:0] _07437_;
  /* cellift = 32'd1 */
  wire [15:0] _07438_;
  wire _07439_;
  /* cellift = 32'd1 */
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire [1:0] _07443_;
  wire [1:0] _07444_;
  wire [1:0] _07445_;
  /* cellift = 32'd1 */
  wire [1:0] _07446_;
  wire [1:0] _07447_;
  /* cellift = 32'd1 */
  wire [1:0] _07448_;
  wire [1:0] _07449_;
  wire [1:0] _07450_;
  /* cellift = 32'd1 */
  wire [1:0] _07451_;
  wire [1:0] _07452_;
  /* cellift = 32'd1 */
  wire [3:0] _07453_;
  wire [3:0] _07454_;
  /* cellift = 32'd1 */
  wire [3:0] _07455_;
  wire [3:0] _07456_;
  /* cellift = 32'd1 */
  wire [3:0] _07457_;
  wire _07458_;
  /* cellift = 32'd1 */
  wire _07459_;
  wire _07460_;
  wire _07461_;
  /* cellift = 32'd1 */
  wire _07462_;
  wire _07463_;
  /* cellift = 32'd1 */
  wire _07464_;
  wire _07465_;
  /* cellift = 32'd1 */
  wire _07466_;
  wire _07467_;
  /* cellift = 32'd1 */
  wire _07468_;
  /* cellift = 32'd1 */
  wire _07469_;
  /* cellift = 32'd1 */
  wire _07470_;
  /* cellift = 32'd1 */
  wire _07471_;
  wire _07472_;
  /* cellift = 32'd1 */
  wire _07473_;
  /* cellift = 32'd1 */
  wire _07474_;
  wire _07475_;
  /* cellift = 32'd1 */
  wire _07476_;
  wire _07477_;
  /* cellift = 32'd1 */
  wire _07478_;
  wire _07479_;
  /* cellift = 32'd1 */
  wire _07480_;
  wire _07481_;
  /* cellift = 32'd1 */
  wire _07482_;
  /* cellift = 32'd1 */
  wire _07483_;
  wire _07484_;
  /* cellift = 32'd1 */
  wire _07485_;
  wire _07486_;
  /* cellift = 32'd1 */
  wire _07487_;
  /* cellift = 32'd1 */
  wire [4:0] _07488_;
  /* cellift = 32'd1 */
  wire [4:0] _07489_;
  wire [4:0] _07490_;
  /* cellift = 32'd1 */
  wire [4:0] _07491_;
  wire [4:0] _07492_;
  /* cellift = 32'd1 */
  wire [4:0] _07493_;
  wire [4:0] _07494_;
  /* cellift = 32'd1 */
  wire [4:0] _07495_;
  wire [4:0] _07496_;
  /* cellift = 32'd1 */
  wire [4:0] _07497_;
  wire [4:0] _07498_;
  /* cellift = 32'd1 */
  wire [4:0] _07499_;
  wire [4:0] _07500_;
  /* cellift = 32'd1 */
  wire [4:0] _07501_;
  wire [4:0] _07502_;
  /* cellift = 32'd1 */
  wire [4:0] _07503_;
  /* cellift = 32'd1 */
  wire [2:0] _07504_;
  /* cellift = 32'd1 */
  wire [2:0] _07505_;
  /* cellift = 32'd1 */
  wire [2:0] _07506_;
  /* cellift = 32'd1 */
  wire [2:0] _07507_;
  wire [2:0] _07508_;
  /* cellift = 32'd1 */
  wire [2:0] _07509_;
  wire [2:0] _07510_;
  /* cellift = 32'd1 */
  wire [2:0] _07511_;
  wire [2:0] _07512_;
  /* cellift = 32'd1 */
  wire [2:0] _07513_;
  /* cellift = 32'd1 */
  wire [2:0] _07514_;
  wire [2:0] _07515_;
  /* cellift = 32'd1 */
  wire [2:0] _07516_;
  wire [2:0] _07517_;
  /* cellift = 32'd1 */
  wire [2:0] _07518_;
  wire [2:0] _07519_;
  /* cellift = 32'd1 */
  wire [2:0] _07520_;
  wire [2:0] _07521_;
  /* cellift = 32'd1 */
  wire [2:0] _07522_;
  wire [2:0] _07523_;
  /* cellift = 32'd1 */
  wire [2:0] _07524_;
  wire [2:0] _07525_;
  /* cellift = 32'd1 */
  wire [2:0] _07526_;
  wire [3:0] _07527_;
  /* cellift = 32'd1 */
  wire [3:0] _07528_;
  wire [3:0] _07529_;
  /* cellift = 32'd1 */
  wire [3:0] _07530_;
  wire [3:0] _07531_;
  /* cellift = 32'd1 */
  wire [3:0] _07532_;
  wire [3:0] _07533_;
  /* cellift = 32'd1 */
  wire [3:0] _07534_;
  /* cellift = 32'd1 */
  wire [5:0] _07535_;
  /* cellift = 32'd1 */
  wire [5:0] _07536_;
  /* cellift = 32'd1 */
  wire [5:0] _07537_;
  /* cellift = 32'd1 */
  wire [5:0] _07538_;
  wire [5:0] _07539_;
  /* cellift = 32'd1 */
  wire [5:0] _07540_;
  wire [5:0] _07541_;
  /* cellift = 32'd1 */
  wire [5:0] _07542_;
  wire [5:0] _07543_;
  /* cellift = 32'd1 */
  wire [5:0] _07544_;
  wire [5:0] _07545_;
  /* cellift = 32'd1 */
  wire [5:0] _07546_;
  wire [5:0] _07547_;
  /* cellift = 32'd1 */
  wire [5:0] _07548_;
  wire [5:0] _07549_;
  /* cellift = 32'd1 */
  wire [5:0] _07550_;
  wire _07551_;
  /* cellift = 32'd1 */
  wire _07552_;
  wire _07553_;
  /* cellift = 32'd1 */
  wire _07554_;
  wire _07555_;
  /* cellift = 32'd1 */
  wire _07556_;
  wire _07557_;
  /* cellift = 32'd1 */
  wire _07558_;
  wire _07559_;
  /* cellift = 32'd1 */
  wire _07560_;
  /* src = "generated/out/vanilla.sv:296.113-296.123" */
  wire _07561_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:296.113-296.123" */
  wire _07562_;
  /* src = "generated/out/vanilla.sv:296.169-296.193" */
  wire _07563_;
  /* src = "generated/out/vanilla.sv:1186.19-1186.57" */
  wire _07564_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1186.19-1186.57" */
  wire _07565_;
  /* src = "generated/out/vanilla.sv:1187.19-1187.57" */
  wire _07566_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1187.19-1187.57" */
  wire _07567_;
  /* src = "generated/out/vanilla.sv:1746.22-1746.53" */
  wire _07568_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1746.22-1746.53" */
  wire _07569_;
  /* src = "generated/out/vanilla.sv:1776.24-1776.46" */
  wire _07570_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1776.24-1776.46" */
  wire _07571_;
  /* src = "generated/out/vanilla.sv:296.44-296.54" */
  wire _07572_;
  /* src = "generated/out/vanilla.sv:795.17-795.96" */
  wire _07573_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:795.17-795.96" */
  wire _07574_;
  /* src = "generated/out/vanilla.sv:827.27-827.51" */
  wire _07575_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:827.27-827.51" */
  wire _07576_;
  /* src = "generated/out/vanilla.sv:994.43-994.254" */
  wire _07577_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:994.43-994.254" */
  wire _07578_;
  /* src = "generated/out/vanilla.sv:995.78-995.259" */
  wire _07579_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:995.78-995.259" */
  wire _07580_;
  /* src = "generated/out/vanilla.sv:330.20-330.43" */
  wire [3:0] _07581_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:330.20-330.43" */
  wire [3:0] _07582_;
  /* src = "generated/out/vanilla.sv:1110.32-1110.49" */
  wire [31:0] _07583_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1110.32-1110.49" */
  wire [31:0] _07584_;
  /* src = "generated/out/vanilla.sv:1216.30-1216.54" */
  /* unused_bits = "4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _07585_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1216.30-1216.54" */
  /* unused_bits = "4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _07586_;
  /* src = "generated/out/vanilla.sv:1591.17-1591.27" */
  /* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _07587_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1591.17-1591.27" */
  /* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _07588_;
  /* src = "generated/out/vanilla.sv:1600.17-1600.27" */
  /* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _07589_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1600.17-1600.27" */
  /* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _07590_;
  /* src = "generated/out/vanilla.sv:1163.33-1163.54" */
  wire [31:0] _07591_;
  /* src = "generated/out/vanilla.sv:1167.24-1167.59" */
  wire [31:0] _07592_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1167.24-1167.59" */
  wire [31:0] _07593_;
  /* src = "generated/out/vanilla.sv:1280.37-1280.109" */
  wire [31:0] _07594_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1280.37-1280.109" */
  wire [31:0] _07595_;
  /* src = "generated/out/vanilla.sv:1323.37-1323.61" */
  wire [31:0] _07596_;
  /* src = "generated/out/vanilla.sv:1405.20-1405.42" */
  wire [31:0] _07597_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1405.20-1405.42" */
  wire [31:0] _07598_;
  /* src = "generated/out/vanilla.sv:1746.22-1746.53" */
  wire [31:0] _07599_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1746.22-1746.53" */
  wire [31:0] _07600_;
  /* src = "generated/out/vanilla.sv:1776.24-1776.46" */
  /* unused_bits = "4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _07601_;
  /* src = "generated/out/vanilla.sv:301.221-301.346" */
  wire [31:0] _07602_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:301.221-301.346" */
  wire [31:0] _07603_;
  /* src = "generated/out/vanilla.sv:301.126-301.347" */
  wire [31:0] _07604_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:301.126-301.347" */
  wire [31:0] _07605_;
  /* src = "generated/out/vanilla.sv:322.21-322.51" */
  wire [3:0] _07606_;
  /* src = "generated/out/vanilla.sv:400.32-400.89" */
  wire [6:0] _07607_;
  /* src = "generated/out/vanilla.sv:512.22-512.58" */
  /* unused_bits = "2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _07608_;
  /* src = "generated/out/vanilla.sv:1135.39-1135.56" */
  wire [31:0] _07609_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1135.39-1135.56" */
  wire [31:0] _07610_;
  /* src = "generated/out/vanilla.sv:1091.13-1091.24" */
  wire [31:0] alu_add_sub;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1091.13-1091.24" */
  wire [31:0] alu_add_sub_t0;
  /* src = "generated/out/vanilla.sv:1094.6-1094.12" */
  wire alu_eq;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1094.6-1094.12" */
  wire alu_eq_t0;
  /* src = "generated/out/vanilla.sv:1096.6-1096.13" */
  wire alu_lts;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1096.6-1096.13" */
  wire alu_lts_t0;
  /* src = "generated/out/vanilla.sv:1095.6-1095.13" */
  wire alu_ltu;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1095.6-1095.13" */
  wire alu_ltu_t0;
  /* src = "generated/out/vanilla.sv:1085.13-1085.20" */
  wire [31:0] alu_out;
  /* src = "generated/out/vanilla.sv:1087.6-1087.15" */
  wire alu_out_0;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1087.6-1087.15" */
  wire alu_out_0_t0;
  /* src = "generated/out/vanilla.sv:1086.13-1086.22" */
  reg [31:0] alu_out_q;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1086.13-1086.22" */
  reg [31:0] alu_out_q_t0;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1085.13-1085.20" */
  wire [31:0] alu_out_t0;
  /* src = "generated/out/vanilla.sv:731.13-731.31" */
  reg [31:0] cached_insn_opcode;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:731.13-731.31" */
  reg [31:0] cached_insn_opcode_t0;
  /* src = "generated/out/vanilla.sv:732.12-732.27" */
  reg [4:0] cached_insn_rs1;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:732.12-732.27" */
  reg [4:0] cached_insn_rs1_t0;
  /* src = "generated/out/vanilla.sv:733.12-733.27" */
  reg [4:0] cached_insn_rs2;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:733.12-733.27" */
  reg [4:0] cached_insn_rs2_t0;
  /* src = "generated/out/vanilla.sv:289.6-289.32" */
  wire clear_prefetched_high_word;
  /* src = "generated/out/vanilla.sv:1142.6-1142.34" */
  reg clear_prefetched_high_word_q;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1142.6-1142.34" */
  reg clear_prefetched_high_word_q_t0;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:289.6-289.32" */
  wire clear_prefetched_high_word_t0;
  /* src = "generated/out/vanilla.sv:85.8-85.11" */
  input clk;
  wire clk;
  /* src = "generated/out/vanilla.sv:593.6-593.22" */
  reg compressed_instr;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:593.6-593.22" */
  reg compressed_instr_t0;
  /* src = "generated/out/vanilla.sv:151.13-151.24" */
  reg [63:0] count_cycle;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:151.13-151.24" */
  reg [63:0] count_cycle_t0;
  /* src = "generated/out/vanilla.sv:152.13-152.24" */
  reg [63:0] count_instr;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:152.13-152.24" */
  reg [63:0] count_instr_t0;
  /* src = "generated/out/vanilla.sv:1045.12-1045.21" */
  reg [7:0] cpu_state;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1045.12-1045.21" */
  reg [7:0] cpu_state_t0;
  reg [31:0] \cpuregs[0] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[0]_t0 ;
  reg [31:0] \cpuregs[10] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[10]_t0 ;
  reg [31:0] \cpuregs[11] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[11]_t0 ;
  reg [31:0] \cpuregs[12] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[12]_t0 ;
  reg [31:0] \cpuregs[13] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[13]_t0 ;
  reg [31:0] \cpuregs[14] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[14]_t0 ;
  reg [31:0] \cpuregs[15] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[15]_t0 ;
  reg [31:0] \cpuregs[16] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[16]_t0 ;
  reg [31:0] \cpuregs[17] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[17]_t0 ;
  reg [31:0] \cpuregs[18] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[18]_t0 ;
  reg [31:0] \cpuregs[19] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[19]_t0 ;
  reg [31:0] \cpuregs[1] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[1]_t0 ;
  reg [31:0] \cpuregs[20] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[20]_t0 ;
  reg [31:0] \cpuregs[21] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[21]_t0 ;
  reg [31:0] \cpuregs[22] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[22]_t0 ;
  reg [31:0] \cpuregs[23] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[23]_t0 ;
  reg [31:0] \cpuregs[24] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[24]_t0 ;
  reg [31:0] \cpuregs[25] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[25]_t0 ;
  reg [31:0] \cpuregs[26] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[26]_t0 ;
  reg [31:0] \cpuregs[27] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[27]_t0 ;
  reg [31:0] \cpuregs[28] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[28]_t0 ;
  reg [31:0] \cpuregs[29] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[29]_t0 ;
  reg [31:0] \cpuregs[2] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[2]_t0 ;
  reg [31:0] \cpuregs[30] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[30]_t0 ;
  reg [31:0] \cpuregs[31] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[31]_t0 ;
  reg [31:0] \cpuregs[3] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[3]_t0 ;
  reg [31:0] \cpuregs[4] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[4]_t0 ;
  reg [31:0] \cpuregs[5] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[5]_t0 ;
  reg [31:0] \cpuregs[6] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[6]_t0 ;
  reg [31:0] \cpuregs[7] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[7]_t0 ;
  reg [31:0] \cpuregs[8] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[8]_t0 ;
  reg [31:0] \cpuregs[9] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[9]_t0 ;
  /* src = "generated/out/vanilla.sv:1153.13-1153.24" */
  wire [31:0] cpuregs_rs1;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1153.13-1153.24" */
  wire [31:0] cpuregs_rs1_t0;
  /* src = "generated/out/vanilla.sv:1154.13-1154.24" */
  wire [31:0] cpuregs_rs2;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1154.13-1154.24" */
  wire [31:0] cpuregs_rs2_t0;
  /* src = "generated/out/vanilla.sv:1152.13-1152.27" */
  wire [31:0] cpuregs_wrdata;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1152.13-1152.27" */
  wire [31:0] cpuregs_wrdata_t0;
  /* src = "generated/out/vanilla.sv:1151.6-1151.19" */
  wire cpuregs_write;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1151.6-1151.19" */
  wire cpuregs_write_t0;
  /* src = "generated/out/vanilla.sv:160.13-160.28" */
  wire [31:0] dbg_insn_opcode;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:160.13-160.28" */
  wire [31:0] dbg_insn_opcode_t0;
  /* src = "generated/out/vanilla.sv:614.12-614.24" */
  wire [4:0] dbg_insn_rs1;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:614.12-614.24" */
  wire [4:0] dbg_insn_rs1_t0;
  /* src = "generated/out/vanilla.sv:615.12-615.24" */
  wire [4:0] dbg_insn_rs2;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:615.12-615.24" */
  wire [4:0] dbg_insn_rs2_t0;
  /* src = "generated/out/vanilla.sv:726.6-726.14" */
  reg dbg_next;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:726.6-726.14" */
  reg dbg_next_t0;
  /* src = "generated/out/vanilla.sv:617.13-617.23" */
  reg [31:0] dbg_rs1val;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:617.13-617.23" */
  reg [31:0] dbg_rs1val_t0;
  /* src = "generated/out/vanilla.sv:619.6-619.22" */
  reg dbg_rs1val_valid;
  /* src = "generated/out/vanilla.sv:618.13-618.23" */
  reg [31:0] dbg_rs2val;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:618.13-618.23" */
  reg [31:0] dbg_rs2val_t0;
  /* src = "generated/out/vanilla.sv:620.6-620.22" */
  reg dbg_rs2val_valid;
  /* src = "generated/out/vanilla.sv:728.6-728.20" */
  reg dbg_valid_insn;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:728.6-728.20" */
  reg dbg_valid_insn_t0;
  /* src = "generated/out/vanilla.sv:587.13-587.24" */
  reg [31:0] decoded_imm;
  /* src = "generated/out/vanilla.sv:588.13-588.26" */
  wire [31:0] decoded_imm_j;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:588.13-588.26" */
  wire [31:0] decoded_imm_j_t0;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:587.13-587.24" */
  reg [31:0] decoded_imm_t0;
  /* src = "generated/out/vanilla.sv:584.28-584.38" */
  reg [4:0] decoded_rd;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:584.28-584.38" */
  reg [4:0] decoded_rd_t0;
  /* src = "generated/out/vanilla.sv:585.28-585.39" */
  reg [4:0] decoded_rs1;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:585.28-585.39" */
  reg [4:0] decoded_rs1_t0;
  /* src = "generated/out/vanilla.sv:586.28-586.39" */
  reg [4:0] decoded_rs2;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:586.28-586.39" */
  reg [4:0] decoded_rs2_t0;
  /* src = "generated/out/vanilla.sv:591.6-591.28" */
  reg decoder_pseudo_trigger;
  /* src = "generated/out/vanilla.sv:592.6-592.30" */
  reg decoder_pseudo_trigger_q;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:592.6-592.30" */
  reg decoder_pseudo_trigger_q_t0;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:591.6-591.28" */
  reg decoder_pseudo_trigger_t0;
  /* src = "generated/out/vanilla.sv:589.6-589.21" */
  reg decoder_trigger;
  /* src = "generated/out/vanilla.sv:590.6-590.23" */
  reg decoder_trigger_q;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:590.6-590.23" */
  reg decoder_trigger_q_t0;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:589.6-589.21" */
  reg decoder_trigger_t0;
  /* src = "generated/out/vanilla.sv:109.20-109.23" */
  output [31:0] eoi;
  wire [31:0] eoi;
  /* cellift = 32'd1 */
  output [31:0] eoi_t0;
  wire [31:0] eoi_t0;
  /* src = "generated/out/vanilla.sv:561.6-561.15" */
  reg instr_add;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:561.6-561.15" */
  reg instr_add_t0;
  /* src = "generated/out/vanilla.sv:552.6-552.16" */
  reg instr_addi;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:552.6-552.16" */
  reg instr_addi_t0;
  /* src = "generated/out/vanilla.sv:570.6-570.15" */
  reg instr_and;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:570.6-570.15" */
  reg instr_and_t0;
  /* src = "generated/out/vanilla.sv:557.6-557.16" */
  reg instr_andi;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:557.6-557.16" */
  reg instr_andi_t0;
  /* src = "generated/out/vanilla.sv:535.6-535.17" */
  reg instr_auipc;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:535.6-535.17" */
  reg instr_auipc_t0;
  /* src = "generated/out/vanilla.sv:538.6-538.15" */
  reg instr_beq;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:538.6-538.15" */
  reg instr_beq_t0;
  /* src = "generated/out/vanilla.sv:541.6-541.15" */
  reg instr_bge;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:541.6-541.15" */
  reg instr_bge_t0;
  /* src = "generated/out/vanilla.sv:543.6-543.16" */
  reg instr_bgeu;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:543.6-543.16" */
  reg instr_bgeu_t0;
  /* src = "generated/out/vanilla.sv:540.6-540.15" */
  reg instr_blt;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:540.6-540.15" */
  reg instr_blt_t0;
  /* src = "generated/out/vanilla.sv:542.6-542.16" */
  reg instr_bltu;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:542.6-542.16" */
  reg instr_bltu_t0;
  /* src = "generated/out/vanilla.sv:539.6-539.15" */
  reg instr_bne;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:539.6-539.15" */
  reg instr_bne_t0;
  /* src = "generated/out/vanilla.sv:575.6-575.24" */
  reg instr_ecall_ebreak;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:575.6-575.24" */
  reg instr_ecall_ebreak_t0;
  /* src = "generated/out/vanilla.sv:576.6-576.17" */
  reg instr_fence;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:576.6-576.17" */
  reg instr_fence_t0;
  /* src = "generated/out/vanilla.sv:536.6-536.15" */
  reg instr_jal;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:536.6-536.15" */
  reg instr_jal_t0;
  /* src = "generated/out/vanilla.sv:537.6-537.16" */
  reg instr_jalr;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:537.6-537.16" */
  reg instr_jalr_t0;
  /* src = "generated/out/vanilla.sv:544.6-544.14" */
  reg instr_lb;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:544.6-544.14" */
  reg instr_lb_t0;
  /* src = "generated/out/vanilla.sv:547.6-547.15" */
  reg instr_lbu;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:547.6-547.15" */
  reg instr_lbu_t0;
  /* src = "generated/out/vanilla.sv:545.6-545.14" */
  reg instr_lh;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:545.6-545.14" */
  reg instr_lh_t0;
  /* src = "generated/out/vanilla.sv:548.6-548.15" */
  reg instr_lhu;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:548.6-548.15" */
  reg instr_lhu_t0;
  /* src = "generated/out/vanilla.sv:534.6-534.15" */
  reg instr_lui;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:534.6-534.15" */
  reg instr_lui_t0;
  /* src = "generated/out/vanilla.sv:546.6-546.14" */
  reg instr_lw;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:546.6-546.14" */
  reg instr_lw_t0;
  /* src = "generated/out/vanilla.sv:569.6-569.14" */
  reg instr_or;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:569.6-569.14" */
  reg instr_or_t0;
  /* src = "generated/out/vanilla.sv:556.6-556.15" */
  reg instr_ori;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:556.6-556.15" */
  reg instr_ori_t0;
  /* src = "generated/out/vanilla.sv:571.6-571.19" */
  reg instr_rdcycle;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:571.6-571.19" */
  reg instr_rdcycle_t0;
  /* src = "generated/out/vanilla.sv:572.6-572.20" */
  reg instr_rdcycleh;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:572.6-572.20" */
  reg instr_rdcycleh_t0;
  /* src = "generated/out/vanilla.sv:573.6-573.19" */
  reg instr_rdinstr;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:573.6-573.19" */
  reg instr_rdinstr_t0;
  /* src = "generated/out/vanilla.sv:574.6-574.20" */
  reg instr_rdinstrh;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:574.6-574.20" */
  reg instr_rdinstrh_t0;
  /* src = "generated/out/vanilla.sv:549.6-549.14" */
  reg instr_sb;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:549.6-549.14" */
  reg instr_sb_t0;
  /* src = "generated/out/vanilla.sv:550.6-550.14" */
  reg instr_sh;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:550.6-550.14" */
  reg instr_sh_t0;
  /* src = "generated/out/vanilla.sv:563.6-563.15" */
  reg instr_sll;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:563.6-563.15" */
  reg instr_sll_t0;
  /* src = "generated/out/vanilla.sv:558.6-558.16" */
  reg instr_slli;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:558.6-558.16" */
  reg instr_slli_t0;
  /* src = "generated/out/vanilla.sv:564.6-564.15" */
  reg instr_slt;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:564.6-564.15" */
  reg instr_slt_t0;
  /* src = "generated/out/vanilla.sv:553.6-553.16" */
  reg instr_slti;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:553.6-553.16" */
  reg instr_slti_t0;
  /* src = "generated/out/vanilla.sv:554.6-554.17" */
  reg instr_sltiu;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:554.6-554.17" */
  reg instr_sltiu_t0;
  /* src = "generated/out/vanilla.sv:565.6-565.16" */
  reg instr_sltu;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:565.6-565.16" */
  reg instr_sltu_t0;
  /* src = "generated/out/vanilla.sv:568.6-568.15" */
  reg instr_sra;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:568.6-568.15" */
  reg instr_sra_t0;
  /* src = "generated/out/vanilla.sv:560.6-560.16" */
  reg instr_srai;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:560.6-560.16" */
  reg instr_srai_t0;
  /* src = "generated/out/vanilla.sv:567.6-567.15" */
  reg instr_srl;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:567.6-567.15" */
  reg instr_srl_t0;
  /* src = "generated/out/vanilla.sv:559.6-559.16" */
  reg instr_srli;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:559.6-559.16" */
  reg instr_srli_t0;
  /* src = "generated/out/vanilla.sv:562.6-562.15" */
  reg instr_sub;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:562.6-562.15" */
  reg instr_sub_t0;
  /* src = "generated/out/vanilla.sv:551.6-551.14" */
  reg instr_sw;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:551.6-551.14" */
  reg instr_sw_t0;
  /* src = "generated/out/vanilla.sv:583.7-583.17" */
  wire instr_trap;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:583.7-583.17" */
  wire instr_trap_t0;
  /* src = "generated/out/vanilla.sv:566.6-566.15" */
  reg instr_xor;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:566.6-566.15" */
  reg instr_xor_t0;
  /* src = "generated/out/vanilla.sv:555.6-555.16" */
  reg instr_xori;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:555.6-555.16" */
  reg instr_xori_t0;
  /* src = "generated/out/vanilla.sv:108.15-108.18" */
  input [31:0] irq;
  wire [31:0] irq;
  /* cellift = 32'd1 */
  input [31:0] irq_t0;
  wire [31:0] irq_t0;
  /* src = "generated/out/vanilla.sv:605.6-605.20" */
  reg is_alu_reg_imm;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:605.6-605.20" */
  reg is_alu_reg_imm_t0;
  /* src = "generated/out/vanilla.sv:606.6-606.20" */
  reg is_alu_reg_reg;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:606.6-606.20" */
  reg is_alu_reg_reg_t0;
  /* src = "generated/out/vanilla.sv:603.6-603.34" */
  reg is_beq_bne_blt_bge_bltu_bgeu;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:603.6-603.34" */
  reg is_beq_bne_blt_bge_bltu_bgeu_t0;
  /* src = "generated/out/vanilla.sv:607.6-607.16" */
  reg is_compare;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:607.6-607.16" */
  reg is_compare_t0;
  /* src = "generated/out/vanilla.sv:597.6-597.43" */
  reg is_jalr_addi_slti_sltiu_xori_ori_andi;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:597.6-597.43" */
  reg is_jalr_addi_slti_sltiu_xori_ori_andi_t0;
  /* src = "generated/out/vanilla.sv:595.6-595.25" */
  reg is_lb_lh_lw_lbu_lhu;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:595.6-595.25" */
  reg is_lb_lh_lw_lbu_lhu_t0;
  /* src = "generated/out/vanilla.sv:594.6-594.22" */
  reg is_lui_auipc_jal;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:594.6-594.22" */
  reg is_lui_auipc_jal_t0;
  /* src = "generated/out/vanilla.sv:609.7-609.43" */
  wire is_rdcycle_rdcycleh_rdinstr_rdinstrh;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:609.7-609.43" */
  wire is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0;
  /* src = "generated/out/vanilla.sv:598.6-598.17" */
  reg is_sb_sh_sw;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:598.6-598.17" */
  reg is_sb_sh_sw_t0;
  /* src = "generated/out/vanilla.sv:599.6-599.20" */
  reg is_sll_srl_sra;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:599.6-599.20" */
  reg is_sll_srl_sra_t0;
  /* src = "generated/out/vanilla.sv:596.6-596.23" */
  reg is_slli_srli_srai;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:596.6-596.23" */
  reg is_slli_srli_srai_t0;
  /* src = "generated/out/vanilla.sv:601.6-601.21" */
  reg is_slti_blt_slt;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:601.6-601.21" */
  reg is_slti_blt_slt_t0;
  /* src = "generated/out/vanilla.sv:602.6-602.24" */
  reg is_sltiu_bltu_sltu;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:602.6-602.24" */
  reg is_sltiu_bltu_sltu_t0;
  /* src = "generated/out/vanilla.sv:285.6-285.20" */
  reg last_mem_valid;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:285.6-285.20" */
  reg last_mem_valid_t0;
  /* src = "generated/out/vanilla.sv:1072.6-1072.20" */
  reg latched_branch;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1072.6-1072.20" */
  reg latched_branch_t0;
  /* src = "generated/out/vanilla.sv:1073.6-1073.19" */
  reg latched_compr;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1073.6-1073.19" */
  reg latched_compr_t0;
  /* src = "generated/out/vanilla.sv:1077.6-1077.19" */
  reg latched_is_lb;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1077.6-1077.19" */
  reg latched_is_lb_t0;
  /* src = "generated/out/vanilla.sv:1076.6-1076.19" */
  reg latched_is_lh;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1076.6-1076.19" */
  reg latched_is_lh_t0;
  /* src = "generated/out/vanilla.sv:1078.28-1078.38" */
  reg [4:0] latched_rd;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1078.28-1078.38" */
  reg [4:0] latched_rd_t0;
  /* src = "generated/out/vanilla.sv:1071.6-1071.19" */
  reg latched_stalu;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1071.6-1071.19" */
  reg latched_stalu_t0;
  /* src = "generated/out/vanilla.sv:1070.6-1070.19" */
  reg latched_store;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1070.6-1070.19" */
  reg latched_store_t0;
  /* src = "generated/out/vanilla.sv:727.7-727.23" */
  wire launch_next_insn;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:727.7-727.23" */
  wire launch_next_insn_t0;
  /* src = "generated/out/vanilla.sv:290.13-290.29" */
  reg [15:0] mem_16bit_buffer;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:290.13-290.29" */
  reg [15:0] mem_16bit_buffer_t0;
  /* src = "generated/out/vanilla.sv:91.20-91.28" */
  output [31:0] mem_addr;
  reg [31:0] mem_addr;
  /* cellift = 32'd1 */
  output [31:0] mem_addr_t0;
  reg [31:0] mem_addr_t0;
  /* src = "generated/out/vanilla.sv:278.6-278.21" */
  reg mem_do_prefetch;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:278.6-278.21" */
  reg mem_do_prefetch_t0;
  /* src = "generated/out/vanilla.sv:280.6-280.18" */
  reg mem_do_rdata;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:280.6-280.18" */
  reg mem_do_rdata_t0;
  /* src = "generated/out/vanilla.sv:279.6-279.18" */
  reg mem_do_rinst;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:279.6-279.18" */
  reg mem_do_rinst_t0;
  /* src = "generated/out/vanilla.sv:281.6-281.18" */
  reg mem_do_wdata;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:281.6-281.18" */
  reg mem_do_wdata_t0;
  /* src = "generated/out/vanilla.sv:296.7-296.15" */
  wire mem_done;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:296.7-296.15" */
  wire mem_done_t0;
  /* src = "generated/out/vanilla.sv:89.13-89.22" */
  output mem_instr;
  reg mem_instr;
  /* cellift = 32'd1 */
  output mem_instr_t0;
  reg mem_instr_t0;
  /* src = "generated/out/vanilla.sv:97.21-97.32" */
  output [31:0] mem_la_addr;
  wire [31:0] mem_la_addr;
  /* cellift = 32'd1 */
  output [31:0] mem_la_addr_t0;
  wire [31:0] mem_la_addr_t0;
  /* src = "generated/out/vanilla.sv:286.7-286.23" */
  wire mem_la_firstword;
  /* src = "generated/out/vanilla.sv:284.6-284.26" */
  reg mem_la_firstword_reg;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:284.6-284.26" */
  reg mem_la_firstword_reg_t0;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:286.7-286.23" */
  wire mem_la_firstword_t0;
  /* src = "generated/out/vanilla.sv:287.7-287.28" */
  wire mem_la_firstword_xfer;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:287.7-287.28" */
  wire mem_la_firstword_xfer_t0;
  /* src = "generated/out/vanilla.sv:95.14-95.25" */
  output mem_la_read;
  wire mem_la_read;
  /* cellift = 32'd1 */
  output mem_la_read_t0;
  wire mem_la_read_t0;
  /* src = "generated/out/vanilla.sv:283.6-283.23" */
  reg mem_la_secondword;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:283.6-283.23" */
  reg mem_la_secondword_t0;
  /* src = "generated/out/vanilla.sv:293.7-293.38" */
  wire mem_la_use_prefetched_high_word;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:293.7-293.38" */
  wire mem_la_use_prefetched_high_word_t0;
  /* src = "generated/out/vanilla.sv:98.20-98.32" */
  output [31:0] mem_la_wdata;
  wire [31:0] mem_la_wdata;
  /* cellift = 32'd1 */
  output [31:0] mem_la_wdata_t0;
  wire [31:0] mem_la_wdata_t0;
  /* src = "generated/out/vanilla.sv:96.14-96.26" */
  output mem_la_write;
  wire mem_la_write;
  /* cellift = 32'd1 */
  output mem_la_write_t0;
  wire mem_la_write_t0;
  /* src = "generated/out/vanilla.sv:99.19-99.31" */
  output [3:0] mem_la_wstrb;
  wire [3:0] mem_la_wstrb;
  /* cellift = 32'd1 */
  output [3:0] mem_la_wstrb_t0;
  wire [3:0] mem_la_wstrb_t0;
  /* src = "generated/out/vanilla.sv:94.15-94.24" */
  input [31:0] mem_rdata;
  wire [31:0] mem_rdata;
  /* src = "generated/out/vanilla.sv:292.14-292.31" */
  wire [31:0] mem_rdata_latched;
  /* src = "generated/out/vanilla.sv:291.14-291.41" */
  wire [31:0] mem_rdata_latched_noshuffle;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:291.14-291.41" */
  wire [31:0] mem_rdata_latched_noshuffle_t0;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:292.14-292.31" */
  wire [31:0] mem_rdata_latched_t0;
  /* src = "generated/out/vanilla.sv:277.13-277.24" */
  reg [31:0] mem_rdata_q;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:277.13-277.24" */
  reg [31:0] mem_rdata_q_t0;
  /* cellift = 32'd1 */
  input [31:0] mem_rdata_t0;
  wire [31:0] mem_rdata_t0;
  /* src = "generated/out/vanilla.sv:276.13-276.27" */
  wire [31:0] mem_rdata_word;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:276.13-276.27" */
  wire [31:0] mem_rdata_word_t0;
  /* src = "generated/out/vanilla.sv:90.8-90.17" */
  input mem_ready;
  wire mem_ready;
  /* cellift = 32'd1 */
  input mem_ready_t0;
  wire mem_ready_t0;
  /* src = "generated/out/vanilla.sv:274.12-274.21" */
  reg [1:0] mem_state;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:274.12-274.21" */
  reg [1:0] mem_state_t0;
  /* src = "generated/out/vanilla.sv:88.13-88.22" */
  output mem_valid;
  reg mem_valid;
  /* cellift = 32'd1 */
  output mem_valid_t0;
  reg mem_valid_t0;
  /* src = "generated/out/vanilla.sv:92.20-92.29" */
  output [31:0] mem_wdata;
  reg [31:0] mem_wdata;
  /* cellift = 32'd1 */
  output [31:0] mem_wdata_t0;
  reg [31:0] mem_wdata_t0;
  /* src = "generated/out/vanilla.sv:275.12-275.24" */
  reg [1:0] mem_wordsize;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:275.12-275.24" */
  reg [1:0] mem_wordsize_t0;
  /* src = "generated/out/vanilla.sv:93.19-93.28" */
  output [3:0] mem_wstrb;
  reg [3:0] mem_wstrb;
  /* cellift = 32'd1 */
  output [3:0] mem_wstrb_t0;
  reg [3:0] mem_wstrb_t0;
  /* src = "generated/out/vanilla.sv:282.7-282.15" */
  wire mem_xfer;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:282.7-282.15" */
  wire mem_xfer_t0;
  /* src = "generated/out/vanilla.sv:159.13-159.29" */
  reg [31:0] next_insn_opcode;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:159.13-159.29" */
  reg [31:0] next_insn_opcode_t0;
  /* src = "generated/out/vanilla.sv:171.14-171.21" */
  /* unused_bits = "0" */
  wire [31:0] next_pc /* verilator public */;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:171.14-171.21" */
  /* unused_bits = "0" */
  wire [31:0] next_pc_t0 /* verilator public */;
  /* src = "generated/out/vanilla.sv:190.14-190.25" */
  wire [31:0] pcpi_div_rd;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:190.14-190.25" */
  wire [31:0] pcpi_div_rd_t0;
  /* src = "generated/out/vanilla.sv:192.7-192.21" */
  wire pcpi_div_ready;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:192.7-192.21" */
  wire pcpi_div_ready_t0;
  /* src = "generated/out/vanilla.sv:191.7-191.20" */
  wire pcpi_div_wait;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:191.7-191.20" */
  /* unused_bits = "0" */
  wire pcpi_div_wait_t0;
  /* src = "generated/out/vanilla.sv:189.7-189.18" */
  wire pcpi_div_wr;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:189.7-189.18" */
  wire pcpi_div_wr_t0;
  /* src = "generated/out/vanilla.sv:101.20-101.29" */
  output [31:0] pcpi_insn;
  reg [31:0] pcpi_insn;
  /* cellift = 32'd1 */
  output [31:0] pcpi_insn_t0;
  reg [31:0] pcpi_insn_t0;
  /* src = "generated/out/vanilla.sv:194.13-194.24" */
  wire [31:0] pcpi_int_rd;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:194.13-194.24" */
  wire [31:0] pcpi_int_rd_t0;
  /* src = "generated/out/vanilla.sv:196.6-196.20" */
  wire pcpi_int_ready;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:196.6-196.20" */
  wire pcpi_int_ready_t0;
  /* src = "generated/out/vanilla.sv:195.6-195.19" */
  wire pcpi_int_wait;
  /* src = "generated/out/vanilla.sv:193.6-193.17" */
  wire pcpi_int_wr;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:193.6-193.17" */
  wire pcpi_int_wr_t0;
  /* src = "generated/out/vanilla.sv:186.14-186.25" */
  wire [31:0] pcpi_mul_rd;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:186.14-186.25" */
  wire [31:0] pcpi_mul_rd_t0;
  /* src = "generated/out/vanilla.sv:188.7-188.21" */
  wire pcpi_mul_ready;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:188.7-188.21" */
  wire pcpi_mul_ready_t0;
  /* src = "generated/out/vanilla.sv:187.7-187.20" */
  wire pcpi_mul_wait;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:187.7-187.20" */
  /* unused_bits = "0" */
  wire pcpi_mul_wait_t0;
  /* src = "generated/out/vanilla.sv:185.7-185.18" */
  wire pcpi_mul_wr;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:185.7-185.18" */
  wire pcpi_mul_wr_t0;
  /* src = "generated/out/vanilla.sv:105.15-105.22" */
  input [31:0] pcpi_rd;
  wire [31:0] pcpi_rd;
  /* cellift = 32'd1 */
  input [31:0] pcpi_rd_t0;
  wire [31:0] pcpi_rd_t0;
  /* src = "generated/out/vanilla.sv:107.8-107.18" */
  input pcpi_ready;
  wire pcpi_ready;
  /* cellift = 32'd1 */
  input pcpi_ready_t0;
  wire pcpi_ready_t0;
  /* src = "generated/out/vanilla.sv:102.21-102.29" */
  output [31:0] pcpi_rs1;
  reg [31:0] pcpi_rs1;
  /* cellift = 32'd1 */
  output [31:0] pcpi_rs1_t0;
  reg [31:0] pcpi_rs1_t0;
  /* src = "generated/out/vanilla.sv:103.21-103.29" */
  output [31:0] pcpi_rs2;
  reg [31:0] pcpi_rs2;
  /* cellift = 32'd1 */
  output [31:0] pcpi_rs2_t0;
  reg [31:0] pcpi_rs2_t0;
  /* src = "generated/out/vanilla.sv:1082.6-1082.18" */
  reg pcpi_timeout;
  /* src = "generated/out/vanilla.sv:1081.12-1081.32" */
  reg [3:0] pcpi_timeout_counter;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1081.12-1081.32" */
  reg [3:0] pcpi_timeout_counter_t0;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1082.6-1082.18" */
  reg pcpi_timeout_t0;
  /* src = "generated/out/vanilla.sv:100.13-100.23" */
  output pcpi_valid;
  reg pcpi_valid;
  /* cellift = 32'd1 */
  output pcpi_valid_t0;
  reg pcpi_valid_t0;
  /* src = "generated/out/vanilla.sv:106.8-106.17" */
  input pcpi_wait;
  wire pcpi_wait;
  /* cellift = 32'd1 */
  input pcpi_wait_t0;
  wire pcpi_wait_t0;
  /* src = "generated/out/vanilla.sv:104.8-104.15" */
  input pcpi_wr;
  wire pcpi_wr;
  /* cellift = 32'd1 */
  input pcpi_wr_t0;
  wire pcpi_wr_t0;
  /* src = "generated/out/vanilla.sv:288.6-288.26" */
  reg prefetched_high_word;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:288.6-288.26" */
  reg prefetched_high_word_t0;
  /* src = "generated/out/vanilla.sv:723.12-723.22" */
  reg [4:0] q_insn_rs1;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:723.12-723.22" */
  reg [4:0] q_insn_rs1_t0;
  /* src = "generated/out/vanilla.sv:724.12-724.22" */
  reg [4:0] q_insn_rs2;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:724.12-724.22" */
  reg [4:0] q_insn_rs2_t0;
  /* src = "generated/out/vanilla.sv:154.13-154.24" */
  reg [31:0] reg_next_pc;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:154.13-154.24" */
  reg [31:0] reg_next_pc_t0;
  /* src = "generated/out/vanilla.sv:157.13-157.20" */
  reg [31:0] reg_out;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:157.13-157.20" */
  reg [31:0] reg_out_t0;
  /* src = "generated/out/vanilla.sv:153.13-153.19" */
  reg [31:0] reg_pc;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:153.13-153.19" */
  reg [31:0] reg_pc_t0;
  /* src = "generated/out/vanilla.sv:158.12-158.18" */
  reg [4:0] reg_sh;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:158.12-158.18" */
  reg [4:0] reg_sh_t0;
  /* src = "generated/out/vanilla.sv:86.8-86.14" */
  input resetn;
  wire resetn;
  /* src = "generated/out/vanilla.sv:133.20-133.41" */
  output [63:0] rvfi_csr_mcycle_rdata;
  wire [63:0] rvfi_csr_mcycle_rdata;
  /* cellift = 32'd1 */
  output [63:0] rvfi_csr_mcycle_rdata_t0;
  wire [63:0] rvfi_csr_mcycle_rdata_t0;
  /* src = "generated/out/vanilla.sv:131.20-131.41" */
  output [63:0] rvfi_csr_mcycle_rmask;
  wire [63:0] rvfi_csr_mcycle_rmask;
  /* cellift = 32'd1 */
  output [63:0] rvfi_csr_mcycle_rmask_t0;
  wire [63:0] rvfi_csr_mcycle_rmask_t0;
  /* src = "generated/out/vanilla.sv:134.20-134.41" */
  output [63:0] rvfi_csr_mcycle_wdata;
  wire [63:0] rvfi_csr_mcycle_wdata;
  /* cellift = 32'd1 */
  output [63:0] rvfi_csr_mcycle_wdata_t0;
  wire [63:0] rvfi_csr_mcycle_wdata_t0;
  /* src = "generated/out/vanilla.sv:132.20-132.41" */
  output [63:0] rvfi_csr_mcycle_wmask;
  wire [63:0] rvfi_csr_mcycle_wmask;
  /* cellift = 32'd1 */
  output [63:0] rvfi_csr_mcycle_wmask_t0;
  wire [63:0] rvfi_csr_mcycle_wmask_t0;
  /* src = "generated/out/vanilla.sv:137.20-137.43" */
  output [63:0] rvfi_csr_minstret_rdata;
  wire [63:0] rvfi_csr_minstret_rdata;
  /* cellift = 32'd1 */
  output [63:0] rvfi_csr_minstret_rdata_t0;
  wire [63:0] rvfi_csr_minstret_rdata_t0;
  /* src = "generated/out/vanilla.sv:135.20-135.43" */
  output [63:0] rvfi_csr_minstret_rmask;
  wire [63:0] rvfi_csr_minstret_rmask;
  /* cellift = 32'd1 */
  output [63:0] rvfi_csr_minstret_rmask_t0;
  wire [63:0] rvfi_csr_minstret_rmask_t0;
  /* src = "generated/out/vanilla.sv:138.20-138.43" */
  output [63:0] rvfi_csr_minstret_wdata;
  wire [63:0] rvfi_csr_minstret_wdata;
  /* cellift = 32'd1 */
  output [63:0] rvfi_csr_minstret_wdata_t0;
  wire [63:0] rvfi_csr_minstret_wdata_t0;
  /* src = "generated/out/vanilla.sv:136.20-136.43" */
  output [63:0] rvfi_csr_minstret_wmask;
  wire [63:0] rvfi_csr_minstret_wmask;
  /* cellift = 32'd1 */
  output [63:0] rvfi_csr_minstret_wmask_t0;
  wire [63:0] rvfi_csr_minstret_wmask_t0;
  /* src = "generated/out/vanilla.sv:114.13-114.22" */
  output rvfi_halt;
  reg rvfi_halt;
  /* cellift = 32'd1 */
  output rvfi_halt_t0;
  reg rvfi_halt_t0;
  /* src = "generated/out/vanilla.sv:112.20-112.29" */
  output [31:0] rvfi_insn;
  wire [31:0] rvfi_insn;
  /* cellift = 32'd1 */
  output [31:0] rvfi_insn_t0;
  wire [31:0] rvfi_insn_t0;
  /* src = "generated/out/vanilla.sv:115.13-115.22" */
  output rvfi_intr;
  wire rvfi_intr;
  /* cellift = 32'd1 */
  output rvfi_intr_t0;
  wire rvfi_intr_t0;
  /* src = "generated/out/vanilla.sv:117.19-117.27" */
  output [1:0] rvfi_ixl;
  wire [1:0] rvfi_ixl;
  /* cellift = 32'd1 */
  output [1:0] rvfi_ixl_t0;
  wire [1:0] rvfi_ixl_t0;
  /* src = "generated/out/vanilla.sv:126.20-126.33" */
  output [31:0] rvfi_mem_addr;
  reg [31:0] rvfi_mem_addr;
  /* cellift = 32'd1 */
  output [31:0] rvfi_mem_addr_t0;
  reg [31:0] rvfi_mem_addr_t0;
  /* src = "generated/out/vanilla.sv:129.20-129.34" */
  output [31:0] rvfi_mem_rdata;
  reg [31:0] rvfi_mem_rdata;
  /* cellift = 32'd1 */
  output [31:0] rvfi_mem_rdata_t0;
  reg [31:0] rvfi_mem_rdata_t0;
  /* src = "generated/out/vanilla.sv:127.19-127.33" */
  output [3:0] rvfi_mem_rmask;
  reg [3:0] rvfi_mem_rmask;
  /* cellift = 32'd1 */
  output [3:0] rvfi_mem_rmask_t0;
  reg [3:0] rvfi_mem_rmask_t0;
  /* src = "generated/out/vanilla.sv:130.20-130.34" */
  output [31:0] rvfi_mem_wdata;
  reg [31:0] rvfi_mem_wdata;
  /* cellift = 32'd1 */
  output [31:0] rvfi_mem_wdata_t0;
  reg [31:0] rvfi_mem_wdata_t0;
  /* src = "generated/out/vanilla.sv:128.19-128.33" */
  output [3:0] rvfi_mem_wmask;
  reg [3:0] rvfi_mem_wmask;
  /* cellift = 32'd1 */
  output [3:0] rvfi_mem_wmask_t0;
  reg [3:0] rvfi_mem_wmask_t0;
  /* src = "generated/out/vanilla.sv:116.19-116.28" */
  output [1:0] rvfi_mode;
  wire [1:0] rvfi_mode;
  /* cellift = 32'd1 */
  output [1:0] rvfi_mode_t0;
  wire [1:0] rvfi_mode_t0;
  /* src = "generated/out/vanilla.sv:111.20-111.30" */
  output [63:0] rvfi_order;
  reg [63:0] rvfi_order;
  /* cellift = 32'd1 */
  output [63:0] rvfi_order_t0;
  reg [63:0] rvfi_order_t0;
  /* src = "generated/out/vanilla.sv:124.20-124.33" */
  output [31:0] rvfi_pc_rdata;
  reg [31:0] rvfi_pc_rdata;
  /* cellift = 32'd1 */
  output [31:0] rvfi_pc_rdata_t0;
  reg [31:0] rvfi_pc_rdata_t0;
  /* src = "generated/out/vanilla.sv:125.20-125.33" */
  output [31:0] rvfi_pc_wdata;
  reg [31:0] rvfi_pc_wdata;
  /* cellift = 32'd1 */
  output [31:0] rvfi_pc_wdata_t0;
  reg [31:0] rvfi_pc_wdata_t0;
  /* src = "generated/out/vanilla.sv:122.19-122.31" */
  output [4:0] rvfi_rd_addr;
  reg [4:0] rvfi_rd_addr;
  /* cellift = 32'd1 */
  output [4:0] rvfi_rd_addr_t0;
  reg [4:0] rvfi_rd_addr_t0;
  /* src = "generated/out/vanilla.sv:123.20-123.33" */
  output [31:0] rvfi_rd_wdata;
  reg [31:0] rvfi_rd_wdata;
  /* cellift = 32'd1 */
  output [31:0] rvfi_rd_wdata_t0;
  reg [31:0] rvfi_rd_wdata_t0;
  /* src = "generated/out/vanilla.sv:118.19-118.32" */
  output [4:0] rvfi_rs1_addr;
  reg [4:0] rvfi_rs1_addr;
  /* cellift = 32'd1 */
  output [4:0] rvfi_rs1_addr_t0;
  reg [4:0] rvfi_rs1_addr_t0;
  /* src = "generated/out/vanilla.sv:120.20-120.34" */
  output [31:0] rvfi_rs1_rdata;
  reg [31:0] rvfi_rs1_rdata;
  /* cellift = 32'd1 */
  output [31:0] rvfi_rs1_rdata_t0;
  reg [31:0] rvfi_rs1_rdata_t0;
  /* src = "generated/out/vanilla.sv:119.19-119.32" */
  output [4:0] rvfi_rs2_addr;
  reg [4:0] rvfi_rs2_addr;
  /* cellift = 32'd1 */
  output [4:0] rvfi_rs2_addr_t0;
  reg [4:0] rvfi_rs2_addr_t0;
  /* src = "generated/out/vanilla.sv:121.20-121.34" */
  output [31:0] rvfi_rs2_rdata;
  reg [31:0] rvfi_rs2_rdata;
  /* cellift = 32'd1 */
  output [31:0] rvfi_rs2_rdata_t0;
  reg [31:0] rvfi_rs2_rdata_t0;
  /* src = "generated/out/vanilla.sv:113.13-113.22" */
  output rvfi_trap;
  wire rvfi_trap;
  /* cellift = 32'd1 */
  output rvfi_trap_t0;
  wire rvfi_trap_t0;
  /* src = "generated/out/vanilla.sv:110.13-110.23" */
  output rvfi_valid;
  reg rvfi_valid;
  /* cellift = 32'd1 */
  output rvfi_valid_t0;
  reg rvfi_valid_t0;
  /* src = "generated/out/vanilla.sv:140.20-140.30" */
  output [35:0] trace_data;
  wire [35:0] trace_data;
  /* cellift = 32'd1 */
  output [35:0] trace_data_t0;
  wire [35:0] trace_data_t0;
  /* src = "generated/out/vanilla.sv:139.13-139.24" */
  output trace_valid;
  wire trace_valid;
  /* cellift = 32'd1 */
  output trace_valid_t0;
  wire trace_valid_t0;
  /* src = "generated/out/vanilla.sv:87.13-87.17" */
  output trap;
  reg trap;
  /* cellift = 32'd1 */
  output trap_t0;
  reg trap_t0;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME _00080_ */
  always_ff @(posedge clk)
    _00080_ <= _06102_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME _00082_ */
  always_ff @(posedge clk)
    _00082_ <= _06104_;
  assign _00084_ = pcpi_rs1 + /* src = "generated/out/vanilla.sv:1110.52-1110.69" */ pcpi_rs2;
  assign _00086_ = reg_pc + /* src = "generated/out/vanilla.sv:1163.23-1163.55" */ _07591_;
  assign _00088_ = count_cycle + /* src = "generated/out/vanilla.sv:1223.29-1223.44" */ 32'd1;
  assign _00090_ = _00060_ + /* src = "generated/out/vanilla.sv:1331.22-1331.61" */ _07596_;
  assign _00092_ = count_instr + /* src = "generated/out/vanilla.sv:1335.23-1335.38" */ 32'd1;
  assign _00094_ = _00060_ + /* src = "generated/out/vanilla.sv:1341.23-1341.49" */ { decoded_imm_j[31:1], 1'h0 };
  assign _00096_ = reg_pc + /* src = "generated/out/vanilla.sv:1554.17-1554.37" */ decoded_imm;
  assign _00098_ = pcpi_rs1 + /* src = "generated/out/vanilla.sv:1645.19-1645.40" */ decoded_imm;
  assign _00100_ = rvfi_order + /* src = "generated/out/vanilla.sv:1716.27-1716.50" */ rvfi_valid;
  assign _00102_ = next_pc[31:2] + /* src = "generated/out/vanilla.sv:299.59-299.96" */ mem_la_firstword_xfer;
  assign _00104_ = 32'd8 + /* src = "generated/out/vanilla.sv:886.25-886.51" */ mem_rdata_latched[4:2];
  assign _00106_ = 32'd8 + /* src = "generated/out/vanilla.sv:897.24-897.50" */ mem_rdata_latched[9:7];
  assign _00108_ = pcpi_rs1 & /* src = "generated/out/vanilla.sv:1137.39-1137.56" */ pcpi_rs2;
  assign _00112_ = mem_la_wstrb & /* src = "generated/out/vanilla.sv:472.18-472.51" */ { mem_la_write, mem_la_write, mem_la_write, mem_la_write };
  assign _00116_ = ~ count_cycle_t0;
  assign _00117_ = ~ _00061_;
  assign _00118_ = ~ count_instr_t0;
  assign _00115_ = ~ reg_pc_t0;
  assign _00114_ = ~ pcpi_rs1_t0;
  assign _00119_ = ~ rvfi_order_t0;
  assign _00120_ = ~ next_pc_t0[31:2];
  assign _00121_ = ~ pcpi_rs2_t0;
  assign _00122_ = ~ { 29'h00000000, latched_compr_t0, latched_compr_t0, 1'h0 };
  assign _00123_ = ~ { 29'h00000000, compressed_instr_t0, compressed_instr_t0, 1'h0 };
  assign _00124_ = ~ { decoded_imm_j_t0[31:1], 1'h0 };
  assign _00125_ = ~ decoded_imm_t0;
  assign _00126_ = ~ { 63'h0000000000000000, rvfi_valid_t0 };
  assign _00127_ = ~ { 29'h00000000, mem_la_firstword_xfer_t0 };
  assign _00128_ = ~ { 29'h00000000, mem_rdata_latched_t0[4:2] };
  assign _00129_ = ~ { 29'h00000000, mem_rdata_latched_t0[9:7] };
  assign _03321_ = pcpi_rs1 & _00114_;
  assign _03458_ = count_cycle & _00116_;
  assign _03459_ = _00060_ & _00117_;
  assign _03461_ = count_instr & _00118_;
  assign _03456_ = reg_pc & _00115_;
  assign _03464_ = rvfi_order & _00119_;
  assign _03466_ = next_pc[31:2] & _00120_;
  assign _03322_ = pcpi_rs2 & _00121_;
  assign _03457_ = _07591_ & _00122_;
  assign _03460_ = _07596_ & _00123_;
  assign _03462_ = { decoded_imm_j[31:1], 1'h0 } & _00124_;
  assign _03463_ = decoded_imm & _00125_;
  assign _03465_ = { 63'h0000000000000000, rvfi_valid } & _00126_;
  assign _03467_ = { 29'h00000000, mem_la_firstword_xfer } & _00127_;
  assign _03468_ = { 29'h00000000, mem_rdata_latched[4:2] } & _00128_;
  assign _03469_ = { 29'h00000000, mem_rdata_latched[9:7] } & _00129_;
  assign _06070_ = _03321_ + _03322_;
  assign _06072_ = _03456_ + _03457_;
  assign _06074_ = _03458_ + 64'h0000000000000001;
  assign _06076_ = _03459_ + _03460_;
  assign _06078_ = _03461_ + 64'h0000000000000001;
  assign _06080_ = _03459_ + _03462_;
  assign _06082_ = _03456_ + _03463_;
  assign _06084_ = _03321_ + _03463_;
  assign _06086_ = _03464_ + _03465_;
  assign _06088_ = _03466_ + _03467_;
  assign _06090_ = 32'd8 + _03468_;
  assign _06092_ = 32'd8 + _03469_;
  assign _05064_ = pcpi_rs1 | pcpi_rs1_t0;
  assign _05140_ = count_cycle | count_cycle_t0;
  assign _05141_ = _00060_ | _00061_;
  assign _05144_ = count_instr | count_instr_t0;
  assign _05137_ = reg_pc | reg_pc_t0;
  assign _05150_ = rvfi_order | rvfi_order_t0;
  assign _05153_ = next_pc[31:2] | next_pc_t0[31:2];
  assign _05065_ = pcpi_rs2 | pcpi_rs2_t0;
  assign _05138_ = _07591_ | { 29'h00000000, latched_compr_t0, latched_compr_t0, 1'h0 };
  assign _05142_ = _07596_ | { 29'h00000000, compressed_instr_t0, compressed_instr_t0, 1'h0 };
  assign _05145_ = { decoded_imm_j[31:1], 1'h0 } | { decoded_imm_j_t0[31:1], 1'h0 };
  assign _05147_ = decoded_imm | decoded_imm_t0;
  assign _05151_ = { 63'h0000000000000000, rvfi_valid } | { 63'h0000000000000000, rvfi_valid_t0 };
  assign _05154_ = { 29'h00000000, mem_la_firstword_xfer } | { 29'h00000000, mem_la_firstword_xfer_t0 };
  assign _05156_ = { 29'h00000000, mem_rdata_latched[4:2] } | { 29'h00000000, mem_rdata_latched_t0[4:2] };
  assign _05158_ = { 29'h00000000, mem_rdata_latched[9:7] } | { 29'h00000000, mem_rdata_latched_t0[9:7] };
  assign _06071_ = _05064_ + _05065_;
  assign _06073_ = _05137_ + _05138_;
  assign _06075_ = _05140_ + 64'h0000000000000001;
  assign _06077_ = _05141_ + _05142_;
  assign _06079_ = _05144_ + 64'h0000000000000001;
  assign _06081_ = _05141_ + _05145_;
  assign _06083_ = _05137_ + _05147_;
  assign _06085_ = _05064_ + _05147_;
  assign _06087_ = _05150_ + _05151_;
  assign _06089_ = _05153_ + _05154_;
  assign _06091_ = 32'd8 + _05156_;
  assign _06093_ = 32'd8 + _05158_;
  assign _05895_ = _06070_ ^ _06071_;
  assign _05896_ = _06072_ ^ _06073_;
  assign _05897_ = _06074_ ^ _06075_;
  assign _05898_ = _06076_ ^ _06077_;
  assign _05899_ = _06078_ ^ _06079_;
  assign _05900_ = _06080_ ^ _06081_;
  assign _05901_ = _06082_ ^ _06083_;
  assign _05902_ = _06084_ ^ _06085_;
  assign _05903_ = _06086_ ^ _06087_;
  assign _05904_ = _06088_ ^ _06089_;
  assign _05157_ = _06090_ ^ _06091_;
  assign _05159_ = _06092_ ^ _06093_;
  assign _05136_ = _05895_ | pcpi_rs1_t0;
  assign _05139_ = _05896_ | reg_pc_t0;
  assign _00089_ = _05897_ | count_cycle_t0;
  assign _05143_ = _05898_ | _00061_;
  assign _00093_ = _05899_ | count_instr_t0;
  assign _05146_ = _05900_ | _00061_;
  assign _05148_ = _05901_ | reg_pc_t0;
  assign _05149_ = _05902_ | pcpi_rs1_t0;
  assign _05152_ = _05903_ | rvfi_order_t0;
  assign _05155_ = _05904_ | next_pc_t0[31:2];
  assign _00085_ = _05136_ | pcpi_rs2_t0;
  assign _00087_ = _05139_ | { 29'h00000000, latched_compr_t0, latched_compr_t0, 1'h0 };
  assign _00091_ = _05143_ | { 29'h00000000, compressed_instr_t0, compressed_instr_t0, 1'h0 };
  assign _00095_ = _05146_ | { decoded_imm_j_t0[31:1], 1'h0 };
  assign _00097_ = _05148_ | decoded_imm_t0;
  assign _00099_ = _05149_ | decoded_imm_t0;
  assign _00101_ = _05152_ | { 63'h0000000000000000, rvfi_valid_t0 };
  assign _00103_ = _05155_ | { 29'h00000000, mem_la_firstword_xfer_t0 };
  assign _00105_ = _05157_ | { 29'h00000000, mem_rdata_latched_t0[4:2] };
  assign _00107_ = _05159_ | { 29'h00000000, mem_rdata_latched_t0[9:7] };
  assign _01333_ = _00001_[0] & _06066_;
  assign _01336_ = _00001_[3] & _06069_;
  assign _01339_ = _00001_[2] & _03362_;
  assign _01342_ = _03361_ & _03364_;
  assign _01346_ = _03369_ & _03364_;
  assign _01350_ = _03373_ & _03364_;
  assign _01349_ = _00001_[0] & _00000_[1];
  assign _01353_ = _03377_ & _03364_;
  assign _01357_ = _03361_ & _03380_;
  assign _01360_ = _03369_ & _03380_;
  assign _01363_ = _03373_ & _03380_;
  assign _01366_ = _03377_ & _03380_;
  assign _01373_ = _03361_ & _03392_;
  assign _01376_ = _03369_ & _03392_;
  assign _01379_ = _03373_ & _03392_;
  assign _01382_ = _03377_ & _03392_;
  assign _01370_ = _00001_[2] & _03390_;
  assign _01386_ = _03361_ & _03402_;
  assign _01389_ = _03369_ & _03402_;
  assign _01392_ = _03373_ & _03402_;
  assign _01395_ = _03377_ & _03402_;
  assign _01399_ = _00001_[2] & _03412_;
  assign _01402_ = _03361_ & _03414_;
  assign _01405_ = _03369_ & _03414_;
  assign _01408_ = _03373_ & _03414_;
  assign _01411_ = _03377_ & _03414_;
  assign _01415_ = _03361_ & _03424_;
  assign _01418_ = _03369_ & _03424_;
  assign _01421_ = _03373_ & _03424_;
  assign _01424_ = _03377_ & _03424_;
  assign _01398_ = _00001_[3] & _00000_[4];
  assign _01427_ = _00001_[2] & _03434_;
  assign _01430_ = _03361_ & _03436_;
  assign _01433_ = _03369_ & _03436_;
  assign _01436_ = _03373_ & _03436_;
  assign _01439_ = _03377_ & _03436_;
  assign _01443_ = _03361_ & _03446_;
  assign _01446_ = _03369_ & _03446_;
  assign _01449_ = _03373_ & _03446_;
  assign _01452_ = _03377_ & _03446_;
  assign _02681_ = _03367_ & _00004_[31];
  assign _02684_ = _03399_ & _00004_[31];
  assign _02687_ = _03401_ & _00004_[31];
  assign _02690_ = _03405_ & _00004_[31];
  assign _02693_ = _03407_ & _00004_[31];
  assign _02696_ = _03409_ & _00004_[31];
  assign _02699_ = _03411_ & _00004_[31];
  assign _02702_ = _03417_ & _00004_[31];
  assign _02705_ = _03419_ & _00004_[31];
  assign _02708_ = _03421_ & _00004_[31];
  assign _02711_ = _03423_ & _00004_[31];
  assign _02714_ = _03371_ & _00004_[31];
  assign _02717_ = _03427_ & _00004_[31];
  assign _02720_ = _03429_ & _00004_[31];
  assign _02723_ = _03431_ & _00004_[31];
  assign _02726_ = _03433_ & _00004_[31];
  assign _02729_ = _03439_ & _00004_[31];
  assign _02732_ = _03441_ & _00004_[31];
  assign _02735_ = _03443_ & _00004_[31];
  assign _02738_ = _03445_ & _00004_[31];
  assign _02741_ = _03449_ & _00004_[31];
  assign _02744_ = _03451_ & _00004_[31];
  assign _02747_ = _03375_ & _00004_[31];
  assign _02750_ = _03453_ & _00004_[31];
  assign _02753_ = _03455_ & _00004_[31];
  assign _02756_ = _03379_ & _00004_[31];
  assign _02759_ = _03383_ & _00004_[31];
  assign _02762_ = _03385_ & _00004_[31];
  assign _02765_ = _03387_ & _00004_[31];
  assign _02768_ = _03389_ & _00004_[31];
  assign _02771_ = _03395_ & _00004_[31];
  assign _02774_ = _03397_ & _00004_[31];
  assign _03470_ = pcpi_rs1_t0 & pcpi_rs2;
  assign _03472_ = mem_la_wstrb_t0 & { mem_la_write, mem_la_write, mem_la_write, mem_la_write };
  assign _01340_ = _03363_ & _06067_;
  assign _01343_ = _03365_ & _03360_;
  assign _01345_ = _00001_[1] & _00000_[0];
  assign _01347_ = _03365_ & _03368_;
  assign _01334_ = _00001_[1] & _06065_;
  assign _01351_ = _03365_ & _03372_;
  assign _01354_ = _03365_ & _03376_;
  assign _01356_ = _03363_ & _00000_[2];
  assign _01358_ = _03381_ & _03360_;
  assign _01361_ = _03381_ & _03368_;
  assign _01364_ = _03381_ & _03372_;
  assign _01367_ = _03381_ & _03376_;
  assign _01369_ = _00001_[4] & _00000_[3];
  assign _01371_ = _03391_ & _06067_;
  assign _01374_ = _03393_ & _03360_;
  assign _01377_ = _03393_ & _03368_;
  assign _01380_ = _03393_ & _03372_;
  assign _01383_ = _03393_ & _03376_;
  assign _01385_ = _03391_ & _00000_[2];
  assign _01387_ = _03403_ & _03360_;
  assign _01390_ = _03403_ & _03368_;
  assign _01393_ = _03403_ & _03372_;
  assign _01396_ = _03403_ & _03376_;
  assign _01337_ = _00001_[4] & _06068_;
  assign _01400_ = _03413_ & _06067_;
  assign _01403_ = _03415_ & _03360_;
  assign _01406_ = _03415_ & _03368_;
  assign _01409_ = _03415_ & _03372_;
  assign _01412_ = _03415_ & _03376_;
  assign _01414_ = _03413_ & _00000_[2];
  assign _01416_ = _03425_ & _03360_;
  assign _01419_ = _03425_ & _03368_;
  assign _01422_ = _03425_ & _03372_;
  assign _01425_ = _03425_ & _03376_;
  assign _01428_ = _03435_ & _06067_;
  assign _01431_ = _03437_ & _03360_;
  assign _01434_ = _03437_ & _03368_;
  assign _01437_ = _03437_ & _03372_;
  assign _01440_ = _03437_ & _03376_;
  assign _01442_ = _03435_ & _00000_[2];
  assign _01444_ = _03447_ & _03360_;
  assign _01447_ = _03447_ & _03368_;
  assign _01450_ = _03447_ & _03372_;
  assign _01453_ = _03447_ & _03376_;
  assign _02682_ = _00005_[31] & _03366_;
  assign _02685_ = _00005_[31] & _03398_;
  assign _02688_ = _00005_[31] & _03400_;
  assign _02691_ = _00005_[31] & _03404_;
  assign _02694_ = _00005_[31] & _03406_;
  assign _02697_ = _00005_[31] & _03408_;
  assign _02700_ = _00005_[31] & _03410_;
  assign _02703_ = _00005_[31] & _03416_;
  assign _02706_ = _00005_[31] & _03418_;
  assign _02709_ = _00005_[31] & _03420_;
  assign _02712_ = _00005_[31] & _03422_;
  assign _02715_ = _00005_[31] & _03370_;
  assign _02718_ = _00005_[31] & _03426_;
  assign _02721_ = _00005_[31] & _03428_;
  assign _02724_ = _00005_[31] & _03430_;
  assign _02727_ = _00005_[31] & _03432_;
  assign _02730_ = _00005_[31] & _03438_;
  assign _02733_ = _00005_[31] & _03440_;
  assign _02736_ = _00005_[31] & _03442_;
  assign _02739_ = _00005_[31] & _03444_;
  assign _02742_ = _00005_[31] & _03448_;
  assign _02745_ = _00005_[31] & _03450_;
  assign _02748_ = _00005_[31] & _03374_;
  assign _02751_ = _00005_[31] & _03452_;
  assign _02754_ = _00005_[31] & _03454_;
  assign _02757_ = _00005_[31] & _03378_;
  assign _02760_ = _00005_[31] & _03382_;
  assign _02763_ = _00005_[31] & _03384_;
  assign _02766_ = _00005_[31] & _03386_;
  assign _02769_ = _00005_[31] & _03388_;
  assign _02772_ = _00005_[31] & _03394_;
  assign _02775_ = _00005_[31] & _03396_;
  assign _03471_ = pcpi_rs2_t0 & pcpi_rs1;
  assign _03473_ = { mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0 } & mem_la_wstrb;
  assign _01335_ = _00001_[0] & _00001_[1];
  assign _01338_ = _00001_[3] & _00001_[4];
  assign _01341_ = _00001_[2] & _03363_;
  assign _01344_ = _03361_ & _03365_;
  assign _01348_ = _03369_ & _03365_;
  assign _01352_ = _03373_ & _03365_;
  assign _01355_ = _03377_ & _03365_;
  assign _01359_ = _03361_ & _03381_;
  assign _01362_ = _03369_ & _03381_;
  assign _01365_ = _03373_ & _03381_;
  assign _01368_ = _03377_ & _03381_;
  assign _01375_ = _03361_ & _03393_;
  assign _01378_ = _03369_ & _03393_;
  assign _01381_ = _03373_ & _03393_;
  assign _01384_ = _03377_ & _03393_;
  assign _01372_ = _00001_[2] & _03391_;
  assign _01388_ = _03361_ & _03403_;
  assign _01391_ = _03369_ & _03403_;
  assign _01394_ = _03373_ & _03403_;
  assign _01397_ = _03377_ & _03403_;
  assign _01401_ = _00001_[2] & _03413_;
  assign _01404_ = _03361_ & _03415_;
  assign _01407_ = _03369_ & _03415_;
  assign _01410_ = _03373_ & _03415_;
  assign _01413_ = _03377_ & _03415_;
  assign _01417_ = _03361_ & _03425_;
  assign _01420_ = _03369_ & _03425_;
  assign _01423_ = _03373_ & _03425_;
  assign _01426_ = _03377_ & _03425_;
  assign _01432_ = _03361_ & _03437_;
  assign _01435_ = _03369_ & _03437_;
  assign _01438_ = _03373_ & _03437_;
  assign _01441_ = _03377_ & _03437_;
  assign _01429_ = _00001_[2] & _03435_;
  assign _01445_ = _03361_ & _03447_;
  assign _01448_ = _03369_ & _03447_;
  assign _01451_ = _03373_ & _03447_;
  assign _01454_ = _03377_ & _03447_;
  assign _02683_ = _03367_ & _00005_[31];
  assign _02686_ = _03399_ & _00005_[31];
  assign _02689_ = _03401_ & _00005_[31];
  assign _02692_ = _03405_ & _00005_[31];
  assign _02695_ = _03407_ & _00005_[31];
  assign _02698_ = _03409_ & _00005_[31];
  assign _02701_ = _03411_ & _00005_[31];
  assign _02704_ = _03417_ & _00005_[31];
  assign _02707_ = _03419_ & _00005_[31];
  assign _02710_ = _03421_ & _00005_[31];
  assign _02713_ = _03423_ & _00005_[31];
  assign _02716_ = _03371_ & _00005_[31];
  assign _02719_ = _03427_ & _00005_[31];
  assign _02722_ = _03429_ & _00005_[31];
  assign _02725_ = _03431_ & _00005_[31];
  assign _02728_ = _03433_ & _00005_[31];
  assign _02731_ = _03439_ & _00005_[31];
  assign _02734_ = _03441_ & _00005_[31];
  assign _02737_ = _03443_ & _00005_[31];
  assign _02740_ = _03445_ & _00005_[31];
  assign _02743_ = _03449_ & _00005_[31];
  assign _02746_ = _03451_ & _00005_[31];
  assign _02749_ = _03375_ & _00005_[31];
  assign _02752_ = _03453_ & _00005_[31];
  assign _02755_ = _03455_ & _00005_[31];
  assign _02758_ = _03379_ & _00005_[31];
  assign _02761_ = _03383_ & _00005_[31];
  assign _02764_ = _03385_ & _00005_[31];
  assign _02767_ = _03387_ & _00005_[31];
  assign _02770_ = _03389_ & _00005_[31];
  assign _02773_ = _03395_ & _00005_[31];
  assign _02776_ = _03397_ & _00005_[31];
  assign _02782_ = pcpi_rs1_t0 & pcpi_rs2_t0;
  assign _03474_ = mem_la_wstrb_t0 & { mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0 };
  assign _03985_ = _01333_ | _01334_;
  assign _03986_ = _01336_ | _01337_;
  assign _03987_ = _01339_ | _01340_;
  assign _03988_ = _01342_ | _01343_;
  assign _03989_ = _01333_ | _01345_;
  assign _03990_ = _01346_ | _01347_;
  assign _03991_ = _01349_ | _01334_;
  assign _03992_ = _01350_ | _01351_;
  assign _03993_ = _01349_ | _01345_;
  assign _03994_ = _01353_ | _01354_;
  assign _03995_ = _01339_ | _01356_;
  assign _03996_ = _01357_ | _01358_;
  assign _03997_ = _01360_ | _01361_;
  assign _03998_ = _01363_ | _01364_;
  assign _03999_ = _01366_ | _01367_;
  assign _04000_ = _01336_ | _01369_;
  assign _04001_ = _01370_ | _01371_;
  assign _04002_ = _01373_ | _01374_;
  assign _04003_ = _01376_ | _01377_;
  assign _04004_ = _01379_ | _01380_;
  assign _04005_ = _01382_ | _01383_;
  assign _04006_ = _01370_ | _01385_;
  assign _04007_ = _01386_ | _01387_;
  assign _04008_ = _01389_ | _01390_;
  assign _04009_ = _01392_ | _01393_;
  assign _04010_ = _01395_ | _01396_;
  assign _04011_ = _01398_ | _01337_;
  assign _04012_ = _01399_ | _01400_;
  assign _04013_ = _01402_ | _01403_;
  assign _04014_ = _01405_ | _01406_;
  assign _04015_ = _01408_ | _01409_;
  assign _04016_ = _01411_ | _01412_;
  assign _04017_ = _01399_ | _01414_;
  assign _04018_ = _01415_ | _01416_;
  assign _04019_ = _01418_ | _01419_;
  assign _04020_ = _01421_ | _01422_;
  assign _04021_ = _01424_ | _01425_;
  assign _04022_ = _01398_ | _01369_;
  assign _04023_ = _01427_ | _01428_;
  assign _04024_ = _01430_ | _01431_;
  assign _04025_ = _01433_ | _01434_;
  assign _04026_ = _01436_ | _01437_;
  assign _04027_ = _01439_ | _01440_;
  assign _04028_ = _01427_ | _01442_;
  assign _04029_ = _01443_ | _01444_;
  assign _04030_ = _01446_ | _01447_;
  assign _04031_ = _01449_ | _01450_;
  assign _04032_ = _01452_ | _01453_;
  assign _04702_ = _02681_ | _02682_;
  assign _04703_ = _02684_ | _02685_;
  assign _04704_ = _02687_ | _02688_;
  assign _04705_ = _02690_ | _02691_;
  assign _04706_ = _02693_ | _02694_;
  assign _04707_ = _02696_ | _02697_;
  assign _04708_ = _02699_ | _02700_;
  assign _04709_ = _02702_ | _02703_;
  assign _04710_ = _02705_ | _02706_;
  assign _04711_ = _02708_ | _02709_;
  assign _04712_ = _02711_ | _02712_;
  assign _04713_ = _02714_ | _02715_;
  assign _04714_ = _02717_ | _02718_;
  assign _04715_ = _02720_ | _02721_;
  assign _04716_ = _02723_ | _02724_;
  assign _04717_ = _02726_ | _02727_;
  assign _04718_ = _02729_ | _02730_;
  assign _04719_ = _02732_ | _02733_;
  assign _04720_ = _02735_ | _02736_;
  assign _04721_ = _02738_ | _02739_;
  assign _04722_ = _02741_ | _02742_;
  assign _04723_ = _02744_ | _02745_;
  assign _04724_ = _02747_ | _02748_;
  assign _04725_ = _02750_ | _02751_;
  assign _04726_ = _02753_ | _02754_;
  assign _04727_ = _02756_ | _02757_;
  assign _04728_ = _02759_ | _02760_;
  assign _04729_ = _02762_ | _02763_;
  assign _04730_ = _02765_ | _02766_;
  assign _04731_ = _02768_ | _02769_;
  assign _04732_ = _02771_ | _02772_;
  assign _04733_ = _02774_ | _02775_;
  assign _05160_ = _03470_ | _03471_;
  assign _05161_ = _03472_ | _03473_;
  assign _03361_ = _03985_ | _01335_;
  assign _03363_ = _03986_ | _01338_;
  assign _03365_ = _03987_ | _01341_;
  assign _03367_ = _03988_ | _01344_;
  assign _03369_ = _03989_ | _01335_;
  assign _03371_ = _03990_ | _01348_;
  assign _03373_ = _03991_ | _01335_;
  assign _03375_ = _03992_ | _01352_;
  assign _03377_ = _03993_ | _01335_;
  assign _03379_ = _03994_ | _01355_;
  assign _03381_ = _03995_ | _01341_;
  assign _03383_ = _03996_ | _01359_;
  assign _03385_ = _03997_ | _01362_;
  assign _03387_ = _03998_ | _01365_;
  assign _03389_ = _03999_ | _01368_;
  assign _03391_ = _04000_ | _01338_;
  assign _03393_ = _04001_ | _01372_;
  assign _03395_ = _04002_ | _01375_;
  assign _03397_ = _04003_ | _01378_;
  assign _03399_ = _04004_ | _01381_;
  assign _03401_ = _04005_ | _01384_;
  assign _03403_ = _04006_ | _01372_;
  assign _03405_ = _04007_ | _01388_;
  assign _03407_ = _04008_ | _01391_;
  assign _03409_ = _04009_ | _01394_;
  assign _03411_ = _04010_ | _01397_;
  assign _03413_ = _04011_ | _01338_;
  assign _03415_ = _04012_ | _01401_;
  assign _03417_ = _04013_ | _01404_;
  assign _03419_ = _04014_ | _01407_;
  assign _03421_ = _04015_ | _01410_;
  assign _03423_ = _04016_ | _01413_;
  assign _03425_ = _04017_ | _01401_;
  assign _03427_ = _04018_ | _01417_;
  assign _03429_ = _04019_ | _01420_;
  assign _03431_ = _04020_ | _01423_;
  assign _03433_ = _04021_ | _01426_;
  assign _03435_ = _04022_ | _01338_;
  assign _03437_ = _04023_ | _01429_;
  assign _03439_ = _04024_ | _01432_;
  assign _03441_ = _04025_ | _01435_;
  assign _03443_ = _04026_ | _01438_;
  assign _03445_ = _04027_ | _01441_;
  assign _03447_ = _04028_ | _01429_;
  assign _03449_ = _04029_ | _01445_;
  assign _03451_ = _04030_ | _01448_;
  assign _03453_ = _04031_ | _01451_;
  assign _03455_ = _04032_ | _01454_;
  assign _07022_ = _04702_ | _02683_;
  assign _07024_ = _04703_ | _02686_;
  assign _07026_ = _04704_ | _02689_;
  assign _07028_ = _04705_ | _02692_;
  assign _07030_ = _04706_ | _02695_;
  assign _07032_ = _04707_ | _02698_;
  assign _07034_ = _04708_ | _02701_;
  assign _07036_ = _04709_ | _02704_;
  assign _07038_ = _04710_ | _02707_;
  assign _07040_ = _04711_ | _02710_;
  assign _07042_ = _04712_ | _02713_;
  assign _07044_ = _04713_ | _02716_;
  assign _07046_ = _04714_ | _02719_;
  assign _07048_ = _04715_ | _02722_;
  assign _07050_ = _04716_ | _02725_;
  assign _07052_ = _04717_ | _02728_;
  assign _07054_ = _04718_ | _02731_;
  assign _07056_ = _04719_ | _02734_;
  assign _07058_ = _04720_ | _02737_;
  assign _07060_ = _04721_ | _02740_;
  assign _07062_ = _04722_ | _02743_;
  assign _07064_ = _04723_ | _02746_;
  assign _07066_ = _04724_ | _02749_;
  assign _07068_ = _04725_ | _02752_;
  assign _07070_ = _04726_ | _02755_;
  assign _07072_ = _04727_ | _02758_;
  assign _07074_ = _04728_ | _02761_;
  assign _07076_ = _04729_ | _02764_;
  assign _07078_ = _04730_ | _02767_;
  assign _07080_ = _04731_ | _02770_;
  assign _07082_ = _04732_ | _02773_;
  assign _07084_ = _04733_ | _02776_;
  assign _00109_ = _05160_ | _02782_;
  assign _00113_ = _05161_ | _03474_;
  reg [23:0] _08119_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME _08119_ */
  always_ff @(posedge clk)
    _08119_ <= { dbg_insn_opcode_t0[31:25], dbg_insn_opcode_t0[19:15], dbg_insn_opcode_t0[11:0] };
  assign { rvfi_insn_t0[31:25], rvfi_insn_t0[19:15], rvfi_insn_t0[11:0] } = _08119_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_valid_t0 */
  always_ff @(posedge clk)
    rvfi_valid_t0 <= _00031_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_halt_t0 */
  always_ff @(posedge clk)
    rvfi_halt_t0 <= trap_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_pc_rdata_t0 */
  always_ff @(posedge clk)
    rvfi_pc_rdata_t0 <= rvfi_pc_wdata_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME reg_out_t0 */
  always_ff @(posedge clk)
    reg_out_t0 <= _00027_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME reg_sh_t0 */
  always_ff @(posedge clk)
    reg_sh_t0 <= _00029_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoder_trigger_t0 */
  always_ff @(posedge clk)
    decoder_trigger_t0 <= _00013_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoder_trigger_q_t0 */
  always_ff @(posedge clk)
    decoder_trigger_q_t0 <= decoder_trigger_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoder_pseudo_trigger_q_t0 */
  always_ff @(posedge clk)
    decoder_pseudo_trigger_q_t0 <= decoder_pseudo_trigger_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_rs1val_t0 */
  always_ff @(posedge clk)
    dbg_rs1val_t0 <= _00007_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_rs2val_t0 */
  always_ff @(posedge clk)
    dbg_rs2val_t0 <= _00010_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME alu_out_q_t0 */
  always_ff @(posedge clk)
    alu_out_q_t0 <= alu_out_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME clear_prefetched_high_word_q_t0 */
  always_ff @(posedge clk)
    clear_prefetched_high_word_q_t0 <= clear_prefetched_high_word_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_lui_auipc_jal_t0 */
  always_ff @(posedge clk)
    is_lui_auipc_jal_t0 <= _00015_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_slti_blt_slt_t0 */
  always_ff @(posedge clk)
    is_slti_blt_slt_t0 <= _00017_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_sltiu_bltu_sltu_t0 */
  always_ff @(posedge clk)
    is_sltiu_bltu_sltu_t0 <= _00019_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME q_insn_rs1_t0 */
  always_ff @(posedge clk)
    q_insn_rs1_t0 <= dbg_insn_rs1_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME q_insn_rs2_t0 */
  always_ff @(posedge clk)
    q_insn_rs2_t0 <= dbg_insn_rs2_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_next_t0 */
  always_ff @(posedge clk)
    dbg_next_t0 <= launch_next_insn_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME _00081_ */
  always_ff @(posedge clk)
    _00081_ <= _06103_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME _00083_ */
  always_ff @(posedge clk)
    _00083_ <= _06105_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_rdata_q_t0[31:7] */
  always_ff @(posedge clk)
    mem_rdata_q_t0[31:7] <= _00021_[31:7];
  assign _05434_ = _06703_ ^ instr_lw;
  assign _05435_ = _06701_ ^ instr_lh;
  assign _05436_ = _06699_ ^ instr_lb;
  assign _05443_ = _07409_ ^ instr_jalr;
  assign _05444_ = _07417_ ^ instr_jal;
  assign _05445_ = _06541_ ^ instr_auipc;
  assign _05446_ = _07427_ ^ instr_lui;
  assign _05447_ = mem_rdata_q ^ pcpi_insn;
  assign _05449_ = _06138_ ^ latched_rd;
  assign _05452_ = compressed_instr ^ latched_compr;
  assign _05461_ = _06224_ ^ pcpi_rs2;
  assign _05462_ = _06234_[31] ^ pcpi_rs1[31];
  assign _05463_ = _06234_[30:0] ^ pcpi_rs1[30:0];
  assign _05465_ = _06220_ ^ mem_wordsize;
  assign _05470_ = { dbg_insn_opcode[24:20], dbg_insn_opcode[14:12] } ^ { rvfi_insn[24:20], rvfi_insn[14:12] };
  assign _05475_ = next_pc[31:1] ^ rvfi_pc_wdata[31:1];
  assign _05476_ = _00002_ ^ \cpuregs[9] ;
  assign _05477_ = _00002_ ^ \cpuregs[8] ;
  assign _05478_ = _00002_ ^ \cpuregs[7] ;
  assign _05479_ = _00002_ ^ \cpuregs[6] ;
  assign _05480_ = _00002_ ^ \cpuregs[5] ;
  assign _05481_ = _00002_ ^ \cpuregs[4] ;
  assign _05482_ = _00002_ ^ \cpuregs[3] ;
  assign _05483_ = _00002_ ^ \cpuregs[31] ;
  assign _05484_ = _00002_ ^ \cpuregs[30] ;
  assign _05485_ = _00002_ ^ \cpuregs[2] ;
  assign _05486_ = _00002_ ^ \cpuregs[29] ;
  assign _05487_ = _00002_ ^ \cpuregs[28] ;
  assign _05488_ = _00002_ ^ \cpuregs[27] ;
  assign _05489_ = _00002_ ^ \cpuregs[26] ;
  assign _05490_ = _00002_ ^ \cpuregs[25] ;
  assign _05491_ = _00002_ ^ \cpuregs[24] ;
  assign _05492_ = _00002_ ^ \cpuregs[23] ;
  assign _05493_ = _00002_ ^ \cpuregs[22] ;
  assign _05494_ = _00002_ ^ \cpuregs[21] ;
  assign _05495_ = _00002_ ^ \cpuregs[20] ;
  assign _05496_ = _00002_ ^ \cpuregs[1] ;
  assign _05497_ = _00002_ ^ \cpuregs[19] ;
  assign _05498_ = _00002_ ^ \cpuregs[18] ;
  assign _05499_ = _00002_ ^ \cpuregs[17] ;
  assign _05500_ = _00002_ ^ \cpuregs[16] ;
  assign _05501_ = _00002_ ^ \cpuregs[15] ;
  assign _05502_ = _00002_ ^ \cpuregs[14] ;
  assign _05503_ = _00002_ ^ \cpuregs[13] ;
  assign _05504_ = _00002_ ^ \cpuregs[12] ;
  assign _05505_ = _00002_ ^ \cpuregs[11] ;
  assign _05506_ = _00002_ ^ \cpuregs[10] ;
  assign _05507_ = _00002_ ^ \cpuregs[0] ;
  assign _05905_ = mem_rdata_latched[6:0] ^ mem_rdata_q[6:0];
  assign _05906_ = mem_rdata_latched ^ next_insn_opcode;
  assign _05907_ = _07437_ ^ mem_16bit_buffer;
  assign _05910_ = _00022_ ^ mem_state;
  assign _05911_ = _07456_ ^ mem_wstrb;
  assign _05913_ = mem_la_addr ^ mem_addr;
  assign _05818_ = _00062_ ^ cached_insn_opcode;
  assign _05914_ = _00024_ ^ mem_valid;
  assign _05816_ = decoded_rs2 ^ cached_insn_rs2;
  assign _05817_ = decoded_rs1 ^ cached_insn_rs1;
  assign _05915_ = _07324_ ^ is_alu_reg_reg;
  assign _05916_ = _07340_ ^ is_alu_reg_imm;
  assign _05918_ = _06897_ ^ instr_ecall_ebreak;
  assign _05920_ = _06817_ ^ is_sll_srl_sra;
  assign _05921_ = _07352_ ^ is_sb_sh_sw;
  assign _05922_ = _06899_ ^ is_jalr_addi_slti_sltiu_xori_ori_andi;
  assign _05923_ = _06813_ ^ is_slli_srli_srai;
  assign _05924_ = _07360_ ^ is_lb_lh_lw_lbu_lhu;
  assign _05925_ = _07362_ ^ compressed_instr;
  assign _05926_ = _07276_ ^ decoded_imm_j[10];
  assign _05927_ = _07278_ ^ decoded_imm_j[7];
  assign _05928_ = _07280_ ^ decoded_imm_j[6];
  assign _05929_ = _07282_ ^ decoded_imm_j[3:1];
  assign _05930_ = _07284_ ^ decoded_imm_j[5];
  assign _05931_ = _07286_ ^ decoded_imm_j[9:8];
  assign _05932_ = _07288_ ^ decoded_imm_j[31:20];
  assign _05933_ = _07290_ ^ decoded_imm_j[4];
  assign _05934_ = _07292_ ^ decoded_imm_j[11];
  assign _05935_ = _07378_ ^ decoded_imm_j[19:12];
  assign _05936_ = _06333_ ^ decoded_imm;
  assign _05508_ = _07376_ ^ decoded_rs2;
  assign _05938_ = mem_la_wdata ^ mem_wdata;
  assign _05939_ = _07274_ ^ decoded_rs1[4];
  assign _05940_ = _07312_ ^ decoded_rs1[3:0];
  assign _05941_ = _07399_ ^ decoded_rd;
  assign _05942_ = _06799_ ^ instr_rdinstrh;
  assign _05943_ = _06795_ ^ instr_rdinstr;
  assign _05944_ = _06791_ ^ instr_rdcycleh;
  assign _05945_ = _06781_ ^ instr_rdcycle;
  assign _05955_ = _06735_ ^ instr_srai;
  assign _05956_ = _06733_ ^ instr_srli;
  assign _05957_ = _06729_ ^ instr_slli;
  assign _05964_ = _06713_ ^ instr_sw;
  assign _05965_ = _06711_ ^ instr_sh;
  assign _05966_ = _06709_ ^ instr_sb;
  assign _05967_ = _06707_ ^ instr_lhu;
  assign _05968_ = _06705_ ^ instr_lbu;
  assign _00132_ = ~ _01045_;
  assign _00133_ = ~ _01049_;
  assign _00134_ = ~ _01057_;
  assign _00135_ = ~ _01059_;
  assign _00136_ = ~ _01061_;
  assign _00137_ = ~ _01063_;
  assign _00138_ = ~ dbg_next;
  assign _00139_ = ~ launch_next_insn;
  assign _00140_ = ~ _07083_;
  assign _00141_ = ~ _07081_;
  assign _00142_ = ~ _07079_;
  assign _00143_ = ~ _07077_;
  assign _00144_ = ~ _07075_;
  assign _00145_ = ~ _07073_;
  assign _00146_ = ~ _07071_;
  assign _00147_ = ~ _07069_;
  assign _00148_ = ~ _07067_;
  assign _00149_ = ~ _07065_;
  assign _00150_ = ~ _07063_;
  assign _00151_ = ~ _07061_;
  assign _00152_ = ~ _07059_;
  assign _00153_ = ~ _07057_;
  assign _00154_ = ~ _07055_;
  assign _00155_ = ~ _07053_;
  assign _00156_ = ~ _07051_;
  assign _00157_ = ~ _07049_;
  assign _00158_ = ~ _07047_;
  assign _00159_ = ~ _07045_;
  assign _00160_ = ~ _07043_;
  assign _00161_ = ~ _07041_;
  assign _00162_ = ~ _07039_;
  assign _00163_ = ~ _07037_;
  assign _00164_ = ~ _07035_;
  assign _00165_ = ~ _07033_;
  assign _00166_ = ~ _07031_;
  assign _00167_ = ~ _07029_;
  assign _00168_ = ~ _07027_;
  assign _00169_ = ~ _07025_;
  assign _00170_ = ~ _07023_;
  assign _00171_ = ~ _07021_;
  assign _00172_ = ~ mem_xfer;
  assign _00173_ = ~ _01029_;
  assign _00174_ = ~ _01035_;
  assign _00175_ = ~ _06888_;
  assign _00176_ = ~ _01039_;
  assign _00178_ = ~ _01041_;
  assign _00177_ = ~ decoder_trigger_q;
  assign _00131_ = ~ _05738_;
  assign _00130_ = ~ _06685_;
  assign _00179_ = ~ _01043_;
  assign _03681_ = _06704_ | instr_lw_t0;
  assign _03685_ = _06702_ | instr_lh_t0;
  assign _03689_ = _06700_ | instr_lb_t0;
  assign _03717_ = _07410_ | instr_jalr_t0;
  assign _03721_ = _07418_ | instr_jal_t0;
  assign _03725_ = _06542_ | instr_auipc_t0;
  assign _03729_ = _07428_ | instr_lui_t0;
  assign _03733_ = mem_rdata_q_t0 | pcpi_insn_t0;
  assign _03741_ = _06139_ | latched_rd_t0;
  assign _03753_ = compressed_instr_t0 | latched_compr_t0;
  assign _03793_ = _06225_ | pcpi_rs2_t0;
  assign _03797_ = _06235_[31] | pcpi_rs1_t0[31];
  assign _03801_ = _06235_[30:0] | pcpi_rs1_t0[30:0];
  assign _03809_ = _06221_ | mem_wordsize_t0;
  assign _03829_ = { dbg_insn_opcode_t0[24:20], dbg_insn_opcode_t0[14:12] } | { rvfi_insn_t0[24:20], rvfi_insn_t0[14:12] };
  assign _03849_ = next_pc_t0[31:1] | rvfi_pc_wdata_t0[31:1];
  assign _03853_ = _00003_ | \cpuregs[9]_t0 ;
  assign _03857_ = _00003_ | \cpuregs[8]_t0 ;
  assign _03861_ = _00003_ | \cpuregs[7]_t0 ;
  assign _03865_ = _00003_ | \cpuregs[6]_t0 ;
  assign _03869_ = _00003_ | \cpuregs[5]_t0 ;
  assign _03873_ = _00003_ | \cpuregs[4]_t0 ;
  assign _03877_ = _00003_ | \cpuregs[3]_t0 ;
  assign _03881_ = _00003_ | \cpuregs[31]_t0 ;
  assign _03885_ = _00003_ | \cpuregs[30]_t0 ;
  assign _03889_ = _00003_ | \cpuregs[2]_t0 ;
  assign _03893_ = _00003_ | \cpuregs[29]_t0 ;
  assign _03897_ = _00003_ | \cpuregs[28]_t0 ;
  assign _03901_ = _00003_ | \cpuregs[27]_t0 ;
  assign _03905_ = _00003_ | \cpuregs[26]_t0 ;
  assign _03909_ = _00003_ | \cpuregs[25]_t0 ;
  assign _03913_ = _00003_ | \cpuregs[24]_t0 ;
  assign _03917_ = _00003_ | \cpuregs[23]_t0 ;
  assign _03921_ = _00003_ | \cpuregs[22]_t0 ;
  assign _03925_ = _00003_ | \cpuregs[21]_t0 ;
  assign _03929_ = _00003_ | \cpuregs[20]_t0 ;
  assign _03933_ = _00003_ | \cpuregs[1]_t0 ;
  assign _03937_ = _00003_ | \cpuregs[19]_t0 ;
  assign _03941_ = _00003_ | \cpuregs[18]_t0 ;
  assign _03945_ = _00003_ | \cpuregs[17]_t0 ;
  assign _03949_ = _00003_ | \cpuregs[16]_t0 ;
  assign _03953_ = _00003_ | \cpuregs[15]_t0 ;
  assign _03957_ = _00003_ | \cpuregs[14]_t0 ;
  assign _03961_ = _00003_ | \cpuregs[13]_t0 ;
  assign _03965_ = _00003_ | \cpuregs[12]_t0 ;
  assign _03969_ = _00003_ | \cpuregs[11]_t0 ;
  assign _03973_ = _00003_ | \cpuregs[10]_t0 ;
  assign _03977_ = _00003_ | \cpuregs[0]_t0 ;
  assign _05162_ = mem_rdata_latched_t0[6:0] | mem_rdata_q_t0[6:0];
  assign _05166_ = mem_rdata_latched_t0 | next_insn_opcode_t0;
  assign _05170_ = _07438_ | mem_16bit_buffer_t0;
  assign _05182_ = _00023_ | mem_state_t0;
  assign _05186_ = _07457_ | mem_wstrb_t0;
  assign _05194_ = mem_la_addr_t0 | mem_addr_t0;
  assign _05198_ = _00063_ | cached_insn_opcode_t0;
  assign _05202_ = _00025_ | mem_valid_t0;
  assign _05206_ = decoded_rs2_t0 | cached_insn_rs2_t0;
  assign _05210_ = decoded_rs1_t0 | cached_insn_rs1_t0;
  assign _05216_ = _07325_ | is_alu_reg_reg_t0;
  assign _05220_ = _07341_ | is_alu_reg_imm_t0;
  assign _05228_ = _06898_ | instr_ecall_ebreak_t0;
  assign _05236_ = _06818_ | is_sll_srl_sra_t0;
  assign _05240_ = _07353_ | is_sb_sh_sw_t0;
  assign _05244_ = _06900_ | is_jalr_addi_slti_sltiu_xori_ori_andi_t0;
  assign _05248_ = _06814_ | is_slli_srli_srai_t0;
  assign _05252_ = _07361_ | is_lb_lh_lw_lbu_lhu_t0;
  assign _05256_ = _06678_ | compressed_instr_t0;
  assign _05260_ = _07277_ | decoded_imm_j_t0[10];
  assign _05264_ = _07279_ | decoded_imm_j_t0[7];
  assign _05268_ = _07281_ | decoded_imm_j_t0[6];
  assign _05272_ = _07283_ | decoded_imm_j_t0[3:1];
  assign _05276_ = _07285_ | decoded_imm_j_t0[5];
  assign _05280_ = _07287_ | decoded_imm_j_t0[9:8];
  assign _05284_ = _07289_ | decoded_imm_j_t0[31:20];
  assign _05288_ = _07291_ | decoded_imm_j_t0[4];
  assign _05292_ = _07293_ | decoded_imm_j_t0[11];
  assign _05296_ = _07379_ | decoded_imm_j_t0[19:12];
  assign _05300_ = _06334_ | decoded_imm_t0;
  assign _05304_ = _07377_ | decoded_rs2_t0;
  assign _05312_ = mem_la_wdata_t0 | mem_wdata_t0;
  assign _05316_ = _07275_ | decoded_rs1_t0[4];
  assign _05320_ = _07313_ | decoded_rs1_t0[3:0];
  assign _05324_ = _07400_ | decoded_rd_t0;
  assign _05328_ = _06800_ | instr_rdinstrh_t0;
  assign _05332_ = _06796_ | instr_rdinstr_t0;
  assign _05336_ = _06792_ | instr_rdcycleh_t0;
  assign _05340_ = _06782_ | instr_rdcycle_t0;
  assign _05380_ = _06736_ | instr_srai_t0;
  assign _05384_ = _06734_ | instr_srli_t0;
  assign _05388_ = _06730_ | instr_slli_t0;
  assign _05416_ = _06714_ | instr_sw_t0;
  assign _05420_ = _06712_ | instr_sh_t0;
  assign _05424_ = _06710_ | instr_sb_t0;
  assign _05428_ = _06708_ | instr_lhu_t0;
  assign _05432_ = _06706_ | instr_lbu_t0;
  assign _03682_ = _05434_ | _03681_;
  assign _03686_ = _05435_ | _03685_;
  assign _03690_ = _05436_ | _03689_;
  assign _03718_ = _05443_ | _03717_;
  assign _03722_ = _05444_ | _03721_;
  assign _03726_ = _05445_ | _03725_;
  assign _03730_ = _05446_ | _03729_;
  assign _03734_ = _05447_ | _03733_;
  assign _03742_ = _05449_ | _03741_;
  assign _03754_ = _05452_ | _03753_;
  assign _03794_ = _05461_ | _03793_;
  assign _03798_ = _05462_ | _03797_;
  assign _03802_ = _05463_ | _03801_;
  assign _03810_ = _05465_ | _03809_;
  assign _03830_ = _05470_ | _03829_;
  assign _03850_ = _05475_ | _03849_;
  assign _03854_ = _05476_ | _03853_;
  assign _03858_ = _05477_ | _03857_;
  assign _03862_ = _05478_ | _03861_;
  assign _03866_ = _05479_ | _03865_;
  assign _03870_ = _05480_ | _03869_;
  assign _03874_ = _05481_ | _03873_;
  assign _03878_ = _05482_ | _03877_;
  assign _03882_ = _05483_ | _03881_;
  assign _03886_ = _05484_ | _03885_;
  assign _03890_ = _05485_ | _03889_;
  assign _03894_ = _05486_ | _03893_;
  assign _03898_ = _05487_ | _03897_;
  assign _03902_ = _05488_ | _03901_;
  assign _03906_ = _05489_ | _03905_;
  assign _03910_ = _05490_ | _03909_;
  assign _03914_ = _05491_ | _03913_;
  assign _03918_ = _05492_ | _03917_;
  assign _03922_ = _05493_ | _03921_;
  assign _03926_ = _05494_ | _03925_;
  assign _03930_ = _05495_ | _03929_;
  assign _03934_ = _05496_ | _03933_;
  assign _03938_ = _05497_ | _03937_;
  assign _03942_ = _05498_ | _03941_;
  assign _03946_ = _05499_ | _03945_;
  assign _03950_ = _05500_ | _03949_;
  assign _03954_ = _05501_ | _03953_;
  assign _03958_ = _05502_ | _03957_;
  assign _03962_ = _05503_ | _03961_;
  assign _03966_ = _05504_ | _03965_;
  assign _03970_ = _05505_ | _03969_;
  assign _03974_ = _05506_ | _03973_;
  assign _03978_ = _05507_ | _03977_;
  assign _05163_ = _05905_ | _05162_;
  assign _05167_ = _05906_ | _05166_;
  assign _05171_ = _05907_ | _05170_;
  assign _05183_ = _05910_ | _05182_;
  assign _05187_ = _05911_ | _05186_;
  assign _05195_ = _05913_ | _05194_;
  assign _05199_ = _05818_ | _05198_;
  assign _05203_ = _05914_ | _05202_;
  assign _05207_ = _05816_ | _05206_;
  assign _05211_ = _05817_ | _05210_;
  assign _05217_ = _05915_ | _05216_;
  assign _05221_ = _05916_ | _05220_;
  assign _05229_ = _05918_ | _05228_;
  assign _05237_ = _05920_ | _05236_;
  assign _05241_ = _05921_ | _05240_;
  assign _05245_ = _05922_ | _05244_;
  assign _05249_ = _05923_ | _05248_;
  assign _05253_ = _05924_ | _05252_;
  assign _05257_ = _05925_ | _05256_;
  assign _05261_ = _05926_ | _05260_;
  assign _05265_ = _05927_ | _05264_;
  assign _05269_ = _05928_ | _05268_;
  assign _05273_ = _05929_ | _05272_;
  assign _05277_ = _05930_ | _05276_;
  assign _05281_ = _05931_ | _05280_;
  assign _05285_ = _05932_ | _05284_;
  assign _05289_ = _05933_ | _05288_;
  assign _05293_ = _05934_ | _05292_;
  assign _05297_ = _05935_ | _05296_;
  assign _05301_ = _05936_ | _05300_;
  assign _05305_ = _05508_ | _05304_;
  assign _05313_ = _05938_ | _05312_;
  assign _05317_ = _05939_ | _05316_;
  assign _05321_ = _05940_ | _05320_;
  assign _05325_ = _05941_ | _05324_;
  assign _05329_ = _05942_ | _05328_;
  assign _05333_ = _05943_ | _05332_;
  assign _05337_ = _05944_ | _05336_;
  assign _05341_ = _05945_ | _05340_;
  assign _05381_ = _05955_ | _05380_;
  assign _05385_ = _05956_ | _05384_;
  assign _05389_ = _05957_ | _05388_;
  assign _05417_ = _05964_ | _05416_;
  assign _05421_ = _05965_ | _05420_;
  assign _05425_ = _05966_ | _05424_;
  assign _05429_ = _05967_ | _05428_;
  assign _05433_ = _05968_ | _05432_;
  assign _01101_ = _06685_ & _06704_;
  assign _01104_ = _06685_ & _06702_;
  assign _01107_ = _06685_ & _06700_;
  assign _01128_ = _05738_ & _07410_;
  assign _01131_ = _05738_ & _07418_;
  assign _01134_ = _05738_ & _06542_;
  assign _01137_ = _05738_ & _07428_;
  assign _01140_ = { _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_ } & mem_rdata_q_t0;
  assign _01146_ = { _01045_, _01045_, _01045_, _01045_, _01045_ } & _06139_;
  assign _01155_ = _01049_ & compressed_instr_t0;
  assign _01186_ = { _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_, _01057_ } & _06225_;
  assign _01189_ = _01059_ & _06235_[31];
  assign _01192_ = { _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_, _01061_ } & _06235_[30:0];
  assign _01198_ = { _01063_, _01063_ } & _06221_;
  assign _01213_ = { dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next } & { dbg_insn_opcode_t0[24:20], dbg_insn_opcode_t0[14:12] };
  assign _01228_ = { launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn } & next_pc_t0[31:1];
  assign _01231_ = { _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_, _07083_ } & _00003_;
  assign _01234_ = { _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_, _07081_ } & _00003_;
  assign _01237_ = { _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_, _07079_ } & _00003_;
  assign _01240_ = { _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_, _07077_ } & _00003_;
  assign _01243_ = { _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_, _07075_ } & _00003_;
  assign _01246_ = { _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_, _07073_ } & _00003_;
  assign _01249_ = { _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_, _07071_ } & _00003_;
  assign _01252_ = { _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_, _07069_ } & _00003_;
  assign _01255_ = { _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_, _07067_ } & _00003_;
  assign _01258_ = { _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_, _07065_ } & _00003_;
  assign _01261_ = { _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_, _07063_ } & _00003_;
  assign _01264_ = { _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_, _07061_ } & _00003_;
  assign _01267_ = { _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_, _07059_ } & _00003_;
  assign _01270_ = { _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_, _07057_ } & _00003_;
  assign _01273_ = { _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_, _07055_ } & _00003_;
  assign _01276_ = { _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_, _07053_ } & _00003_;
  assign _01279_ = { _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_, _07051_ } & _00003_;
  assign _01282_ = { _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_, _07049_ } & _00003_;
  assign _01285_ = { _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_, _07047_ } & _00003_;
  assign _01288_ = { _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_, _07045_ } & _00003_;
  assign _01291_ = { _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_, _07043_ } & _00003_;
  assign _01294_ = { _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_, _07041_ } & _00003_;
  assign _01297_ = { _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_, _07039_ } & _00003_;
  assign _01300_ = { _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_, _07037_ } & _00003_;
  assign _01303_ = { _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_, _07035_ } & _00003_;
  assign _01306_ = { _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_, _07033_ } & _00003_;
  assign _01309_ = { _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_, _07031_ } & _00003_;
  assign _01312_ = { _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_, _07029_ } & _00003_;
  assign _01315_ = { _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_, _07027_ } & _00003_;
  assign _01318_ = { _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_, _07025_ } & _00003_;
  assign _01321_ = { _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_, _07023_ } & _00003_;
  assign _01324_ = { _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_, _07021_ } & _00003_;
  assign _03475_ = { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer } & mem_rdata_latched_t0[6:0];
  assign _03478_ = { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer } & mem_rdata_latched_t0;
  assign _03481_ = { _01029_, _01029_, _01029_, _01029_, _01029_, _01029_, _01029_, _01029_, _01029_, _01029_, _01029_, _01029_, _01029_, _01029_, _01029_, _01029_ } & _07438_;
  assign _03490_ = { _01035_, _01035_ } & _00023_;
  assign _03493_ = { _00175_, _00175_, _00175_, _00175_ } & _07457_;
  assign _03499_ = { _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_, _01039_ } & mem_la_addr_t0;
  assign _03502_ = { decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q } & _00063_;
  assign _03505_ = _01041_ & _00025_;
  assign _03508_ = { decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q } & decoded_rs2_t0;
  assign _03511_ = { decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q } & decoded_rs1_t0;
  assign _03516_ = _05738_ & _07325_;
  assign _03519_ = _05738_ & _07341_;
  assign _03525_ = _06685_ & _06898_;
  assign _03531_ = _06685_ & _06818_;
  assign _03534_ = _05738_ & _07353_;
  assign _03537_ = _06685_ & _06900_;
  assign _03540_ = _06685_ & _06814_;
  assign _03543_ = _05738_ & _07361_;
  assign _03546_ = _05738_ & _06678_;
  assign _03549_ = _05738_ & _07277_;
  assign _03552_ = _05738_ & _07279_;
  assign _03555_ = _05738_ & _07281_;
  assign _03558_ = { _05738_, _05738_, _05738_ } & _07283_;
  assign _03561_ = _05738_ & _07285_;
  assign _03564_ = { _05738_, _05738_ } & _07287_;
  assign _03567_ = { _05738_, _05738_, _05738_, _05738_, _05738_, _05738_, _05738_, _05738_, _05738_, _05738_, _05738_, _05738_ } & _07289_;
  assign _03570_ = _05738_ & _07291_;
  assign _03573_ = _05738_ & _07293_;
  assign _03576_ = { _05738_, _05738_, _05738_, _05738_, _05738_, _05738_, _05738_, _05738_ } & _07379_;
  assign _03579_ = { _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_, _06685_ } & _06334_;
  assign _03582_ = { _05738_, _05738_, _05738_, _05738_, _05738_ } & _07377_;
  assign _03588_ = { _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_, _01043_ } & mem_la_wdata_t0;
  assign _03591_ = _05738_ & _07275_;
  assign _03594_ = { _05738_, _05738_, _05738_, _05738_ } & _07313_;
  assign _03597_ = { _05738_, _05738_, _05738_, _05738_, _05738_ } & _07400_;
  assign _03600_ = _06685_ & _06800_;
  assign _03603_ = _06685_ & _06796_;
  assign _03606_ = _06685_ & _06792_;
  assign _03609_ = _06685_ & _06782_;
  assign _03639_ = _06685_ & _06736_;
  assign _03642_ = _06685_ & _06734_;
  assign _03645_ = _06685_ & _06730_;
  assign _03666_ = _06685_ & _06714_;
  assign _03669_ = _06685_ & _06712_;
  assign _03672_ = _06685_ & _06710_;
  assign _03675_ = _06685_ & _06708_;
  assign _03678_ = _06685_ & _06706_;
  assign _01099_ = _00130_ & instr_lbu_t0;
  assign _01102_ = _00130_ & instr_lw_t0;
  assign _01105_ = _00130_ & instr_lh_t0;
  assign _01108_ = _00130_ & instr_lb_t0;
  assign _01129_ = _00131_ & instr_jalr_t0;
  assign _01132_ = _00131_ & instr_jal_t0;
  assign _01135_ = _00131_ & instr_auipc_t0;
  assign _01138_ = _00131_ & instr_lui_t0;
  assign _01141_ = { _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_ } & pcpi_insn_t0;
  assign _01147_ = { _00132_, _00132_, _00132_, _00132_, _00132_ } & latched_rd_t0;
  assign _01156_ = _00133_ & latched_compr_t0;
  assign _01187_ = { _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_, _00134_ } & pcpi_rs2_t0;
  assign _01190_ = _00135_ & pcpi_rs1_t0[31];
  assign _01193_ = { _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_, _00136_ } & pcpi_rs1_t0[30:0];
  assign _01199_ = { _00137_, _00137_ } & mem_wordsize_t0;
  assign _01214_ = { _00138_, _00138_, _00138_, _00138_, _00138_, _00138_, _00138_, _00138_ } & { rvfi_insn_t0[24:20], rvfi_insn_t0[14:12] };
  assign _01229_ = { _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_, _00139_ } & rvfi_pc_wdata_t0[31:1];
  assign _01232_ = { _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_, _00140_ } & \cpuregs[9]_t0 ;
  assign _01235_ = { _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_, _00141_ } & \cpuregs[8]_t0 ;
  assign _01238_ = { _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_, _00142_ } & \cpuregs[7]_t0 ;
  assign _01241_ = { _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_, _00143_ } & \cpuregs[6]_t0 ;
  assign _01244_ = { _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_, _00144_ } & \cpuregs[5]_t0 ;
  assign _01247_ = { _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_, _00145_ } & \cpuregs[4]_t0 ;
  assign _01250_ = { _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_, _00146_ } & \cpuregs[3]_t0 ;
  assign _01253_ = { _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_, _00147_ } & \cpuregs[31]_t0 ;
  assign _01256_ = { _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_, _00148_ } & \cpuregs[30]_t0 ;
  assign _01259_ = { _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_, _00149_ } & \cpuregs[2]_t0 ;
  assign _01262_ = { _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_, _00150_ } & \cpuregs[29]_t0 ;
  assign _01265_ = { _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_, _00151_ } & \cpuregs[28]_t0 ;
  assign _01268_ = { _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_, _00152_ } & \cpuregs[27]_t0 ;
  assign _01271_ = { _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_, _00153_ } & \cpuregs[26]_t0 ;
  assign _01274_ = { _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_, _00154_ } & \cpuregs[25]_t0 ;
  assign _01277_ = { _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_, _00155_ } & \cpuregs[24]_t0 ;
  assign _01280_ = { _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_, _00156_ } & \cpuregs[23]_t0 ;
  assign _01283_ = { _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_, _00157_ } & \cpuregs[22]_t0 ;
  assign _01286_ = { _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_, _00158_ } & \cpuregs[21]_t0 ;
  assign _01289_ = { _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_, _00159_ } & \cpuregs[20]_t0 ;
  assign _01292_ = { _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_, _00160_ } & \cpuregs[1]_t0 ;
  assign _01295_ = { _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_, _00161_ } & \cpuregs[19]_t0 ;
  assign _01298_ = { _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_, _00162_ } & \cpuregs[18]_t0 ;
  assign _01301_ = { _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_, _00163_ } & \cpuregs[17]_t0 ;
  assign _01304_ = { _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_, _00164_ } & \cpuregs[16]_t0 ;
  assign _01307_ = { _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_, _00165_ } & \cpuregs[15]_t0 ;
  assign _01310_ = { _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_, _00166_ } & \cpuregs[14]_t0 ;
  assign _01313_ = { _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_, _00167_ } & \cpuregs[13]_t0 ;
  assign _01316_ = { _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_, _00168_ } & \cpuregs[12]_t0 ;
  assign _01319_ = { _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_, _00169_ } & \cpuregs[11]_t0 ;
  assign _01322_ = { _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_, _00170_ } & \cpuregs[10]_t0 ;
  assign _01325_ = { _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_, _00171_ } & \cpuregs[0]_t0 ;
  assign _03476_ = { _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_ } & mem_rdata_q_t0[6:0];
  assign _03479_ = { _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_, _00172_ } & next_insn_opcode_t0;
  assign _03482_ = { _00173_, _00173_, _00173_, _00173_, _00173_, _00173_, _00173_, _00173_, _00173_, _00173_, _00173_, _00173_, _00173_, _00173_, _00173_, _00173_ } & mem_16bit_buffer_t0;
  assign _03491_ = { _00174_, _00174_ } & mem_state_t0;
  assign _03494_ = { _06888_, _06888_, _06888_, _06888_ } & mem_wstrb_t0;
  assign _03500_ = { _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_, _00176_ } & mem_addr_t0;
  assign _03503_ = { _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_, _00177_ } & cached_insn_opcode_t0;
  assign _03506_ = _00178_ & mem_valid_t0;
  assign _03509_ = { _00177_, _00177_, _00177_, _00177_, _00177_ } & cached_insn_rs2_t0;
  assign _03512_ = { _00177_, _00177_, _00177_, _00177_, _00177_ } & cached_insn_rs1_t0;
  assign _03517_ = _00131_ & is_alu_reg_reg_t0;
  assign _03520_ = _00131_ & is_alu_reg_imm_t0;
  assign _03526_ = _00130_ & instr_ecall_ebreak_t0;
  assign _03532_ = _00130_ & is_sll_srl_sra_t0;
  assign _03535_ = _00131_ & is_sb_sh_sw_t0;
  assign _03538_ = _00130_ & is_jalr_addi_slti_sltiu_xori_ori_andi_t0;
  assign _03541_ = _00130_ & is_slli_srli_srai_t0;
  assign _03544_ = _00131_ & is_lb_lh_lw_lbu_lhu_t0;
  assign _03547_ = _00131_ & compressed_instr_t0;
  assign _03550_ = _00131_ & decoded_imm_j_t0[10];
  assign _03553_ = _00131_ & decoded_imm_j_t0[7];
  assign _03556_ = _00131_ & decoded_imm_j_t0[6];
  assign _03559_ = { _00131_, _00131_, _00131_ } & decoded_imm_j_t0[3:1];
  assign _03562_ = _00131_ & decoded_imm_j_t0[5];
  assign _03565_ = { _00131_, _00131_ } & decoded_imm_j_t0[9:8];
  assign _03568_ = { _00131_, _00131_, _00131_, _00131_, _00131_, _00131_, _00131_, _00131_, _00131_, _00131_, _00131_, _00131_ } & decoded_imm_j_t0[31:20];
  assign _03571_ = _00131_ & decoded_imm_j_t0[4];
  assign _03574_ = _00131_ & decoded_imm_j_t0[11];
  assign _03577_ = { _00131_, _00131_, _00131_, _00131_, _00131_, _00131_, _00131_, _00131_ } & decoded_imm_j_t0[19:12];
  assign _03580_ = { _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_, _00130_ } & decoded_imm_t0;
  assign _03583_ = { _00131_, _00131_, _00131_, _00131_, _00131_ } & decoded_rs2_t0;
  assign _03589_ = { _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_, _00179_ } & mem_wdata_t0;
  assign _03592_ = _00131_ & decoded_rs1_t0[4];
  assign _03595_ = { _00131_, _00131_, _00131_, _00131_ } & decoded_rs1_t0[3:0];
  assign _03598_ = { _00131_, _00131_, _00131_, _00131_, _00131_ } & decoded_rd_t0;
  assign _03601_ = _00130_ & instr_rdinstrh_t0;
  assign _03604_ = _00130_ & instr_rdinstr_t0;
  assign _03607_ = _00130_ & instr_rdcycleh_t0;
  assign _03610_ = _00130_ & instr_rdcycle_t0;
  assign _03640_ = _00130_ & instr_srai_t0;
  assign _03643_ = _00130_ & instr_srli_t0;
  assign _03646_ = _00130_ & instr_slli_t0;
  assign _03667_ = _00130_ & instr_sw_t0;
  assign _03670_ = _00130_ & instr_sh_t0;
  assign _03673_ = _00130_ & instr_sb_t0;
  assign _03676_ = _00130_ & instr_lhu_t0;
  assign _01100_ = _05433_ & _06686_;
  assign _01103_ = _03682_ & _06686_;
  assign _01106_ = _03686_ & _06686_;
  assign _01109_ = _03690_ & _06686_;
  assign _01130_ = _03718_ & _06608_;
  assign _01133_ = _03722_ & _06608_;
  assign _01136_ = _03726_ & _06608_;
  assign _01139_ = _03730_ & _06608_;
  assign _01142_ = _03734_ & { _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_ };
  assign _01148_ = _03742_ & { _01046_, _01046_, _01046_, _01046_, _01046_ };
  assign _01157_ = _03754_ & _01050_;
  assign _01188_ = _03794_ & { _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_, _01058_ };
  assign _01191_ = _03798_ & _01060_;
  assign _01194_ = _03802_ & { _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_, _01062_ };
  assign _01200_ = _03810_ & { _01064_, _01064_ };
  assign _01215_ = _03830_ & { dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0 };
  assign _01230_ = _03850_ & { launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0 };
  assign _01233_ = _03854_ & { _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_, _07084_ };
  assign _01236_ = _03858_ & { _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_, _07082_ };
  assign _01239_ = _03862_ & { _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_, _07080_ };
  assign _01242_ = _03866_ & { _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_, _07078_ };
  assign _01245_ = _03870_ & { _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_, _07076_ };
  assign _01248_ = _03874_ & { _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_, _07074_ };
  assign _01251_ = _03878_ & { _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_, _07072_ };
  assign _01254_ = _03882_ & { _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_, _07070_ };
  assign _01257_ = _03886_ & { _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_, _07068_ };
  assign _01260_ = _03890_ & { _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_, _07066_ };
  assign _01263_ = _03894_ & { _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_, _07064_ };
  assign _01266_ = _03898_ & { _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_, _07062_ };
  assign _01269_ = _03902_ & { _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_, _07060_ };
  assign _01272_ = _03906_ & { _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_, _07058_ };
  assign _01275_ = _03910_ & { _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_, _07056_ };
  assign _01278_ = _03914_ & { _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_, _07054_ };
  assign _01281_ = _03918_ & { _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_, _07052_ };
  assign _01284_ = _03922_ & { _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_, _07050_ };
  assign _01287_ = _03926_ & { _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_, _07048_ };
  assign _01290_ = _03930_ & { _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_, _07046_ };
  assign _01293_ = _03934_ & { _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_, _07044_ };
  assign _01296_ = _03938_ & { _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_, _07042_ };
  assign _01299_ = _03942_ & { _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_, _07040_ };
  assign _01302_ = _03946_ & { _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_, _07038_ };
  assign _01305_ = _03950_ & { _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_, _07036_ };
  assign _01308_ = _03954_ & { _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_, _07034_ };
  assign _01311_ = _03958_ & { _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_, _07032_ };
  assign _01314_ = _03962_ & { _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_, _07030_ };
  assign _01317_ = _03966_ & { _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_, _07028_ };
  assign _01320_ = _03970_ & { _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_, _07026_ };
  assign _01323_ = _03974_ & { _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_, _07024_ };
  assign _01326_ = _03978_ & { _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_, _07022_ };
  assign _03477_ = _05163_ & { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 };
  assign _03480_ = _05167_ & { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 };
  assign _03483_ = _05171_ & { _01030_, _01030_, _01030_, _01030_, _01030_, _01030_, _01030_, _01030_, _01030_, _01030_, _01030_, _01030_, _01030_, _01030_, _01030_, _01030_ };
  assign _03492_ = _05183_ & { _01036_, _01036_ };
  assign _03495_ = _05187_ & { _00797_, _00797_, _00797_, _00797_ };
  assign _03501_ = _05195_ & { _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_, _01040_ };
  assign _03504_ = _05199_ & { decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0 };
  assign _03507_ = _05203_ & _01042_;
  assign _03510_ = _05207_ & { decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0 };
  assign _03513_ = _05211_ & { decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0, decoder_trigger_q_t0 };
  assign _03518_ = _05217_ & _06608_;
  assign _03521_ = _05221_ & _06608_;
  assign _03527_ = _05229_ & _06686_;
  assign _03533_ = _05237_ & _06686_;
  assign _03536_ = _05241_ & _06608_;
  assign _03539_ = _05245_ & _06686_;
  assign _03542_ = _05249_ & _06686_;
  assign _03545_ = _05253_ & _06608_;
  assign _03548_ = _05257_ & _06608_;
  assign _03551_ = _05261_ & _06608_;
  assign _03554_ = _05265_ & _06608_;
  assign _03557_ = _05269_ & _06608_;
  assign _03560_ = _05273_ & { _06608_, _06608_, _06608_ };
  assign _03563_ = _05277_ & _06608_;
  assign _03566_ = _05281_ & { _06608_, _06608_ };
  assign _03569_ = _05285_ & { _06608_, _06608_, _06608_, _06608_, _06608_, _06608_, _06608_, _06608_, _06608_, _06608_, _06608_, _06608_ };
  assign _03572_ = _05289_ & _06608_;
  assign _03575_ = _05293_ & _06608_;
  assign _03578_ = _05297_ & { _06608_, _06608_, _06608_, _06608_, _06608_, _06608_, _06608_, _06608_ };
  assign _03581_ = _05301_ & { _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_, _06686_ };
  assign _03584_ = _05305_ & { _06608_, _06608_, _06608_, _06608_, _06608_ };
  assign _03590_ = _05313_ & { _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_, _01044_ };
  assign _03593_ = _05317_ & _06608_;
  assign _03596_ = _05321_ & { _06608_, _06608_, _06608_, _06608_ };
  assign _03599_ = _05325_ & { _06608_, _06608_, _06608_, _06608_, _06608_ };
  assign _03602_ = _05329_ & _06686_;
  assign _03605_ = _05333_ & _06686_;
  assign _03608_ = _05337_ & _06686_;
  assign _03611_ = _05341_ & _06686_;
  assign _03641_ = _05381_ & _06686_;
  assign _03644_ = _05385_ & _06686_;
  assign _03647_ = _05389_ & _06686_;
  assign _03668_ = _05417_ & _06686_;
  assign _03671_ = _05421_ & _06686_;
  assign _03674_ = _05425_ & _06686_;
  assign _03677_ = _05429_ & _06686_;
  assign _03679_ = _03678_ | _01099_;
  assign _03683_ = _01101_ | _01102_;
  assign _03687_ = _01104_ | _01105_;
  assign _03691_ = _01107_ | _01108_;
  assign _03719_ = _01128_ | _01129_;
  assign _03723_ = _01131_ | _01132_;
  assign _03727_ = _01134_ | _01135_;
  assign _03731_ = _01137_ | _01138_;
  assign _03735_ = _01140_ | _01141_;
  assign _03743_ = _01146_ | _01147_;
  assign _03755_ = _01155_ | _01156_;
  assign _03795_ = _01186_ | _01187_;
  assign _03799_ = _01189_ | _01190_;
  assign _03803_ = _01192_ | _01193_;
  assign _03811_ = _01198_ | _01199_;
  assign _03831_ = _01213_ | _01214_;
  assign _03851_ = _01228_ | _01229_;
  assign _03855_ = _01231_ | _01232_;
  assign _03859_ = _01234_ | _01235_;
  assign _03863_ = _01237_ | _01238_;
  assign _03867_ = _01240_ | _01241_;
  assign _03871_ = _01243_ | _01244_;
  assign _03875_ = _01246_ | _01247_;
  assign _03879_ = _01249_ | _01250_;
  assign _03883_ = _01252_ | _01253_;
  assign _03887_ = _01255_ | _01256_;
  assign _03891_ = _01258_ | _01259_;
  assign _03895_ = _01261_ | _01262_;
  assign _03899_ = _01264_ | _01265_;
  assign _03903_ = _01267_ | _01268_;
  assign _03907_ = _01270_ | _01271_;
  assign _03911_ = _01273_ | _01274_;
  assign _03915_ = _01276_ | _01277_;
  assign _03919_ = _01279_ | _01280_;
  assign _03923_ = _01282_ | _01283_;
  assign _03927_ = _01285_ | _01286_;
  assign _03931_ = _01288_ | _01289_;
  assign _03935_ = _01291_ | _01292_;
  assign _03939_ = _01294_ | _01295_;
  assign _03943_ = _01297_ | _01298_;
  assign _03947_ = _01300_ | _01301_;
  assign _03951_ = _01303_ | _01304_;
  assign _03955_ = _01306_ | _01307_;
  assign _03959_ = _01309_ | _01310_;
  assign _03963_ = _01312_ | _01313_;
  assign _03967_ = _01315_ | _01316_;
  assign _03971_ = _01318_ | _01319_;
  assign _03975_ = _01321_ | _01322_;
  assign _03979_ = _01324_ | _01325_;
  assign _05164_ = _03475_ | _03476_;
  assign _05168_ = _03478_ | _03479_;
  assign _05172_ = _03481_ | _03482_;
  assign _05184_ = _03490_ | _03491_;
  assign _05188_ = _03493_ | _03494_;
  assign _05196_ = _03499_ | _03500_;
  assign _05200_ = _03502_ | _03503_;
  assign _05204_ = _03505_ | _03506_;
  assign _05208_ = _03508_ | _03509_;
  assign _05212_ = _03511_ | _03512_;
  assign _05218_ = _03516_ | _03517_;
  assign _05222_ = _03519_ | _03520_;
  assign _05230_ = _03525_ | _03526_;
  assign _05238_ = _03531_ | _03532_;
  assign _05242_ = _03534_ | _03535_;
  assign _05246_ = _03537_ | _03538_;
  assign _05250_ = _03540_ | _03541_;
  assign _05254_ = _03543_ | _03544_;
  assign _05258_ = _03546_ | _03547_;
  assign _05262_ = _03549_ | _03550_;
  assign _05266_ = _03552_ | _03553_;
  assign _05270_ = _03555_ | _03556_;
  assign _05274_ = _03558_ | _03559_;
  assign _05278_ = _03561_ | _03562_;
  assign _05282_ = _03564_ | _03565_;
  assign _05286_ = _03567_ | _03568_;
  assign _05290_ = _03570_ | _03571_;
  assign _05294_ = _03573_ | _03574_;
  assign _05298_ = _03576_ | _03577_;
  assign _05302_ = _03579_ | _03580_;
  assign _05306_ = _03582_ | _03583_;
  assign _05314_ = _03588_ | _03589_;
  assign _05318_ = _03591_ | _03592_;
  assign _05322_ = _03594_ | _03595_;
  assign _05326_ = _03597_ | _03598_;
  assign _05330_ = _03600_ | _03601_;
  assign _05334_ = _03603_ | _03604_;
  assign _05338_ = _03606_ | _03607_;
  assign _05342_ = _03609_ | _03610_;
  assign _05382_ = _03639_ | _03640_;
  assign _05386_ = _03642_ | _03643_;
  assign _05390_ = _03645_ | _03646_;
  assign _05418_ = _03666_ | _03667_;
  assign _05422_ = _03669_ | _03670_;
  assign _05426_ = _03672_ | _03673_;
  assign _05430_ = _03675_ | _03676_;
  assign _03680_ = _03679_ | _01100_;
  assign _03684_ = _03683_ | _01103_;
  assign _03688_ = _03687_ | _01106_;
  assign _03692_ = _03691_ | _01109_;
  assign _03720_ = _03719_ | _01130_;
  assign _03724_ = _03723_ | _01133_;
  assign _03728_ = _03727_ | _01136_;
  assign _03732_ = _03731_ | _01139_;
  assign _03736_ = _03735_ | _01142_;
  assign _03744_ = _03743_ | _01148_;
  assign _03756_ = _03755_ | _01157_;
  assign _03796_ = _03795_ | _01188_;
  assign _03800_ = _03799_ | _01191_;
  assign _03804_ = _03803_ | _01194_;
  assign _03812_ = _03811_ | _01200_;
  assign _03832_ = _03831_ | _01215_;
  assign _03852_ = _03851_ | _01230_;
  assign _03856_ = _03855_ | _01233_;
  assign _03860_ = _03859_ | _01236_;
  assign _03864_ = _03863_ | _01239_;
  assign _03868_ = _03867_ | _01242_;
  assign _03872_ = _03871_ | _01245_;
  assign _03876_ = _03875_ | _01248_;
  assign _03880_ = _03879_ | _01251_;
  assign _03884_ = _03883_ | _01254_;
  assign _03888_ = _03887_ | _01257_;
  assign _03892_ = _03891_ | _01260_;
  assign _03896_ = _03895_ | _01263_;
  assign _03900_ = _03899_ | _01266_;
  assign _03904_ = _03903_ | _01269_;
  assign _03908_ = _03907_ | _01272_;
  assign _03912_ = _03911_ | _01275_;
  assign _03916_ = _03915_ | _01278_;
  assign _03920_ = _03919_ | _01281_;
  assign _03924_ = _03923_ | _01284_;
  assign _03928_ = _03927_ | _01287_;
  assign _03932_ = _03931_ | _01290_;
  assign _03936_ = _03935_ | _01293_;
  assign _03940_ = _03939_ | _01296_;
  assign _03944_ = _03943_ | _01299_;
  assign _03948_ = _03947_ | _01302_;
  assign _03952_ = _03951_ | _01305_;
  assign _03956_ = _03955_ | _01308_;
  assign _03960_ = _03959_ | _01311_;
  assign _03964_ = _03963_ | _01314_;
  assign _03968_ = _03967_ | _01317_;
  assign _03972_ = _03971_ | _01320_;
  assign _03976_ = _03975_ | _01323_;
  assign _03980_ = _03979_ | _01326_;
  assign _05165_ = _05164_ | _03477_;
  assign _05169_ = _05168_ | _03480_;
  assign _05173_ = _05172_ | _03483_;
  assign _05185_ = _05184_ | _03492_;
  assign _05189_ = _05188_ | _03495_;
  assign _05197_ = _05196_ | _03501_;
  assign _05201_ = _05200_ | _03504_;
  assign _05205_ = _05204_ | _03507_;
  assign _05209_ = _05208_ | _03510_;
  assign _05213_ = _05212_ | _03513_;
  assign _05219_ = _05218_ | _03518_;
  assign _05223_ = _05222_ | _03521_;
  assign _05231_ = _05230_ | _03527_;
  assign _05239_ = _05238_ | _03533_;
  assign _05243_ = _05242_ | _03536_;
  assign _05247_ = _05246_ | _03539_;
  assign _05251_ = _05250_ | _03542_;
  assign _05255_ = _05254_ | _03545_;
  assign _05259_ = _05258_ | _03548_;
  assign _05263_ = _05262_ | _03551_;
  assign _05267_ = _05266_ | _03554_;
  assign _05271_ = _05270_ | _03557_;
  assign _05275_ = _05274_ | _03560_;
  assign _05279_ = _05278_ | _03563_;
  assign _05283_ = _05282_ | _03566_;
  assign _05287_ = _05286_ | _03569_;
  assign _05291_ = _05290_ | _03572_;
  assign _05295_ = _05294_ | _03575_;
  assign _05299_ = _05298_ | _03578_;
  assign _05303_ = _05302_ | _03581_;
  assign _05307_ = _05306_ | _03584_;
  assign _05315_ = _05314_ | _03590_;
  assign _05319_ = _05318_ | _03593_;
  assign _05323_ = _05322_ | _03596_;
  assign _05327_ = _05326_ | _03599_;
  assign _05331_ = _05330_ | _03602_;
  assign _05335_ = _05334_ | _03605_;
  assign _05339_ = _05338_ | _03608_;
  assign _05343_ = _05342_ | _03611_;
  assign _05383_ = _05382_ | _03641_;
  assign _05387_ = _05386_ | _03644_;
  assign _05391_ = _05390_ | _03647_;
  assign _05419_ = _05418_ | _03668_;
  assign _05423_ = _05422_ | _03671_;
  assign _05427_ = _05426_ | _03674_;
  assign _05431_ = _05430_ | _03677_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lbu_t0 */
  always_ff @(posedge clk)
    instr_lbu_t0 <= _03680_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lw_t0 */
  always_ff @(posedge clk)
    instr_lw_t0 <= _03684_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lh_t0 */
  always_ff @(posedge clk)
    instr_lh_t0 <= _03688_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lb_t0 */
  always_ff @(posedge clk)
    instr_lb_t0 <= _03692_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_jalr_t0 */
  always_ff @(posedge clk)
    instr_jalr_t0 <= _03720_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_jal_t0 */
  always_ff @(posedge clk)
    instr_jal_t0 <= _03724_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_auipc_t0 */
  always_ff @(posedge clk)
    instr_auipc_t0 <= _03728_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lui_t0 */
  always_ff @(posedge clk)
    instr_lui_t0 <= _03732_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_insn_t0 */
  always_ff @(posedge clk)
    pcpi_insn_t0 <= _03736_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_rd_t0 */
  always_ff @(posedge clk)
    latched_rd_t0 <= _03744_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_compr_t0 */
  always_ff @(posedge clk)
    latched_compr_t0 <= _03756_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_rs2_t0 */
  always_ff @(posedge clk)
    pcpi_rs2_t0 <= _03796_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_rs1_t0[31] */
  always_ff @(posedge clk)
    pcpi_rs1_t0[31] <= _03800_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_rs1_t0[30:0] */
  always_ff @(posedge clk)
    pcpi_rs1_t0[30:0] <= _03804_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_wordsize_t0 */
  always_ff @(posedge clk)
    mem_wordsize_t0 <= _03812_;
  reg [7:0] _08966_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME _08966_ */
  always_ff @(posedge clk)
    _08966_ <= _03832_;
  assign { rvfi_insn_t0[24:20], rvfi_insn_t0[14:12] } = _08966_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_pc_wdata_t0[31:1] */
  always_ff @(posedge clk)
    rvfi_pc_wdata_t0[31:1] <= _03852_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[9]_t0  */
  always_ff @(posedge clk)
    \cpuregs[9]_t0  <= _03856_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[8]_t0  */
  always_ff @(posedge clk)
    \cpuregs[8]_t0  <= _03860_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[7]_t0  */
  always_ff @(posedge clk)
    \cpuregs[7]_t0  <= _03864_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[6]_t0  */
  always_ff @(posedge clk)
    \cpuregs[6]_t0  <= _03868_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[5]_t0  */
  always_ff @(posedge clk)
    \cpuregs[5]_t0  <= _03872_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[4]_t0  */
  always_ff @(posedge clk)
    \cpuregs[4]_t0  <= _03876_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[3]_t0  */
  always_ff @(posedge clk)
    \cpuregs[3]_t0  <= _03880_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[31]_t0  */
  always_ff @(posedge clk)
    \cpuregs[31]_t0  <= _03884_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[30]_t0  */
  always_ff @(posedge clk)
    \cpuregs[30]_t0  <= _03888_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[2]_t0  */
  always_ff @(posedge clk)
    \cpuregs[2]_t0  <= _03892_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[29]_t0  */
  always_ff @(posedge clk)
    \cpuregs[29]_t0  <= _03896_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[28]_t0  */
  always_ff @(posedge clk)
    \cpuregs[28]_t0  <= _03900_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[27]_t0  */
  always_ff @(posedge clk)
    \cpuregs[27]_t0  <= _03904_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[26]_t0  */
  always_ff @(posedge clk)
    \cpuregs[26]_t0  <= _03908_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[25]_t0  */
  always_ff @(posedge clk)
    \cpuregs[25]_t0  <= _03912_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[24]_t0  */
  always_ff @(posedge clk)
    \cpuregs[24]_t0  <= _03916_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[23]_t0  */
  always_ff @(posedge clk)
    \cpuregs[23]_t0  <= _03920_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[22]_t0  */
  always_ff @(posedge clk)
    \cpuregs[22]_t0  <= _03924_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[21]_t0  */
  always_ff @(posedge clk)
    \cpuregs[21]_t0  <= _03928_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[20]_t0  */
  always_ff @(posedge clk)
    \cpuregs[20]_t0  <= _03932_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[1]_t0  */
  always_ff @(posedge clk)
    \cpuregs[1]_t0  <= _03936_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[19]_t0  */
  always_ff @(posedge clk)
    \cpuregs[19]_t0  <= _03940_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[18]_t0  */
  always_ff @(posedge clk)
    \cpuregs[18]_t0  <= _03944_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[17]_t0  */
  always_ff @(posedge clk)
    \cpuregs[17]_t0  <= _03948_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[16]_t0  */
  always_ff @(posedge clk)
    \cpuregs[16]_t0  <= _03952_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[15]_t0  */
  always_ff @(posedge clk)
    \cpuregs[15]_t0  <= _03956_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[14]_t0  */
  always_ff @(posedge clk)
    \cpuregs[14]_t0  <= _03960_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[13]_t0  */
  always_ff @(posedge clk)
    \cpuregs[13]_t0  <= _03964_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[12]_t0  */
  always_ff @(posedge clk)
    \cpuregs[12]_t0  <= _03968_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[11]_t0  */
  always_ff @(posedge clk)
    \cpuregs[11]_t0  <= _03972_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[10]_t0  */
  always_ff @(posedge clk)
    \cpuregs[10]_t0  <= _03976_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[0]_t0  */
  always_ff @(posedge clk)
    \cpuregs[0]_t0  <= _03980_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_rdata_q_t0[6:0] */
  always_ff @(posedge clk)
    mem_rdata_q_t0[6:0] <= _05165_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME next_insn_opcode_t0 */
  always_ff @(posedge clk)
    next_insn_opcode_t0 <= _05169_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_16bit_buffer_t0 */
  always_ff @(posedge clk)
    mem_16bit_buffer_t0 <= _05173_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_state_t0 */
  always_ff @(posedge clk)
    mem_state_t0 <= _05185_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_wstrb_t0 */
  always_ff @(posedge clk)
    mem_wstrb_t0 <= _05189_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_addr_t0 */
  always_ff @(posedge clk)
    mem_addr_t0 <= _05197_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME cached_insn_opcode_t0 */
  always_ff @(posedge clk)
    cached_insn_opcode_t0 <= _05201_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_valid_t0 */
  always_ff @(posedge clk)
    mem_valid_t0 <= _05205_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME cached_insn_rs2_t0 */
  always_ff @(posedge clk)
    cached_insn_rs2_t0 <= _05209_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME cached_insn_rs1_t0 */
  always_ff @(posedge clk)
    cached_insn_rs1_t0 <= _05213_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_alu_reg_reg_t0 */
  always_ff @(posedge clk)
    is_alu_reg_reg_t0 <= _05219_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_alu_reg_imm_t0 */
  always_ff @(posedge clk)
    is_alu_reg_imm_t0 <= _05223_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_ecall_ebreak_t0 */
  always_ff @(posedge clk)
    instr_ecall_ebreak_t0 <= _05231_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_sll_srl_sra_t0 */
  always_ff @(posedge clk)
    is_sll_srl_sra_t0 <= _05239_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_sb_sh_sw_t0 */
  always_ff @(posedge clk)
    is_sb_sh_sw_t0 <= _05243_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_jalr_addi_slti_sltiu_xori_ori_andi_t0 */
  always_ff @(posedge clk)
    is_jalr_addi_slti_sltiu_xori_ori_andi_t0 <= _05247_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_slli_srli_srai_t0 */
  always_ff @(posedge clk)
    is_slli_srli_srai_t0 <= _05251_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_lb_lh_lw_lbu_lhu_t0 */
  always_ff @(posedge clk)
    is_lb_lh_lw_lbu_lhu_t0 <= _05255_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME compressed_instr_t0 */
  always_ff @(posedge clk)
    compressed_instr_t0 <= _05259_;
  reg \decoded_imm_j_t0_reg[10] ;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_t0_reg[10]  */
  always_ff @(posedge clk)
    \decoded_imm_j_t0_reg[10]  <= _05263_;
  assign decoded_imm_j_t0[10] = \decoded_imm_j_t0_reg[10] ;
  reg \decoded_imm_j_t0_reg[7] ;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_t0_reg[7]  */
  always_ff @(posedge clk)
    \decoded_imm_j_t0_reg[7]  <= _05267_;
  assign decoded_imm_j_t0[7] = \decoded_imm_j_t0_reg[7] ;
  reg \decoded_imm_j_t0_reg[6] ;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_t0_reg[6]  */
  always_ff @(posedge clk)
    \decoded_imm_j_t0_reg[6]  <= _05271_;
  assign decoded_imm_j_t0[6] = \decoded_imm_j_t0_reg[6] ;
  reg [2:0] _09022_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME _09022_ */
  always_ff @(posedge clk)
    _09022_ <= _05275_;
  assign decoded_imm_j_t0[3:1] = _09022_;
  reg \decoded_imm_j_t0_reg[5] ;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_t0_reg[5]  */
  always_ff @(posedge clk)
    \decoded_imm_j_t0_reg[5]  <= _05279_;
  assign decoded_imm_j_t0[5] = \decoded_imm_j_t0_reg[5] ;
  reg [1:0] _09024_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME _09024_ */
  always_ff @(posedge clk)
    _09024_ <= _05283_;
  assign decoded_imm_j_t0[9:8] = _09024_;
  reg [11:0] _09025_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME _09025_ */
  always_ff @(posedge clk)
    _09025_ <= _05287_;
  assign decoded_imm_j_t0[31:20] = _09025_;
  reg \decoded_imm_j_t0_reg[4] ;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_t0_reg[4]  */
  always_ff @(posedge clk)
    \decoded_imm_j_t0_reg[4]  <= _05291_;
  assign decoded_imm_j_t0[4] = \decoded_imm_j_t0_reg[4] ;
  reg \decoded_imm_j_t0_reg[11] ;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_t0_reg[11]  */
  always_ff @(posedge clk)
    \decoded_imm_j_t0_reg[11]  <= _05295_;
  assign decoded_imm_j_t0[11] = \decoded_imm_j_t0_reg[11] ;
  reg [7:0] _09028_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME _09028_ */
  always_ff @(posedge clk)
    _09028_ <= _05299_;
  assign decoded_imm_j_t0[19:12] = _09028_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_imm_t0 */
  always_ff @(posedge clk)
    decoded_imm_t0 <= _05303_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_rs2_t0 */
  always_ff @(posedge clk)
    decoded_rs2_t0 <= _05307_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_wdata_t0 */
  always_ff @(posedge clk)
    mem_wdata_t0 <= _05315_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_rs1_t0[4] */
  always_ff @(posedge clk)
    decoded_rs1_t0[4] <= _05319_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_rs1_t0[3:0] */
  always_ff @(posedge clk)
    decoded_rs1_t0[3:0] <= _05323_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_rd_t0 */
  always_ff @(posedge clk)
    decoded_rd_t0 <= _05327_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_rdinstrh_t0 */
  always_ff @(posedge clk)
    instr_rdinstrh_t0 <= _05331_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_rdinstr_t0 */
  always_ff @(posedge clk)
    instr_rdinstr_t0 <= _05335_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_rdcycleh_t0 */
  always_ff @(posedge clk)
    instr_rdcycleh_t0 <= _05339_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_rdcycle_t0 */
  always_ff @(posedge clk)
    instr_rdcycle_t0 <= _05343_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_srai_t0 */
  always_ff @(posedge clk)
    instr_srai_t0 <= _05383_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_srli_t0 */
  always_ff @(posedge clk)
    instr_srli_t0 <= _05387_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_slli_t0 */
  always_ff @(posedge clk)
    instr_slli_t0 <= _05391_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sw_t0 */
  always_ff @(posedge clk)
    instr_sw_t0 <= _05419_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sh_t0 */
  always_ff @(posedge clk)
    instr_sh_t0 <= _05423_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sb_t0 */
  always_ff @(posedge clk)
    instr_sb_t0 <= _05427_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lhu_t0 */
  always_ff @(posedge clk)
    instr_lhu_t0 <= _05431_;
  assign _00180_ = | { mem_do_rdata_t0, mem_la_read_t0 };
  assign _00181_ = | { mem_la_use_prefetched_high_word_t0, mem_la_read_t0 };
  assign _00182_ = | { _00797_, _06538_, mem_do_rinst_t0 };
  assign _00183_ = | { _00797_, _06837_, _06885_, mem_do_wdata_t0 };
  assign _00184_ = | { _00797_, _07440_, mem_xfer_t0 };
  assign _00185_ = | { _00797_, _06536_, mem_xfer_t0 };
  assign _00186_ = | { _00797_, _07440_, mem_la_read_t0, mem_xfer_t0 };
  assign _00187_ = | { _00797_, _06890_ };
  assign _00188_ = | { _06492_, is_beq_bne_blt_bge_bltu_bgeu_t0 };
  assign _00189_ = | { _06498_, _06866_, mem_do_rdata_t0 };
  assign _00190_ = | { _06498_, _06866_ };
  assign _00191_ = | { is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, instr_trap_t0, _06488_ };
  assign _00192_ = | { instr_trap_t0, _06490_ };
  assign _00193_ = | { _01081_, _01093_, _06614_, instr_trap_t0, _06488_, _06873_, is_sll_srl_sra_t0 };
  assign _00194_ = | { _06490_, _06873_, is_sll_srl_sra_t0 };
  assign _00195_ = | { _06494_, _06500_, _06873_ };
  assign _00196_ = | { _01093_, _06488_, _06873_ };
  assign _00197_ = | { _06494_, _06488_, _06490_, _06873_, _06486_ };
  assign _00198_ = | { _06496_, _06866_, mem_do_wdata_t0 };
  assign _00199_ = | { _06850_, _06860_, _06858_, _06598_, _06494_, _06500_ };
  assign _00200_ = | { _06850_, _06598_, _06494_, _06500_ };
  assign _00201_ = | { _06494_, _06500_ };
  assign _00202_ = | { _06496_, _06866_ };
  assign _00203_ = | { _06215_[1], _06868_, _06498_, _06866_, mem_do_rdata_t0, instr_lw_t0 };
  assign _00204_ = | { _06496_, _06866_, instr_sb_t0, instr_sh_t0, instr_sw_t0, mem_do_wdata_t0 };
  assign _00205_ = | { _00858_, instr_trap_t0 };
  assign _00206_ = | { pcpi_rs2_t0, pcpi_rs1_t0 };
  assign _00207_ = | rvfi_insn_t0[6:0];
  assign _00208_ = | rvfi_insn_t0[13:12];
  assign _00209_ = | rvfi_insn_t0[31:20];
  assign _00212_ = | mem_rdata_latched_t0[6:0];
  assign _00214_ = | mem_rdata_latched_t0[12:10];
  assign _00215_ = | mem_rdata_q_t0[31:20];
  assign _00216_ = | mem_rdata_q_t0[6:0];
  assign _00217_ = | mem_rdata_q_t0[15:0];
  assign _00221_ = | cpu_state_t0;
  assign _07610_ = pcpi_rs1_t0 | pcpi_rs2_t0;
  assign _00226_ = ~ { mem_la_read_t0, mem_do_rdata_t0 };
  assign _00227_ = ~ { mem_la_read_t0, mem_la_use_prefetched_high_word_t0 };
  assign _00228_ = ~ { _00797_, 1'h0 };
  assign _00229_ = ~ { _06538_, _00797_, mem_do_rinst_t0 };
  assign _00230_ = ~ { _06837_, _00797_, _06885_, mem_do_wdata_t0 };
  assign _00231_ = ~ { _07440_, _00797_, mem_xfer_t0 };
  assign _00232_ = ~ { _06536_, _00797_, mem_xfer_t0 };
  assign _00233_ = ~ { _07440_, _00797_, mem_la_read_t0, mem_xfer_t0 };
  assign _00234_ = ~ { _00797_, _06890_ };
  assign _00235_ = ~ { _06492_, is_beq_bne_blt_bge_bltu_bgeu_t0 };
  assign _00236_ = ~ { _06498_, _06866_, mem_do_rdata_t0 };
  assign _00237_ = ~ { _06498_, _06866_ };
  assign _00238_ = ~ { _06488_, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, instr_trap_t0 };
  assign _00239_ = ~ { _06490_, instr_trap_t0 };
  assign _00240_ = ~ { _01081_, _06488_, _01093_, _06873_, _06614_, instr_trap_t0, is_sll_srl_sra_t0, 1'h0 };
  assign _00241_ = ~ { _06490_, _06873_, is_sll_srl_sra_t0, 1'h0 };
  assign _00242_ = ~ { _06494_, _06873_, _06500_, 1'h0 };
  assign _00243_ = ~ { _06488_, _01093_, _06873_, 1'h0 };
  assign _00244_ = ~ { _06488_, _06490_, _06486_, _06494_, _06873_, 1'h0 };
  assign _00245_ = ~ { _06496_, _06866_, mem_do_wdata_t0 };
  assign _00246_ = ~ { _06494_, _06850_, _06860_, _06858_, _06598_, _06500_ };
  assign _00247_ = ~ { _06494_, _06850_, _06598_, _06500_ };
  assign _00248_ = ~ { _06494_, _06500_ };
  assign _00249_ = ~ { _06496_, _06866_ };
  assign _00250_ = ~ { _06498_, _06215_[1], _06868_, _06866_, instr_lw_t0, mem_do_rdata_t0 };
  assign _00251_ = ~ { _06496_, _06866_, instr_sw_t0, instr_sh_t0, instr_sb_t0, mem_do_wdata_t0 };
  assign _00252_ = ~ { _00858_, instr_trap_t0 };
  assign _00253_ = ~ _07610_;
  assign _00254_ = ~ rvfi_insn_t0[6:0];
  assign _00255_ = ~ rvfi_insn_t0[13:12];
  assign _00256_ = ~ rvfi_insn_t0[31:20];
  assign _00257_ = ~ mem_rdata_latched_t0[11:10];
  assign _00258_ = ~ mem_rdata_latched_t0[6:5];
  assign _00259_ = ~ mem_rdata_latched_t0[6:0];
  assign _00260_ = ~ mem_rdata_latched_t0[11:7];
  assign _00261_ = ~ mem_rdata_latched_t0[12:10];
  assign _00262_ = ~ mem_rdata_q_t0[31:20];
  assign _00263_ = ~ mem_rdata_q_t0[6:0];
  assign _00264_ = ~ mem_rdata_q_t0[15:0];
  assign _00265_ = ~ mem_rdata_q_t0[14:12];
  assign _00266_ = ~ mem_rdata_q_t0[31:25];
  assign _00267_ = ~ mem_rdata_latched_t0[1:0];
  assign _00268_ = ~ cpu_state_t0;
  assign _00269_ = ~ mem_rdata_latched_t0[15:13];
  assign _00270_ = ~ mem_state_t0;
  assign _00271_ = ~ pcpi_rs1_t0[1:0];
  assign _00272_ = ~ mem_wordsize_t0;
  assign _01456_ = { mem_la_read, mem_do_rdata } & _00226_;
  assign _01457_ = { mem_la_read, mem_la_use_prefetched_high_word } & _00227_;
  assign _01458_ = { _06888_, resetn } & _00228_;
  assign _01459_ = { _06537_, _06888_, mem_do_rinst } & _00229_;
  assign _01460_ = { _06836_, _06888_, _06884_, mem_do_wdata } & _00230_;
  assign _01461_ = { _07439_, _06888_, mem_xfer } & _00231_;
  assign _01462_ = { _06535_, _06888_, mem_xfer } & _00232_;
  assign _01463_ = { _07439_, _06888_, mem_la_read, mem_xfer } & _00233_;
  assign _01466_ = { _06888_, _06889_ } & _00234_;
  assign _01470_ = { _06491_, is_beq_bne_blt_bge_bltu_bgeu } & _00235_;
  assign _01472_ = { _06497_, _06865_, mem_do_rdata } & _00236_;
  assign _01473_ = { _06497_, _06865_ } & _00237_;
  assign _01475_ = { _06487_, is_rdcycle_rdcycleh_rdinstr_rdinstrh, instr_trap } & _00238_;
  assign _01476_ = { _06489_, instr_trap } & _00239_;
  assign _01479_ = { _01080_, _06487_, _01092_, _06872_, _06613_, instr_trap, is_sll_srl_sra, resetn } & _00240_;
  assign _01480_ = { _06489_, _06872_, is_sll_srl_sra, resetn } & _00241_;
  assign _01481_ = { _06493_, _06872_, _06499_, resetn } & _00242_;
  assign _01482_ = { _06487_, _01092_, _06872_, resetn } & _00243_;
  assign _01483_ = { _06487_, _06489_, _06485_, _06493_, _06872_, resetn } & _00244_;
  assign _01484_ = { _06495_, _06865_, mem_do_wdata } & _00245_;
  assign _01485_ = { _06493_, _06849_, _06859_, _06857_, _06597_, _06499_ } & _00246_;
  assign _01486_ = { _06493_, _06849_, _06597_, _06499_ } & _00247_;
  assign _01487_ = { _06493_, _06499_ } & _00248_;
  assign _01488_ = { _06495_, _06865_ } & _00249_;
  assign _01490_ = { _06497_, _06869_, _06867_, _06865_, instr_lw, mem_do_rdata } & _00250_;
  assign _01491_ = { _06495_, _06865_, instr_sw, instr_sh, instr_sb, mem_do_wdata } & _00251_;
  assign _01494_ = { _00857_, instr_trap } & _00252_;
  assign _02085_ = pcpi_rs1 & _00253_;
  assign _02088_ = rvfi_insn[6:0] & _00254_;
  assign _02089_ = rvfi_insn[13:12] & _00255_;
  assign _02090_ = rvfi_insn[31:20] & _00256_;
  assign _02091_ = mem_rdata_latched[11:10] & _00257_;
  assign _02092_ = mem_rdata_latched[6:5] & _00258_;
  assign _02093_ = mem_rdata_latched[6:0] & _00259_;
  assign _02095_ = mem_rdata_latched[11:7] & _00260_;
  assign _02096_ = mem_rdata_latched[12:10] & _00261_;
  assign _02098_ = mem_rdata_q[31:20] & _00262_;
  assign _02099_ = mem_rdata_q[6:0] & _00263_;
  assign _02100_ = mem_rdata_q[15:0] & _00264_;
  assign _02101_ = mem_rdata_q[14:12] & _00265_;
  assign _02102_ = mem_rdata_q[31:25] & _00266_;
  assign _02778_ = mem_rdata_latched[1:0] & _00267_;
  assign _02814_ = cpu_state & _00268_;
  assign _03043_ = mem_rdata_latched[15:13] & _00269_;
  assign _03135_ = mem_state & _00270_;
  assign _02777_ = pcpi_rs1[1:0] & _00271_;
  assign _03291_ = mem_wordsize & _00272_;
  assign _02086_ = pcpi_rs2 & _00253_;
  assign _05969_ = _01456_ == { 1'h0, _00226_[0] };
  assign _05970_ = _01457_ == _00227_;
  assign _05971_ = _01458_ == _00228_;
  assign _05972_ = _01459_ == { _00229_[2], 2'h0 };
  assign _05973_ = _01460_ == { _00230_[3], 3'h0 };
  assign _05974_ = _01461_ == { _00231_[2], 2'h0 };
  assign _05975_ = _01462_ == { _00232_[2], 2'h0 };
  assign _05976_ = _01463_ == { _00233_[3], 1'h0, _00233_[1:0] };
  assign _05977_ = _01466_ == { _00234_[1], 1'h0 };
  assign _05978_ = _01470_ == { _00235_[1], 1'h0 };
  assign _05979_ = _01472_ == _00236_;
  assign _05980_ = _01473_ == { _00237_[1], 1'h0 };
  assign _05981_ = _01470_ == _00235_;
  assign _05982_ = _01475_ == { _00238_[2], 2'h0 };
  assign _05983_ = _01476_ == { _00239_[1], 1'h0 };
  assign _05984_ = _01479_ == { 1'h0, _00240_[6], 4'h0, _00240_[1:0] };
  assign _05985_ = _01480_ == { _00241_[3], 1'h0, _00241_[1:0] };
  assign _05986_ = _01481_ == { _00242_[3], 2'h0, _00242_[0] };
  assign _05987_ = _01482_ == { _00243_[3:2], 1'h0, _00243_[0] };
  assign _05988_ = _01483_ == { 5'h00, _00244_[0] };
  assign _05989_ = _01484_ == _00245_;
  assign _05990_ = _01485_ == { _00246_[5], 5'h00 };
  assign _05991_ = _01486_ == { _00247_[3:2], 2'h0 };
  assign _05992_ = _01485_ == { _00246_[5], 3'h0, _00246_[1], 1'h0 };
  assign _05993_ = _01486_ == { _00247_[3:1], 1'h0 };
  assign _05994_ = _01487_ == _00248_;
  assign _05995_ = _01488_ == { _00249_[1], 1'h0 };
  assign _05996_ = _01490_ == { _00250_[5], 2'h0, _00250_[2], 2'h0 };
  assign _05997_ = _01491_ == { _00251_[5:4], 4'h0 };
  assign _05998_ = _01494_ == { _00252_[1], 1'h0 };
  assign _05999_ = _02085_ == _02086_;
  assign _06000_ = _02088_ == { _00254_[6:4], 2'h0, _00254_[1:0] };
  assign _06001_ = _02089_ == { _00255_[1], 1'h0 };
  assign _06002_ = _02090_ == { _00256_[11:10], 10'h000 };
  assign _06003_ = _02090_ == { _00256_[11:10], 2'h0, _00256_[7], 7'h00 };
  assign _06004_ = _02090_ == { _00256_[11:10], 8'h00, _00256_[1], 1'h0 };
  assign _06005_ = _02090_ == { _00256_[11:10], 2'h0, _00256_[7], 5'h00, _00256_[1], 1'h0 };
  assign _06006_ = _02091_ == { 1'h0, _00257_[0] };
  assign _06007_ = _02092_ == { 1'h0, _00258_[0] };
  assign _06008_ = _02092_ == { _00258_[1], 1'h0 };
  assign _06009_ = _02092_ == _00258_;
  assign _06010_ = _02093_ == { 1'h0, _00259_[5:4], 1'h0, _00259_[2:0] };
  assign _06011_ = _02093_ == { 2'h0, _00259_[4], 1'h0, _00259_[2:0] };
  assign _06012_ = _02093_ == { _00259_[6:5], 1'h0, _00259_[3:0] };
  assign _06013_ = _02093_ == { _00259_[6:5], 2'h0, _00259_[2:0] };
  assign _06014_ = _02093_ == { _00259_[6:5], 3'h0, _00259_[1:0] };
  assign _06015_ = _02093_ == { 5'h00, _00259_[1:0] };
  assign _06016_ = _02093_ == { 1'h0, _00259_[5], 3'h0, _00259_[1:0] };
  assign _06017_ = _02093_ == { 2'h0, _00259_[4], 2'h0, _00259_[1:0] };
  assign _06018_ = _02093_ == { 1'h0, _00259_[5:4], 2'h0, _00259_[1:0] };
  assign _06019_ = _02095_ == { 3'h0, _00260_[1], 1'h0 };
  assign _06020_ = _02091_ == { _00257_[1], 1'h0 };
  assign _06021_ = _02096_ == { 1'h0, _00261_[1:0] };
  assign _06022_ = _02098_ == { _00262_[11], 1'h0, _00262_[9:8], 8'h00 };
  assign _06023_ = _02098_ == { _00262_[11], 1'h0, _00262_[9:8], 7'h00, _00262_[0] };
  assign _06024_ = _02098_ == { _00262_[11], 1'h0, _00262_[9:7], 7'h00 };
  assign _06025_ = _02098_ == { _00262_[11], 1'h0, _00262_[9:7], 6'h00, _00262_[0] };
  assign _06026_ = _02098_ == { _00262_[11], 1'h0, _00262_[9:8], 6'h00, _00262_[1], 1'h0 };
  assign _06027_ = _02098_ == { _00262_[11], 1'h0, _00262_[9:7], 5'h00, _00262_[1], 1'h0 };
  assign _06028_ = _02099_ == { _00263_[6:4], 2'h0, _00263_[1:0] };
  assign _06029_ = _02100_ == { _00264_[15], 2'h0, _00264_[12], 10'h000, _00264_[1], 1'h0 };
  assign _06030_ = _02099_ == { 3'h0, _00263_[3:0] };
  assign _06031_ = _02101_ == _00265_;
  assign _06032_ = _02101_ == { _00265_[2:1], 1'h0 };
  assign _06033_ = _02101_ == { _00265_[2], 2'h0 };
  assign _06034_ = _02101_ == { 1'h0, _00265_[1:0] };
  assign _06035_ = _02101_ == { 1'h0, _00265_[1], 1'h0 };
  assign _06036_ = _02102_ == { 1'h0, _00266_[5], 5'h00 };
  assign _06037_ = _02101_ == { _00265_[2], 1'h0, _00265_[0] };
  assign _06038_ = _02101_ == { 2'h0, _00265_[0] };
  assign _06039_ = _02778_ == _00267_;
  assign _06040_ = _02814_ == { _00268_[7], 7'h00 };
  assign _06041_ = _02814_ == { 4'h0, _00268_[3], 3'h0 };
  assign _06042_ = _02814_ == { 7'h00, _00268_[0] };
  assign _06043_ = _02814_ == { 6'h00, _00268_[1], 1'h0 };
  assign _06044_ = _02814_ == { 5'h00, _00268_[2], 2'h0 };
  assign _06045_ = _02814_ == { 1'h0, _00268_[6], 6'h00 };
  assign _06046_ = _02814_ == { 3'h0, _00268_[4], 4'h0 };
  assign _06047_ = _02814_ == { 2'h0, _00268_[5], 5'h00 };
  assign _06048_ = _03043_ == { _00269_[2:1], 1'h0 };
  assign _06049_ = _03043_ == { 1'h0, _00269_[1], 1'h0 };
  assign _06050_ = _03043_ == { _00269_[2], 2'h0 };
  assign _06051_ = _02778_ == { _00267_[1], 1'h0 };
  assign _06052_ = _03043_ == { _00269_[2], 1'h0, _00269_[0] };
  assign _06053_ = _03043_ == { 2'h0, _00269_[0] };
  assign _06054_ = _03043_ == { 1'h0, _00269_[1:0] };
  assign _06055_ = _02778_ == { 1'h0, _00267_[0] };
  assign _06056_ = _03135_ == { 1'h0, _00270_[0] };
  assign _06057_ = _03135_ == _00270_;
  assign _06058_ = _03135_ == { _00270_[1], 1'h0 };
  assign _06059_ = _03043_ == _00269_;
  assign _06060_ = _02777_ == _00271_;
  assign _06061_ = _02777_ == { _00271_[1], 1'h0 };
  assign _06062_ = _02777_ == { 1'h0, _00271_[0] };
  assign _06063_ = _03291_ == { _00272_[1], 1'h0 };
  assign _06064_ = _03291_ == { 1'h0, _00272_[0] };
  assign _00946_ = _05969_ & _00180_;
  assign _00948_ = _05970_ & _00181_;
  assign _00950_ = _05971_ & _00797_;
  assign _00952_ = _05972_ & _00182_;
  assign _00954_ = _05973_ & _00183_;
  assign _00956_ = _05974_ & _00184_;
  assign _00958_ = _05975_ & _00185_;
  assign _00960_ = _05976_ & _00186_;
  assign _00966_ = _05977_ & _00187_;
  assign _00974_ = _05978_ & _00188_;
  assign _00978_ = _05979_ & _00189_;
  assign _00980_ = _05980_ & _00190_;
  assign _00984_ = _05981_ & _00188_;
  assign _00986_ = _05982_ & _00191_;
  assign _00988_ = _05983_ & _00192_;
  assign _00994_ = _05984_ & _00193_;
  assign _00996_ = _05985_ & _00194_;
  assign _00998_ = _05986_ & _00195_;
  assign _01000_ = _05987_ & _00196_;
  assign _01002_ = _05988_ & _00197_;
  assign _01004_ = _05989_ & _00198_;
  assign _01006_ = _05990_ & _00199_;
  assign _01008_ = _05991_ & _00200_;
  assign _01010_ = _05992_ & _00199_;
  assign _01012_ = _05993_ & _00200_;
  assign _01014_ = _05994_ & _00201_;
  assign _01016_ = _05995_ & _00202_;
  assign _01020_ = _05996_ & _00203_;
  assign _01022_ = _05997_ & _00204_;
  assign _01028_ = _05998_ & _00205_;
  assign alu_eq_t0 = _05999_ & _00206_;
  assign _06506_ = _06000_ & _00207_;
  assign _06508_ = _06001_ & _00208_;
  assign _00052_[31] = _06002_ & _00209_;
  assign _06511_ = _06003_ & _00209_;
  assign _00056_[31] = _06004_ & _00209_;
  assign _06514_ = _06005_ & _00209_;
  assign _06520_ = _06006_ & _00210_;
  assign _06528_ = _06007_ & _00211_;
  assign _06530_ = _06008_ & _00211_;
  assign _06532_ = _06009_ & _00211_;
  assign _06540_ = _06010_ & _00212_;
  assign _06542_ = _06011_ & _00212_;
  assign _06544_ = _06012_ & _00212_;
  assign _06546_ = _06013_ & _00212_;
  assign _06550_ = _06014_ & _00212_;
  assign _06552_ = _06015_ & _00212_;
  assign _06554_ = _06016_ & _00212_;
  assign _06556_ = _06017_ & _00212_;
  assign _06558_ = _06018_ & _00212_;
  assign _06516_ = _06019_ & _00213_;
  assign _06522_ = _06020_ & _00210_;
  assign _06524_ = _06021_ & _00214_;
  assign _06582_ = _06022_ & _00215_;
  assign _06584_ = _06023_ & _00215_;
  assign _06586_ = _06024_ & _00215_;
  assign _06588_ = _06025_ & _00215_;
  assign _06590_ = _06026_ & _00215_;
  assign _06592_ = _06027_ & _00215_;
  assign _06580_ = _06028_ & _00216_;
  assign _06594_ = _06029_ & _00217_;
  assign _06596_ = _06030_ & _00216_;
  assign _06570_ = _06031_ & _00218_;
  assign _06568_ = _06032_ & _00218_;
  assign _06564_ = _06033_ & _00218_;
  assign _06574_ = _06034_ & _00218_;
  assign _06572_ = _06035_ & _00218_;
  assign _06578_ = _06036_ & _00219_;
  assign _06566_ = _06037_ & _00218_;
  assign _06562_ = _06038_ & _00218_;
  assign _06678_ = _06039_ & _00220_;
  assign _06484_ = _06040_ & _00221_;
  assign _06492_ = _06041_ & _00221_;
  assign _06498_ = _06042_ & _00221_;
  assign _06496_ = _06043_ & _00221_;
  assign _06494_ = _06044_ & _00221_;
  assign _06486_ = _06045_ & _00221_;
  assign _06490_ = _06046_ & _00221_;
  assign _06488_ = _06047_ & _00221_;
  assign _07255_ = _06048_ & _00222_;
  assign _07271_ = _06049_ & _00222_;
  assign _07248_ = _06050_ & _00222_;
  assign _07252_ = _06051_ & _00220_;
  assign _07414_ = _06052_ & _00222_;
  assign _06362_[0] = _06053_ & _00222_;
  assign _07266_ = _06054_ & _00222_;
  assign _07268_ = _06055_ & _00220_;
  assign _07440_ = _06056_ & _00223_;
  assign _06538_ = _06057_ & _00223_;
  assign _06536_ = _06058_ & _00223_;
  assign _06427_[0] = _06059_ & _00222_;
  assign _07552_ = _06060_ & _00224_;
  assign _07554_ = _06061_ & _00224_;
  assign _07556_ = _06062_ & _00224_;
  assign _07558_ = _06063_ & _00225_;
  assign _06504_ = _06064_ & _00225_;
  /* src = "generated/out/vanilla.sv:302.2-311.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME last_mem_valid */
  always_ff @(posedge clk)
    if (!resetn) last_mem_valid <= 1'h0;
    else last_mem_valid <= _06661_;
  /* src = "generated/out/vanilla.sv:302.2-311.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_la_firstword_reg */
  always_ff @(posedge clk)
    if (!resetn) mem_la_firstword_reg <= 1'h0;
    else mem_la_firstword_reg <= _07559_;
  /* src = "generated/out/vanilla.sv:339.2-446.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_rdata_q[6:0] */
  always_ff @(posedge clk)
    if (mem_xfer) mem_rdata_q[6:0] <= mem_rdata_latched[6:0];
  /* src = "generated/out/vanilla.sv:339.2-446.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_rdata_q[31:7] */
  always_ff @(posedge clk)
    mem_rdata_q[31:7] <= _00020_[31:7];
  /* src = "generated/out/vanilla.sv:339.2-446.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME next_insn_opcode */
  always_ff @(posedge clk)
    if (mem_xfer) next_insn_opcode <= mem_rdata_latched;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_16bit_buffer */
  always_ff @(posedge clk)
    if (_01029_) mem_16bit_buffer <= _07437_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME prefetched_high_word */
  always_ff @(posedge clk)
    if (_01071_) prefetched_high_word <= 1'h0;
    else if (_01031_) prefetched_high_word <= _07441_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_la_secondword */
  always_ff @(posedge clk)
    if (_06888_) mem_la_secondword <= 1'h0;
    else if (_01033_) mem_la_secondword <= _07442_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_state */
  always_ff @(posedge clk)
    if (_01035_) mem_state <= _00022_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_wstrb */
  always_ff @(posedge clk)
    if (!_06888_) mem_wstrb <= _07456_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_instr */
  always_ff @(posedge clk)
    if (_01037_)
      if (mem_do_wdata) mem_instr <= 1'h0;
      else mem_instr <= _07458_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_addr */
  always_ff @(posedge clk)
    if (_01039_) mem_addr <= mem_la_addr;
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME cached_insn_opcode */
  always_ff @(posedge clk)
    if (decoder_trigger_q) cached_insn_opcode <= _00062_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_valid */
  always_ff @(posedge clk)
    if (_01041_) mem_valid <= _00024_;
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME cached_insn_rs2 */
  always_ff @(posedge clk)
    if (decoder_trigger_q) cached_insn_rs2 <= decoded_rs2;
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME cached_insn_rs1 */
  always_ff @(posedge clk)
    if (decoder_trigger_q) cached_insn_rs1 <= decoded_rs1;
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_valid_insn */
  always_ff @(posedge clk)
    if (_06888_) dbg_valid_insn <= 1'h0;
    else if (launch_next_insn) dbg_valid_insn <= 1'h1;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_compare */
  always_ff @(posedge clk)
    if (_01072_) is_compare <= 1'h0;
    else is_compare <= _07573_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_alu_reg_reg */
  always_ff @(posedge clk)
    if (_05738_) is_alu_reg_reg <= _07324_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_alu_reg_imm */
  always_ff @(posedge clk)
    if (_05738_) is_alu_reg_imm <= _07340_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_fence */
  always_ff @(posedge clk)
    if (!resetn) instr_fence <= 1'h0;
    else if (_06685_) instr_fence <= _06805_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_ecall_ebreak */
  always_ff @(posedge clk)
    if (_06685_) instr_ecall_ebreak <= _06897_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_beq_bne_blt_bge_bltu_bgeu */
  always_ff @(posedge clk)
    if (!resetn) is_beq_bne_blt_bge_bltu_bgeu <= 1'h0;
    else if (_05738_) is_beq_bne_blt_bge_bltu_bgeu <= _07346_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_sll_srl_sra */
  always_ff @(posedge clk)
    if (_06685_) is_sll_srl_sra <= _06817_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_sb_sh_sw */
  always_ff @(posedge clk)
    if (_05738_) is_sb_sh_sw <= _07352_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_jalr_addi_slti_sltiu_xori_ori_andi */
  always_ff @(posedge clk)
    if (_06685_) is_jalr_addi_slti_sltiu_xori_ori_andi <= _06899_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_slli_srli_srai */
  always_ff @(posedge clk)
    if (_06685_) is_slli_srli_srai <= _06813_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_lb_lh_lw_lbu_lhu */
  always_ff @(posedge clk)
    if (_05738_) is_lb_lh_lw_lbu_lhu <= _07360_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME compressed_instr */
  always_ff @(posedge clk)
    if (_05738_) compressed_instr <= _07362_;
  reg \decoded_imm_j_reg[10] ;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_reg[10]  */
  always_ff @(posedge clk)
    if (_05738_) \decoded_imm_j_reg[10]  <= _07276_;
  assign decoded_imm_j[10] = \decoded_imm_j_reg[10] ;
  reg \decoded_imm_j_reg[7] ;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_reg[7]  */
  always_ff @(posedge clk)
    if (_05738_) \decoded_imm_j_reg[7]  <= _07278_;
  assign decoded_imm_j[7] = \decoded_imm_j_reg[7] ;
  reg \decoded_imm_j_reg[6] ;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_reg[6]  */
  always_ff @(posedge clk)
    if (_05738_) \decoded_imm_j_reg[6]  <= _07280_;
  assign decoded_imm_j[6] = \decoded_imm_j_reg[6] ;
  reg [2:0] _09402_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME _09402_ */
  always_ff @(posedge clk)
    if (_05738_) _09402_ <= _07282_;
  assign decoded_imm_j[3:1] = _09402_;
  reg \decoded_imm_j_reg[5] ;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_reg[5]  */
  always_ff @(posedge clk)
    if (_05738_) \decoded_imm_j_reg[5]  <= _07284_;
  assign decoded_imm_j[5] = \decoded_imm_j_reg[5] ;
  reg [1:0] _09404_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME _09404_ */
  always_ff @(posedge clk)
    if (_05738_) _09404_ <= _07286_;
  assign decoded_imm_j[9:8] = _09404_;
  reg [11:0] _09405_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME _09405_ */
  always_ff @(posedge clk)
    if (_05738_) _09405_ <= _07288_;
  assign decoded_imm_j[31:20] = _09405_;
  reg \decoded_imm_j_reg[4] ;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_reg[4]  */
  always_ff @(posedge clk)
    if (_05738_) \decoded_imm_j_reg[4]  <= _07290_;
  assign decoded_imm_j[4] = \decoded_imm_j_reg[4] ;
  reg \decoded_imm_j_reg[11] ;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_reg[11]  */
  always_ff @(posedge clk)
    if (_05738_) \decoded_imm_j_reg[11]  <= _07292_;
  assign decoded_imm_j[11] = \decoded_imm_j_reg[11] ;
  reg [7:0] _09408_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME _09408_ */
  always_ff @(posedge clk)
    if (_05738_) _09408_ <= _07378_;
  assign decoded_imm_j[19:12] = _09408_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_imm */
  always_ff @(posedge clk)
    if (_06685_) decoded_imm <= _06333_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_rs2 */
  always_ff @(posedge clk)
    if (_05738_) decoded_rs2 <= _07376_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME trap */
  always_ff @(posedge clk)
    if (!resetn) trap <= 1'h0;
    else trap <= _07142_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_wdata */
  always_ff @(posedge clk)
    if (_00971_)
      if (mem_instr) rvfi_mem_wdata <= 32'd0;
      else rvfi_mem_wdata <= _07098_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_wdata */
  always_ff @(posedge clk)
    if (_01043_) mem_wdata <= mem_la_wdata;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_rs1[4] */
  always_ff @(posedge clk)
    if (_05738_) decoded_rs1[4] <= _07274_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_rs1[3:0] */
  always_ff @(posedge clk)
    if (_05738_) decoded_rs1[3:0] <= _07312_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_rd */
  always_ff @(posedge clk)
    if (_05738_) decoded_rd <= _07399_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_rdinstrh */
  always_ff @(posedge clk)
    if (_06685_) instr_rdinstrh <= _06799_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_rdinstr */
  always_ff @(posedge clk)
    if (_06685_) instr_rdinstr <= _06795_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_rdcycleh */
  always_ff @(posedge clk)
    if (_06685_) instr_rdcycleh <= _06791_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_rdcycle */
  always_ff @(posedge clk)
    if (_06685_) instr_rdcycle <= _06781_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_and */
  always_ff @(posedge clk)
    if (!resetn) instr_and <= 1'h0;
    else if (_06685_) instr_and <= _06771_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_or */
  always_ff @(posedge clk)
    if (!resetn) instr_or <= 1'h0;
    else if (_06685_) instr_or <= _06767_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sra */
  always_ff @(posedge clk)
    if (!resetn) instr_sra <= 1'h0;
    else if (_06685_) instr_sra <= _06763_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_srl */
  always_ff @(posedge clk)
    if (!resetn) instr_srl <= 1'h0;
    else if (_06685_) instr_srl <= _06761_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_xor */
  always_ff @(posedge clk)
    if (!resetn) instr_xor <= 1'h0;
    else if (_06685_) instr_xor <= _06757_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sltu */
  always_ff @(posedge clk)
    if (!resetn) instr_sltu <= 1'h0;
    else if (_06685_) instr_sltu <= _06753_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_slt */
  always_ff @(posedge clk)
    if (!resetn) instr_slt <= 1'h0;
    else if (_06685_) instr_slt <= _06749_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sub */
  always_ff @(posedge clk)
    if (!resetn) instr_sub <= 1'h0;
    else if (_06685_) instr_sub <= _06741_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_add */
  always_ff @(posedge clk)
    if (!resetn) instr_add <= 1'h0;
    else if (_06685_) instr_add <= _06739_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_srai */
  always_ff @(posedge clk)
    if (_06685_) instr_srai <= _06735_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_srli */
  always_ff @(posedge clk)
    if (_06685_) instr_srli <= _06733_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_slli */
  always_ff @(posedge clk)
    if (_06685_) instr_slli <= _06729_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_andi */
  always_ff @(posedge clk)
    if (!resetn) instr_andi <= 1'h0;
    else if (_06685_) instr_andi <= _06725_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_ori */
  always_ff @(posedge clk)
    if (!resetn) instr_ori <= 1'h0;
    else if (_06685_) instr_ori <= _06723_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_xori */
  always_ff @(posedge clk)
    if (!resetn) instr_xori <= 1'h0;
    else if (_06685_) instr_xori <= _06721_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sltiu */
  always_ff @(posedge clk)
    if (!resetn) instr_sltiu <= 1'h0;
    else if (_06685_) instr_sltiu <= _06719_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_slti */
  always_ff @(posedge clk)
    if (!resetn) instr_slti <= 1'h0;
    else if (_06685_) instr_slti <= _06717_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_addi */
  always_ff @(posedge clk)
    if (!resetn) instr_addi <= 1'h0;
    else if (_06685_) instr_addi <= _06715_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sw */
  always_ff @(posedge clk)
    if (_06685_) instr_sw <= _06713_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sh */
  always_ff @(posedge clk)
    if (_06685_) instr_sh <= _06711_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sb */
  always_ff @(posedge clk)
    if (_06685_) instr_sb <= _06709_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lhu */
  always_ff @(posedge clk)
    if (_06685_) instr_lhu <= _06707_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lbu */
  always_ff @(posedge clk)
    if (_06685_) instr_lbu <= _06705_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lw */
  always_ff @(posedge clk)
    if (_06685_) instr_lw <= _06703_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lh */
  always_ff @(posedge clk)
    if (_06685_) instr_lh <= _06701_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lb */
  always_ff @(posedge clk)
    if (_06685_) instr_lb <= _06699_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_bgeu */
  always_ff @(posedge clk)
    if (!resetn) instr_bgeu <= 1'h0;
    else if (_06685_) instr_bgeu <= _06697_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_bltu */
  always_ff @(posedge clk)
    if (!resetn) instr_bltu <= 1'h0;
    else if (_06685_) instr_bltu <= _06695_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_bge */
  always_ff @(posedge clk)
    if (!resetn) instr_bge <= 1'h0;
    else if (_06685_) instr_bge <= _06693_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_blt */
  always_ff @(posedge clk)
    if (!resetn) instr_blt <= 1'h0;
    else if (_06685_) instr_blt <= _06691_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_bne */
  always_ff @(posedge clk)
    if (!resetn) instr_bne <= 1'h0;
    else if (_06685_) instr_bne <= _06689_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_beq */
  always_ff @(posedge clk)
    if (!resetn) instr_beq <= 1'h0;
    else if (_06685_) instr_beq <= _06687_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_jalr */
  always_ff @(posedge clk)
    if (_05738_) instr_jalr <= _07409_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_jal */
  always_ff @(posedge clk)
    if (_05738_) instr_jal <= _07417_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_auipc */
  always_ff @(posedge clk)
    if (_05738_) instr_auipc <= _06541_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lui */
  always_ff @(posedge clk)
    if (_05738_) instr_lui <= _07427_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_insn */
  always_ff @(posedge clk)
    if (_06685_) pcpi_insn <= mem_rdata_q;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_timeout */
  always_ff @(posedge clk)
    if (!resetn) pcpi_timeout <= 1'h0;
    else pcpi_timeout <= _06829_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_timeout_counter */
  always_ff @(posedge clk)
    if (!_06607_) pcpi_timeout_counter <= 4'hf;
    else if (_07143_) pcpi_timeout_counter <= _07585_[3:0];
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_rd */
  always_ff @(posedge clk)
    if (_01045_) latched_rd <= _06138_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_is_lb */
  always_ff @(posedge clk)
    if (!resetn) latched_is_lb <= 1'h0;
    else if (_01047_) latched_is_lb <= _06140_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_is_lh */
  always_ff @(posedge clk)
    if (!resetn) latched_is_lh <= 1'h0;
    else if (_01047_) latched_is_lh <= _06142_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_compr */
  always_ff @(posedge clk)
    if (_01049_) latched_compr <= compressed_instr;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_branch */
  always_ff @(posedge clk)
    if (!resetn) latched_branch <= 1'h0;
    else if (_00975_) latched_branch <= _06144_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_stalu */
  always_ff @(posedge clk)
    if (!resetn) latched_stalu <= 1'h0;
    else if (_01051_) latched_stalu <= _06146_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_store */
  always_ff @(posedge clk)
    if (!resetn) latched_store <= 1'h0;
    else if (_01053_) latched_store <= _06154_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME count_cycle */
  always_ff @(posedge clk)
    if (!resetn) count_cycle <= 64'h0000000000000000;
    else count_cycle <= _00088_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME reg_pc */
  always_ff @(posedge clk)
    if (!resetn) reg_pc <= 32'd2147483648;
    else if (_06485_) reg_pc <= _00060_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME reg_next_pc */
  always_ff @(posedge clk)
    if (!resetn) reg_next_pc <= 32'd2147483648;
    else if (_06485_) reg_next_pc <= _07232_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_wmask */
  always_ff @(posedge clk)
    if (_00971_)
      if (mem_instr) rvfi_mem_wmask <= 4'h0;
      else rvfi_mem_wmask <= _07102_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_rmask */
  always_ff @(posedge clk)
    if (_00971_)
      if (mem_instr) rvfi_mem_rmask <= 4'h0;
      else rvfi_mem_rmask <= _07104_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_do_wdata */
  always_ff @(posedge clk)
    if (_00034_) mem_do_wdata <= 1'h1;
    else if (_06872_) mem_do_wdata <= 1'h0;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_do_rdata */
  always_ff @(posedge clk)
    if (_00032_) mem_do_rdata <= 1'h1;
    else if (_06872_) mem_do_rdata <= 1'h0;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_do_rinst */
  always_ff @(posedge clk)
    if (_00033_) mem_do_rinst <= 1'h1;
    else if (_01055_) mem_do_rinst <= _07209_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_rs2 */
  always_ff @(posedge clk)
    if (_01057_) pcpi_rs2 <= _06224_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_rs1[31] */
  always_ff @(posedge clk)
    if (_01059_) pcpi_rs1[31] <= _06234_[31];
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_rs1[30:0] */
  always_ff @(posedge clk)
    if (_01061_) pcpi_rs1[30:0] <= _06234_[30:0];
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_rdata */
  always_ff @(posedge clk)
    if (_00971_)
      if (mem_instr) rvfi_mem_rdata <= 32'd0;
      else rvfi_mem_rdata <= _07100_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_wordsize */
  always_ff @(posedge clk)
    if (_01063_) mem_wordsize <= _06220_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sll */
  always_ff @(posedge clk)
    if (!resetn) instr_sll <= 1'h0;
    else if (_06685_) instr_sll <= _06745_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_addr */
  always_ff @(posedge clk)
    if (_00971_)
      if (mem_instr) rvfi_mem_addr <= 32'd0;
      else rvfi_mem_addr <= _07106_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rd_wdata */
  always_ff @(posedge clk)
    if (_01073_) rvfi_rd_wdata <= 32'd0;
    else if (_01025_) rvfi_rd_wdata <= _07109_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rd_addr */
  always_ff @(posedge clk)
    if (_01073_) rvfi_rd_addr <= 5'h00;
    else if (_01025_) rvfi_rd_addr <= _07113_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rs2_rdata */
  always_ff @(posedge clk)
    if (!dbg_rs2val_valid) rvfi_rs2_rdata <= 32'd0;
    else rvfi_rs2_rdata <= dbg_rs2val;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rs1_rdata */
  always_ff @(posedge clk)
    if (_01074_) rvfi_rs1_rdata <= 32'd0;
    else rvfi_rs1_rdata <= dbg_rs1val;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rs2_addr */
  always_ff @(posedge clk)
    if (!dbg_rs2val_valid) rvfi_rs2_addr <= 5'h00;
    else rvfi_rs2_addr <= dbg_insn_rs2;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rs1_addr */
  always_ff @(posedge clk)
    if (_01074_) rvfi_rs1_addr <= 5'h00;
    else rvfi_rs1_addr <= dbg_insn_rs1;
  reg [7:0] _09488_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME _09488_ */
  always_ff @(posedge clk)
    if (dbg_next) _09488_ <= { dbg_insn_opcode[24:20], dbg_insn_opcode[14:12] };
  assign { rvfi_insn[24:20], rvfi_insn[14:12] } = _09488_;
  reg [23:0] _09489_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME _09489_ */
  always_ff @(posedge clk)
    _09489_ <= { dbg_insn_opcode[31:25], dbg_insn_opcode[19:15], dbg_insn_opcode[11:0] };
  assign { rvfi_insn[31:25], rvfi_insn[19:15], rvfi_insn[11:0] } = _09489_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_order */
  always_ff @(posedge clk)
    if (!resetn) rvfi_order <= 64'h0000000000000000;
    else rvfi_order <= _00100_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME cpu_state */
  always_ff @(posedge clk)
    if (_06624_) cpu_state <= 8'h80;
    else cpu_state <= _07185_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_do_prefetch */
  always_ff @(posedge clk)
    if (_06872_) mem_do_prefetch <= 1'h0;
    else if (_01065_) mem_do_prefetch <= _06610_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoder_pseudo_trigger */
  always_ff @(posedge clk)
    if (!_01075_) decoder_pseudo_trigger <= 1'h0;
    else decoder_pseudo_trigger <= _07119_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME count_instr */
  always_ff @(posedge clk)
    if (!resetn) count_instr <= 64'h0000000000000000;
    else if (_01067_) count_instr <= _00092_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_valid */
  always_ff @(posedge clk)
    if (!resetn) pcpi_valid <= 1'h0;
    else if (_01069_) pcpi_valid <= _07238_;
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_pc_wdata[0] */
  always_ff @(posedge clk)
    if (launch_next_insn)
      if (_06599_) rvfi_pc_wdata[0] <= 1'h0;
      else rvfi_pc_wdata[0] <= reg_next_pc[0];
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_pc_wdata[31:1] */
  always_ff @(posedge clk)
    if (launch_next_insn) rvfi_pc_wdata[31:1] <= next_pc[31:1];
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[9]  */
  always_ff @(posedge clk)
    if (_07083_) \cpuregs[9]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[8]  */
  always_ff @(posedge clk)
    if (_07081_) \cpuregs[8]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[7]  */
  always_ff @(posedge clk)
    if (_07079_) \cpuregs[7]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[6]  */
  always_ff @(posedge clk)
    if (_07077_) \cpuregs[6]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[5]  */
  always_ff @(posedge clk)
    if (_07075_) \cpuregs[5]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[4]  */
  always_ff @(posedge clk)
    if (_07073_) \cpuregs[4]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[3]  */
  always_ff @(posedge clk)
    if (_07071_) \cpuregs[3]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[31]  */
  always_ff @(posedge clk)
    if (_07069_) \cpuregs[31]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[30]  */
  always_ff @(posedge clk)
    if (_07067_) \cpuregs[30]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[2]  */
  always_ff @(posedge clk)
    if (_07065_) \cpuregs[2]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[29]  */
  always_ff @(posedge clk)
    if (_07063_) \cpuregs[29]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[28]  */
  always_ff @(posedge clk)
    if (_07061_) \cpuregs[28]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[27]  */
  always_ff @(posedge clk)
    if (_07059_) \cpuregs[27]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[26]  */
  always_ff @(posedge clk)
    if (_07057_) \cpuregs[26]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[25]  */
  always_ff @(posedge clk)
    if (_07055_) \cpuregs[25]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[24]  */
  always_ff @(posedge clk)
    if (_07053_) \cpuregs[24]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[23]  */
  always_ff @(posedge clk)
    if (_07051_) \cpuregs[23]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[22]  */
  always_ff @(posedge clk)
    if (_07049_) \cpuregs[22]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[21]  */
  always_ff @(posedge clk)
    if (_07047_) \cpuregs[21]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[20]  */
  always_ff @(posedge clk)
    if (_07045_) \cpuregs[20]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[1]  */
  always_ff @(posedge clk)
    if (_07043_) \cpuregs[1]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[19]  */
  always_ff @(posedge clk)
    if (_07041_) \cpuregs[19]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[18]  */
  always_ff @(posedge clk)
    if (_07039_) \cpuregs[18]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[17]  */
  always_ff @(posedge clk)
    if (_07037_) \cpuregs[17]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[16]  */
  always_ff @(posedge clk)
    if (_07035_) \cpuregs[16]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[15]  */
  always_ff @(posedge clk)
    if (_07033_) \cpuregs[15]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[14]  */
  always_ff @(posedge clk)
    if (_07031_) \cpuregs[14]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[13]  */
  always_ff @(posedge clk)
    if (_07029_) \cpuregs[13]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[12]  */
  always_ff @(posedge clk)
    if (_07027_) \cpuregs[12]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[11]  */
  always_ff @(posedge clk)
    if (_07025_) \cpuregs[11]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[10]  */
  always_ff @(posedge clk)
    if (_07023_) \cpuregs[10]  <= _00002_;
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[0]  */
  always_ff @(posedge clk)
    if (_07021_) \cpuregs[0]  <= _00002_;
  assign _06102_ = _05738_ ? _07376_ : decoded_rs2;
  assign _06104_ = _05738_ ? { _07274_, _07312_ } : decoded_rs1;
  assign _04481_ = { 26'h0000000, reg_sh } | { 26'h0000000, reg_sh_t0 };
  assign _00937_ = { 1'h0, _02103_ } >= 32'd4;
  assign _00938_ = { 1'h0, _04481_ } >= 32'd4;
  assign _06598_ = _00937_ ^ _00938_;
  assign _00273_ = ~ { 26'h0000000, reg_sh_t0 };
  assign _02103_ = { 26'h0000000, reg_sh } & _00273_;
  assign _02104_ = latched_store_t0 & latched_branch;
  assign _02110_ = _06486_ & decoder_trigger;
  assign _02113_ = mem_do_rinst_t0 & mem_done;
  assign _02116_ = latched_store_t0 & _06827_;
  assign _02117_ = is_lb_lh_lw_lbu_lhu_t0 & _06831_;
  assign _02120_ = mem_do_prefetch_t0 & mem_done;
  assign _02123_ = _06502_ & _07087_;
  assign _02126_ = _06504_ & pcpi_rs1[0];
  assign _02129_ = _06626_ & dbg_valid_insn;
  assign _02132_ = mem_valid_t0 & mem_ready;
  assign _02135_ = rvfi_valid_t0 & _06505_;
  assign _02138_ = _06630_ & _06507_;
  assign _02141_ = _06634_ & next_pc[1];
  assign _02144_ = _06636_ & _06833_;
  assign _02147_ = mem_la_firstword_t0 & prefetched_high_word;
  assign _02150_ = _06638_ & _06834_;
  assign _02153_ = mem_la_use_prefetched_high_word_t0 & mem_do_rinst;
  assign _02156_ = mem_xfer_t0 & _07572_;
  assign _02159_ = _06642_ & _06878_;
  assign _02162_ = _07562_ & mem_do_rinst;
  assign _02165_ = _06822_ & mem_xfer;
  assign _02168_ = _06648_ & _06882_;
  assign _02171_ = _06652_ & mem_do_wdata;
  assign _02174_ = mem_la_use_prefetched_high_word_t0 & _06836_;
  assign _02177_ = _06654_ & _06884_;
  assign _02180_ = mem_xfer_t0 & _07559_;
  assign _02183_ = mem_la_firstword_xfer_t0 & _06833_;
  assign _02186_ = _06658_ & _07563_;
  assign _02189_ = mem_valid_t0 & _06839_;
  assign _02190_ = mem_done_t0 & _06633_;
  assign _02193_ = mem_rdata_latched_t0[12] & _06533_;
  assign _02196_ = _06546_ & _06547_;
  assign _02199_ = mem_rdata_latched_t0[11] & _06841_;
  assign _02202_ = mem_rdata_latched_t0[12] & _07090_;
  assign _02205_ = _06682_ & _06533_;
  assign _02208_ = mem_rdata_latched_t0[12] & _07089_;
  assign _02210_ = _06670_ & _06533_;
  assign _02214_ = decoder_trigger_t0 & _06842_;
  assign _02217_ = is_beq_bne_blt_bge_bltu_bgeu_t0 & _06559_;
  assign _02220_ = is_beq_bne_blt_bge_bltu_bgeu_t0 & _06561_;
  assign _02223_ = is_beq_bne_blt_bge_bltu_bgeu_t0 & _06563_;
  assign _02226_ = is_beq_bne_blt_bge_bltu_bgeu_t0 & _06565_;
  assign _02229_ = is_beq_bne_blt_bge_bltu_bgeu_t0 & _06567_;
  assign _02232_ = is_beq_bne_blt_bge_bltu_bgeu_t0 & _06569_;
  assign _02235_ = is_lb_lh_lw_lbu_lhu_t0 & _06559_;
  assign _02238_ = is_lb_lh_lw_lbu_lhu_t0 & _06561_;
  assign _02241_ = is_lb_lh_lw_lbu_lhu_t0 & _06571_;
  assign _02244_ = is_lb_lh_lw_lbu_lhu_t0 & _06563_;
  assign _02247_ = is_lb_lh_lw_lbu_lhu_t0 & _06565_;
  assign _02250_ = is_sb_sh_sw_t0 & _06559_;
  assign _02253_ = is_sb_sh_sw_t0 & _06561_;
  assign _02256_ = is_sb_sh_sw_t0 & _06571_;
  assign _02259_ = is_alu_reg_imm_t0 & _06559_;
  assign _02262_ = is_alu_reg_imm_t0 & _06571_;
  assign _02265_ = is_alu_reg_imm_t0 & _06573_;
  assign _02268_ = is_alu_reg_imm_t0 & _06563_;
  assign _02271_ = is_alu_reg_imm_t0 & _06567_;
  assign _02274_ = is_alu_reg_imm_t0 & _06569_;
  assign _02277_ = is_alu_reg_imm_t0 & _06561_;
  assign _02280_ = _06728_ & _06575_;
  assign _02283_ = _06732_ & _06575_;
  assign _02286_ = is_alu_reg_imm_t0 & _06565_;
  assign _02289_ = _06732_ & _06577_;
  assign _02292_ = _06738_ & _06575_;
  assign _02295_ = is_alu_reg_reg_t0 & _06559_;
  assign _02298_ = _06738_ & _06577_;
  assign _02301_ = is_alu_reg_reg_t0 & _06561_;
  assign _02304_ = _06744_ & _06575_;
  assign _02307_ = is_alu_reg_reg_t0 & _06571_;
  assign _02310_ = _06748_ & _06575_;
  assign _02313_ = is_alu_reg_reg_t0 & _06573_;
  assign _02316_ = _06752_ & _06575_;
  assign _02319_ = is_alu_reg_reg_t0 & _06563_;
  assign _02322_ = _06756_ & _06575_;
  assign _02325_ = _06760_ & _06575_;
  assign _02328_ = is_alu_reg_reg_t0 & _06565_;
  assign _02331_ = _06760_ & _06577_;
  assign _02334_ = is_alu_reg_reg_t0 & _06567_;
  assign _02337_ = _06766_ & _06575_;
  assign _02340_ = is_alu_reg_reg_t0 & _06569_;
  assign _02343_ = _06770_ & _06575_;
  assign _02346_ = _06580_ & _06581_;
  assign _02349_ = _06774_ & _07092_;
  assign _02352_ = _06580_ & _06583_;
  assign _02355_ = _06778_ & _07092_;
  assign _02358_ = _06580_ & _06585_;
  assign _02361_ = _06784_ & _07092_;
  assign _02364_ = _06580_ & _06587_;
  assign _02367_ = _06788_ & _07092_;
  assign _02370_ = _06580_ & _06589_;
  assign _02373_ = _06794_ & _07092_;
  assign _02376_ = _06580_ & _06591_;
  assign _02379_ = _06798_ & _07092_;
  assign _02382_ = _06580_ & _06843_;
  assign _02385_ = _06802_ & _06845_;
  assign _02388_ = _06596_ & _06847_;
  assign _02391_ = is_alu_reg_imm_t0 & _07577_;
  assign _02394_ = is_alu_reg_imm_t0 & _07579_;
  assign _02397_ = _06566_ & _06577_;
  assign _02400_ = _06566_ & _06575_;
  assign _02403_ = _06562_ & _06575_;
  assign _02406_ = is_alu_reg_reg_t0 & _07577_;
  assign _02105_ = latched_branch_t0 & latched_store;
  assign _06604_ = cpuregs_write_t0 & resetn;
  assign _02111_ = decoder_trigger_t0 & _06485_;
  assign _02114_ = mem_done_t0 & mem_do_rinst;
  assign _02118_ = instr_trap_t0 & is_lb_lh_lw_lbu_lhu;
  assign _02121_ = mem_done_t0 & _06832_;
  assign _06618_ = _06871_ & resetn;
  assign _02124_ = _07088_ & _06501_;
  assign _02127_ = pcpi_rs1_t0[0] & _06503_;
  assign _06626_ = _06875_ & resetn;
  assign _02130_ = dbg_valid_insn_t0 & _06625_;
  assign _02133_ = mem_ready_t0 & mem_valid;
  assign _02136_ = _06506_ & rvfi_valid;
  assign _02139_ = _06508_ & _06629_;
  assign _02142_ = next_pc_t0[1] & _06633_;
  assign _02145_ = mem_la_secondword_t0 & _06635_;
  assign _02148_ = prefetched_high_word_t0 & mem_la_firstword;
  assign _02151_ = clear_prefetched_high_word_t0 & _06637_;
  assign _02154_ = mem_do_rinst_t0 & mem_la_use_prefetched_high_word;
  assign _02157_ = _06837_ & mem_xfer;
  assign _02160_ = _06879_ & _06641_;
  assign _02163_ = mem_do_rinst_t0 & _07561_;
  assign _06648_ = _06881_ & resetn;
  assign _02166_ = mem_xfer_t0 & _06821_;
  assign _02169_ = _06883_ & _06647_;
  assign _06652_ = _06837_ & resetn;
  assign _02172_ = mem_do_wdata_t0 & _06651_;
  assign _02175_ = _06837_ & _06838_;
  assign _02178_ = _06885_ & _06653_;
  assign _02181_ = _07560_ & mem_xfer;
  assign _02184_ = mem_la_secondword_t0 & mem_la_firstword_xfer;
  assign _02187_ = _06822_ & _06657_;
  assign mem_la_read_t0 = _06887_ & resetn;
  assign _02191_ = _06634_ & mem_done;
  assign _02194_ = _06534_ & _00704_;
  assign _02197_ = _06548_ & _06545_;
  assign _02200_ = mem_rdata_latched_t0[12] & _06840_;
  assign _02203_ = _07091_ & _00704_;
  assign _02206_ = _06534_ & _06681_;
  assign _02209_ = _07091_ & mem_rdata_latched[12];
  assign _02211_ = _06534_ & _06669_;
  assign _02213_ = _06534_ & mem_rdata_latched[12];
  assign _02215_ = decoder_pseudo_trigger_t0 & decoder_trigger;
  assign _02218_ = _06560_ & is_beq_bne_blt_bge_bltu_bgeu;
  assign _02221_ = _06562_ & is_beq_bne_blt_bge_bltu_bgeu;
  assign _02224_ = _06564_ & is_beq_bne_blt_bge_bltu_bgeu;
  assign _02227_ = _06566_ & is_beq_bne_blt_bge_bltu_bgeu;
  assign _02230_ = _06568_ & is_beq_bne_blt_bge_bltu_bgeu;
  assign _02233_ = _06570_ & is_beq_bne_blt_bge_bltu_bgeu;
  assign _02236_ = _06560_ & is_lb_lh_lw_lbu_lhu;
  assign _02239_ = _06562_ & is_lb_lh_lw_lbu_lhu;
  assign _02242_ = _06572_ & is_lb_lh_lw_lbu_lhu;
  assign _02245_ = _06564_ & is_lb_lh_lw_lbu_lhu;
  assign _02248_ = _06566_ & is_lb_lh_lw_lbu_lhu;
  assign _02251_ = _06560_ & is_sb_sh_sw;
  assign _02254_ = _06562_ & is_sb_sh_sw;
  assign _02257_ = _06572_ & is_sb_sh_sw;
  assign _02260_ = _06560_ & is_alu_reg_imm;
  assign _02263_ = _06572_ & is_alu_reg_imm;
  assign _02266_ = _06574_ & is_alu_reg_imm;
  assign _02269_ = _06564_ & is_alu_reg_imm;
  assign _02272_ = _06568_ & is_alu_reg_imm;
  assign _02275_ = _06570_ & is_alu_reg_imm;
  assign _02278_ = _06562_ & is_alu_reg_imm;
  assign _02281_ = _06576_ & _06727_;
  assign _02284_ = _06576_ & _06731_;
  assign _02287_ = _06566_ & is_alu_reg_imm;
  assign _02290_ = _06578_ & _06731_;
  assign _02293_ = _06576_ & _06737_;
  assign _02296_ = _06560_ & is_alu_reg_reg;
  assign _02299_ = _06578_ & _06737_;
  assign _02302_ = _06562_ & is_alu_reg_reg;
  assign _02305_ = _06576_ & _06743_;
  assign _02308_ = _06572_ & is_alu_reg_reg;
  assign _02311_ = _06576_ & _06747_;
  assign _02314_ = _06574_ & is_alu_reg_reg;
  assign _02317_ = _06576_ & _06751_;
  assign _02320_ = _06564_ & is_alu_reg_reg;
  assign _02323_ = _06576_ & _06755_;
  assign _02326_ = _06576_ & _06759_;
  assign _02329_ = _06566_ & is_alu_reg_reg;
  assign _02332_ = _06578_ & _06759_;
  assign _02335_ = _06568_ & is_alu_reg_reg;
  assign _02338_ = _06576_ & _06765_;
  assign _02341_ = _06570_ & is_alu_reg_reg;
  assign _02344_ = _06576_ & _06769_;
  assign _02347_ = _06582_ & _06579_;
  assign _02350_ = _07093_ & _06773_;
  assign _02353_ = _06584_ & _06579_;
  assign _02356_ = _07093_ & _06777_;
  assign _02359_ = _06586_ & _06579_;
  assign _02362_ = _07093_ & _06783_;
  assign _02365_ = _06588_ & _06579_;
  assign _02368_ = _07093_ & _06787_;
  assign _02371_ = _06590_ & _06579_;
  assign _02374_ = _07093_ & _06793_;
  assign _02377_ = _06592_ & _06579_;
  assign _02380_ = _07093_ & _06797_;
  assign _02383_ = _06844_ & _06579_;
  assign _02386_ = _06846_ & _06801_;
  assign _02389_ = _06848_ & _06595_;
  assign _02392_ = _07578_ & is_alu_reg_imm;
  assign _02395_ = _07580_ & is_alu_reg_imm;
  assign _02398_ = _06578_ & _06565_;
  assign _02401_ = _06576_ & _06565_;
  assign _02404_ = _06576_ & _06561_;
  assign _02407_ = _07578_ & is_alu_reg_reg;
  assign _02106_ = latched_store_t0 & latched_branch_t0;
  assign _02112_ = _06486_ & decoder_trigger_t0;
  assign _02115_ = mem_do_rinst_t0 & mem_done_t0;
  assign _02119_ = is_lb_lh_lw_lbu_lhu_t0 & instr_trap_t0;
  assign _02122_ = mem_do_prefetch_t0 & mem_done_t0;
  assign _02125_ = _06502_ & _07088_;
  assign _02128_ = _06504_ & pcpi_rs1_t0[0];
  assign _02131_ = _06626_ & dbg_valid_insn_t0;
  assign _02134_ = mem_valid_t0 & mem_ready_t0;
  assign _02137_ = rvfi_valid_t0 & _06506_;
  assign _02140_ = _06630_ & _06508_;
  assign _02143_ = _06634_ & next_pc_t0[1];
  assign _02146_ = _06636_ & mem_la_secondword_t0;
  assign _02149_ = mem_la_firstword_t0 & prefetched_high_word_t0;
  assign _02152_ = _06638_ & clear_prefetched_high_word_t0;
  assign _02155_ = mem_la_use_prefetched_high_word_t0 & mem_do_rinst_t0;
  assign _02158_ = mem_xfer_t0 & _06837_;
  assign _02161_ = _06642_ & _06879_;
  assign _02164_ = _07562_ & mem_do_rinst_t0;
  assign _02167_ = _06822_ & mem_xfer_t0;
  assign _02170_ = _06648_ & _06883_;
  assign _02173_ = _06652_ & mem_do_wdata_t0;
  assign _02176_ = mem_la_use_prefetched_high_word_t0 & _06837_;
  assign _02179_ = _06654_ & _06885_;
  assign _02182_ = mem_xfer_t0 & _07560_;
  assign _02185_ = mem_la_firstword_xfer_t0 & mem_la_secondword_t0;
  assign _02188_ = _06658_ & _06822_;
  assign _02192_ = mem_done_t0 & _06634_;
  assign _02195_ = mem_rdata_latched_t0[12] & _06534_;
  assign _02198_ = _06546_ & _06548_;
  assign _02201_ = mem_rdata_latched_t0[11] & mem_rdata_latched_t0[12];
  assign _02204_ = mem_rdata_latched_t0[12] & _07091_;
  assign _02207_ = _06682_ & _06534_;
  assign _02212_ = _06670_ & _06534_;
  assign _02216_ = decoder_trigger_t0 & decoder_pseudo_trigger_t0;
  assign _02219_ = is_beq_bne_blt_bge_bltu_bgeu_t0 & _06560_;
  assign _02222_ = is_beq_bne_blt_bge_bltu_bgeu_t0 & _06562_;
  assign _02225_ = is_beq_bne_blt_bge_bltu_bgeu_t0 & _06564_;
  assign _02228_ = is_beq_bne_blt_bge_bltu_bgeu_t0 & _06566_;
  assign _02231_ = is_beq_bne_blt_bge_bltu_bgeu_t0 & _06568_;
  assign _02234_ = is_beq_bne_blt_bge_bltu_bgeu_t0 & _06570_;
  assign _02237_ = is_lb_lh_lw_lbu_lhu_t0 & _06560_;
  assign _02240_ = is_lb_lh_lw_lbu_lhu_t0 & _06562_;
  assign _02243_ = is_lb_lh_lw_lbu_lhu_t0 & _06572_;
  assign _02246_ = is_lb_lh_lw_lbu_lhu_t0 & _06564_;
  assign _02249_ = is_lb_lh_lw_lbu_lhu_t0 & _06566_;
  assign _02252_ = is_sb_sh_sw_t0 & _06560_;
  assign _02255_ = is_sb_sh_sw_t0 & _06562_;
  assign _02258_ = is_sb_sh_sw_t0 & _06572_;
  assign _02261_ = is_alu_reg_imm_t0 & _06560_;
  assign _02264_ = is_alu_reg_imm_t0 & _06572_;
  assign _02267_ = is_alu_reg_imm_t0 & _06574_;
  assign _02270_ = is_alu_reg_imm_t0 & _06564_;
  assign _02273_ = is_alu_reg_imm_t0 & _06568_;
  assign _02276_ = is_alu_reg_imm_t0 & _06570_;
  assign _02279_ = is_alu_reg_imm_t0 & _06562_;
  assign _02282_ = _06728_ & _06576_;
  assign _02285_ = _06732_ & _06576_;
  assign _02288_ = is_alu_reg_imm_t0 & _06566_;
  assign _02291_ = _06732_ & _06578_;
  assign _02294_ = _06738_ & _06576_;
  assign _02297_ = is_alu_reg_reg_t0 & _06560_;
  assign _02300_ = _06738_ & _06578_;
  assign _02303_ = is_alu_reg_reg_t0 & _06562_;
  assign _02306_ = _06744_ & _06576_;
  assign _02309_ = is_alu_reg_reg_t0 & _06572_;
  assign _02312_ = _06748_ & _06576_;
  assign _02315_ = is_alu_reg_reg_t0 & _06574_;
  assign _02318_ = _06752_ & _06576_;
  assign _02321_ = is_alu_reg_reg_t0 & _06564_;
  assign _02324_ = _06756_ & _06576_;
  assign _02327_ = _06760_ & _06576_;
  assign _02330_ = is_alu_reg_reg_t0 & _06566_;
  assign _02333_ = _06760_ & _06578_;
  assign _02336_ = is_alu_reg_reg_t0 & _06568_;
  assign _02339_ = _06766_ & _06576_;
  assign _02342_ = is_alu_reg_reg_t0 & _06570_;
  assign _02345_ = _06770_ & _06576_;
  assign _02348_ = _06580_ & _06582_;
  assign _02351_ = _06774_ & _07093_;
  assign _02354_ = _06580_ & _06584_;
  assign _02357_ = _06778_ & _07093_;
  assign _02360_ = _06580_ & _06586_;
  assign _02363_ = _06784_ & _07093_;
  assign _02366_ = _06580_ & _06588_;
  assign _02369_ = _06788_ & _07093_;
  assign _02372_ = _06580_ & _06590_;
  assign _02375_ = _06794_ & _07093_;
  assign _02378_ = _06580_ & _06592_;
  assign _02381_ = _06798_ & _07093_;
  assign _02384_ = _06580_ & _06844_;
  assign _02387_ = _06802_ & _06846_;
  assign _02390_ = _06596_ & _06848_;
  assign _02393_ = is_alu_reg_imm_t0 & _07578_;
  assign _02396_ = is_alu_reg_imm_t0 & _07580_;
  assign _02399_ = _06566_ & _06578_;
  assign _02402_ = _06566_ & _06576_;
  assign _02405_ = _06562_ & _06576_;
  assign _02408_ = is_alu_reg_reg_t0 & _07578_;
  assign _04482_ = _02104_ | _02105_;
  assign _04484_ = _02110_ | _02111_;
  assign _04485_ = _02113_ | _02114_;
  assign _04486_ = _02116_ | _02105_;
  assign _04487_ = _02117_ | _02118_;
  assign _04488_ = _02120_ | _02121_;
  assign _04489_ = _02123_ | _02124_;
  assign _04490_ = _02126_ | _02127_;
  assign _04491_ = _02129_ | _02130_;
  assign _04492_ = _02132_ | _02133_;
  assign _04493_ = _02135_ | _02136_;
  assign _04494_ = _02138_ | _02139_;
  assign _04495_ = _02141_ | _02142_;
  assign _04496_ = _02144_ | _02145_;
  assign _04497_ = _02147_ | _02148_;
  assign _04498_ = _02150_ | _02151_;
  assign _04499_ = _02153_ | _02154_;
  assign _04500_ = _02156_ | _02157_;
  assign _04501_ = _02159_ | _02160_;
  assign _04502_ = _02162_ | _02163_;
  assign _04503_ = _02165_ | _02166_;
  assign _04504_ = _02168_ | _02169_;
  assign _04505_ = _02171_ | _02172_;
  assign _04506_ = _02174_ | _02175_;
  assign _04507_ = _02177_ | _02178_;
  assign _04508_ = _02180_ | _02181_;
  assign _04509_ = _02183_ | _02184_;
  assign _04510_ = _02186_ | _02187_;
  assign _04511_ = _02189_ | _02133_;
  assign _04512_ = _02190_ | _02191_;
  assign _04513_ = _02193_ | _02194_;
  assign _04514_ = _02196_ | _02197_;
  assign _04515_ = _02199_ | _02200_;
  assign _04516_ = _02202_ | _02203_;
  assign _04517_ = _02205_ | _02206_;
  assign _04518_ = _02208_ | _02194_;
  assign _04519_ = _02202_ | _02209_;
  assign _04520_ = _02210_ | _02211_;
  assign _04521_ = _02208_ | _02213_;
  assign _04522_ = _02214_ | _02215_;
  assign _04523_ = _02217_ | _02218_;
  assign _04524_ = _02220_ | _02221_;
  assign _04525_ = _02223_ | _02224_;
  assign _04526_ = _02226_ | _02227_;
  assign _04527_ = _02229_ | _02230_;
  assign _04528_ = _02232_ | _02233_;
  assign _04529_ = _02235_ | _02236_;
  assign _04530_ = _02238_ | _02239_;
  assign _04531_ = _02241_ | _02242_;
  assign _04532_ = _02244_ | _02245_;
  assign _04533_ = _02247_ | _02248_;
  assign _04534_ = _02250_ | _02251_;
  assign _04535_ = _02253_ | _02254_;
  assign _04536_ = _02256_ | _02257_;
  assign _04537_ = _02259_ | _02260_;
  assign _04538_ = _02262_ | _02263_;
  assign _04539_ = _02265_ | _02266_;
  assign _04540_ = _02268_ | _02269_;
  assign _04541_ = _02271_ | _02272_;
  assign _04542_ = _02274_ | _02275_;
  assign _04543_ = _02277_ | _02278_;
  assign _04544_ = _02280_ | _02281_;
  assign _04545_ = _02283_ | _02284_;
  assign _04546_ = _02286_ | _02287_;
  assign _04547_ = _02289_ | _02290_;
  assign _04548_ = _02292_ | _02293_;
  assign _04549_ = _02295_ | _02296_;
  assign _04550_ = _02298_ | _02299_;
  assign _04551_ = _02301_ | _02302_;
  assign _04552_ = _02304_ | _02305_;
  assign _04553_ = _02307_ | _02308_;
  assign _04554_ = _02310_ | _02311_;
  assign _04555_ = _02313_ | _02314_;
  assign _04556_ = _02316_ | _02317_;
  assign _04557_ = _02319_ | _02320_;
  assign _04558_ = _02322_ | _02323_;
  assign _04559_ = _02325_ | _02326_;
  assign _04560_ = _02328_ | _02329_;
  assign _04561_ = _02331_ | _02332_;
  assign _04562_ = _02334_ | _02335_;
  assign _04563_ = _02337_ | _02338_;
  assign _04564_ = _02340_ | _02341_;
  assign _04565_ = _02343_ | _02344_;
  assign _04566_ = _02346_ | _02347_;
  assign _04567_ = _02349_ | _02350_;
  assign _04568_ = _02352_ | _02353_;
  assign _04569_ = _02355_ | _02356_;
  assign _04570_ = _02358_ | _02359_;
  assign _04571_ = _02361_ | _02362_;
  assign _04572_ = _02364_ | _02365_;
  assign _04573_ = _02367_ | _02368_;
  assign _04574_ = _02370_ | _02371_;
  assign _04575_ = _02373_ | _02374_;
  assign _04576_ = _02376_ | _02377_;
  assign _04577_ = _02379_ | _02380_;
  assign _04578_ = _02382_ | _02383_;
  assign _04579_ = _02385_ | _02386_;
  assign _04580_ = _02388_ | _02389_;
  assign _04581_ = _02391_ | _02392_;
  assign _04582_ = _02394_ | _02395_;
  assign _04583_ = _02397_ | _02398_;
  assign _04584_ = _02400_ | _02401_;
  assign _04585_ = _02403_ | _02404_;
  assign _04586_ = _02406_ | _02407_;
  assign _06600_ = _04482_ | _02106_;
  assign launch_next_insn_t0 = _04484_ | _02112_;
  assign _06608_ = _04485_ | _02115_;
  assign _06602_ = _04486_ | _02106_;
  assign _06614_ = _04487_ | _02119_;
  assign _06616_ = _04488_ | _02122_;
  assign _06620_ = _04489_ | _02125_;
  assign _06622_ = _04490_ | _02128_;
  assign _00031_ = _04491_ | _02131_;
  assign _06628_ = _04492_ | _02134_;
  assign _06630_ = _04493_ | _02137_;
  assign _06632_ = _04494_ | _02140_;
  assign _06636_ = _04495_ | _02143_;
  assign mem_la_firstword_t0 = _04496_ | _02146_;
  assign _06638_ = _04497_ | _02149_;
  assign mem_la_use_prefetched_high_word_t0 = _04498_ | _02152_;
  assign _06640_ = _04499_ | _02155_;
  assign _06642_ = _04500_ | _02158_;
  assign _06644_ = _04501_ | _02161_;
  assign _06646_ = _04502_ | _02164_;
  assign _06650_ = _04503_ | _02167_;
  assign mem_done_t0 = _04504_ | _02170_;
  assign mem_la_write_t0 = _04505_ | _02173_;
  assign _06654_ = _04506_ | _02176_;
  assign _06656_ = _04507_ | _02179_;
  assign mem_la_firstword_xfer_t0 = _04508_ | _02182_;
  assign _06658_ = _04509_ | _02185_;
  assign _06660_ = _04510_ | _02188_;
  assign _06662_ = _04511_ | _02134_;
  assign _06664_ = _04512_ | _02192_;
  assign _06666_ = _04513_ | _02195_;
  assign _06676_ = _04514_ | _02198_;
  assign _06680_ = _04515_ | _02201_;
  assign _06682_ = _04516_ | _02204_;
  assign _06684_ = _04517_ | _02207_;
  assign _06668_ = _04518_ | _02195_;
  assign _06670_ = _04519_ | _02204_;
  assign _06672_ = _04520_ | _02212_;
  assign _06674_ = _04521_ | _02195_;
  assign _06686_ = _04522_ | _02216_;
  assign _06688_ = _04523_ | _02219_;
  assign _06690_ = _04524_ | _02222_;
  assign _06692_ = _04525_ | _02225_;
  assign _06694_ = _04526_ | _02228_;
  assign _06696_ = _04527_ | _02231_;
  assign _06698_ = _04528_ | _02234_;
  assign _06700_ = _04529_ | _02237_;
  assign _06702_ = _04530_ | _02240_;
  assign _06704_ = _04531_ | _02243_;
  assign _06706_ = _04532_ | _02246_;
  assign _06708_ = _04533_ | _02249_;
  assign _06710_ = _04534_ | _02252_;
  assign _06712_ = _04535_ | _02255_;
  assign _06714_ = _04536_ | _02258_;
  assign _06716_ = _04537_ | _02261_;
  assign _06718_ = _04538_ | _02264_;
  assign _06720_ = _04539_ | _02267_;
  assign _06722_ = _04540_ | _02270_;
  assign _06724_ = _04541_ | _02273_;
  assign _06726_ = _04542_ | _02276_;
  assign _06728_ = _04543_ | _02279_;
  assign _06730_ = _04544_ | _02282_;
  assign _06734_ = _04545_ | _02285_;
  assign _06732_ = _04546_ | _02288_;
  assign _06736_ = _04547_ | _02291_;
  assign _06740_ = _04548_ | _02294_;
  assign _06738_ = _04549_ | _02297_;
  assign _06742_ = _04550_ | _02300_;
  assign _06744_ = _04551_ | _02303_;
  assign _06746_ = _04552_ | _02306_;
  assign _06748_ = _04553_ | _02309_;
  assign _06750_ = _04554_ | _02312_;
  assign _06752_ = _04555_ | _02315_;
  assign _06754_ = _04556_ | _02318_;
  assign _06756_ = _04557_ | _02321_;
  assign _06758_ = _04558_ | _02324_;
  assign _06762_ = _04559_ | _02327_;
  assign _06760_ = _04560_ | _02330_;
  assign _06764_ = _04561_ | _02333_;
  assign _06766_ = _04562_ | _02336_;
  assign _06768_ = _04563_ | _02339_;
  assign _06770_ = _04564_ | _02342_;
  assign _06772_ = _04565_ | _02345_;
  assign _06774_ = _04566_ | _02348_;
  assign _06776_ = _04567_ | _02351_;
  assign _06778_ = _04568_ | _02354_;
  assign _06780_ = _04569_ | _02357_;
  assign _06784_ = _04570_ | _02360_;
  assign _06786_ = _04571_ | _02363_;
  assign _06788_ = _04572_ | _02366_;
  assign _06790_ = _04573_ | _02369_;
  assign _06794_ = _04574_ | _02372_;
  assign _06796_ = _04575_ | _02375_;
  assign _06798_ = _04576_ | _02378_;
  assign _06800_ = _04577_ | _02381_;
  assign _06802_ = _04578_ | _02384_;
  assign _06804_ = _04579_ | _02387_;
  assign _06806_ = _04580_ | _02390_;
  assign _06814_ = _04581_ | _02393_;
  assign _06816_ = _04582_ | _02396_;
  assign _06808_ = _04583_ | _02399_;
  assign _06810_ = _04584_ | _02402_;
  assign _06812_ = _04585_ | _02405_;
  assign _06818_ = _04586_ | _02408_;
  assign _00274_ = ~ _06604_;
  assign _00275_ = ~ latched_rd_t0;
  assign _00276_ = _06603_ & _00274_;
  assign _00277_ = _06603_ | _06604_;
  assign _02107_ = latched_rd & _00275_;
  assign _04483_ = latched_rd | latched_rd_t0;
  assign _00278_ = | _02107_;
  assign _00279_ = | _04483_;
  assign _02108_ = _00276_ & _00278_;
  assign _02109_ = _00277_ & _00279_;
  assign _00005_[31] = _02108_ ^ _02109_;
  assign _00280_ = | { _06894_, mem_do_rdata_t0, mem_la_read_t0 };
  assign _00281_ = | { _00797_, _06536_, _07440_, _06837_, _06538_ };
  assign _00282_ = | { _06885_, mem_do_wdata_t0 };
  assign _00283_ = | { _00797_, _06536_, _07440_, _06837_ };
  assign _00284_ = | { _06488_, _06490_ };
  assign _00285_ = | { _06628_, mem_instr_t0 };
  assign _00286_ = | { _06492_, _06486_ };
  assign _00287_ = | { _06498_, _06486_ };
  assign _00288_ = | { _01083_, _06492_, _06488_, _06490_, _06486_ };
  assign _00289_ = | { _06496_, _06494_, _06498_, _06488_ };
  assign _00290_ = | { _06496_, _06498_, _06486_ };
  assign _00291_ = | { cpuregs_write_t0, rvfi_valid_t0 };
  assign _00292_ = | { is_lui_auipc_jal_t0, is_jalr_addi_slti_sltiu_xori_ori_andi_t0 };
  assign _00293_ = | { _06494_, _06498_ };
  assign _00294_ = | { is_lui_auipc_jal_t0, _06614_, instr_rdcycle_t0, instr_rdcycleh_t0, instr_rdinstr_t0, instr_rdinstrh_t0, is_jalr_addi_slti_sltiu_xori_ori_andi_t0 };
  assign _00295_ = | { _06362_[0], _07414_ };
  assign _00296_ = | { _07271_, _07255_ };
  assign _00297_ = | { _06427_[0], _07255_ };
  assign _00298_ = | { _06427_[0], _06303_[1], _07266_, _07271_, _07255_ };
  assign _00299_ = | { instr_rdcycle_t0, instr_rdcycleh_t0, instr_rdinstr_t0, instr_rdinstrh_t0, is_slli_srli_srai_t0 };
  assign _00300_ = | { _06602_, latched_branch_t0 };
  assign _00301_ = | { _06614_, instr_rdcycle_t0, instr_rdcycleh_t0, instr_rdinstr_t0, instr_rdinstrh_t0, is_slli_srli_srai_t0 };
  assign _00302_ = | { _06496_, _06498_ };
  assign _00303_ = | { is_lui_auipc_jal_t0, _06614_, instr_rdcycle_t0, instr_rdcycleh_t0, instr_rdinstr_t0, instr_rdinstrh_t0, is_jalr_addi_slti_sltiu_xori_ori_andi_t0, is_slli_srli_srai_t0 };
  assign _00304_ = | { is_lui_auipc_jal_t0, instr_rdcycle_t0, instr_rdcycleh_t0, instr_rdinstr_t0, instr_rdinstrh_t0 };
  assign _00305_ = | { _07273_, _07252_ };
  assign _00306_ = | { _06303_[1], _07271_ };
  assign _00307_ = | { _06303_[1], _07271_, _07255_ };
  assign _00308_ = | { pcpi_div_ready_t0, pcpi_mul_ready_t0 };
  assign _00309_ = | { _06496_, _06494_, _06498_, _06492_ };
  assign _00310_ = | { is_lui_auipc_jal_t0, _06614_, is_jalr_addi_slti_sltiu_xori_ori_andi_t0, is_slli_srli_srai_t0 };
  assign _00311_ = | { is_sltiu_bltu_sltu_t0, is_slti_blt_slt_t0, instr_bgeu_t0 };
  assign _00312_ = | { instr_jalr_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_sb_sh_sw_t0, is_lb_lh_lw_lbu_lhu_t0, is_alu_reg_imm_t0 };
  assign _00313_ = | reg_sh_t0;
  assign _00210_ = | mem_rdata_latched_t0[11:10];
  assign _00211_ = | mem_rdata_latched_t0[6:5];
  assign _00314_ = | mem_rdata_latched_t0[14:12];
  assign _00315_ = | mem_rdata_latched_t0[6:2];
  assign _00218_ = | mem_rdata_q_t0[14:12];
  assign _00219_ = | mem_rdata_q_t0[31:25];
  assign _00316_ = | pcpi_timeout_counter_t0;
  assign _00317_ = | { instr_sll_t0, instr_lui_t0, instr_auipc_t0, instr_jal_t0, instr_jalr_t0, instr_beq_t0, instr_bne_t0, instr_blt_t0, instr_bge_t0, instr_bltu_t0, instr_bgeu_t0, instr_lb_t0, instr_lh_t0, instr_lw_t0, instr_lbu_t0, instr_lhu_t0, instr_sb_t0, instr_sh_t0, instr_sw_t0, instr_addi_t0, instr_slti_t0, instr_sltiu_t0, instr_xori_t0, instr_ori_t0, instr_andi_t0, instr_slli_t0, instr_srli_t0, instr_srai_t0, instr_add_t0, instr_sub_t0, instr_slt_t0, instr_sltu_t0, instr_xor_t0, instr_srl_t0, instr_sra_t0, instr_or_t0, instr_and_t0, instr_rdcycle_t0, instr_rdcycleh_t0, instr_rdinstr_t0, instr_rdinstrh_t0, instr_fence_t0 };
  assign _00318_ = | mem_rdata_q_t0[31:21];
  assign _00319_ = | mem_rdata_q_t0[19:7];
  assign _00320_ = | mem_rdata_q_t0[15:12];
  assign _00224_ = | pcpi_rs1_t0[1:0];
  assign _00213_ = | mem_rdata_latched_t0[11:7];
  assign _00321_ = | mem_rdata_q_t0[13:12];
  assign _00222_ = | mem_rdata_latched_t0[15:13];
  assign _00220_ = | mem_rdata_latched_t0[1:0];
  assign _00223_ = | mem_state_t0;
  assign _00225_ = | mem_wordsize_t0;
  assign _00322_ = | decoded_rs1_t0;
  assign _00323_ = | decoded_rs2_t0;
  assign _00324_ = | latched_rd_t0;
  assign _00325_ = | mem_wstrb_t0;
  assign _00326_ = | { instr_lui_t0, instr_auipc_t0 };
  assign _00327_ = | { instr_rdcycle_t0, instr_rdcycleh_t0, instr_rdinstr_t0, instr_rdinstrh_t0 };
  assign _00328_ = | { instr_lui_t0, instr_auipc_t0, instr_jal_t0 };
  assign _00329_ = | { instr_blt_t0, instr_slti_t0, instr_slt_t0 };
  assign _00330_ = | { instr_bltu_t0, instr_sltiu_t0, instr_sltu_t0 };
  assign _00331_ = | { instr_slti_t0, instr_sltiu_t0, instr_slt_t0, instr_sltu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0 };
  assign _00332_ = | mem_rdata_latched_t0[12:5];
  assign _00333_ = | { _06560_, _06572_, _06574_, _06564_, _06568_, _06570_ };
  assign _00334_ = | { _06812_, _06810_, _06808_ };
  assign _00335_ = ~ { _06894_, mem_la_read_t0, mem_do_rdata_t0 };
  assign _00336_ = ~ { _06837_, _06536_, _06538_, _07440_, _00797_ };
  assign _00337_ = ~ { _06885_, mem_do_wdata_t0 };
  assign _00338_ = ~ { _06837_, _06536_, _07440_, _00797_ };
  assign _00339_ = ~ { _06488_, _06490_ };
  assign _00340_ = ~ { _06628_, mem_instr_t0 };
  assign _00341_ = ~ { _06486_, _06492_ };
  assign _00342_ = ~ { _06486_, _06498_ };
  assign _00343_ = ~ { _06488_, _06490_, _06486_, _06492_, _01083_ };
  assign _00344_ = ~ { _06873_, 1'h0 };
  assign _00345_ = ~ { _06488_, _06494_, _06496_, _06498_ };
  assign _00346_ = ~ { _06486_, _06496_, _06498_ };
  assign _00347_ = ~ { cpuregs_write_t0, rvfi_valid_t0 };
  assign _00348_ = ~ { is_jalr_addi_slti_sltiu_xori_ori_andi_t0, is_lui_auipc_jal_t0 };
  assign _00349_ = ~ { _06498_, _06494_ };
  assign _00350_ = ~ { _06614_, is_jalr_addi_slti_sltiu_xori_ori_andi_t0, is_lui_auipc_jal_t0, instr_rdinstrh_t0, instr_rdinstr_t0, instr_rdcycleh_t0, instr_rdcycle_t0 };
  assign _00351_ = ~ { _07414_, _06362_[0] };
  assign _00352_ = ~ { _07271_, _07255_ };
  assign _00353_ = ~ { _07255_, _06427_[0] };
  assign _00354_ = ~ { _07271_, _07266_, _07255_, _06427_[0], _06303_[1] };
  assign _00355_ = ~ { is_slli_srli_srai_t0, instr_rdinstrh_t0, instr_rdinstr_t0, instr_rdcycleh_t0, instr_rdcycle_t0 };
  assign _00356_ = ~ { _06602_, latched_branch_t0 };
  assign _00357_ = ~ { _06614_, is_slli_srli_srai_t0, instr_rdinstrh_t0, instr_rdinstr_t0, instr_rdcycleh_t0, instr_rdcycle_t0 };
  assign _00358_ = ~ { _06498_, _06496_ };
  assign _00359_ = ~ { _06490_, _06488_ };
  assign _00360_ = ~ { _06614_, is_jalr_addi_slti_sltiu_xori_ori_andi_t0, is_slli_srli_srai_t0, is_lui_auipc_jal_t0, instr_rdinstrh_t0, instr_rdinstr_t0, instr_rdcycleh_t0, instr_rdcycle_t0 };
  assign _00361_ = ~ { is_lui_auipc_jal_t0, instr_rdinstrh_t0, instr_rdinstr_t0, instr_rdcycleh_t0, instr_rdcycle_t0 };
  assign _00362_ = ~ { _07273_, _07252_ };
  assign _00363_ = ~ { _07271_, _06303_[1] };
  assign _00364_ = ~ { _07271_, _07255_, _06303_[1] };
  assign _00365_ = ~ { pcpi_div_ready_t0, pcpi_mul_ready_t0 };
  assign _00366_ = ~ { _06498_, _06496_, _06494_, _06492_ };
  assign _00367_ = ~ { _06614_, is_jalr_addi_slti_sltiu_xori_ori_andi_t0, is_slli_srli_srai_t0, is_lui_auipc_jal_t0 };
  assign _00368_ = ~ { is_sltiu_bltu_sltu_t0, is_slti_blt_slt_t0, instr_bgeu_t0 };
  assign _00369_ = ~ { is_alu_reg_imm_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_sb_sh_sw_t0, is_lb_lh_lw_lbu_lhu_t0, instr_jalr_t0 };
  assign _00370_ = ~ reg_sh_t0;
  assign _00371_ = ~ mem_rdata_latched_t0[14:12];
  assign _00372_ = ~ mem_rdata_latched_t0[6:2];
  assign _00373_ = ~ pcpi_timeout_counter_t0;
  assign _00374_ = ~ { instr_lui_t0, instr_auipc_t0, instr_jal_t0, instr_jalr_t0, instr_beq_t0, instr_bne_t0, instr_blt_t0, instr_bge_t0, instr_bltu_t0, instr_bgeu_t0, instr_lb_t0, instr_lh_t0, instr_lw_t0, instr_lbu_t0, instr_lhu_t0, instr_sb_t0, instr_sh_t0, instr_sw_t0, instr_addi_t0, instr_slti_t0, instr_sltiu_t0, instr_xori_t0, instr_ori_t0, instr_andi_t0, instr_slli_t0, instr_srli_t0, instr_srai_t0, instr_add_t0, instr_sub_t0, instr_sll_t0, instr_slt_t0, instr_sltu_t0, instr_xor_t0, instr_srl_t0, instr_sra_t0, instr_or_t0, instr_and_t0, instr_rdcycle_t0, instr_rdcycleh_t0, instr_rdinstr_t0, instr_rdinstrh_t0, instr_fence_t0, 6'h00 };
  assign _00375_ = ~ mem_rdata_q_t0[31:21];
  assign _00376_ = ~ mem_rdata_q_t0[19:7];
  assign _00377_ = ~ mem_rdata_q_t0[15:12];
  assign _00378_ = ~ mem_rdata_q_t0[13:12];
  assign _00379_ = ~ decoded_rs1_t0;
  assign _00380_ = ~ decoded_rs2_t0;
  assign _00381_ = ~ mem_wstrb_t0;
  assign _00382_ = ~ { instr_auipc_t0, instr_lui_t0 };
  assign _00383_ = ~ { instr_rdinstrh_t0, instr_rdinstr_t0, instr_rdcycleh_t0, instr_rdcycle_t0 };
  assign _00384_ = ~ { instr_jal_t0, instr_auipc_t0, instr_lui_t0 };
  assign _00385_ = ~ { instr_slt_t0, instr_slti_t0, instr_blt_t0 };
  assign _00386_ = ~ { instr_sltu_t0, instr_sltiu_t0, instr_bltu_t0 };
  assign _00387_ = ~ { is_beq_bne_blt_bge_bltu_bgeu_t0, instr_sltu_t0, instr_slt_t0, instr_sltiu_t0, instr_slti_t0 };
  assign _00388_ = ~ mem_rdata_latched_t0[12:5];
  assign _00389_ = ~ { _06574_, _06572_, _06570_, _06568_, _06564_, _06560_ };
  assign _00390_ = ~ { _06812_, _06810_, _06808_ };
  assign _01455_ = { _06893_, mem_la_read, mem_do_rdata } & _00335_;
  assign _01464_ = { _06836_, _06535_, _06537_, _07439_, _06888_ } & _00336_;
  assign _01465_ = { _06884_, mem_do_wdata } & _00337_;
  assign _01467_ = { _06836_, _06535_, _07439_, _06888_ } & _00338_;
  assign _01468_ = { _06487_, _06489_ } & _00339_;
  assign _01469_ = { _06627_, mem_instr } & _00340_;
  assign _01471_ = { _06485_, _06491_ } & _00341_;
  assign _01474_ = { _06485_, _06497_ } & _00342_;
  assign _01477_ = { _06487_, _06489_, _06485_, _06491_, _01082_ } & _00343_;
  assign _01478_ = { _06872_, resetn } & _00344_;
  assign _01489_ = { _06487_, _06493_, _06495_, _06497_ } & _00345_;
  assign _01492_ = { _06485_, _06495_, _06497_ } & _00346_;
  assign _01493_ = { cpuregs_write, rvfi_valid } & _00347_;
  assign _01495_ = { is_jalr_addi_slti_sltiu_xori_ori_andi, is_lui_auipc_jal } & _00348_;
  assign _01496_ = { _06497_, _06493_ } & _00349_;
  assign _01497_ = { _06613_, is_jalr_addi_slti_sltiu_xori_ori_andi, is_lui_auipc_jal, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle } & _00350_;
  assign _01498_ = { _07413_, _07397_ } & _00351_;
  assign _01499_ = { _07270_, _07254_ } & _00352_;
  assign _01500_ = { _07254_, _07253_ } & _00353_;
  assign _01501_ = { _07270_, _07265_, _07254_, _07253_, _07250_ } & _00354_;
  assign _01502_ = { is_slli_srli_srai, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle } & _00355_;
  assign _01503_ = { _06601_, latched_branch } & _00356_;
  assign _01504_ = { _06613_, is_slli_srli_srai, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle } & _00357_;
  assign _01505_ = { _06497_, _06495_ } & _00358_;
  assign _01506_ = { _06489_, _06487_ } & _00359_;
  assign _01507_ = { _06613_, is_jalr_addi_slti_sltiu_xori_ori_andi, is_slli_srli_srai, is_lui_auipc_jal, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle } & _00360_;
  assign _01508_ = { is_lui_auipc_jal, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle } & _00361_;
  assign _01509_ = { _07272_, _07251_ } & _00362_;
  assign _01510_ = { _07270_, _07250_ } & _00363_;
  assign _01511_ = { _07270_, _07254_, _07250_ } & _00364_;
  assign _01512_ = { pcpi_div_ready, pcpi_mul_ready } & _00365_;
  assign _01567_ = { _06497_, _06495_, _06493_, _06491_ } & _00366_;
  assign _01568_ = { _06613_, is_jalr_addi_slti_sltiu_xori_ori_andi, is_slli_srli_srai, is_lui_auipc_jal } & _00367_;
  assign _01569_ = { is_sltiu_bltu_sltu, is_slti_blt_slt, instr_bgeu } & _00368_;
  assign _01570_ = { is_alu_reg_imm, is_beq_bne_blt_bge_bltu_bgeu, is_sb_sh_sw, is_lb_lh_lw_lbu_lhu, instr_jalr } & _00369_;
  assign _02087_ = reg_sh & _00370_;
  assign _02094_ = mem_rdata_latched[14:12] & _00371_;
  assign _02097_ = mem_rdata_latched[6:2] & _00372_;
  assign _02409_ = pcpi_timeout_counter & _00373_;
  assign _02410_ = { instr_lui, instr_auipc, instr_jal, instr_jalr, instr_beq, instr_bne, instr_blt, instr_bge, instr_bltu, instr_bgeu, instr_lb, instr_lh, instr_lw, instr_lbu, instr_lhu, instr_sb, instr_sh, instr_sw, instr_addi, instr_slti, instr_sltiu, instr_xori, instr_ori, instr_andi, instr_slli, instr_srli, instr_srai, instr_add, instr_sub, instr_sll, instr_slt, instr_sltu, instr_xor, instr_srl, instr_sra, instr_or, instr_and, instr_rdcycle, instr_rdcycleh, instr_rdinstr, instr_rdinstrh, instr_fence, 6'h00 } & _00374_;
  assign _02411_ = mem_rdata_q[31:21] & _00375_;
  assign _02412_ = mem_rdata_q[19:7] & _00376_;
  assign _02413_ = mem_rdata_q[15:12] & _00377_;
  assign _02779_ = mem_rdata_q[13:12] & _00378_;
  assign _03309_ = decoded_rs1 & _00379_;
  assign _03310_ = decoded_rs2 & _00380_;
  assign _03311_ = mem_wstrb & _00381_;
  assign _03312_ = { instr_auipc, instr_lui } & _00382_;
  assign _03313_ = { instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle } & _00383_;
  assign _03314_ = { instr_jal, instr_auipc, instr_lui } & _00384_;
  assign _03315_ = { instr_slt, instr_slti, instr_blt } & _00385_;
  assign _03316_ = { instr_sltu, instr_sltiu, instr_bltu } & _00386_;
  assign _03317_ = { is_beq_bne_blt_bge_bltu_bgeu, instr_sltu, instr_slt, instr_sltiu, instr_slti } & _00387_;
  assign _03318_ = mem_rdata_latched[12:5] & _00388_;
  assign _03319_ = { _06573_, _06571_, _06569_, _06567_, _06563_, _06559_ } & _00389_;
  assign _03320_ = { _06811_, _06809_, _06807_ } & _00390_;
  assign _00391_ = ! _01455_;
  assign _00392_ = ! _01464_;
  assign _00393_ = ! _01465_;
  assign _00394_ = ! _01467_;
  assign _00395_ = ! _01468_;
  assign _00396_ = ! _01469_;
  assign _00397_ = ! _01471_;
  assign _00398_ = ! _01474_;
  assign _00399_ = ! _01477_;
  assign _00400_ = ! _01478_;
  assign _00401_ = ! _01489_;
  assign _00402_ = ! _01492_;
  assign _00403_ = ! _01493_;
  assign _00404_ = ! _01495_;
  assign _00405_ = ! _01496_;
  assign _00406_ = ! _01497_;
  assign _00407_ = ! _01498_;
  assign _00408_ = ! _01499_;
  assign _00409_ = ! _01500_;
  assign _00410_ = ! _01501_;
  assign _00411_ = ! _01502_;
  assign _00412_ = ! _01503_;
  assign _00413_ = ! _01504_;
  assign _00414_ = ! _01505_;
  assign _00415_ = ! _01506_;
  assign _00416_ = ! _01507_;
  assign _00417_ = ! _01508_;
  assign _00418_ = ! _01509_;
  assign _00419_ = ! _01510_;
  assign _00420_ = ! _01511_;
  assign _00421_ = ! _01512_;
  assign _00422_ = ! _01567_;
  assign _00423_ = ! _01568_;
  assign _00424_ = ! _01569_;
  assign _00425_ = ! _01570_;
  assign _00426_ = ! _02087_;
  assign _00427_ = ! _02091_;
  assign _00428_ = ! _02092_;
  assign _00429_ = ! _02094_;
  assign _00430_ = ! _02097_;
  assign _00431_ = ! _02101_;
  assign _00432_ = ! _02102_;
  assign _00433_ = ! _02409_;
  assign _00434_ = ! _02410_;
  assign _00435_ = ! _02411_;
  assign _00436_ = ! _02412_;
  assign _00437_ = ! _02413_;
  assign _00438_ = ! _02777_;
  assign _00439_ = ! _02095_;
  assign _00440_ = ! _02779_;
  assign _00441_ = ! _03043_;
  assign _00442_ = ! _02778_;
  assign _00443_ = ! _03135_;
  assign _00444_ = ! _03291_;
  assign _00445_ = ! _03309_;
  assign _00446_ = ! _03310_;
  assign _00447_ = ! _02107_;
  assign _00448_ = ! _03311_;
  assign _00449_ = ! _03312_;
  assign _00450_ = ! _03313_;
  assign _00451_ = ! _03314_;
  assign _00452_ = ! _03315_;
  assign _00453_ = ! _03316_;
  assign _00454_ = ! _03317_;
  assign _00455_ = ! _03318_;
  assign _00456_ = ! _03319_;
  assign _00457_ = ! _03320_;
  assign _00944_ = _00391_ & _00280_;
  assign _00962_ = _00392_ & _00281_;
  assign _00964_ = _00393_ & _00282_;
  assign _00968_ = _00394_ & _00283_;
  assign _00970_ = _00395_ & _00284_;
  assign _00972_ = _00396_ & _00285_;
  assign _00976_ = _00397_ & _00286_;
  assign _00982_ = _00398_ & _00287_;
  assign _00990_ = _00399_ & _00288_;
  assign _00992_ = _00400_ & _06873_;
  assign _01018_ = _00401_ & _00289_;
  assign _01024_ = _00402_ & _00290_;
  assign _01026_ = _00403_ & _00291_;
  assign _01081_ = _00404_ & _00292_;
  assign _01083_ = _00405_ & _00293_;
  assign _01085_ = _00406_ & _00294_;
  assign _01089_ = _00407_ & _00295_;
  assign _01077_ = _00408_ & _00296_;
  assign _01079_ = _00409_ & _00297_;
  assign _01091_ = _00410_ & _00298_;
  assign _01093_ = _00411_ & _00299_;
  assign _00040_ = _00412_ & _00300_;
  assign _01096_ = _00413_ & _00301_;
  assign _01098_ = _00414_ & _00302_;
  assign _00858_ = _00415_ & _00284_;
  assign _00856_ = _00416_ & _00303_;
  assign _00860_ = _00417_ & _00304_;
  assign _00864_ = _00418_ & _00305_;
  assign _00866_ = _00419_ & _00306_;
  assign _00862_ = _00420_ & _00307_;
  assign pcpi_int_ready_t0 = _00421_ & _00308_;
  assign _00868_ = _00422_ & _00309_;
  assign _00870_ = _00423_ & _00310_;
  assign _00872_ = _00424_ & _00311_;
  assign _00874_ = _00425_ & _00312_;
  assign _06500_ = _00426_ & _00313_;
  assign _06518_ = _00427_ & _00210_;
  assign _06526_ = _00428_ & _00211_;
  assign _06548_ = _00429_ & _00314_;
  assign _06534_ = _00430_ & _00315_;
  assign _06560_ = _00431_ & _00218_;
  assign _06576_ = _00432_ & _00219_;
  assign _06830_ = _00433_ & _00316_;
  assign instr_trap_t0 = _00434_ & _00317_;
  assign _06844_ = _00435_ & _00318_;
  assign _06846_ = _00436_ & _00319_;
  assign _06848_ = _00437_ & _00320_;
  assign _07088_ = _00438_ & _00224_;
  assign _07091_ = _00439_ & _00213_;
  assign _07093_ = _00440_ & _00321_;
  assign _06303_[1] = _00441_ & _00222_;
  assign _07273_ = _00442_ & _00220_;
  assign _06837_ = _00443_ & _00223_;
  assign _06502_ = _00444_ & _00225_;
  assign _07565_ = _00445_ & _00322_;
  assign _07567_ = _00446_ & _00323_;
  assign _07569_ = _00447_ & _00324_;
  assign _07571_ = _00448_ & _00325_;
  assign _07364_ = _00449_ & _00326_;
  assign is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0 = _00450_ & _00327_;
  assign _00015_ = _00451_ & _00328_;
  assign _00017_ = _00452_ & _00329_;
  assign _00019_ = _00453_ & _00330_;
  assign _07574_ = _00454_ & _00331_;
  assign _07576_ = _00455_ & _00332_;
  assign _07580_ = _00456_ & _00333_;
  assign _07578_ = _00457_ & _00334_;
  assign _00458_ = ~ instr_sra;
  assign _00459_ = ~ instr_xori;
  assign _00460_ = ~ instr_ori;
  assign _00461_ = ~ instr_andi;
  assign _00462_ = ~ pcpi_timeout;
  assign _00463_ = ~ instr_slli;
  assign _00464_ = ~ instr_srli;
  assign _00465_ = ~ instr_lb;
  assign _00466_ = ~ instr_lh;
  assign _00467_ = ~ mem_do_rdata;
  assign _00468_ = ~ _06627_;
  assign _00469_ = ~ _06876_;
  assign _00470_ = ~ _06643_;
  assign _00471_ = ~ _06655_;
  assign _00472_ = ~ mem_la_read;
  assign _00473_ = ~ _06633_;
  assign _00474_ = ~ mem_do_prefetch;
  assign _00476_ = ~ mem_do_rinst;
  assign _00477_ = ~ _06775_;
  assign _00478_ = ~ _06785_;
  assign _00479_ = ~ _06803_;
  assign _00480_ = ~ instr_jalr;
  assign _00481_ = ~ instr_srai;
  assign _00482_ = ~ instr_xor;
  assign _00483_ = ~ instr_or;
  assign _00484_ = ~ instr_and;
  assign _00485_ = ~ instr_ecall_ebreak;
  assign _00486_ = ~ instr_sll;
  assign _00487_ = ~ instr_srl;
  assign _00488_ = ~ mem_done;
  assign _00489_ = ~ instr_lbu;
  assign _00490_ = ~ instr_lhu;
  assign _00491_ = ~ mem_do_wdata;
  assign _00492_ = ~ trap;
  assign _00493_ = ~ _06639_;
  assign _00494_ = ~ _06645_;
  assign _00495_ = ~ _06649_;
  assign _00496_ = ~ _06659_;
  assign _00497_ = ~ mem_la_write;
  assign _00498_ = ~ mem_la_secondword;
  assign _00499_ = ~ _06779_;
  assign _00500_ = ~ _06789_;
  assign _00501_ = ~ _06593_;
  assign _00502_ = ~ _06815_;
  assign _02414_ = instr_sra_t0 & _00481_;
  assign _02417_ = instr_xori_t0 & _00482_;
  assign _02420_ = instr_ori_t0 & _00483_;
  assign _02423_ = instr_andi_t0 & _00484_;
  assign _06864_ = _06862_ & resetn;
  assign _02426_ = pcpi_timeout_t0 & _00485_;
  assign _02429_ = instr_slli_t0 & _00486_;
  assign _02432_ = instr_srli_t0 & _00487_;
  assign _02435_ = mem_do_prefetch_t0 & _00488_;
  assign _02437_ = instr_lb_t0 & _00489_;
  assign _02440_ = instr_lh_t0 & _00490_;
  assign _02443_ = mem_do_rdata_t0 & _00491_;
  assign _02446_ = launch_next_insn_t0 & _00492_;
  assign _02449_ = _06628_ & _00493_;
  assign _02452_ = _06877_ & _00491_;
  assign _02455_ = _06644_ & _00494_;
  assign _02458_ = mem_la_firstword_t0 & _00495_;
  assign _02461_ = _06656_ & _00496_;
  assign _02464_ = mem_la_read_t0 & _00497_;
  assign _02467_ = _06634_ & _00467_;
  assign _02470_ = mem_do_prefetch_t0 & _00476_;
  assign _02473_ = _06820_ & _00498_;
  assign _02476_ = mem_do_rinst_t0 & _00467_;
  assign _02479_ = _06776_ & _00499_;
  assign _02482_ = _06786_ & _00500_;
  assign _02485_ = _06804_ & _00501_;
  assign _02488_ = instr_jalr_t0 & _00502_;
  assign _02415_ = instr_srai_t0 & _00458_;
  assign _02418_ = instr_xor_t0 & _00459_;
  assign _02421_ = instr_or_t0 & _00460_;
  assign _02424_ = instr_and_t0 & _00461_;
  assign _02427_ = instr_ecall_ebreak_t0 & _00462_;
  assign _02430_ = instr_sll_t0 & _00463_;
  assign _02433_ = instr_srl_t0 & _00464_;
  assign _02436_ = mem_done_t0 & mem_do_prefetch;
  assign _02438_ = instr_lbu_t0 & _00465_;
  assign _02441_ = instr_lhu_t0 & _00466_;
  assign _02444_ = mem_do_wdata_t0 & _00467_;
  assign _06873_ = mem_done_t0 & resetn;
  assign _02447_ = trap_t0 & _00139_;
  assign _02450_ = _06640_ & _00468_;
  assign _02453_ = mem_do_wdata_t0 & _00469_;
  assign _02456_ = _06646_ & _00470_;
  assign _02459_ = _06650_ & mem_la_firstword;
  assign _02462_ = _06660_ & _00471_;
  assign _06890_ = mem_ready_t0 & resetn;
  assign _02465_ = mem_la_write_t0 & _00472_;
  assign _02468_ = mem_do_rdata_t0 & _00473_;
  assign _02471_ = mem_do_rinst_t0 & _00474_;
  assign _02474_ = mem_la_secondword_t0 & _00475_;
  assign _02477_ = mem_do_rdata_t0 & _00476_;
  assign _00797_ = trap_t0 & resetn;
  assign _02480_ = _06780_ & _00477_;
  assign _02483_ = _06790_ & _00478_;
  assign _02486_ = _06594_ & _00479_;
  assign _02489_ = _06816_ & _00480_;
  assign _02416_ = instr_sra_t0 & instr_srai_t0;
  assign _02419_ = instr_xori_t0 & instr_xor_t0;
  assign _02422_ = instr_ori_t0 & instr_or_t0;
  assign _02425_ = instr_andi_t0 & instr_and_t0;
  assign _02428_ = pcpi_timeout_t0 & instr_ecall_ebreak_t0;
  assign _02431_ = instr_slli_t0 & instr_sll_t0;
  assign _02434_ = instr_srli_t0 & instr_srl_t0;
  assign _02439_ = instr_lb_t0 & instr_lbu_t0;
  assign _02442_ = instr_lh_t0 & instr_lhu_t0;
  assign _02445_ = mem_do_rdata_t0 & mem_do_wdata_t0;
  assign _02448_ = launch_next_insn_t0 & trap_t0;
  assign _02451_ = _06628_ & _06640_;
  assign _02454_ = _06877_ & mem_do_wdata_t0;
  assign _02457_ = _06644_ & _06646_;
  assign _02460_ = mem_la_firstword_t0 & _06650_;
  assign _02463_ = _06656_ & _06660_;
  assign _02466_ = mem_la_read_t0 & mem_la_write_t0;
  assign _02469_ = _06634_ & mem_do_rdata_t0;
  assign _02472_ = mem_do_prefetch_t0 & mem_do_rinst_t0;
  assign _02475_ = _06820_ & mem_la_secondword_t0;
  assign _02478_ = mem_do_rinst_t0 & mem_do_rdata_t0;
  assign _02481_ = _06776_ & _06780_;
  assign _02484_ = _06786_ & _06790_;
  assign _02487_ = _06804_ & _06594_;
  assign _02490_ = instr_jalr_t0 & _06816_;
  assign _04587_ = _02414_ | _02415_;
  assign _04588_ = _02417_ | _02418_;
  assign _04589_ = _02420_ | _02421_;
  assign _04590_ = _02423_ | _02424_;
  assign _04591_ = _02426_ | _02427_;
  assign _04592_ = _02429_ | _02430_;
  assign _04593_ = _02432_ | _02433_;
  assign _04594_ = _02435_ | _02436_;
  assign _04595_ = _02437_ | _02438_;
  assign _04596_ = _02440_ | _02441_;
  assign _04597_ = _02443_ | _02444_;
  assign _04598_ = _02446_ | _02447_;
  assign _04599_ = _02449_ | _02450_;
  assign _04600_ = _02452_ | _02453_;
  assign _04601_ = _02455_ | _02456_;
  assign _04602_ = _02458_ | _02459_;
  assign _04603_ = _02461_ | _02462_;
  assign _04604_ = _02464_ | _02465_;
  assign _04605_ = _02467_ | _02468_;
  assign _04606_ = _02470_ | _02471_;
  assign _04607_ = _02473_ | _02474_;
  assign _04608_ = _02476_ | _02477_;
  assign _04612_ = _02479_ | _02480_;
  assign _04613_ = _02482_ | _02483_;
  assign _04614_ = _02485_ | _02486_;
  assign _04615_ = _02488_ | _02489_;
  assign _06850_ = _04587_ | _02416_;
  assign _06852_ = _04588_ | _02419_;
  assign _06854_ = _04589_ | _02422_;
  assign _06856_ = _04590_ | _02425_;
  assign _06612_ = _04591_ | _02428_;
  assign _06858_ = _04592_ | _02431_;
  assign _06860_ = _04593_ | _02434_;
  assign _06866_ = _04594_ | _02122_;
  assign _06868_ = _04595_ | _02439_;
  assign _06215_[1] = _04596_ | _02442_;
  assign _06871_ = _04597_ | _02445_;
  assign _06875_ = _04598_ | _02448_;
  assign mem_xfer_t0 = _04599_ | _02451_;
  assign _06879_ = _04600_ | _02454_;
  assign _06881_ = _04601_ | _02457_;
  assign _06883_ = _04602_ | _02460_;
  assign _06887_ = _04603_ | _02463_;
  assign _06892_ = _04604_ | _02466_;
  assign _06885_ = _04605_ | _02469_;
  assign _06634_ = _04606_ | _02472_;
  assign _06894_ = _04607_ | _02475_;
  assign _06877_ = _04608_ | _02478_;
  assign _06782_ = _04612_ | _02481_;
  assign _06792_ = _04613_ | _02484_;
  assign _06898_ = _04614_ | _02487_;
  assign _06900_ = _04615_ | _02490_;
  assign _00503_ = ~ latched_branch_t0;
  assign _00504_ = ~ mem_rdata_latched_t0[12];
  assign _00505_ = latched_branch & _00503_;
  assign _00506_ = mem_rdata_latched[12] & _00504_;
  assign _00507_ = latched_branch | latched_branch_t0;
  assign _00508_ = mem_rdata_latched[12] | mem_rdata_latched_t0[12];
  assign _04609_ = mem_rdata_latched[6:2] | mem_rdata_latched_t0[6:2];
  assign _00509_ = | _02097_;
  assign _00510_ = | _04609_;
  assign _04610_ = _00506_ | _00509_;
  assign _04611_ = _00508_ | _00510_;
  assign _06862_ = _00505_ ^ _00507_;
  assign _06896_ = _04610_ ^ _04611_;
  assign _00939_ = $signed({ _04616_, _02493_ }) < $signed({ _02492_, _04619_ });
  assign _00940_ = { _02491_, _02493_ } < { _04617_, _04619_ };
  assign _00941_ = $signed({ _02491_, _04618_ }) < $signed({ _04617_, _02494_ });
  assign _00942_ = { _04616_, _04618_ } < { _02492_, _02494_ };
  assign alu_lts_t0 = _00939_ ^ _00941_;
  assign alu_ltu_t0 = _00940_ ^ _00942_;
  assign _00511_ = ~ pcpi_rs1_t0[30:0];
  assign _00512_ = ~ pcpi_rs1_t0[31];
  assign _00513_ = ~ pcpi_rs2_t0[30:0];
  assign _00514_ = ~ pcpi_rs2_t0[31];
  assign _04616_ = pcpi_rs1[31] | pcpi_rs1_t0[31];
  assign _04617_ = pcpi_rs2[31] | pcpi_rs2_t0[31];
  assign _02491_ = pcpi_rs1[31] & _00512_;
  assign _02492_ = pcpi_rs2[31] & _00514_;
  assign _02493_ = pcpi_rs1[30:0] & _00511_;
  assign _02494_ = pcpi_rs2[30:0] & _00513_;
  assign _04618_ = pcpi_rs1[30:0] | pcpi_rs1_t0[30:0];
  assign _04619_ = pcpi_rs2[30:0] | pcpi_rs2_t0[30:0];
  assign _06065_ = ~ _00000_[0];
  assign _06066_ = ~ _00000_[1];
  assign _06067_ = ~ _00000_[2];
  assign _06068_ = ~ _00000_[3];
  assign _06069_ = ~ _00000_[4];
  assign _03360_ = _06065_ & _06066_;
  assign _03362_ = _06068_ & _06069_;
  assign _03364_ = _06067_ & _03362_;
  assign _03366_ = _03360_ & _03364_;
  assign _03368_ = _00000_[0] & _06066_;
  assign _03370_ = _03368_ & _03364_;
  assign _03372_ = _06065_ & _00000_[1];
  assign _03374_ = _03372_ & _03364_;
  assign _03376_ = _00000_[0] & _00000_[1];
  assign _03378_ = _03376_ & _03364_;
  assign _03380_ = _00000_[2] & _03362_;
  assign _03382_ = _03360_ & _03380_;
  assign _03384_ = _03368_ & _03380_;
  assign _03386_ = _03372_ & _03380_;
  assign _03388_ = _03376_ & _03380_;
  assign _03390_ = _00000_[3] & _06069_;
  assign _03392_ = _06067_ & _03390_;
  assign _03394_ = _03360_ & _03392_;
  assign _03396_ = _03368_ & _03392_;
  assign _03398_ = _03372_ & _03392_;
  assign _03400_ = _03376_ & _03392_;
  assign _03402_ = _00000_[2] & _03390_;
  assign _03404_ = _03360_ & _03402_;
  assign _03406_ = _03368_ & _03402_;
  assign _03408_ = _03372_ & _03402_;
  assign _03410_ = _03376_ & _03402_;
  assign _03412_ = _06068_ & _00000_[4];
  assign _03414_ = _06067_ & _03412_;
  assign _03416_ = _03360_ & _03414_;
  assign _03418_ = _03368_ & _03414_;
  assign _03420_ = _03372_ & _03414_;
  assign _03422_ = _03376_ & _03414_;
  assign _03424_ = _00000_[2] & _03412_;
  assign _03426_ = _03360_ & _03424_;
  assign _03428_ = _03368_ & _03424_;
  assign _03430_ = _03372_ & _03424_;
  assign _03432_ = _03376_ & _03424_;
  assign _03434_ = _00000_[3] & _00000_[4];
  assign _03436_ = _06067_ & _03434_;
  assign _03438_ = _03360_ & _03436_;
  assign _03440_ = _03368_ & _03436_;
  assign _03442_ = _03372_ & _03436_;
  assign _03444_ = _03376_ & _03436_;
  assign _03446_ = _00000_[2] & _03434_;
  assign _03448_ = _03360_ & _03446_;
  assign _03450_ = _03368_ & _03446_;
  assign _03452_ = _03372_ & _03446_;
  assign _03454_ = _03376_ & _03446_;
  assign _00515_ = ~ { _05738_, _05738_, _05738_, _05738_, _05738_ };
  assign _00516_ = ~ _06497_;
  assign _00517_ = ~ _06491_;
  assign _00518_ = ~ _01097_;
  assign _00519_ = ~ { latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh };
  assign _00520_ = ~ { latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb };
  assign _00521_ = ~ { _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_ };
  assign _00522_ = ~ { _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_ };
  assign _00523_ = ~ { _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_ };
  assign _00524_ = ~ { _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_ };
  assign _00525_ = ~ { is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh };
  assign _00526_ = ~ { instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh };
  assign _00527_ = ~ { instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh };
  assign _00528_ = ~ { _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_ };
  assign _00529_ = ~ { _06489_, _06489_, _06489_, _06489_, _06489_ };
  assign _00530_ = ~ { _06493_, _06493_, _06493_, _06493_, _06493_ };
  assign _00531_ = ~ { is_slli_srli_srai, is_slli_srli_srai, is_slli_srli_srai, is_slli_srli_srai, is_slli_srli_srai };
  assign _00532_ = ~ { _01084_, _01084_, _01084_, _01084_, _01084_ };
  assign _00533_ = ~ { _06491_, _06491_, _06491_, _06491_, _06491_ };
  assign _00534_ = ~ _01082_;
  assign _00535_ = ~ _06487_;
  assign _00536_ = ~ _06489_;
  assign _00537_ = ~ _05104_;
  assign _00538_ = ~ is_rdcycle_rdcycleh_rdinstr_rdinstrh;
  assign _00539_ = ~ { _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_ };
  assign _00540_ = ~ { _01097_, _01097_, _01097_, _01097_, _01097_, _01097_, _01097_, _01097_ };
  assign _00541_ = ~ { _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_ };
  assign _00542_ = ~ { _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_ };
  assign _00543_ = ~ { _05106_, _05106_, _05106_, _05106_, _05106_, _05106_, _05106_, _05106_ };
  assign _00544_ = ~ { _00867_, _00867_, _00867_, _00867_, _00867_, _00867_, _00867_, _00867_ };
  assign _00545_ = ~ { is_sll_srl_sra, is_sll_srl_sra, is_sll_srl_sra, is_sll_srl_sra, is_sll_srl_sra, is_sll_srl_sra, is_sll_srl_sra, is_sll_srl_sra };
  assign _00546_ = ~ { instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap };
  assign _00547_ = ~ { _05108_, _05108_, _05108_, _05108_, _05108_, _05108_, _05108_, _05108_ };
  assign _00548_ = ~ { _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_ };
  assign _00549_ = ~ { is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh };
  assign _00550_ = ~ { _00869_, _00869_, _00869_, _00869_, _00869_, _00869_, _00869_, _00869_ };
  assign _00551_ = ~ { _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_ };
  assign _00552_ = ~ _06493_;
  assign _00553_ = ~ _05110_;
  assign _00554_ = ~ is_sll_srl_sra;
  assign _00555_ = ~ instr_trap;
  assign _00556_ = ~ _05108_;
  assign _00557_ = ~ is_sb_sh_sw;
  assign _00558_ = ~ _01080_;
  assign _00559_ = ~ _06613_;
  assign _00560_ = ~ _05112_;
  assign _00561_ = ~ { instr_lw, instr_lw };
  assign _00562_ = ~ { _06497_, _06497_ };
  assign _00563_ = ~ { instr_sw, instr_sw };
  assign _00564_ = ~ { _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_, _01095_ };
  assign _00565_ = ~ { _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_ };
  assign _00566_ = ~ { _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_ };
  assign _00567_ = ~ { _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_ };
  assign _00568_ = ~ { _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_ };
  assign _00569_ = ~ { _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_ };
  assign _00570_ = ~ { is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal };
  assign _00571_ = ~ { _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_ };
  assign _00572_ = ~ { _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_ };
  assign _00573_ = ~ { is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare };
  assign _00574_ = ~ { _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_ };
  assign _00575_ = ~ { _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_ };
  assign _00576_ = ~ is_slti_blt_slt;
  assign _00577_ = ~ is_sltiu_bltu_sltu;
  assign _00578_ = ~ instr_bne;
  assign _00579_ = ~ instr_bge;
  assign _00580_ = ~ _00871_;
  assign _00581_ = ~ _07250_;
  assign _00582_ = ~ _07247_;
  assign _00583_ = ~ _07251_;
  assign _00584_ = ~ _07272_;
  assign _00585_ = ~ _05118_;
  assign _00586_ = ~ _01078_;
  assign _00587_ = ~ _07265_;
  assign _00588_ = ~ _05120_;
  assign _00589_ = ~ { _07254_, _07254_, _07254_, _07254_ };
  assign _00590_ = ~ { _07270_, _07270_, _07270_, _07270_ };
  assign _00591_ = ~ { _05122_, _05122_, _05122_, _05122_ };
  assign _00592_ = ~ { _07251_, _07251_, _07251_, _07251_ };
  assign _00593_ = ~ { _07272_, _07272_, _07272_, _07272_ };
  assign _00594_ = ~ { _05118_, _05118_, _05118_, _05118_ };
  assign _00595_ = ~ { _01078_, _01078_, _01078_, _01078_ };
  assign _00596_ = ~ { _07265_, _07265_, _07265_, _07265_ };
  assign _00597_ = ~ { _05120_, _05120_, _05120_, _05120_ };
  assign _00598_ = ~ { _01076_, _01076_, _01076_, _01076_ };
  assign _00599_ = ~ _07267_;
  assign _00600_ = ~ _00865_;
  assign _00601_ = ~ _05124_;
  assign _00602_ = ~ { is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu };
  assign _00603_ = ~ { is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw };
  assign _00604_ = ~ { instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal };
  assign _00605_ = ~ { _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_ };
  assign _00606_ = ~ { _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_ };
  assign _00607_ = ~ { _07254_, _07254_, _07254_, _07254_, _07254_ };
  assign _00608_ = ~ { _07250_, _07250_, _07250_, _07250_, _07250_ };
  assign _00609_ = ~ { _05122_, _05122_, _05122_, _05122_, _05122_ };
  assign _00610_ = ~ { _07251_, _07251_, _07251_, _07251_, _07251_ };
  assign _00611_ = ~ { _07272_, _07272_, _07272_, _07272_, _07272_ };
  assign _00612_ = ~ { _05118_, _05118_, _05118_, _05118_, _05118_ };
  assign _00613_ = ~ { _07247_, _07247_, _07247_, _07247_, _07247_ };
  assign _00614_ = ~ { _05126_, _05126_, _05126_, _05126_, _05126_ };
  assign _00615_ = ~ { _00865_, _00865_, _00865_, _00865_, _00865_ };
  assign _00616_ = ~ { _05124_, _05124_, _05124_, _05124_, _05124_ };
  assign _00617_ = ~ { _07439_, _07439_ };
  assign _00618_ = ~ { _05128_, _05128_ };
  assign _00619_ = ~ _07439_;
  assign _00620_ = ~ _06535_;
  assign _00621_ = ~ _00861_;
  assign _00622_ = ~ _01090_;
  assign _00623_ = ~ _00863_;
  assign _00624_ = ~ { _07270_, _07270_, _07270_, _07270_, _07270_ };
  assign _00625_ = ~ { _01076_, _01076_, _01076_ };
  assign _00626_ = ~ { _07250_, _07250_, _07250_ };
  assign _00627_ = ~ { _05130_, _05130_, _05130_ };
  assign _00628_ = ~ { _07251_, _07251_, _07251_ };
  assign _00629_ = ~ { _07272_, _07272_, _07272_ };
  assign _00630_ = ~ { _05118_, _05118_, _05118_ };
  assign _00631_ = ~ { _07265_, _07265_, _07265_ };
  assign _00632_ = ~ { _07247_, _07247_, _07247_ };
  assign _00633_ = ~ { _05132_, _05132_, _05132_ };
  assign _00634_ = ~ { _07254_, _07254_, _07254_, _07254_, _07254_, _07254_ };
  assign _00635_ = ~ { _07250_, _07250_, _07250_, _07250_, _07250_, _07250_ };
  assign _00636_ = ~ { _07270_, _07270_, _07270_, _07270_, _07270_, _07270_ };
  assign _00637_ = ~ { _05122_, _05122_, _05122_, _05122_, _05122_, _05122_ };
  assign _00638_ = ~ { _07251_, _07251_, _07251_, _07251_, _07251_, _07251_ };
  assign _00639_ = ~ { _07272_, _07272_, _07272_, _07272_, _07272_, _07272_ };
  assign _00640_ = ~ { _05118_, _05118_, _05118_, _05118_, _05118_, _05118_ };
  assign _00641_ = ~ { _01078_, _01078_, _01078_, _01078_, _01078_, _01078_ };
  assign _00642_ = ~ { _00865_, _00865_, _00865_, _00865_, _00865_, _00865_ };
  assign _00643_ = ~ { _07265_, _07265_, _07265_, _07265_, _07265_, _07265_ };
  assign _00644_ = ~ { _05120_, _05120_, _05120_, _05120_, _05120_, _05120_ };
  assign _00645_ = ~ { _01076_, _01076_, _01076_, _01076_, _01076_, _01076_ };
  assign _00646_ = ~ { _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_ };
  assign _00647_ = ~ { _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_ };
  assign _00648_ = ~ { _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_ };
  assign _00649_ = ~ { pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1] };
  assign _00650_ = ~ { _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_ };
  assign _00651_ = ~ { _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_ };
  assign _00652_ = ~ { _07557_, _07557_, _07557_, _07557_ };
  assign _00653_ = ~ { pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready };
  assign _00654_ = ~ pcpi_div_ready;
  assign _00655_ = ~ { _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4] };
  assign _00656_ = ~ { _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3] };
  assign _00657_ = ~ { _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2] };
  assign _00658_ = ~ { _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1] };
  assign _00659_ = ~ { _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0] };
  assign _00660_ = ~ { _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4] };
  assign _00661_ = ~ { _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3] };
  assign _00662_ = ~ { _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2] };
  assign _00663_ = ~ { _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1] };
  assign _00664_ = ~ { _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0] };
  assign _00665_ = ~ _06865_;
  assign _00666_ = ~ is_beq_bne_blt_bge_bltu_bgeu;
  assign _00667_ = ~ alu_out_0;
  assign _00668_ = ~ { latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch };
  assign _00669_ = ~ { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn };
  assign _00670_ = ~ resetn;
  assign _00671_ = ~ _06615_;
  assign _00672_ = ~ { _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_ };
  assign _00673_ = ~ { _06597_, _06597_, _06597_, _06597_, _06597_ };
  assign _00674_ = ~ { _06499_, _06499_, _06499_, _06499_, _06499_ };
  assign _00675_ = ~ instr_jal;
  assign _00676_ = ~ decoder_trigger;
  assign _00677_ = ~ pcpi_int_ready;
  assign _00678_ = ~ { _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_ };
  assign _00679_ = ~ { _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_ };
  assign _00680_ = ~ { _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_ };
  assign _00681_ = ~ { mem_done, mem_done, mem_done, mem_done, mem_done, mem_done, mem_done, mem_done };
  assign _00682_ = ~ { _06611_, _06611_, _06611_, _06611_, _06611_, _06611_, _06611_, _06611_ };
  assign _00683_ = ~ { pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready };
  assign _00684_ = ~ { decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger };
  assign _00685_ = ~ { _06619_, _06619_, _06619_, _06619_, _06619_, _06619_, _06619_, _06619_ };
  assign _00686_ = ~ { _06621_, _06621_, _06621_, _06621_, _06621_, _06621_, _06621_, _06621_ };
  assign _00687_ = ~ { _06617_, _06617_, _06617_, _06617_, _06617_, _06617_, _06617_, _06617_ };
  assign _00688_ = ~ { launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn };
  assign _00689_ = ~ { _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_ };
  assign _00690_ = ~ { _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_ };
  assign _00691_ = ~ _06872_;
  assign _00692_ = ~ { mem_do_rdata, mem_do_rdata };
  assign _00693_ = ~ { mem_do_wdata, mem_do_wdata };
  assign _00694_ = ~ { mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata };
  assign _00695_ = ~ { mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata };
  assign _00696_ = ~ { _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_ };
  assign _00697_ = ~ { decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger };
  assign _00698_ = ~ _06485_;
  assign _00699_ = ~ _06863_;
  assign _00700_ = ~ _06683_;
  assign _00701_ = ~ _06667_;
  assign _00702_ = ~ _06671_;
  assign _00703_ = ~ _06673_;
  assign _00704_ = ~ mem_rdata_latched[12];
  assign _00705_ = ~ _06679_;
  assign _00706_ = ~ _06521_;
  assign _00707_ = ~ _06523_;
  assign _00708_ = ~ _06515_;
  assign _00709_ = ~ _06895_;
  assign _00710_ = ~ _01076_;
  assign _00711_ = ~ _06677_;
  assign _00712_ = ~ { _06677_, _06677_, _06677_ };
  assign _00713_ = ~ { _06677_, _06677_ };
  assign _00714_ = ~ { _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_ };
  assign _00715_ = ~ { _06667_, _06667_, _06667_, _06667_ };
  assign _00716_ = ~ { _06671_, _06671_, _06671_, _06671_ };
  assign _00717_ = ~ { _06673_, _06673_, _06673_, _06673_ };
  assign _00718_ = ~ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] };
  assign _00719_ = ~ { _06521_, _06521_, _06521_, _06521_ };
  assign _00720_ = ~ { _06523_, _06523_, _06523_, _06523_ };
  assign _00721_ = ~ { _06677_, _06677_, _06677_, _06677_ };
  assign _00722_ = ~ _07254_;
  assign _00723_ = ~ _07090_;
  assign _00724_ = ~ _07270_;
  assign _00725_ = ~ { _06673_, _06673_, _06673_, _06673_, _06673_ };
  assign _00726_ = ~ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] };
  assign _00727_ = ~ { _06523_, _06523_, _06523_, _06523_, _06523_ };
  assign _00728_ = ~ { _06677_, _06677_, _06677_, _06677_, _06677_ };
  assign _00729_ = ~ { _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_ };
  assign _00730_ = ~ { _06671_, _06671_, _06671_, _06671_, _06671_ };
  assign _00731_ = ~ { _06521_, _06521_, _06521_, _06521_, _06521_ };
  assign _00732_ = ~ _01088_;
  assign _00733_ = ~ { decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q };
  assign _00734_ = ~ { decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q };
  assign _00735_ = ~ { dbg_next, dbg_next, dbg_next, dbg_next, dbg_next };
  assign _00736_ = ~ { dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next };
  assign _00737_ = ~ { _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_ };
  assign _00738_ = ~ { mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata };
  assign _00739_ = ~ { mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word };
  assign _00740_ = ~ { mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read };
  assign _00741_ = ~ { mem_la_read, mem_la_read };
  assign _00742_ = ~ { _06888_, _06888_ };
  assign _00743_ = ~ { _06891_, _06891_, _06891_, _06891_ };
  assign _00744_ = ~ { _06884_, _06884_, _06884_, _06884_ };
  assign _00745_ = ~ { _06836_, _06836_, _06836_, _06836_ };
  assign _00746_ = ~ _06665_;
  assign _00747_ = ~ _06517_;
  assign _00748_ = ~ _06519_;
  assign _00749_ = ~ _06663_;
  assign _00750_ = ~ { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer };
  assign _00751_ = ~ { _06665_, _06665_, _06665_, _06665_, _06665_ };
  assign _00752_ = ~ { _06515_, _06515_, _06515_, _06515_, _06515_ };
  assign _00753_ = ~ { _06663_, _06663_, _06663_, _06663_, _06663_ };
  assign _00754_ = ~ { _07265_, _07265_, _07265_, _07265_, _07265_ };
  assign _00755_ = ~ { _07267_, _07267_, _07267_, _07267_, _07267_ };
  assign _00756_ = ~ { mem_xfer, mem_xfer, mem_xfer };
  assign _00757_ = ~ { _06665_, _06665_, _06665_ };
  assign _00758_ = ~ { _06667_, _06667_, _06667_ };
  assign _00759_ = ~ { _06671_, _06671_, _06671_ };
  assign _00760_ = ~ { _06673_, _06673_, _06673_ };
  assign _00761_ = ~ { _06517_, _06517_, _06517_ };
  assign _00762_ = ~ { _06519_, _06519_, _06519_ };
  assign _00763_ = ~ { _06521_, _06521_, _06521_ };
  assign _00764_ = ~ { _06525_, _06525_, _06525_ };
  assign _00765_ = ~ { _06527_, _06527_, _06527_ };
  assign _00766_ = ~ { _06529_, _06529_, _06529_ };
  assign _00767_ = ~ { _06531_, _06531_, _06531_ };
  assign _00768_ = ~ { _06523_, _06523_, _06523_ };
  assign _00769_ = ~ { _06515_, _06515_, _06515_ };
  assign _00770_ = ~ { _06663_, _06663_, _06663_ };
  assign _00771_ = ~ { mem_xfer, mem_xfer, mem_xfer, mem_xfer };
  assign _00772_ = ~ { _06663_, _06663_, _06663_, _06663_ };
  assign _00773_ = ~ { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer };
  assign _00774_ = ~ { _06665_, _06665_, _06665_, _06665_, _06665_, _06665_ };
  assign _00775_ = ~ { _06667_, _06667_, _06667_, _06667_, _06667_, _06667_ };
  assign _00776_ = ~ { _06671_, _06671_, _06671_, _06671_, _06671_, _06671_ };
  assign _00777_ = ~ { _06673_, _06673_, _06673_, _06673_, _06673_, _06673_ };
  assign _00778_ = ~ { _06517_, _06517_, _06517_, _06517_, _06517_, _06517_ };
  assign _00779_ = ~ { _06519_, _06519_, _06519_, _06519_, _06519_, _06519_ };
  assign _00780_ = ~ { _06521_, _06521_, _06521_, _06521_, _06521_, _06521_ };
  assign _00781_ = ~ { _06523_, _06523_, _06523_, _06523_, _06523_, _06523_ };
  assign _00782_ = ~ { _06515_, _06515_, _06515_, _06515_, _06515_, _06515_ };
  assign _00783_ = ~ { _06663_, _06663_, _06663_, _06663_, _06663_, _06663_ };
  assign _00784_ = ~ last_mem_valid;
  assign _00785_ = ~ { _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_ };
  assign _00786_ = ~ { _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_ };
  assign _00787_ = ~ { _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_ };
  assign _00788_ = ~ { instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub };
  assign _00789_ = ~ { latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store };
  assign _00790_ = ~ { latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu };
  assign _00791_ = ~ { instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui };
  assign _00792_ = ~ { _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_ };
  assign _00793_ = ~ { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer };
  assign _00794_ = ~ { mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word };
  assign _00795_ = ~ { mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword };
  assign _00796_ = ~ { mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword };
  assign _03981_ = { _06608_, _06608_, _06608_, _06608_, _06608_ } | _00515_;
  assign _04073_ = _06492_ | _00517_;
  assign _04076_ = _01098_ | _00518_;
  assign _04079_ = { latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0 } | _00519_;
  assign _04082_ = { latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0 } | _00520_;
  assign _04085_ = { _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_ } | _00521_;
  assign _04088_ = { _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_ } | _00522_;
  assign _04091_ = { _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_ } | _00523_;
  assign _04094_ = { _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_ } | _00524_;
  assign _04097_ = { is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0 } | _00525_;
  assign _04100_ = { instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0 } | _00526_;
  assign _04103_ = { instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0 } | _00527_;
  assign _04106_ = { _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_ } | _00528_;
  assign _04109_ = { _06490_, _06490_, _06490_, _06490_, _06490_ } | _00529_;
  assign _04112_ = { _06494_, _06494_, _06494_, _06494_, _06494_ } | _00530_;
  assign _04115_ = { is_slli_srli_srai_t0, is_slli_srli_srai_t0, is_slli_srli_srai_t0, is_slli_srli_srai_t0, is_slli_srli_srai_t0 } | _00531_;
  assign _04118_ = { _01085_, _01085_, _01085_, _01085_, _01085_ } | _00532_;
  assign _04119_ = { _06492_, _06492_, _06492_, _06492_, _06492_ } | _00533_;
  assign _04121_ = _01083_ | _00534_;
  assign _04122_ = _06488_ | _00535_;
  assign _04124_ = _06490_ | _00536_;
  assign _04127_ = _05105_ | _00537_;
  assign _04130_ = is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0 | _00538_;
  assign _04131_ = { _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_ } | _00539_;
  assign _04134_ = { _01098_, _01098_, _01098_, _01098_, _01098_, _01098_, _01098_, _01098_ } | _00540_;
  assign _04137_ = { _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_ } | _00541_;
  assign _04140_ = { _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_ } | _00542_;
  assign _04143_ = { _05107_, _05107_, _05107_, _05107_, _05107_, _05107_, _05107_, _05107_ } | _00543_;
  assign _04146_ = { _00868_, _00868_, _00868_, _00868_, _00868_, _00868_, _00868_, _00868_ } | _00544_;
  assign _04149_ = { is_sll_srl_sra_t0, is_sll_srl_sra_t0, is_sll_srl_sra_t0, is_sll_srl_sra_t0, is_sll_srl_sra_t0, is_sll_srl_sra_t0, is_sll_srl_sra_t0, is_sll_srl_sra_t0 } | _00545_;
  assign _04150_ = { instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0 } | _00546_;
  assign _04152_ = { _05109_, _05109_, _05109_, _05109_, _05109_, _05109_, _05109_, _05109_ } | _00547_;
  assign _04155_ = { _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_ } | _00548_;
  assign _04157_ = { is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0 } | _00549_;
  assign _04158_ = { _00870_, _00870_, _00870_, _00870_, _00870_, _00870_, _00870_, _00870_ } | _00550_;
  assign _04161_ = { _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_ } | _00551_;
  assign _04165_ = _06494_ | _00552_;
  assign _04169_ = _05111_ | _00553_;
  assign _04172_ = is_sll_srl_sra_t0 | _00554_;
  assign _04173_ = instr_trap_t0 | _00555_;
  assign _04176_ = _05109_ | _00556_;
  assign _04177_ = is_sb_sh_sw_t0 | _00557_;
  assign _04180_ = _06614_ | _00559_;
  assign _04181_ = _05113_ | _00560_;
  assign _04184_ = { instr_lw_t0, instr_lw_t0 } | _00561_;
  assign _04186_ = { _06498_, _06498_ } | _00562_;
  assign _04189_ = { instr_sw_t0, instr_sw_t0 } | _00563_;
  assign _04191_ = { _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_, _01096_ } | _00564_;
  assign _04192_ = { _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_ } | _00565_;
  assign _04196_ = { _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_ } | _00566_;
  assign _04199_ = { _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_ } | _00567_;
  assign _04202_ = { _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_ } | _00568_;
  assign _04205_ = { _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_ } | _00569_;
  assign _04210_ = { is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0 } | _00570_;
  assign _04213_ = { _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_ } | _00571_;
  assign _04216_ = { _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_ } | _00572_;
  assign _04219_ = { is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0 } | _00573_;
  assign _04222_ = { _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_ } | _00574_;
  assign _04225_ = { _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_ } | _00575_;
  assign _04228_ = is_slti_blt_slt_t0 | _00576_;
  assign _04231_ = is_sltiu_bltu_sltu_t0 | _00577_;
  assign _04234_ = instr_bne_t0 | _00578_;
  assign _04237_ = instr_bge_t0 | _00579_;
  assign _04240_ = _00872_ | _00580_;
  assign _04243_ = _06303_[1] | _00581_;
  assign _04245_ = _07248_ | _00582_;
  assign _04248_ = _07252_ | _00583_;
  assign _04251_ = _07273_ | _00584_;
  assign _04253_ = _05119_ | _00585_;
  assign _04256_ = _01079_ | _00586_;
  assign _04259_ = _07266_ | _00587_;
  assign _04262_ = _05121_ | _00588_;
  assign _04265_ = { _07255_, _07255_, _07255_, _07255_ } | _00589_;
  assign _04268_ = { _07271_, _07271_, _07271_, _07271_ } | _00590_;
  assign _04271_ = { _05123_, _05123_, _05123_, _05123_ } | _00591_;
  assign _04274_ = { _07252_, _07252_, _07252_, _07252_ } | _00592_;
  assign _04277_ = { _07273_, _07273_, _07273_, _07273_ } | _00593_;
  assign _04279_ = { _05119_, _05119_, _05119_, _05119_ } | _00594_;
  assign _04282_ = { _01079_, _01079_, _01079_, _01079_ } | _00595_;
  assign _04285_ = { _07266_, _07266_, _07266_, _07266_ } | _00596_;
  assign _04288_ = { _05121_, _05121_, _05121_, _05121_ } | _00597_;
  assign _04291_ = { _01077_, _01077_, _01077_, _01077_ } | _00598_;
  assign _04294_ = _07268_ | _00599_;
  assign _04302_ = _00866_ | _00600_;
  assign _04303_ = _05125_ | _00601_;
  assign _04308_ = { is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0 } | _00602_;
  assign _04311_ = { is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0 } | _00603_;
  assign _04314_ = { instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0 } | _00604_;
  assign _04316_ = { _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_ } | _00605_;
  assign _04319_ = { _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_ } | _00606_;
  assign _04322_ = { _07255_, _07255_, _07255_, _07255_, _07255_ } | _00607_;
  assign _04325_ = { _06303_[1], _06303_[1], _06303_[1], _06303_[1], _06303_[1] } | _00608_;
  assign _04327_ = { _05123_, _05123_, _05123_, _05123_, _05123_ } | _00609_;
  assign _04330_ = { _07252_, _07252_, _07252_, _07252_, _07252_ } | _00610_;
  assign _04333_ = { _07273_, _07273_, _07273_, _07273_, _07273_ } | _00611_;
  assign _04335_ = { _05119_, _05119_, _05119_, _05119_, _05119_ } | _00612_;
  assign _04338_ = { _07248_, _07248_, _07248_, _07248_, _07248_ } | _00613_;
  assign _04341_ = { _05127_, _05127_, _05127_, _05127_, _05127_ } | _00614_;
  assign _04347_ = { _00866_, _00866_, _00866_, _00866_, _00866_ } | _00615_;
  assign _04350_ = { _05125_, _05125_, _05125_, _05125_, _05125_ } | _00616_;
  assign _04353_ = { _07440_, _07440_ } | _00617_;
  assign _04356_ = { _05129_, _05129_ } | _00618_;
  assign _04359_ = _07440_ | _00619_;
  assign _04362_ = _06536_ | _00620_;
  assign _04364_ = _00862_ | _00621_;
  assign _04369_ = _01091_ | _00622_;
  assign _04373_ = _00864_ | _00623_;
  assign _04376_ = { _07271_, _07271_, _07271_, _07271_, _07271_ } | _00624_;
  assign _04388_ = { _01077_, _01077_, _01077_ } | _00625_;
  assign _04389_ = { _06303_[1], _06303_[1], _06303_[1] } | _00626_;
  assign _04390_ = { _05131_, _05131_, _05131_ } | _00627_;
  assign _04393_ = { _07252_, _07252_, _07252_ } | _00628_;
  assign _04396_ = { _07273_, _07273_, _07273_ } | _00629_;
  assign _04399_ = { _05119_, _05119_, _05119_ } | _00630_;
  assign _04402_ = { _07266_, _07266_, _07266_ } | _00631_;
  assign _04405_ = { _07248_, _07248_, _07248_ } | _00632_;
  assign _04408_ = { _05133_, _05133_, _05133_ } | _00633_;
  assign _04414_ = { _07255_, _07255_, _07255_, _07255_, _07255_, _07255_ } | _00634_;
  assign _04417_ = { _06303_[1], _06303_[1], _06303_[1], _06303_[1], _06303_[1], _06303_[1] } | _00635_;
  assign _04419_ = { _07271_, _07271_, _07271_, _07271_, _07271_, _07271_ } | _00636_;
  assign _04422_ = { _05123_, _05123_, _05123_, _05123_, _05123_, _05123_ } | _00637_;
  assign _04425_ = { _07252_, _07252_, _07252_, _07252_, _07252_, _07252_ } | _00638_;
  assign _04428_ = { _07273_, _07273_, _07273_, _07273_, _07273_, _07273_ } | _00639_;
  assign _04431_ = { _05119_, _05119_, _05119_, _05119_, _05119_, _05119_ } | _00640_;
  assign _04434_ = { _01079_, _01079_, _01079_, _01079_, _01079_, _01079_ } | _00641_;
  assign _04437_ = { _00866_, _00866_, _00866_, _00866_, _00866_, _00866_ } | _00642_;
  assign _04440_ = { _07266_, _07266_, _07266_, _07266_, _07266_, _07266_ } | _00643_;
  assign _04443_ = { _05121_, _05121_, _05121_, _05121_, _05121_, _05121_ } | _00644_;
  assign _04447_ = { _01077_, _01077_, _01077_, _01077_, _01077_, _01077_ } | _00645_;
  assign _04450_ = { _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_ } | _00646_;
  assign _04453_ = { _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_ } | _00647_;
  assign _04456_ = { _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_ } | _00648_;
  assign _04459_ = { pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1] } | _00649_;
  assign _04462_ = { _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_ } | _00650_;
  assign _04465_ = { _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_ } | _00651_;
  assign _04469_ = { _07558_, _07558_, _07558_, _07558_ } | _00652_;
  assign _04474_ = { pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0 } | _00653_;
  assign _04478_ = pcpi_div_ready_t0 | _00654_;
  assign _04620_ = { _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4] } | _00655_;
  assign _04623_ = { _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3] } | _00656_;
  assign _04627_ = { _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2] } | _00657_;
  assign _04633_ = { _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1] } | _00658_;
  assign _04643_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } | _00659_;
  assign _04661_ = { _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4] } | _00660_;
  assign _04664_ = { _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3] } | _00661_;
  assign _04668_ = { _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2] } | _00662_;
  assign _04674_ = { _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1] } | _00663_;
  assign _04684_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } | _00664_;
  assign _04741_ = _06866_ | _00665_;
  assign _04743_ = is_beq_bne_blt_bge_bltu_bgeu_t0 | _00666_;
  assign _04745_ = mem_do_wdata_t0 | _00491_;
  assign _04746_ = mem_do_rdata_t0 | _00467_;
  assign _04747_ = alu_out_0_t0 | _00667_;
  assign _04748_ = { latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0 } | _00668_;
  assign _04752_ = _06616_ | _00671_;
  assign _04757_ = { _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_ } | _00672_;
  assign _04761_ = { _06598_, _06598_, _06598_, _06598_, _06598_ } | _00673_;
  assign _04764_ = { _06500_, _06500_, _06500_, _06500_, _06500_ } | _00674_;
  assign _04766_ = decoder_trigger_t0 | _00676_;
  assign _04768_ = pcpi_int_ready_t0 | _00677_;
  assign _04771_ = { _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_ } | _00678_;
  assign _04772_ = { _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_ } | _00679_;
  assign _04775_ = { _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_ } | _00680_;
  assign _04776_ = { mem_done_t0, mem_done_t0, mem_done_t0, mem_done_t0, mem_done_t0, mem_done_t0, mem_done_t0, mem_done_t0 } | _00681_;
  assign _04778_ = { _06612_, _06612_, _06612_, _06612_, _06612_, _06612_, _06612_, _06612_ } | _00682_;
  assign _04779_ = { pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0 } | _00683_;
  assign _04781_ = { decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0 } | _00684_;
  assign _04784_ = { _06620_, _06620_, _06620_, _06620_, _06620_, _06620_, _06620_, _06620_ } | _00685_;
  assign _04785_ = { _06622_, _06622_, _06622_, _06622_, _06622_, _06622_, _06622_, _06622_ } | _00686_;
  assign _04786_ = { _06618_, _06618_, _06618_, _06618_, _06618_, _06618_, _06618_, _06618_ } | _00687_;
  assign _04789_ = { launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0, launch_next_insn_t0 } | _00688_;
  assign _04790_ = { _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_ } | _00689_;
  assign _04793_ = { _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_ } | _00690_;
  assign _04799_ = _06873_ | _00691_;
  assign _04800_ = { mem_do_rdata_t0, mem_do_rdata_t0 } | _00692_;
  assign _04802_ = { mem_do_wdata_t0, mem_do_wdata_t0 } | _00693_;
  assign _04803_ = { mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0 } | _00694_;
  assign _04804_ = { mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0, mem_do_wdata_t0 } | _00695_;
  assign _04805_ = { _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_ } | _00696_;
  assign _04809_ = { decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0 } | _00697_;
  assign _04816_ = _06864_ | _00699_;
  assign _04818_ = _06684_ | _00700_;
  assign _04820_ = _06668_ | _00701_;
  assign _04821_ = _06672_ | _00702_;
  assign _04824_ = _06674_ | _00703_;
  assign _04827_ = mem_rdata_latched_t0[12] | _00704_;
  assign _04828_ = _06680_ | _00705_;
  assign _04830_ = _06522_ | _00706_;
  assign _04833_ = _06524_ | _00707_;
  assign _04836_ = _06516_ | _00708_;
  assign _04838_ = _06896_ | _00709_;
  assign _04841_ = _06678_ | _00711_;
  assign _04847_ = { _06678_, _06678_, _06678_ } | _00712_;
  assign _04851_ = { _06678_, _06678_ } | _00713_;
  assign _04854_ = { _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_ } | _00714_;
  assign _04860_ = { _06668_, _06668_, _06668_, _06668_ } | _00715_;
  assign _04861_ = { _06672_, _06672_, _06672_, _06672_ } | _00716_;
  assign _04864_ = { _06674_, _06674_, _06674_, _06674_ } | _00717_;
  assign _04867_ = { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] } | _00718_;
  assign _04869_ = { _06522_, _06522_, _06522_, _06522_ } | _00719_;
  assign _04872_ = { _06524_, _06524_, _06524_, _06524_ } | _00720_;
  assign _04877_ = { _06678_, _06678_, _06678_, _06678_ } | _00721_;
  assign _04890_ = _07255_ | _00722_;
  assign _04892_ = _07091_ | _00723_;
  assign _04893_ = _07271_ | _00724_;
  assign _04898_ = { _06674_, _06674_, _06674_, _06674_, _06674_ } | _00725_;
  assign _04901_ = { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] } | _00726_;
  assign _04903_ = { _06524_, _06524_, _06524_, _06524_, _06524_ } | _00727_;
  assign _04906_ = { _06678_, _06678_, _06678_, _06678_, _06678_ } | _00728_;
  assign _04909_ = { _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_ } | _00729_;
  assign _04912_ = { _06672_, _06672_, _06672_, _06672_, _06672_ } | _00730_;
  assign _04915_ = { _06522_, _06522_, _06522_, _06522_, _06522_ } | _00731_;
  assign _04924_ = _01089_ | _00732_;
  assign _04931_ = { decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0 } | _00733_;
  assign _04935_ = { decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0 } | _00734_;
  assign _04938_ = { dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0 } | _00735_;
  assign _04942_ = { dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0 } | _00736_;
  assign _04945_ = { _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_ } | _00737_;
  assign _04949_ = { mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0, mem_do_rdata_t0 } | _00738_;
  assign _04950_ = { mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0 } | _00739_;
  assign _04951_ = { mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0 } | _00740_;
  assign _04955_ = { mem_la_read_t0, mem_la_read_t0 } | _00741_;
  assign _04956_ = { _00797_, _00797_ } | _00742_;
  assign _04957_ = { _06892_, _06892_, _06892_, _06892_ } | _00743_;
  assign _04960_ = { _06885_, _06885_, _06885_, _06885_ } | _00744_;
  assign _04961_ = { _06837_, _06837_, _06837_, _06837_ } | _00745_;
  assign _04965_ = mem_xfer_t0 | _00172_;
  assign _04967_ = _00797_ | _00175_;
  assign _04969_ = _06666_ | _00746_;
  assign _04970_ = _06518_ | _00747_;
  assign _04971_ = _06520_ | _00748_;
  assign _04973_ = _06664_ | _00749_;
  assign _04979_ = { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 } | _00750_;
  assign _04982_ = { _06666_, _06666_, _06666_, _06666_, _06666_ } | _00751_;
  assign _04984_ = { _06516_, _06516_, _06516_, _06516_, _06516_ } | _00752_;
  assign _04987_ = { _06664_, _06664_, _06664_, _06664_, _06664_ } | _00753_;
  assign _04992_ = { _07266_, _07266_, _07266_, _07266_, _07266_ } | _00754_;
  assign _04995_ = { _07268_, _07268_, _07268_, _07268_, _07268_ } | _00755_;
  assign _04999_ = { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 } | _00756_;
  assign _05002_ = { _06666_, _06666_, _06666_ } | _00757_;
  assign _05003_ = { _06668_, _06668_, _06668_ } | _00758_;
  assign _05004_ = { _06672_, _06672_, _06672_ } | _00759_;
  assign _05005_ = { _06674_, _06674_, _06674_ } | _00760_;
  assign _05006_ = { _06518_, _06518_, _06518_ } | _00761_;
  assign _05007_ = { _06520_, _06520_, _06520_ } | _00762_;
  assign _05008_ = { _06522_, _06522_, _06522_ } | _00763_;
  assign _05009_ = { _06526_, _06526_, _06526_ } | _00764_;
  assign _05010_ = { _06528_, _06528_, _06528_ } | _00765_;
  assign _05011_ = { _06530_, _06530_, _06530_ } | _00766_;
  assign _05012_ = { _06532_, _06532_, _06532_ } | _00767_;
  assign _05013_ = { _06524_, _06524_, _06524_ } | _00768_;
  assign _05016_ = { _06516_, _06516_, _06516_ } | _00769_;
  assign _05017_ = { _06664_, _06664_, _06664_ } | _00770_;
  assign _05020_ = { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 } | _00771_;
  assign _05026_ = { _06664_, _06664_, _06664_, _06664_ } | _00772_;
  assign _05029_ = { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 } | _00773_;
  assign _05032_ = { _06666_, _06666_, _06666_, _06666_, _06666_, _06666_ } | _00774_;
  assign _05033_ = { _06668_, _06668_, _06668_, _06668_, _06668_, _06668_ } | _00775_;
  assign _05034_ = { _06672_, _06672_, _06672_, _06672_, _06672_, _06672_ } | _00776_;
  assign _05035_ = { _06674_, _06674_, _06674_, _06674_, _06674_, _06674_ } | _00777_;
  assign _05036_ = { _06518_, _06518_, _06518_, _06518_, _06518_, _06518_ } | _00778_;
  assign _05037_ = { _06520_, _06520_, _06520_, _06520_, _06520_, _06520_ } | _00779_;
  assign _05038_ = { _06522_, _06522_, _06522_, _06522_, _06522_, _06522_ } | _00780_;
  assign _05041_ = { _06524_, _06524_, _06524_, _06524_, _06524_, _06524_ } | _00781_;
  assign _05044_ = { _06516_, _06516_, _06516_, _06516_, _06516_, _06516_ } | _00782_;
  assign _05047_ = { _06664_, _06664_, _06664_, _06664_, _06664_, _06664_ } | _00783_;
  assign _05050_ = last_mem_valid_t0 | _00784_;
  assign _05053_ = { _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_ } | _00785_;
  assign _05057_ = { _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_ } | _00786_;
  assign _05069_ = { _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_ } | _00787_;
  assign _05072_ = { instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0 } | _00788_;
  assign _05077_ = { latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0 } | _00789_;
  assign _05080_ = { latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0 } | _00790_;
  assign _05083_ = { instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0 } | _00791_;
  assign _05085_ = { _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_ } | _00792_;
  assign _05088_ = { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 } | _00793_;
  assign _05091_ = { mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0 } | _00794_;
  assign _05094_ = { mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0 } | _00795_;
  assign _05097_ = { mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0 } | _00796_;
  assign _03982_ = { _06608_, _06608_, _06608_, _06608_, _06608_ } | { _05738_, _05738_, _05738_, _05738_, _05738_ };
  assign _04072_ = _06498_ | _06497_;
  assign _04074_ = _06492_ | _06491_;
  assign _04077_ = _01098_ | _01097_;
  assign _04080_ = { latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0 } | { latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh };
  assign _04083_ = { latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0 } | { latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb };
  assign _04086_ = { _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_ } | { _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_, _06497_ };
  assign _04089_ = { _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_ } | { _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_ };
  assign _04092_ = { _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_ } | { _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_, _06491_ };
  assign _04095_ = { _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_ } | { _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_, _05100_ };
  assign _04098_ = { is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0 } | { is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh };
  assign _04101_ = { instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0 } | { instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh };
  assign _04104_ = { instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0 } | { instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh };
  assign _04107_ = { _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_ } | { _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_, _05102_ };
  assign _04110_ = { _06490_, _06490_, _06490_, _06490_, _06490_ } | { _06489_, _06489_, _06489_, _06489_, _06489_ };
  assign _04113_ = { _06494_, _06494_, _06494_, _06494_, _06494_ } | { _06493_, _06493_, _06493_, _06493_, _06493_ };
  assign _04116_ = { is_slli_srli_srai_t0, is_slli_srli_srai_t0, is_slli_srli_srai_t0, is_slli_srli_srai_t0, is_slli_srli_srai_t0 } | { is_slli_srli_srai, is_slli_srli_srai, is_slli_srli_srai, is_slli_srli_srai, is_slli_srli_srai };
  assign _04123_ = _06488_ | _06487_;
  assign _04125_ = _06490_ | _06489_;
  assign _04128_ = _05105_ | _05104_;
  assign _04132_ = { _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_ } | { _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_ };
  assign _04135_ = { _01098_, _01098_, _01098_, _01098_, _01098_, _01098_, _01098_, _01098_ } | { _01097_, _01097_, _01097_, _01097_, _01097_, _01097_, _01097_, _01097_ };
  assign _04138_ = { _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_ } | { _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_, _06489_ };
  assign _04141_ = { _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_ } | { _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_ };
  assign _04144_ = { _05107_, _05107_, _05107_, _05107_, _05107_, _05107_, _05107_, _05107_ } | { _05106_, _05106_, _05106_, _05106_, _05106_, _05106_, _05106_, _05106_ };
  assign _04147_ = { _00868_, _00868_, _00868_, _00868_, _00868_, _00868_, _00868_, _00868_ } | { _00867_, _00867_, _00867_, _00867_, _00867_, _00867_, _00867_, _00867_ };
  assign _04151_ = { instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0 } | { instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap };
  assign _04153_ = { _05109_, _05109_, _05109_, _05109_, _05109_, _05109_, _05109_, _05109_ } | { _05108_, _05108_, _05108_, _05108_, _05108_, _05108_, _05108_, _05108_ };
  assign _04159_ = { _00870_, _00870_, _00870_, _00870_, _00870_, _00870_, _00870_, _00870_ } | { _00869_, _00869_, _00869_, _00869_, _00869_, _00869_, _00869_, _00869_ };
  assign _04162_ = { _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_ } | { _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_, _06487_ };
  assign _04166_ = _06494_ | _06493_;
  assign _04170_ = _05111_ | _05110_;
  assign _04174_ = instr_trap_t0 | instr_trap;
  assign _04178_ = _01081_ | _01080_;
  assign _04182_ = _05113_ | _05112_;
  assign _04185_ = { _06496_, _06496_ } | { _06495_, _06495_ };
  assign _04187_ = { _06498_, _06498_ } | { _06497_, _06497_ };
  assign _04193_ = { _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_ } | { _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_, _01080_ };
  assign _04197_ = { _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_ } | { _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_, _06493_ };
  assign _04200_ = { _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_ } | { _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_, _05114_ };
  assign _04203_ = { _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_ } | { _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_, _06859_ };
  assign _04206_ = { _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_ } | { _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_, _06849_ };
  assign _04211_ = { is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0 } | { is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal };
  assign _04214_ = { _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_ } | { _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_, _06601_ };
  assign _04217_ = { _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_ } | { _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_, _06855_ };
  assign _04220_ = { is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0 } | { is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare };
  assign _04223_ = { _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_ } | { _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_, _06851_ };
  assign _04226_ = { _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_ } | { _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_, _05116_ };
  assign _04229_ = is_slti_blt_slt_t0 | is_slti_blt_slt;
  assign _04232_ = is_sltiu_bltu_sltu_t0 | is_sltiu_bltu_sltu;
  assign _04235_ = instr_bne_t0 | instr_bne;
  assign _04238_ = instr_bge_t0 | instr_bge;
  assign _04241_ = _00872_ | _00871_;
  assign _04244_ = _06303_[1] | _07250_;
  assign _04246_ = _07248_ | _07247_;
  assign _04249_ = _07252_ | _07251_;
  assign _04252_ = _07273_ | _07272_;
  assign _04254_ = _05119_ | _05118_;
  assign _04257_ = _01079_ | _01078_;
  assign _04260_ = _07266_ | _07265_;
  assign _04263_ = _05121_ | _05120_;
  assign _04266_ = { _07255_, _07255_, _07255_, _07255_ } | { _07254_, _07254_, _07254_, _07254_ };
  assign _04267_ = { _06303_[1], _06303_[1], _06303_[1], _06303_[1] } | { _07250_, _07250_, _07250_, _07250_ };
  assign _04269_ = { _07271_, _07271_, _07271_, _07271_ } | { _07270_, _07270_, _07270_, _07270_ };
  assign _04272_ = { _05123_, _05123_, _05123_, _05123_ } | { _05122_, _05122_, _05122_, _05122_ };
  assign _04275_ = { _07252_, _07252_, _07252_, _07252_ } | { _07251_, _07251_, _07251_, _07251_ };
  assign _04278_ = { _07273_, _07273_, _07273_, _07273_ } | { _07272_, _07272_, _07272_, _07272_ };
  assign _04280_ = { _05119_, _05119_, _05119_, _05119_ } | { _05118_, _05118_, _05118_, _05118_ };
  assign _04283_ = { _01079_, _01079_, _01079_, _01079_ } | { _01078_, _01078_, _01078_, _01078_ };
  assign _04286_ = { _07266_, _07266_, _07266_, _07266_ } | { _07265_, _07265_, _07265_, _07265_ };
  assign _04289_ = { _05121_, _05121_, _05121_, _05121_ } | { _05120_, _05120_, _05120_, _05120_ };
  assign _04292_ = { _01077_, _01077_, _01077_, _01077_ } | { _01076_, _01076_, _01076_, _01076_ };
  assign _04295_ = _07268_ | _07267_;
  assign _04304_ = _05125_ | _05124_;
  assign _04309_ = { is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0 } | { is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu };
  assign _04312_ = { is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0 } | { is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw };
  assign _04315_ = { instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0 } | { instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal };
  assign _04317_ = { _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_ } | { _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_, _07363_ };
  assign _04320_ = { _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_ } | { _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_, _00873_ };
  assign _04323_ = { _07255_, _07255_, _07255_, _07255_, _07255_ } | { _07254_, _07254_, _07254_, _07254_, _07254_ };
  assign _04326_ = { _06303_[1], _06303_[1], _06303_[1], _06303_[1], _06303_[1] } | { _07250_, _07250_, _07250_, _07250_, _07250_ };
  assign _04328_ = { _05123_, _05123_, _05123_, _05123_, _05123_ } | { _05122_, _05122_, _05122_, _05122_, _05122_ };
  assign _04331_ = { _07252_, _07252_, _07252_, _07252_, _07252_ } | { _07251_, _07251_, _07251_, _07251_, _07251_ };
  assign _04334_ = { _07273_, _07273_, _07273_, _07273_, _07273_ } | { _07272_, _07272_, _07272_, _07272_, _07272_ };
  assign _04336_ = { _05119_, _05119_, _05119_, _05119_, _05119_ } | { _05118_, _05118_, _05118_, _05118_, _05118_ };
  assign _04339_ = { _07248_, _07248_, _07248_, _07248_, _07248_ } | { _07247_, _07247_, _07247_, _07247_, _07247_ };
  assign _04342_ = { _05127_, _05127_, _05127_, _05127_, _05127_ } | { _05126_, _05126_, _05126_, _05126_, _05126_ };
  assign _04348_ = { _00866_, _00866_, _00866_, _00866_, _00866_ } | { _00865_, _00865_, _00865_, _00865_, _00865_ };
  assign _04351_ = { _05125_, _05125_, _05125_, _05125_, _05125_ } | { _05124_, _05124_, _05124_, _05124_, _05124_ };
  assign _04354_ = { _07440_, _07440_ } | { _07439_, _07439_ };
  assign _04357_ = { _05129_, _05129_ } | { _05128_, _05128_ };
  assign _04360_ = _07440_ | _07439_;
  assign _04370_ = _01091_ | _01090_;
  assign _04374_ = _00864_ | _00863_;
  assign _04377_ = { _07271_, _07271_, _07271_, _07271_, _07271_ } | { _07270_, _07270_, _07270_, _07270_, _07270_ };
  assign _04391_ = { _05131_, _05131_, _05131_ } | { _05130_, _05130_, _05130_ };
  assign _04394_ = { _07252_, _07252_, _07252_ } | { _07251_, _07251_, _07251_ };
  assign _04397_ = { _07273_, _07273_, _07273_ } | { _07272_, _07272_, _07272_ };
  assign _04400_ = { _05119_, _05119_, _05119_ } | { _05118_, _05118_, _05118_ };
  assign _04403_ = { _07266_, _07266_, _07266_ } | { _07265_, _07265_, _07265_ };
  assign _04406_ = { _07248_, _07248_, _07248_ } | { _07247_, _07247_, _07247_ };
  assign _04409_ = { _05133_, _05133_, _05133_ } | { _05132_, _05132_, _05132_ };
  assign _04415_ = { _07255_, _07255_, _07255_, _07255_, _07255_, _07255_ } | { _07254_, _07254_, _07254_, _07254_, _07254_, _07254_ };
  assign _04418_ = { _06303_[1], _06303_[1], _06303_[1], _06303_[1], _06303_[1], _06303_[1] } | { _07250_, _07250_, _07250_, _07250_, _07250_, _07250_ };
  assign _04420_ = { _07271_, _07271_, _07271_, _07271_, _07271_, _07271_ } | { _07270_, _07270_, _07270_, _07270_, _07270_, _07270_ };
  assign _04423_ = { _05123_, _05123_, _05123_, _05123_, _05123_, _05123_ } | { _05122_, _05122_, _05122_, _05122_, _05122_, _05122_ };
  assign _04426_ = { _07252_, _07252_, _07252_, _07252_, _07252_, _07252_ } | { _07251_, _07251_, _07251_, _07251_, _07251_, _07251_ };
  assign _04429_ = { _07273_, _07273_, _07273_, _07273_, _07273_, _07273_ } | { _07272_, _07272_, _07272_, _07272_, _07272_, _07272_ };
  assign _04432_ = { _05119_, _05119_, _05119_, _05119_, _05119_, _05119_ } | { _05118_, _05118_, _05118_, _05118_, _05118_, _05118_ };
  assign _04435_ = { _01079_, _01079_, _01079_, _01079_, _01079_, _01079_ } | { _01078_, _01078_, _01078_, _01078_, _01078_, _01078_ };
  assign _04438_ = { _00866_, _00866_, _00866_, _00866_, _00866_, _00866_ } | { _00865_, _00865_, _00865_, _00865_, _00865_, _00865_ };
  assign _04441_ = { _07266_, _07266_, _07266_, _07266_, _07266_, _07266_ } | { _07265_, _07265_, _07265_, _07265_, _07265_, _07265_ };
  assign _04444_ = { _05121_, _05121_, _05121_, _05121_, _05121_, _05121_ } | { _05120_, _05120_, _05120_, _05120_, _05120_, _05120_ };
  assign _04448_ = { _01077_, _01077_, _01077_, _01077_, _01077_, _01077_ } | { _01076_, _01076_, _01076_, _01076_, _01076_, _01076_ };
  assign _04451_ = { _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_ } | { _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_, _07551_ };
  assign _04454_ = { _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_ } | { _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_, _07555_ };
  assign _04457_ = { _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_ } | { _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_, _05134_ };
  assign _04460_ = { pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1] } | { pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1] };
  assign _04463_ = { _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_ } | { _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_, _06503_ };
  assign _04466_ = { _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_ } | { _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_, _07557_ };
  assign _04468_ = { _06504_, _06504_, _06504_, _06504_ } | { _06503_, _06503_, _06503_, _06503_ };
  assign _04470_ = { _07558_, _07558_, _07558_, _07558_ } | { _07557_, _07557_, _07557_, _07557_ };
  assign _04475_ = { pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0 } | { pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready };
  assign _04477_ = pcpi_mul_ready_t0 | pcpi_mul_ready;
  assign _04479_ = pcpi_div_ready_t0 | pcpi_div_ready;
  assign _04621_ = { _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4] } | { _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4], _00080_[4] };
  assign _04624_ = { _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3] } | { _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3], _00080_[3] };
  assign _04628_ = { _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2] } | { _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2], _00080_[2] };
  assign _04634_ = { _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1] } | { _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1], _00080_[1] };
  assign _04644_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } | { _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0], _00080_[0] };
  assign _04662_ = { _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4] } | { _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4], _00082_[4] };
  assign _04665_ = { _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3] } | { _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3], _00082_[3] };
  assign _04669_ = { _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2] } | { _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2], _00082_[2] };
  assign _04675_ = { _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1] } | { _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1], _00082_[1] };
  assign _04685_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } | { _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0], _00082_[0] };
  assign _04735_ = { _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31] } | { _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_, _06509_ };
  assign _04736_ = { _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_ } | { _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_, _06631_ };
  assign _04737_ = { _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_, _06628_ } | { _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_, _06627_ };
  assign _04738_ = { _06628_, _06628_, _06628_, _06628_ } | { _06627_, _06627_, _06627_, _06627_ };
  assign _04739_ = { cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0 } | { cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write };
  assign _04740_ = { cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0 } | { cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write };
  assign _04742_ = _06866_ | _06865_;
  assign _04744_ = is_beq_bne_blt_bge_bltu_bgeu_t0 | is_beq_bne_blt_bge_bltu_bgeu;
  assign _03785_ = mem_do_wdata_t0 | mem_do_wdata;
  assign _03787_ = mem_do_rdata_t0 | mem_do_rdata;
  assign _04749_ = { latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0 } | { latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch };
  assign _04751_ = { _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_ } | { _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_ };
  assign _04755_ = { _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_ } | { _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_, _06615_ };
  assign _04756_ = { _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_ } | { _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_ };
  assign _04758_ = { _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_ } | { _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_, _06499_ };
  assign _04759_ = { instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0 } | { instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap };
  assign _04760_ = { pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0 } | { pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready };
  assign _04762_ = { _06598_, _06598_, _06598_, _06598_, _06598_ } | { _06597_, _06597_, _06597_, _06597_, _06597_ };
  assign _04767_ = decoder_trigger_t0 | decoder_trigger;
  assign _04769_ = pcpi_int_ready_t0 | pcpi_int_ready;
  assign _04773_ = { _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_ } | { _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_, _06865_ };
  assign _04777_ = { is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0 } | { is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu };
  assign _04780_ = { instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0 } | { instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal };
  assign _04782_ = { decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0 } | { decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger };
  assign _04787_ = { _06618_, _06618_, _06618_, _06618_, _06618_, _06618_, _06618_, _06618_ } | { _06617_, _06617_, _06617_, _06617_, _06617_, _06617_, _06617_, _06617_ };
  assign _04791_ = { _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_ } | { _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_, _00855_ };
  assign _04794_ = { _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_ } | { _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_, _00859_ };
  assign _04797_ = _06500_ | _06499_;
  assign _04801_ = { _06866_, _06866_ } | { _06865_, _06865_ };
  assign _04806_ = { _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_ } | { _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_, _06597_ };
  assign _04810_ = { decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0 } | { decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger };
  assign _04812_ = _00858_ | _00857_;
  assign _04813_ = { _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31] } | { _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_, _06605_ };
  assign _04814_ = { _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31] } | { _06605_, _06605_, _06605_, _06605_, _06605_ };
  assign _04815_ = _06486_ | _06485_;
  assign _04817_ = prefetched_high_word_t0 | prefetched_high_word;
  assign _04819_ = _06684_ | _06683_;
  assign _04822_ = _06672_ | _06671_;
  assign _04825_ = _06674_ | _06673_;
  assign _04829_ = _06680_ | _06679_;
  assign _04831_ = _06522_ | _06521_;
  assign _04834_ = _06524_ | _06523_;
  assign _04837_ = _06516_ | _06515_;
  assign _04839_ = _06896_ | _06895_;
  assign _04840_ = _01077_ | _01076_;
  assign _04842_ = _06678_ | _06677_;
  assign _04848_ = { _06678_, _06678_, _06678_ } | { _06677_, _06677_, _06677_ };
  assign _04852_ = { _06678_, _06678_ } | { _06677_, _06677_ };
  assign _04855_ = { _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_ } | { _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_ };
  assign _04859_ = { _06684_, _06684_, _06684_, _06684_ } | { _06683_, _06683_, _06683_, _06683_ };
  assign _04862_ = { _06672_, _06672_, _06672_, _06672_ } | { _06671_, _06671_, _06671_, _06671_ };
  assign _04865_ = { _06674_, _06674_, _06674_, _06674_ } | { _06673_, _06673_, _06673_, _06673_ };
  assign _04868_ = { _06680_, _06680_, _06680_, _06680_ } | { _06679_, _06679_, _06679_, _06679_ };
  assign _04870_ = { _06522_, _06522_, _06522_, _06522_ } | { _06521_, _06521_, _06521_, _06521_ };
  assign _04873_ = { _06524_, _06524_, _06524_, _06524_ } | { _06523_, _06523_, _06523_, _06523_ };
  assign _04875_ = { _06516_, _06516_, _06516_, _06516_ } | { _06515_, _06515_, _06515_, _06515_ };
  assign _04876_ = { _06896_, _06896_, _06896_, _06896_ } | { _06895_, _06895_, _06895_, _06895_ };
  assign _04878_ = { _06678_, _06678_, _06678_, _06678_ } | { _06677_, _06677_, _06677_, _06677_ };
  assign _04894_ = _07271_ | _07270_;
  assign _04897_ = { _06668_, _06668_, _06668_, _06668_, _06668_ } | { _06667_, _06667_, _06667_, _06667_, _06667_ };
  assign _04899_ = { _06674_, _06674_, _06674_, _06674_, _06674_ } | { _06673_, _06673_, _06673_, _06673_, _06673_ };
  assign _04902_ = { _06680_, _06680_, _06680_, _06680_, _06680_ } | { _06679_, _06679_, _06679_, _06679_, _06679_ };
  assign _04904_ = { _06524_, _06524_, _06524_, _06524_, _06524_ } | { _06523_, _06523_, _06523_, _06523_, _06523_ };
  assign _04907_ = { _06678_, _06678_, _06678_, _06678_, _06678_ } | { _06677_, _06677_, _06677_, _06677_, _06677_ };
  assign _04910_ = { _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_ } | { _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_, _06677_ };
  assign _04914_ = { _07091_, _07091_, _07091_, _07091_, _07091_ } | { _07090_, _07090_, _07090_, _07090_, _07090_ };
  assign _04916_ = { _06522_, _06522_, _06522_, _06522_, _06522_ } | { _06521_, _06521_, _06521_, _06521_, _06521_ };
  assign _04919_ = { _06896_, _06896_, _06896_, _06896_, _06896_ } | { _06895_, _06895_, _06895_, _06895_, _06895_ };
  assign _04932_ = { decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0 } | { decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q };
  assign _04936_ = { decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0 } | { decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q };
  assign _04939_ = { dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0 } | { dbg_next, dbg_next, dbg_next, dbg_next, dbg_next };
  assign _04943_ = { dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0 } | { dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next };
  assign _04946_ = { _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_ } | { _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_, _07429_ };
  assign _04948_ = { _06894_, _06894_, _06894_, _06894_, _06894_, _06894_, _06894_, _06894_, _06894_, _06894_, _06894_, _06894_, _06894_, _06894_, _06894_, _06894_ } | { _06893_, _06893_, _06893_, _06893_, _06893_, _06893_, _06893_, _06893_, _06893_, _06893_, _06893_, _06893_, _06893_, _06893_, _06893_, _06893_ };
  assign _04952_ = { mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0 } | { mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read };
  assign _04954_ = { mem_xfer_t0, mem_xfer_t0 } | { mem_xfer, mem_xfer };
  assign _04958_ = { _06892_, _06892_, _06892_, _06892_ } | { _06891_, _06891_, _06891_, _06891_ };
  assign _04962_ = { _06837_, _06837_, _06837_, _06837_ } | { _06836_, _06836_, _06836_, _06836_ };
  assign _04964_ = _06885_ | _06884_;
  assign _04966_ = mem_xfer_t0 | mem_xfer;
  assign _04974_ = _06664_ | _06663_;
  assign _04980_ = { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 } | { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer };
  assign _04985_ = { _06516_, _06516_, _06516_, _06516_, _06516_ } | { _06515_, _06515_, _06515_, _06515_, _06515_ };
  assign _04988_ = { _06664_, _06664_, _06664_, _06664_, _06664_ } | { _06663_, _06663_, _06663_, _06663_, _06663_ };
  assign _04993_ = { _07266_, _07266_, _07266_, _07266_, _07266_ } | { _07265_, _07265_, _07265_, _07265_, _07265_ };
  assign _04996_ = { _07268_, _07268_, _07268_, _07268_, _07268_ } | { _07267_, _07267_, _07267_, _07267_, _07267_ };
  assign _05000_ = { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 } | { mem_xfer, mem_xfer, mem_xfer };
  assign _05014_ = { _06524_, _06524_, _06524_ } | { _06523_, _06523_, _06523_ };
  assign _05018_ = { _06664_, _06664_, _06664_ } | { _06663_, _06663_, _06663_ };
  assign _05021_ = { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 } | { mem_xfer, mem_xfer, mem_xfer, mem_xfer };
  assign _05027_ = { _06664_, _06664_, _06664_, _06664_ } | { _06663_, _06663_, _06663_, _06663_ };
  assign _05030_ = { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 } | { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer };
  assign _05039_ = { _06522_, _06522_, _06522_, _06522_, _06522_, _06522_ } | { _06521_, _06521_, _06521_, _06521_, _06521_, _06521_ };
  assign _05042_ = { _06524_, _06524_, _06524_, _06524_, _06524_, _06524_ } | { _06523_, _06523_, _06523_, _06523_, _06523_, _06523_ };
  assign _05045_ = { _06516_, _06516_, _06516_, _06516_, _06516_, _06516_ } | { _06515_, _06515_, _06515_, _06515_, _06515_, _06515_ };
  assign _05048_ = { _06664_, _06664_, _06664_, _06664_, _06664_, _06664_ } | { _06663_, _06663_, _06663_, _06663_, _06663_, _06663_ };
  assign _05051_ = last_mem_valid_t0 | last_mem_valid;
  assign _05054_ = { _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_ } | { _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_, _06513_ };
  assign _05056_ = { _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31] } | { _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_, _06512_ };
  assign _05058_ = { _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_ } | { _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_, _06510_ };
  assign _05070_ = { _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_ } | { _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_, _06599_ };
  assign _05073_ = { instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0 } | { instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub };
  assign _05075_ = { _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_ } | { _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_, _07564_ };
  assign _05076_ = { _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_ } | { _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_, _07566_ };
  assign _05078_ = { latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0 } | { latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store };
  assign _05081_ = { latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0 } | { latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu };
  assign _05084_ = { _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_ } | { _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_, _07568_ };
  assign _05086_ = { _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_ } | { _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_, _06633_ };
  assign _05089_ = { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 } | { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer };
  assign _05092_ = { mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0 } | { mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word };
  assign _05095_ = { mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0 } | { mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword };
  assign _05098_ = { mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0 } | { mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword };
  assign _01327_ = decoded_rs2_t0 & _03981_;
  assign _01330_ = decoded_rs1_t0 & _03981_;
  assign _01571_ = _06608_ & _04073_;
  assign _01574_ = _06107_ & _04076_;
  assign _01577_ = mem_rdata_word_t0 & _04079_;
  assign _01580_ = _06111_ & _04082_;
  assign _01583_ = _07133_ & _04085_;
  assign _01586_ = _06123_ & _04088_;
  assign _01589_ = _06117_ & _04091_;
  assign _01592_ = _06119_ & _04094_;
  assign _01595_ = _07135_ & _04097_;
  assign _01598_ = count_instr_t0[31:0] & _04100_;
  assign _01601_ = count_cycle_t0[31:0] & _04103_;
  assign _01604_ = _06127_ & _04106_;
  assign _01607_ = _06137_ & _04109_;
  assign _01610_ = _06131_ & _04112_;
  assign _01613_ = cpuregs_rs2_t0[4:0] & _04115_;
  assign _06137_ = _06135_ & _04118_;
  assign _01616_ = decoded_rd_t0 & _04119_;
  assign _01622_ = _07154_ & _04073_;
  assign _01625_ = _07156_ & _04121_;
  assign _01629_ = _06151_ & _04124_;
  assign _01632_ = _06153_ & _04127_;
  assign _01635_ = _07158_ & _04130_;
  assign _01637_ = _07170_ & _04131_;
  assign _01640_ = _06158_ & _04134_;
  assign _01643_ = _06185_ & _04137_;
  assign _01646_ = cpu_state_t0 & _04140_;
  assign _01649_ = _06164_ & _04143_;
  assign _01652_ = _06166_ & _04146_;
  assign _01657_ = _06171_ & _04152_;
  assign _01660_ = { 4'h0, is_sb_sh_sw_t0, 1'h0, is_sb_sh_sw_t0, 1'h0 } & _04149_;
  assign _01662_ = { 5'h00, is_slli_srli_srai_t0, 1'h0, is_slli_srli_srai_t0 } & _04155_;
  assign _01664_ = _06176_ & _04150_;
  assign _01666_ = _06181_ & _04157_;
  assign _01668_ = _06183_ & _04158_;
  assign _01671_ = _07193_ & _04161_;
  assign _01674_ = _06189_ & _04088_;
  assign _01677_ = _06202_ & _04165_;
  assign _01680_ = _07207_ & _04122_;
  assign _01683_ = _06195_ & _04169_;
  assign _01686_ = mem_do_prefetch_t0 & _04173_;
  assign _01689_ = _06200_ & _04176_;
  assign _01691_ = mem_do_prefetch_t0 & _04177_;
  assign _06206_ = _06204_ & _04172_;
  assign _01693_ = _06206_ & _04173_;
  assign _01695_ = _06210_ & _04180_;
  assign _01697_ = _06212_ & _04181_;
  assign _01700_ = { _06215_[1], _06215_[1] } & _04184_;
  assign _01704_ = _06219_ & _04186_;
  assign _01707_ = { instr_sh_t0, instr_sh_t0 } & _04189_;
  assign _01709_ = _06229_ & _04088_;
  assign _06227_ = cpuregs_rs2_t0 & _04191_;
  assign _01711_ = _06227_ & _04192_;
  assign _01714_ = _07225_ & _04085_;
  assign _01717_ = _06247_ & _04196_;
  assign _01720_ = _06233_ & _04199_;
  assign _01723_ = { pcpi_rs1_t0[30:0], 1'h0 } & _04202_;
  assign _01726_ = _06237_ & _04205_;
  assign _01729_ = { pcpi_rs1_t0[27:0], 4'h0 } & _04202_;
  assign _01732_ = _06241_ & _04205_;
  assign _06245_ = cpuregs_rs1_t0 & _04097_;
  assign _01735_ = _06245_ & _04210_;
  assign _01738_ = _00087_ & _04213_;
  assign _01741_ = _07095_ & _04216_;
  assign _01744_ = alu_add_sub_t0 & _04219_;
  assign _01747_ = _06251_ & _04222_;
  assign _01750_ = _06253_ & _04225_;
  assign _01753_ = alu_ltu_t0 & _04228_;
  assign _01756_ = _06255_ & _04231_;
  assign _01759_ = alu_eq_t0 & _04234_;
  assign _01762_ = _06259_ & _04237_;
  assign _01765_ = _06261_ & _04240_;
  assign _01770_ = _06263_ & _04245_;
  assign _01773_ = _06279_ & _04248_;
  assign _01778_ = _06269_ & _04253_;
  assign _01781_ = _07261_ & _04256_;
  assign _01786_ = _06275_ & _04259_;
  assign _01789_ = _06277_ & _04262_;
  assign _01792_ = _07300_ & _04265_;
  assign _01796_ = _06283_ & _04268_;
  assign _01799_ = _06285_ & _04271_;
  assign _01802_ = _06301_ & _04274_;
  assign _01807_ = _06291_ & _04279_;
  assign _01810_ = _07308_ & _04282_;
  assign _01815_ = _06297_ & _04285_;
  assign _01818_ = _06299_ & _04288_;
  assign _01821_ = { 2'h0, _06303_[1], 1'h0 } & _04291_;
  assign _01824_ = _06558_ & _04294_;
  assign _01827_ = _06306_ & _04248_;
  assign _01830_ = _06320_ & _04248_;
  assign _01833_ = _06556_ & _04251_;
  assign _01836_ = _06312_ & _04253_;
  assign _01839_ = _07337_ & _04245_;
  assign _01842_ = _06556_ & _04302_;
  assign _01844_ = _06318_ & _04303_;
  assign _01847_ = _06552_ & _04251_;
  assign _01850_ = _06322_ & _04248_;
  assign _01853_ = { mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31:20] } & _04308_;
  assign _01856_ = _06326_ & _04311_;
  assign _01861_ = _06330_ & _04316_;
  assign _01864_ = _06332_ & _04319_;
  assign _01867_ = _07368_ & _04322_;
  assign _01872_ = _06338_ & _04327_;
  assign _01875_ = _07374_ & _04330_;
  assign _01880_ = _06344_ & _04335_;
  assign _01883_ = _07387_ & _04338_;
  assign _01888_ = _06350_ & _04341_;
  assign _01891_ = _06366_ & _04330_;
  assign _01896_ = _06356_ & _04335_;
  assign _01899_ = _07396_ & _04338_;
  assign _01902_ = { 4'h0, _06362_[0] } & _04347_;
  assign _01905_ = _06364_ & _04350_;
  assign _01908_ = _07451_ & _04353_;
  assign _01911_ = _06370_ & _04356_;
  assign _01914_ = _07466_ & _04359_;
  assign _01917_ = _06374_ & _04362_;
  assign _01919_ = _07468_ & _04245_;
  assign _01922_ = _06377_ & _04364_;
  assign _01924_ = _06389_ & _04248_;
  assign _01927_ = _07468_ & _04251_;
  assign _01930_ = _06383_ & _04253_;
  assign _01935_ = _06387_ & _04369_;
  assign _01938_ = _07483_ & _04294_;
  assign _01941_ = _06391_ & _04373_;
  assign _01944_ = _07488_ & _04376_;
  assign _01947_ = _06395_ & _04338_;
  assign _01950_ = _06409_ & _04330_;
  assign _01953_ = _07488_ & _04333_;
  assign _01956_ = _06401_ & _04335_;
  assign _01959_ = _07495_ & _04338_;
  assign _01962_ = _07488_ & _04347_;
  assign _01965_ = _06407_ & _04350_;
  assign _01968_ = _07488_ & _04325_;
  assign _01971_ = _06411_ & _04376_;
  assign _01974_ = _07509_ & _04388_;
  assign _01976_ = _07504_ & _04389_;
  assign _01978_ = _06417_ & _04390_;
  assign _01981_ = _06433_ & _04393_;
  assign _01984_ = _07504_ & _04396_;
  assign _01987_ = _06423_ & _04399_;
  assign _01990_ = _07504_ & _04402_;
  assign _01993_ = _06429_ & _04405_;
  assign _01996_ = _06431_ & _04408_;
  assign _02000_ = _06435_ & _04388_;
  assign _02002_ = _07532_ & _04274_;
  assign _02005_ = _07528_ & _04277_;
  assign _02008_ = _06441_ & _04279_;
  assign _02011_ = _07540_ & _04414_;
  assign _02014_ = _07535_ & _04417_;
  assign _02016_ = _06447_ & _04419_;
  assign _02019_ = _06449_ & _04422_;
  assign _02022_ = _06465_ & _04425_;
  assign _02025_ = _07535_ & _04428_;
  assign _02028_ = _06455_ & _04431_;
  assign _02031_ = _07548_ & _04434_;
  assign _02034_ = _07535_ & _04437_;
  assign _02037_ = _06461_ & _04440_;
  assign _02040_ = _06463_ & _04443_;
  assign _02045_ = _06467_ & _04447_;
  assign _02048_ = { 24'h000000, mem_rdata_t0[23:16] } & _04450_;
  assign _02051_ = { 24'h000000, mem_rdata_t0[7:0] } & _04453_;
  assign _02054_ = _06473_ & _04456_;
  assign _02057_ = { 16'h0000, mem_rdata_t0[15:0] } & _04459_;
  assign _02060_ = mem_rdata_t0 & _04462_;
  assign _02063_ = _06475_ & _04465_;
  assign _02068_ = _06477_ & _04469_;
  assign _02071_ = pcpi_rs2_t0 & _04462_;
  assign _02074_ = _06479_ & _04465_;
  assign _02077_ = pcpi_mul_rd_t0 & _04474_;
  assign _02082_ = _06481_ & _04478_;
  assign _02495_ = _06902_ & _04620_;
  assign _02498_ = _06906_ & _04623_;
  assign _02501_ = _06910_ & _04623_;
  assign _02504_ = _06914_ & _04627_;
  assign _02507_ = _06918_ & _04627_;
  assign _02510_ = _06922_ & _04627_;
  assign _02513_ = _06926_ & _04627_;
  assign _02516_ = _06930_ & _04633_;
  assign _02519_ = _06934_ & _04633_;
  assign _02522_ = _06938_ & _04633_;
  assign _02525_ = _06942_ & _04633_;
  assign _02528_ = _06946_ & _04633_;
  assign _02531_ = _06950_ & _04633_;
  assign _02534_ = _06954_ & _04633_;
  assign _02537_ = _06958_ & _04633_;
  assign _02540_ = \cpuregs[0]_t0  & _04643_;
  assign _02543_ = \cpuregs[20]_t0  & _04643_;
  assign _02546_ = \cpuregs[22]_t0  & _04643_;
  assign _02549_ = \cpuregs[24]_t0  & _04643_;
  assign _02552_ = \cpuregs[26]_t0  & _04643_;
  assign _02555_ = \cpuregs[28]_t0  & _04643_;
  assign _02558_ = \cpuregs[30]_t0  & _04643_;
  assign _02561_ = \cpuregs[2]_t0  & _04643_;
  assign _02564_ = \cpuregs[4]_t0  & _04643_;
  assign _02567_ = \cpuregs[6]_t0  & _04643_;
  assign _02570_ = \cpuregs[8]_t0  & _04643_;
  assign _02573_ = \cpuregs[10]_t0  & _04643_;
  assign _02576_ = \cpuregs[12]_t0  & _04643_;
  assign _02579_ = \cpuregs[14]_t0  & _04643_;
  assign _02582_ = \cpuregs[16]_t0  & _04643_;
  assign _02585_ = \cpuregs[18]_t0  & _04643_;
  assign _02588_ = _06962_ & _04661_;
  assign _02591_ = _06966_ & _04664_;
  assign _02594_ = _06970_ & _04664_;
  assign _02597_ = _06974_ & _04668_;
  assign _02600_ = _06978_ & _04668_;
  assign _02603_ = _06982_ & _04668_;
  assign _02606_ = _06986_ & _04668_;
  assign _02609_ = _06990_ & _04674_;
  assign _02612_ = _06994_ & _04674_;
  assign _02615_ = _06998_ & _04674_;
  assign _02618_ = _07002_ & _04674_;
  assign _02621_ = _07006_ & _04674_;
  assign _02624_ = _07010_ & _04674_;
  assign _02627_ = _07014_ & _04674_;
  assign _02630_ = _07018_ & _04674_;
  assign _02633_ = \cpuregs[0]_t0  & _04684_;
  assign _02636_ = \cpuregs[20]_t0  & _04684_;
  assign _02639_ = \cpuregs[22]_t0  & _04684_;
  assign _02642_ = \cpuregs[24]_t0  & _04684_;
  assign _02645_ = \cpuregs[26]_t0  & _04684_;
  assign _02648_ = \cpuregs[28]_t0  & _04684_;
  assign _02651_ = \cpuregs[30]_t0  & _04684_;
  assign _02654_ = \cpuregs[2]_t0  & _04684_;
  assign _02657_ = \cpuregs[4]_t0  & _04684_;
  assign _02660_ = \cpuregs[6]_t0  & _04684_;
  assign _02663_ = \cpuregs[8]_t0  & _04684_;
  assign _02666_ = \cpuregs[10]_t0  & _04684_;
  assign _02669_ = \cpuregs[12]_t0  & _04684_;
  assign _02672_ = \cpuregs[14]_t0  & _04684_;
  assign _02675_ = \cpuregs[16]_t0  & _04684_;
  assign _02678_ = \cpuregs[18]_t0  & _04684_;
  assign _02796_ = reg_next_pc_t0 & _04748_;
  assign _02799_ = _06608_ & _04752_;
  assign _02801_ = _06608_ & _04741_;
  assign _02804_ = _06608_ & _04747_;
  assign _02806_ = _06608_ & _04743_;
  assign _02809_ = _06608_ & _00670_;
  assign _02811_ = _07590_[4:0] & _04761_;
  assign _07141_ = _07139_ & _04764_;
  assign _07146_ = instr_lb_t0 & _04746_;
  assign _07149_ = instr_lh_t0 & _04746_;
  assign _02815_ = instr_jalr_t0 & _04743_;
  assign _02820_ = latched_store_t0 & _04768_;
  assign _02823_ = cpu_state_t0 & _04771_;
  assign _02825_ = cpu_state_t0 & _04772_;
  assign _02828_ = cpu_state_t0 & _04775_;
  assign _02830_ = cpu_state_t0 & _04776_;
  assign _02834_ = cpu_state_t0 & _04778_;
  assign _02836_ = _07172_ & _04779_;
  assign _02840_ = cpu_state_t0 & _04781_;
  assign _02843_ = _07180_ & _04784_;
  assign _02845_ = _07182_ & _04785_;
  assign _02847_ = _07180_ & _04786_;
  assign _07193_ = dbg_rs2val_t0 & _04789_;
  assign _02850_ = cpuregs_rs2_t0 & _04790_;
  assign _02853_ = _07193_ & _00669_;
  assign _07197_ = dbg_rs1val_t0 & _04789_;
  assign _02855_ = cpuregs_rs1_t0 & _04793_;
  assign _02858_ = _07197_ & _04161_;
  assign _02861_ = _07197_ & _00669_;
  assign _02863_ = mem_do_rinst_t0 & _04768_;
  assign _02865_ = decoder_trigger_t0 & _04766_;
  assign _02867_ = _07208_ & _04799_;
  assign _07212_ = _06217_ & _04800_;
  assign _07216_ = _06223_ & _04802_;
  assign _07219_ = _00099_ & _04803_;
  assign _07223_ = _00099_ & _04804_;
  assign _02869_ = _06239_ & _04805_;
  assign _07229_ = _07227_ & _04757_;
  assign _02872_ = _00091_ & _04314_;
  assign _02875_ = _00061_ & _04809_;
  assign _02878_ = _06612_ & _04768_;
  assign _02882_ = _00036_ & _04816_;
  assign _02888_ = _07240_ & _04820_;
  assign _02890_ = _07242_ & _04821_;
  assign _02893_ = _07244_ & _04824_;
  assign _02896_ = mem_rdata_latched_t0[11] & _04827_;
  assign _02900_ = _07257_ & _04830_;
  assign _02903_ = _07259_ & _04833_;
  assign _02912_ = mem_rdata_latched_t0[19] & _04841_;
  assign _02915_ = mem_rdata_latched_t0[30] & _04841_;
  assign _02918_ = mem_rdata_latched_t0[27] & _04841_;
  assign _02921_ = mem_rdata_latched_t0[26] & _04841_;
  assign _02924_ = mem_rdata_latched_t0[23:21] & _04847_;
  assign _02927_ = mem_rdata_latched_t0[25] & _04841_;
  assign _02930_ = mem_rdata_latched_t0[29:28] & _04851_;
  assign _02933_ = { mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31] } & _04854_;
  assign _02936_ = mem_rdata_latched_t0[24] & _04841_;
  assign _02939_ = mem_rdata_latched_t0[20] & _04841_;
  assign _02944_ = _07294_ & _04860_;
  assign _02946_ = _07296_ & _04861_;
  assign _02949_ = _07298_ & _04864_;
  assign _02952_ = mem_rdata_latched_t0[10:7] & _04867_;
  assign _02956_ = _07304_ & _04869_;
  assign _02959_ = _07306_ & _04872_;
  assign _02966_ = mem_rdata_latched_t0[18:15] & _04877_;
  assign _02969_ = _06558_ & _04820_;
  assign _02971_ = _07315_ & _04824_;
  assign _02973_ = _06558_ & _04245_;
  assign _02976_ = _06558_ & _04833_;
  assign _02980_ = _06558_ & _04841_;
  assign _02985_ = _06556_ & _04243_;
  assign _02988_ = _06556_ & _04828_;
  assign _02990_ = _07331_ & _04830_;
  assign _02992_ = _06556_ & _04836_;
  assign _02994_ = _06556_ & _04838_;
  assign _02999_ = _06556_ & _04841_;
  assign _03002_ = _06550_ & _04256_;
  assign _03004_ = _06550_ & _04294_;
  assign _03007_ = _06550_ & _04841_;
  assign _03010_ = _06554_ & _04373_;
  assign _03013_ = _06554_ & _04890_;
  assign _03015_ = _06554_ & _04841_;
  assign _03018_ = _06552_ & _04892_;
  assign _03020_ = _06552_ & _04893_;
  assign _03024_ = _06552_ & _04841_;
  assign _03029_ = _07366_ & _04898_;
  assign _03032_ = mem_rdata_latched_t0[6:2] & _04901_;
  assign _03036_ = _07371_ & _04903_;
  assign _03044_ = mem_rdata_latched_t0[24:20] & _04906_;
  assign _03047_ = mem_rdata_latched_t0[19:12] & _04909_;
  assign _03052_ = _07381_ & _04912_;
  assign _03054_ = _07383_ & _04898_;
  assign _03059_ = mem_rdata_latched_t0[11:7] & _04901_;
  assign _03063_ = _07390_ & _04915_;
  assign _03066_ = _07392_ & _04903_;
  assign _03073_ = mem_rdata_latched_t0[11:7] & _04906_;
  assign _03076_ = _06676_ & _04818_;
  assign _03078_ = _07402_ & _04821_;
  assign _03080_ = _06676_ & _04245_;
  assign _03083_ = _06676_ & _04248_;
  assign _03086_ = _06676_ & _04841_;
  assign _03089_ = _06544_ & _04924_;
  assign _03091_ = _06544_ & _04294_;
  assign _03094_ = _06544_ & _04841_;
  assign _03099_ = _06540_ & _04838_;
  assign _03102_ = _06540_ & _04259_;
  assign _03105_ = _06540_ & _04294_;
  assign _03108_ = _06540_ & _04841_;
  assign _03111_ = decoded_rs2_t0 & _04931_;
  assign _03114_ = decoded_rs1_t0 & _04931_;
  assign _03117_ = _00063_ & _04935_;
  assign _03120_ = q_insn_rs2_t0 & _04938_;
  assign _03123_ = q_insn_rs1_t0 & _04938_;
  assign _03126_ = { rvfi_insn_t0[31:25], 5'h00, rvfi_insn_t0[19:15], 3'h0, rvfi_insn_t0[11:0] } & _04942_;
  assign _03129_ = { 16'h0000, next_insn_opcode_t0[15:0] } & _04945_;
  assign _07434_ = _07432_ & _04949_;
  assign _07436_ = mem_rdata_t0[31:16] & _04950_;
  assign _03132_ = _07434_ & _04951_;
  assign _07446_ = { _06877_, _06877_ } & _04955_;
  assign _03136_ = _06372_ & _04956_;
  assign _03138_ = mem_wstrb_t0 & _04957_;
  assign _03141_ = _07453_ & _04960_;
  assign _03143_ = _07453_ & _04961_;
  assign _03146_ = _07464_ & _04745_;
  assign _03148_ = _06376_ & _04967_;
  assign _03150_ = mem_rdata_q_t0[31] & _04965_;
  assign _03153_ = _07468_ & _04969_;
  assign _03155_ = _07469_ & _04820_;
  assign _03157_ = _07470_ & _04821_;
  assign _03159_ = _07471_ & _04824_;
  assign _03161_ = _07468_ & _04970_;
  assign _03163_ = _07474_ & _04971_;
  assign _03165_ = _07476_ & _04830_;
  assign _03168_ = _07478_ & _04833_;
  assign _03170_ = _07468_ & _04364_;
  assign _03172_ = _07468_ & _04973_;
  assign _03175_ = mem_rdata_q_t0[7] & _04965_;
  assign _03178_ = _07483_ & _04890_;
  assign _03180_ = _07483_ & _04256_;
  assign _03183_ = _07483_ & _04973_;
  assign _03186_ = mem_rdata_q_t0[24:20] & _04979_;
  assign _03189_ = _07488_ & _04982_;
  assign _03191_ = _07489_ & _04912_;
  assign _03193_ = _07488_ & _04915_;
  assign _03196_ = { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] } & _04984_;
  assign _03199_ = _07488_ & _04987_;
  assign _03202_ = mem_rdata_q_t0[19:15] & _04979_;
  assign _03205_ = { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[6:5] } & _04984_;
  assign _03208_ = _07497_ & _04992_;
  assign _03211_ = _07497_ & _04995_;
  assign _03214_ = _07497_ & _04987_;
  assign _03217_ = mem_rdata_q_t0[14:12] & _04999_;
  assign _03220_ = _07504_ & _05002_;
  assign _03222_ = _07505_ & _05003_;
  assign _03224_ = _07506_ & _05004_;
  assign _03226_ = _07507_ & _05005_;
  assign _03228_ = _07504_ & _05006_;
  assign _03230_ = _07511_ & _05007_;
  assign _03232_ = _07513_ & _05008_;
  assign _03234_ = _07514_ & _05009_;
  assign _03236_ = _07516_ & _05010_;
  assign _03238_ = _07518_ & _05011_;
  assign _03240_ = _07520_ & _05012_;
  assign _03242_ = _07514_ & _05013_;
  assign _03245_ = mem_rdata_latched_t0[4:2] & _05016_;
  assign _03247_ = _07504_ & _05017_;
  assign _03250_ = mem_rdata_q_t0[11:8] & _05020_;
  assign _03253_ = _07528_ & _04265_;
  assign _03256_ = _07528_ & _04282_;
  assign _03261_ = _07528_ & _05026_;
  assign _03264_ = mem_rdata_q_t0[30:25] & _05029_;
  assign _03267_ = _07535_ & _05032_;
  assign _03269_ = _07536_ & _05033_;
  assign _03271_ = _07537_ & _05034_;
  assign _03273_ = _07538_ & _05035_;
  assign _03275_ = _07535_ & _05036_;
  assign _03277_ = _07542_ & _05037_;
  assign _03279_ = _07544_ & _05038_;
  assign _03282_ = _07546_ & _05041_;
  assign _03285_ = { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] } & _05044_;
  assign _03288_ = _07535_ & _05047_;
  assign _03292_ = mem_la_firstword_t0 & _05050_;
  assign _03295_ = _00054_ & _05053_;
  assign _03298_ = { 32'h00000000, _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31] } & _05053_;
  assign _03302_ = _00050_ & _05057_;
  assign _03305_ = { 32'h00000000, _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31] } & _05057_;
  assign _03325_ = reg_next_pc_t0 & _05069_;
  assign _03328_ = _00085_ & _05072_;
  assign _03335_ = reg_next_pc_t0 & _05077_;
  assign _03338_ = reg_out_t0 & _05080_;
  assign _03341_ = reg_pc_t0 & _05083_;
  assign _03345_ = { pcpi_rs1_t0[31:2], 2'h0 } & _05085_;
  assign _03348_ = mem_rdata_q_t0 & _05088_;
  assign _03351_ = _07605_ & _05091_;
  assign _03354_ = mem_rdata_latched_noshuffle_t0 & _05094_;
  assign _03357_ = _07603_ & _05097_;
  assign _01328_ = _07377_ & _03982_;
  assign _01331_ = { _07275_, _07313_ } & _03982_;
  assign _01572_ = _07127_ & _04074_;
  assign _01575_ = _07123_ & _04077_;
  assign _01578_ = { mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15:0] } & _04080_;
  assign _01581_ = { mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7:0] } & _04083_;
  assign _01584_ = _07131_ & _04086_;
  assign _01587_ = _07137_ & _04089_;
  assign _01590_ = _00097_ & _04092_;
  assign _01593_ = _06115_ & _04095_;
  assign _01596_ = _06129_ & _04098_;
  assign _01599_ = count_instr_t0[63:32] & _04101_;
  assign _01602_ = count_cycle_t0[63:32] & _04104_;
  assign _01605_ = _06125_ & _04107_;
  assign _01608_ = cpuregs_rs2_t0[4:0] & _04110_;
  assign _01611_ = _07141_ & _04113_;
  assign _01614_ = decoded_rs2_t0 & _04116_;
  assign _01618_ = _07147_ & _04072_;
  assign _01620_ = _07150_ & _04072_;
  assign _01623_ = _07152_ & _04074_;
  assign _01627_ = _06156_ & _04123_;
  assign _01630_ = _07160_ & _04125_;
  assign _01633_ = _06149_ & _04128_;
  assign _01638_ = _07166_ & _04132_;
  assign _01641_ = _07164_ & _04135_;
  assign _01644_ = _06173_ & _04138_;
  assign _01647_ = _07178_ & _04141_;
  assign _01650_ = _06162_ & _04144_;
  assign _01653_ = _06160_ & _04147_;
  assign _01655_ = _07174_ & _04151_;
  assign _01658_ = { 5'h00, is_sll_srl_sra_t0, is_sll_srl_sra_t0, 1'h0 } & _04153_;
  assign _01669_ = _06179_ & _04159_;
  assign _01672_ = _07195_ & _04162_;
  assign _01675_ = cpuregs_rs2_t0 & _04089_;
  assign _01678_ = _07203_ & _04166_;
  assign _01681_ = _06214_ & _04123_;
  assign _01684_ = _06193_ & _04170_;
  assign _01687_ = _07205_ & _04174_;
  assign _06208_ = mem_do_prefetch_t0 & _04178_;
  assign _01698_ = _06208_ & _04182_;
  assign _01702_ = _07217_ & _04185_;
  assign _01705_ = _07214_ & _04187_;
  assign _01712_ = decoded_imm_t0 & _04193_;
  assign _01715_ = _07221_ & _04086_;
  assign _01718_ = _07229_ & _04197_;
  assign _01721_ = _06231_ & _04200_;
  assign _01724_ = { 1'h0, pcpi_rs1_t0[31:1] } & _04203_;
  assign _01727_ = { 1'h0, pcpi_rs1_t0[31:1] } & _04206_;
  assign _01730_ = { 4'h0, pcpi_rs1_t0[31:4] } & _04203_;
  assign _01733_ = { 1'h0, pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31:4] } & _04206_;
  assign _01736_ = _07598_ & _04211_;
  assign _01739_ = { _00111_[31:1], _07593_[0] } & _04214_;
  assign _01742_ = _00109_ & _04217_;
  assign _01745_ = { 31'h00000000, alu_out_0_t0 } & _04220_;
  assign _01748_ = _07610_ & _04223_;
  assign _01751_ = _06249_ & _04226_;
  assign _01754_ = alu_lts_t0 & _04229_;
  assign _01757_ = alu_ltu_t0 & _04232_;
  assign _01760_ = alu_eq_t0 & _04235_;
  assign _01763_ = alu_lts_t0 & _04238_;
  assign _01766_ = _06257_ & _04241_;
  assign _01768_ = _07249_ & _04244_;
  assign _01771_ = _07246_ & _04246_;
  assign _01774_ = _06265_ & _04249_;
  assign _01776_ = _07269_ & _04252_;
  assign _01779_ = _06267_ & _04254_;
  assign _01782_ = _00107_[4] & _04257_;
  assign _01784_ = mem_rdata_latched_t0[11] & _04244_;
  assign _01787_ = _07264_ & _04260_;
  assign _01790_ = _06273_ & _04263_;
  assign _01794_ = _07302_ & _04267_;
  assign _01797_ = { 2'h0, _07091_, 1'h0 } & _04269_;
  assign _01800_ = _06281_ & _04272_;
  assign _01803_ = _06287_ & _04275_;
  assign _01805_ = _06304_ & _04278_;
  assign _01808_ = _06289_ & _04280_;
  assign _01811_ = _00107_[3:0] & _04283_;
  assign _01813_ = mem_rdata_latched_t0[10:7] & _04267_;
  assign _01816_ = _07311_ & _04286_;
  assign _01819_ = _06295_ & _04289_;
  assign _01822_ = _00107_[3:0] & _04292_;
  assign _01825_ = _07323_ & _04295_;
  assign _01828_ = _07319_ & _04249_;
  assign _01831_ = _07329_ & _04249_;
  assign _01834_ = _07339_ & _04252_;
  assign _01837_ = _06310_ & _04254_;
  assign _01840_ = _07333_ & _04246_;
  assign _01845_ = _06316_ & _04304_;
  assign _01848_ = _07359_ & _04252_;
  assign _01851_ = _07357_ & _04249_;
  assign _01854_ = { mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[7], mem_rdata_q_t0[30:25], mem_rdata_q_t0[11:8], 1'h0 } & _04309_;
  assign _01857_ = { mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31:25], mem_rdata_q_t0[11:7] } & _04312_;
  assign _01859_ = { decoded_imm_j_t0[31:1], 1'h0 } & _04315_;
  assign _01862_ = { mem_rdata_q_t0[31:12], 12'h000 } & _04317_;
  assign _01865_ = _06328_ & _04320_;
  assign _01868_ = mem_rdata_latched_t0[6:2] & _04323_;
  assign _01870_ = _07369_ & _04326_;
  assign _01873_ = _06336_ & _04328_;
  assign _01876_ = _06340_ & _04331_;
  assign _01878_ = _07375_ & _04334_;
  assign _01881_ = _06342_ & _04336_;
  assign _01884_ = _07385_ & _04339_;
  assign _01886_ = _07388_ & _04326_;
  assign _01889_ = _06348_ & _04342_;
  assign _01892_ = _06352_ & _04331_;
  assign _01894_ = _07398_ & _04334_;
  assign _01897_ = _06354_ & _04336_;
  assign _01900_ = _07394_ & _04339_;
  assign _01903_ = mem_rdata_latched_t0[11:7] & _04348_;
  assign _01906_ = _06360_ & _04351_;
  assign _01909_ = _07448_ & _04354_;
  assign _01912_ = _06368_ & _04357_;
  assign _01915_ = _07462_ & _04360_;
  assign _01920_ = _07473_ & _04246_;
  assign _01925_ = _06379_ & _04249_;
  assign _01928_ = _07482_ & _04252_;
  assign _01931_ = _06381_ & _04254_;
  assign _01933_ = _07480_ & _04246_;
  assign _01936_ = mem_rdata_latched_t0[12] & _04370_;
  assign _01939_ = _07487_ & _04295_;
  assign _01942_ = _07485_ & _04374_;
  assign _01945_ = { mem_rdata_latched_t0[6:4], 2'h0 } & _04377_;
  assign _01948_ = _07491_ & _04339_;
  assign _01951_ = _06397_ & _04331_;
  assign _01954_ = _06413_ & _04334_;
  assign _01957_ = _06399_ & _04336_;
  assign _01960_ = _07493_ & _04339_;
  assign _01963_ = mem_rdata_latched_t0[6:2] & _04348_;
  assign _01966_ = _06405_ & _04351_;
  assign _01969_ = { mem_rdata_latched_t0[11], mem_rdata_latched_t0[5], mem_rdata_latched_t0[6], 2'h0 } & _04326_;
  assign _01972_ = { mem_rdata_latched_t0[11:10], mem_rdata_latched_t0[6], 2'h0 } & _04377_;
  assign _01979_ = _06415_ & _04391_;
  assign _01982_ = _06419_ & _04394_;
  assign _01985_ = _06437_ & _04397_;
  assign _01988_ = _06421_ & _04400_;
  assign _01991_ = _07526_ & _04403_;
  assign _01994_ = _07524_ & _04406_;
  assign _01997_ = { 2'h0, _06427_[0] } & _04409_;
  assign _02003_ = _07530_ & _04275_;
  assign _02006_ = _07534_ & _04278_;
  assign _02009_ = _06439_ & _04280_;
  assign _02012_ = { 3'h0, mem_rdata_latched_t0[8:7], mem_rdata_latched_t0[12] } & _04415_;
  assign _02017_ = { 3'h0, mem_rdata_latched_t0[3:2], mem_rdata_latched_t0[12] } & _04420_;
  assign _02020_ = _06445_ & _04423_;
  assign _02023_ = _06451_ & _04426_;
  assign _02026_ = _06469_ & _04429_;
  assign _02029_ = _06453_ & _04432_;
  assign _02032_ = { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[6:5], mem_rdata_latched_t0[2] } & _04435_;
  assign _02035_ = { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] } & _04438_;
  assign _02038_ = _07550_ & _04441_;
  assign _02041_ = _06459_ & _04444_;
  assign _02043_ = { 1'h0, mem_rdata_latched_t0[10:7], mem_rdata_latched_t0[12] } & _04418_;
  assign _02046_ = { 4'h0, mem_rdata_latched_t0[5], mem_rdata_latched_t0[12] } & _04448_;
  assign _02049_ = { 24'h000000, mem_rdata_t0[31:24] } & _04451_;
  assign _02052_ = { 24'h000000, mem_rdata_t0[15:8] } & _04454_;
  assign _02055_ = _06471_ & _04457_;
  assign _02058_ = { 16'h0000, mem_rdata_t0[31:16] } & _04460_;
  assign _02061_ = _00048_ & _04463_;
  assign _02064_ = _00065_ & _04466_;
  assign _02066_ = { pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1] } & _04468_;
  assign _02069_ = _07582_ & _04470_;
  assign _02072_ = { pcpi_rs2_t0[15:0], pcpi_rs2_t0[15:0] } & _04463_;
  assign _02075_ = { pcpi_rs2_t0[7:0], pcpi_rs2_t0[7:0], pcpi_rs2_t0[7:0], pcpi_rs2_t0[7:0] } & _04466_;
  assign _02078_ = pcpi_div_rd_t0 & _04475_;
  assign _02080_ = pcpi_mul_wr_t0 & _04477_;
  assign _02083_ = pcpi_div_wr_t0 & _04479_;
  assign _02496_ = _06904_ & _04621_;
  assign _02499_ = _06908_ & _04624_;
  assign _02502_ = _06912_ & _04624_;
  assign _02505_ = _06916_ & _04628_;
  assign _02508_ = _06920_ & _04628_;
  assign _02511_ = _06924_ & _04628_;
  assign _02514_ = _06928_ & _04628_;
  assign _02517_ = _06932_ & _04634_;
  assign _02520_ = _06936_ & _04634_;
  assign _02523_ = _06940_ & _04634_;
  assign _02526_ = _06944_ & _04634_;
  assign _02529_ = _06948_ & _04634_;
  assign _02532_ = _06952_ & _04634_;
  assign _02535_ = _06956_ & _04634_;
  assign _02538_ = _06960_ & _04634_;
  assign _02541_ = \cpuregs[1]_t0  & _04644_;
  assign _02544_ = \cpuregs[21]_t0  & _04644_;
  assign _02547_ = \cpuregs[23]_t0  & _04644_;
  assign _02550_ = \cpuregs[25]_t0  & _04644_;
  assign _02553_ = \cpuregs[27]_t0  & _04644_;
  assign _02556_ = \cpuregs[29]_t0  & _04644_;
  assign _02559_ = \cpuregs[31]_t0  & _04644_;
  assign _02562_ = \cpuregs[3]_t0  & _04644_;
  assign _02565_ = \cpuregs[5]_t0  & _04644_;
  assign _02568_ = \cpuregs[7]_t0  & _04644_;
  assign _02571_ = \cpuregs[9]_t0  & _04644_;
  assign _02574_ = \cpuregs[11]_t0  & _04644_;
  assign _02577_ = \cpuregs[13]_t0  & _04644_;
  assign _02580_ = \cpuregs[15]_t0  & _04644_;
  assign _02583_ = \cpuregs[17]_t0  & _04644_;
  assign _02586_ = \cpuregs[19]_t0  & _04644_;
  assign _02589_ = _06964_ & _04662_;
  assign _02592_ = _06968_ & _04665_;
  assign _02595_ = _06972_ & _04665_;
  assign _02598_ = _06976_ & _04669_;
  assign _02601_ = _06980_ & _04669_;
  assign _02604_ = _06984_ & _04669_;
  assign _02607_ = _06988_ & _04669_;
  assign _02610_ = _06992_ & _04675_;
  assign _02613_ = _06996_ & _04675_;
  assign _02616_ = _07000_ & _04675_;
  assign _02619_ = _07004_ & _04675_;
  assign _02622_ = _07008_ & _04675_;
  assign _02625_ = _07012_ & _04675_;
  assign _02628_ = _07016_ & _04675_;
  assign _02631_ = _07020_ & _04675_;
  assign _02634_ = \cpuregs[1]_t0  & _04685_;
  assign _02637_ = \cpuregs[21]_t0  & _04685_;
  assign _02640_ = \cpuregs[23]_t0  & _04685_;
  assign _02643_ = \cpuregs[25]_t0  & _04685_;
  assign _02646_ = \cpuregs[27]_t0  & _04685_;
  assign _02649_ = \cpuregs[29]_t0  & _04685_;
  assign _02652_ = \cpuregs[31]_t0  & _04685_;
  assign _02655_ = \cpuregs[3]_t0  & _04685_;
  assign _02658_ = \cpuregs[5]_t0  & _04685_;
  assign _02661_ = \cpuregs[7]_t0  & _04685_;
  assign _02664_ = \cpuregs[9]_t0  & _04685_;
  assign _02667_ = \cpuregs[11]_t0  & _04685_;
  assign _02670_ = \cpuregs[13]_t0  & _04685_;
  assign _02673_ = \cpuregs[15]_t0  & _04685_;
  assign _02676_ = \cpuregs[17]_t0  & _04685_;
  assign _02679_ = \cpuregs[19]_t0  & _04685_;
  assign _02783_ = _00071_ & _04736_;
  assign _02785_ = _00073_ & _04736_;
  assign _02787_ = _00067_ & _04736_;
  assign _02789_ = _00069_ & _04736_;
  assign _07099_ = mem_wdata_t0 & _04737_;
  assign _07101_ = mem_rdata_t0 & _04737_;
  assign _07103_ = mem_wstrb_t0 & _04738_;
  assign _07105_ = { _07571_, _07571_, _07571_, _07571_ } & _04738_;
  assign _07107_ = mem_addr_t0 & _04737_;
  assign _02791_ = _07600_ & _04739_;
  assign _02793_ = latched_rd_t0 & _04740_;
  assign _02795_ = alu_out_0_t0 & _04744_;
  assign _02797_ = _07595_ & _04749_;
  assign _07118_ = _07116_ & _04751_;
  assign _00061_ = _07118_ & { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn };
  assign _02802_ = _07121_ & _04742_;
  assign _02807_ = _07125_ & _04744_;
  assign _02810_ = _06109_ & resetn;
  assign _07129_ = _06113_ & _04755_;
  assign _07131_ = _07129_ & _04756_;
  assign _07133_ = pcpi_rs1_t0 & _04758_;
  assign _07137_ = _07135_ & _04759_;
  assign _07135_ = pcpi_int_rd_t0 & _04760_;
  assign _00027_ = _06121_ & { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn };
  assign _02812_ = _07588_[4:0] & _04762_;
  assign _00029_ = _06133_ & { resetn, resetn, resetn, resetn, resetn };
  assign _07147_ = _07146_ & _04742_;
  assign _07150_ = _07149_ & _04742_;
  assign _02817_ = instr_jal_t0 & _04767_;
  assign _07160_ = _07158_ & _04174_;
  assign _02821_ = pcpi_int_wr_t0 & _04769_;
  assign _02826_ = _07162_ & _04773_;
  assign _02832_ = _07168_ & _04777_;
  assign _02838_ = cpu_state_t0 & _04780_;
  assign _02841_ = _07176_ & _04782_;
  assign _07180_ = _06168_ & { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn };
  assign _02848_ = _07184_ & _04787_;
  assign _02851_ = _07193_ & _04791_;
  assign _02854_ = _06191_ & { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn };
  assign _02856_ = _07197_ & _04794_;
  assign _02859_ = _07199_ & _04162_;
  assign _02862_ = _07201_ & { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn };
  assign _07203_ = mem_do_prefetch_t0 & _04797_;
  assign _07208_ = _06197_ & resetn;
  assign _07214_ = _07212_ & _04801_;
  assign _07217_ = _07216_ & _04801_;
  assign _07221_ = _07219_ & _04756_;
  assign _07225_ = _07223_ & _04756_;
  assign _02870_ = _06243_ & _04806_;
  assign _02873_ = _00095_ & _04315_;
  assign _02876_ = _07231_ & _04810_;
  assign _07239_ = _07237_ & _04812_;
  assign _07237_ = _07235_ & _04174_;
  assign _00003_ = cpuregs_wrdata_t0 & _04813_;
  assign _00001_ = latched_rd_t0 & _04814_;
  assign cpuregs_wrdata_t0 = _00038_ & _04751_;
  assign _02880_ = _00040_ & _04815_;
  assign _02884_ = clear_prefetched_high_word_q_t0 & _04817_;
  assign _02886_ = mem_rdata_latched_t0[11] & _04819_;
  assign _02891_ = mem_rdata_latched_t0[11] & _04822_;
  assign _02894_ = mem_rdata_latched_t0[11] & _04825_;
  assign _02898_ = _00107_[4] & _04829_;
  assign _02901_ = _00107_[4] & _04831_;
  assign _02904_ = _00107_[4] & _04834_;
  assign _02906_ = mem_rdata_latched_t0[11] & _04837_;
  assign _02908_ = _07262_ & _04839_;
  assign _02910_ = _00107_[4] & _04840_;
  assign _02913_ = _06271_ & _04842_;
  assign _02916_ = mem_rdata_latched_t0[8] & _04842_;
  assign _02919_ = mem_rdata_latched_t0[6] & _04842_;
  assign _02922_ = mem_rdata_latched_t0[7] & _04842_;
  assign _02925_ = mem_rdata_latched_t0[5:3] & _04848_;
  assign _02928_ = mem_rdata_latched_t0[2] & _04842_;
  assign _02931_ = mem_rdata_latched_t0[10:9] & _04852_;
  assign _02934_ = { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] } & _04855_;
  assign _02937_ = mem_rdata_latched_t0[11] & _04842_;
  assign _02940_ = mem_rdata_latched_t0[12] & _04842_;
  assign _02942_ = mem_rdata_latched_t0[10:7] & _04859_;
  assign _02947_ = mem_rdata_latched_t0[10:7] & _04862_;
  assign _02950_ = mem_rdata_latched_t0[10:7] & _04865_;
  assign _02954_ = _00107_[3:0] & _04868_;
  assign _02957_ = _00107_[3:0] & _04870_;
  assign _02960_ = _00107_[3:0] & _04873_;
  assign _02962_ = mem_rdata_latched_t0[10:7] & _04875_;
  assign _02964_ = _07309_ & _04876_;
  assign _02967_ = _06293_ & _04878_;
  assign _02974_ = _07317_ & _04246_;
  assign _02978_ = _07321_ & _04246_;
  assign _02981_ = _06308_ & _04842_;
  assign _02983_ = _06556_ & _00508_;
  assign _02986_ = _07327_ & _04244_;
  assign _02995_ = _07335_ & _04839_;
  assign _02997_ = _07576_ & _04244_;
  assign _03000_ = _06314_ & _04842_;
  assign _03005_ = _07343_ & _04295_;
  assign _03008_ = _07345_ & _04842_;
  assign _03011_ = _07349_ & _04374_;
  assign _03016_ = _07351_ & _04842_;
  assign _03021_ = _07355_ & _04894_;
  assign _03025_ = _06324_ & _04842_;
  assign _03027_ = mem_rdata_latched_t0[6:2] & _04897_;
  assign _03030_ = mem_rdata_latched_t0[6:2] & _04899_;
  assign _03034_ = mem_rdata_latched_t0[6:2] & _04902_;
  assign _03037_ = _00105_[4:0] & _04904_;
  assign _03039_ = _07372_ & _04339_;
  assign _03041_ = _00105_[4:0] & _04323_;
  assign _03045_ = _06346_ & _04907_;
  assign _03048_ = { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] } & _04910_;
  assign _03050_ = mem_rdata_latched_t0[11:7] & _04897_;
  assign _03055_ = mem_rdata_latched_t0[11:7] & _04899_;
  assign _03057_ = mem_rdata_latched_t0[11:7] & _04914_;
  assign _03061_ = _00107_[4:0] & _04902_;
  assign _03064_ = _00107_[4:0] & _04916_;
  assign _03067_ = _00107_[4:0] & _04904_;
  assign _03069_ = mem_rdata_latched_t0[11:7] & _04919_;
  assign _03071_ = _00105_[4:0] & _04348_;
  assign _03074_ = _06358_ & _04907_;
  assign _03081_ = _07404_ & _04246_;
  assign _03084_ = _07406_ & _04249_;
  assign _03087_ = _07408_ & _04842_;
  assign _03092_ = _07412_ & _04295_;
  assign _03095_ = _07416_ & _04842_;
  assign _03097_ = _06540_ & _04837_;
  assign _03100_ = _07420_ & _04839_;
  assign _03103_ = _07422_ & _04260_;
  assign _03106_ = _07424_ & _04295_;
  assign _03109_ = _07426_ & _04842_;
  assign _03112_ = cached_insn_rs2_t0 & _04932_;
  assign _03115_ = cached_insn_rs1_t0 & _04932_;
  assign _03118_ = cached_insn_opcode_t0 & _04936_;
  assign _03121_ = _00046_ & _04939_;
  assign _03124_ = _00044_ & _04939_;
  assign _03127_ = _00042_ & _04943_;
  assign _03130_ = next_insn_opcode_t0 & _04946_;
  assign _07432_ = mem_rdata_t0[31:16] & _04948_;
  assign _03133_ = _07436_ & _04952_;
  assign _07448_ = _07446_ & _04954_;
  assign _03139_ = _00113_ & _04958_;
  assign _03144_ = _07455_ & _04962_;
  assign _07459_ = _06634_ & _04964_;
  assign _07462_ = mem_la_read_t0 & _04966_;
  assign _07464_ = mem_la_use_prefetched_high_word_t0 & _04964_;
  assign _03151_ = mem_rdata_latched_t0[31] & _04966_;
  assign _03166_ = mem_rdata_latched_t0[12] & _04831_;
  assign _03173_ = _06385_ & _04974_;
  assign _03176_ = mem_rdata_latched_t0[7] & _04966_;
  assign _03181_ = mem_rdata_latched_t0[12] & _04257_;
  assign _03184_ = _06393_ & _04974_;
  assign _03187_ = mem_rdata_latched_t0[24:20] & _04980_;
  assign _03194_ = mem_rdata_latched_t0[6:2] & _04916_;
  assign _03197_ = { mem_rdata_latched_t0[6], 4'h0 } & _04985_;
  assign _03200_ = _06403_ & _04988_;
  assign _03203_ = mem_rdata_latched_t0[19:15] & _04980_;
  assign _03206_ = _07497_ & _04985_;
  assign _03209_ = _07499_ & _04993_;
  assign _03212_ = _07501_ & _04996_;
  assign _03215_ = _07503_ & _04988_;
  assign _03218_ = mem_rdata_latched_t0[14:12] & _05000_;
  assign _03243_ = _07522_ & _05014_;
  assign _03248_ = _06425_ & _05018_;
  assign _03251_ = mem_rdata_latched_t0[11:8] & _05021_;
  assign _03254_ = { mem_rdata_latched_t0[11:9], 1'h0 } & _04266_;
  assign _03257_ = { mem_rdata_latched_t0[11:10], mem_rdata_latched_t0[4:3] } & _04283_;
  assign _03259_ = { mem_rdata_latched_t0[11:10], mem_rdata_latched_t0[6], 1'h0 } & _04266_;
  assign _03262_ = _06443_ & _05027_;
  assign _03265_ = mem_rdata_latched_t0[30:25] & _05030_;
  assign _03280_ = { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] } & _05039_;
  assign _03283_ = { _06526_, 5'h00 } & _05042_;
  assign _03286_ = { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[4:3], mem_rdata_latched_t0[5], mem_rdata_latched_t0[2] } & _05045_;
  assign _03289_ = _06457_ & _05048_;
  assign _03293_ = mem_la_firstword_reg_t0 & _05051_;
  assign _03296_ = { rvfi_rd_wdata_t0, 32'h00000000 } & _05054_;
  assign _03300_ = { 32'h00000000, rvfi_rd_wdata_t0 } & _05056_;
  assign _03303_ = { rvfi_rd_wdata_t0, 32'h00000000 } & _05058_;
  assign _03307_ = { 32'h00000000, rvfi_rd_wdata_t0 } & _04735_;
  assign _03326_ = { reg_out_t0[31:1], 1'h0 } & _05070_;
  assign _03329_ = _07584_ & _05073_;
  assign _03331_ = _07085_ & _05075_;
  assign _03333_ = _07086_ & _05076_;
  assign _03336_ = { _00111_[31:1], 1'h0 } & _05078_;
  assign _03339_ = alu_out_q_t0 & _05081_;
  assign _03343_ = cpuregs_wrdata_t0 & _05084_;
  assign _03346_ = { _00103_, 2'h0 } & _05086_;
  assign _03349_ = mem_rdata_t0 & _05089_;
  assign _03352_ = { 16'h0000, mem_16bit_buffer_t0 } & _05092_;
  assign _03355_ = { 16'h0000, mem_rdata_latched_noshuffle_t0[31:16] } & _05095_;
  assign _03358_ = { mem_rdata_latched_noshuffle_t0[15:0], mem_16bit_buffer_t0 } & _05098_;
  assign _03983_ = _01327_ | _01328_;
  assign _03984_ = _01330_ | _01331_;
  assign _04075_ = _01571_ | _01572_;
  assign _04078_ = _01574_ | _01575_;
  assign _04081_ = _01577_ | _01578_;
  assign _04084_ = _01580_ | _01581_;
  assign _04087_ = _01583_ | _01584_;
  assign _04090_ = _01586_ | _01587_;
  assign _04093_ = _01589_ | _01590_;
  assign _04096_ = _01592_ | _01593_;
  assign _04099_ = _01595_ | _01596_;
  assign _04102_ = _01598_ | _01599_;
  assign _04105_ = _01601_ | _01602_;
  assign _04108_ = _01604_ | _01605_;
  assign _04111_ = _01607_ | _01608_;
  assign _04114_ = _01610_ | _01611_;
  assign _04117_ = _01613_ | _01614_;
  assign _04120_ = _01622_ | _01623_;
  assign _04126_ = _01629_ | _01630_;
  assign _04129_ = _01632_ | _01633_;
  assign _04133_ = _01637_ | _01638_;
  assign _04136_ = _01640_ | _01641_;
  assign _04139_ = _01643_ | _01644_;
  assign _04142_ = _01646_ | _01647_;
  assign _04145_ = _01649_ | _01650_;
  assign _04148_ = _01652_ | _01653_;
  assign _04154_ = _01657_ | _01658_;
  assign _04156_ = _01664_ | _01655_;
  assign _04160_ = _01668_ | _01669_;
  assign _04163_ = _01671_ | _01672_;
  assign _04164_ = _01674_ | _01675_;
  assign _04167_ = _01677_ | _01678_;
  assign _04168_ = _01680_ | _01681_;
  assign _04171_ = _01683_ | _01684_;
  assign _04175_ = _01686_ | _01687_;
  assign _04179_ = _01693_ | _01687_;
  assign _04183_ = _01697_ | _01698_;
  assign _04188_ = _01704_ | _01705_;
  assign _04190_ = _01709_ | _01675_;
  assign _04194_ = _01711_ | _01712_;
  assign _04195_ = _01714_ | _01715_;
  assign _04198_ = _01717_ | _01718_;
  assign _04201_ = _01720_ | _01721_;
  assign _04204_ = _01723_ | _01724_;
  assign _04207_ = _01726_ | _01727_;
  assign _04208_ = _01729_ | _01730_;
  assign _04209_ = _01732_ | _01733_;
  assign _04212_ = _01735_ | _01736_;
  assign _04215_ = _01738_ | _01739_;
  assign _04218_ = _01741_ | _01742_;
  assign _04221_ = _01744_ | _01745_;
  assign _04224_ = _01747_ | _01748_;
  assign _04227_ = _01750_ | _01751_;
  assign _04230_ = _01753_ | _01754_;
  assign _04233_ = _01756_ | _01757_;
  assign _04236_ = _01759_ | _01760_;
  assign _04239_ = _01762_ | _01763_;
  assign _04242_ = _01765_ | _01766_;
  assign _04247_ = _01770_ | _01771_;
  assign _04250_ = _01773_ | _01774_;
  assign _04255_ = _01778_ | _01779_;
  assign _04258_ = _01781_ | _01782_;
  assign _04261_ = _01786_ | _01787_;
  assign _04264_ = _01789_ | _01790_;
  assign _04270_ = _01796_ | _01797_;
  assign _04273_ = _01799_ | _01800_;
  assign _04276_ = _01802_ | _01803_;
  assign _04281_ = _01807_ | _01808_;
  assign _04284_ = _01810_ | _01811_;
  assign _04287_ = _01815_ | _01816_;
  assign _04290_ = _01818_ | _01819_;
  assign _04293_ = _01821_ | _01822_;
  assign _04296_ = _01824_ | _01825_;
  assign _04297_ = _01827_ | _01828_;
  assign _04298_ = _01830_ | _01831_;
  assign _04299_ = _01833_ | _01834_;
  assign _04300_ = _01836_ | _01837_;
  assign _04301_ = _01839_ | _01840_;
  assign _04305_ = _01844_ | _01845_;
  assign _04306_ = _01847_ | _01848_;
  assign _04307_ = _01850_ | _01851_;
  assign _04310_ = _01853_ | _01854_;
  assign _04313_ = _01856_ | _01857_;
  assign _04318_ = _01861_ | _01862_;
  assign _04321_ = _01864_ | _01865_;
  assign _04324_ = _01867_ | _01868_;
  assign _04329_ = _01872_ | _01873_;
  assign _04332_ = _01875_ | _01876_;
  assign _04337_ = _01880_ | _01881_;
  assign _04340_ = _01883_ | _01884_;
  assign _04343_ = _01888_ | _01889_;
  assign _04344_ = _01891_ | _01892_;
  assign _04345_ = _01896_ | _01897_;
  assign _04346_ = _01899_ | _01900_;
  assign _04349_ = _01902_ | _01903_;
  assign _04352_ = _01905_ | _01906_;
  assign _04355_ = _01908_ | _01909_;
  assign _04358_ = _01911_ | _01912_;
  assign _04361_ = _01914_ | _01915_;
  assign _04363_ = _01919_ | _01920_;
  assign _04365_ = _01924_ | _01925_;
  assign _04366_ = _01927_ | _01928_;
  assign _04367_ = _01930_ | _01931_;
  assign _04368_ = _01919_ | _01933_;
  assign _04371_ = _01935_ | _01936_;
  assign _04372_ = _01938_ | _01939_;
  assign _04375_ = _01941_ | _01942_;
  assign _04378_ = _01944_ | _01945_;
  assign _04379_ = _01947_ | _01948_;
  assign _04380_ = _01950_ | _01951_;
  assign _04381_ = _01953_ | _01954_;
  assign _04382_ = _01956_ | _01957_;
  assign _04383_ = _01959_ | _01960_;
  assign _04384_ = _01962_ | _01963_;
  assign _04385_ = _01965_ | _01966_;
  assign _04386_ = _01968_ | _01969_;
  assign _04387_ = _01971_ | _01972_;
  assign _04392_ = _01978_ | _01979_;
  assign _04395_ = _01981_ | _01982_;
  assign _04398_ = _01984_ | _01985_;
  assign _04401_ = _01987_ | _01988_;
  assign _04404_ = _01990_ | _01991_;
  assign _04407_ = _01993_ | _01994_;
  assign _04410_ = _01996_ | _01997_;
  assign _04411_ = _02002_ | _02003_;
  assign _04412_ = _02005_ | _02006_;
  assign _04413_ = _02008_ | _02009_;
  assign _04416_ = _02011_ | _02012_;
  assign _04421_ = _02016_ | _02017_;
  assign _04424_ = _02019_ | _02020_;
  assign _04427_ = _02022_ | _02023_;
  assign _04430_ = _02025_ | _02026_;
  assign _04433_ = _02028_ | _02029_;
  assign _04436_ = _02031_ | _02032_;
  assign _04439_ = _02034_ | _02035_;
  assign _04442_ = _02037_ | _02038_;
  assign _04445_ = _02040_ | _02041_;
  assign _04446_ = _02014_ | _02043_;
  assign _04449_ = _02045_ | _02046_;
  assign _04452_ = _02048_ | _02049_;
  assign _04455_ = _02051_ | _02052_;
  assign _04458_ = _02054_ | _02055_;
  assign _04461_ = _02057_ | _02058_;
  assign _04464_ = _02060_ | _02061_;
  assign _04467_ = _02063_ | _02064_;
  assign _04471_ = _02068_ | _02069_;
  assign _04472_ = _02071_ | _02072_;
  assign _04473_ = _02074_ | _02075_;
  assign _04476_ = _02077_ | _02078_;
  assign _04480_ = _02082_ | _02083_;
  assign _04622_ = _02495_ | _02496_;
  assign _04625_ = _02498_ | _02499_;
  assign _04626_ = _02501_ | _02502_;
  assign _04629_ = _02504_ | _02505_;
  assign _04630_ = _02507_ | _02508_;
  assign _04631_ = _02510_ | _02511_;
  assign _04632_ = _02513_ | _02514_;
  assign _04635_ = _02516_ | _02517_;
  assign _04636_ = _02519_ | _02520_;
  assign _04637_ = _02522_ | _02523_;
  assign _04638_ = _02525_ | _02526_;
  assign _04639_ = _02528_ | _02529_;
  assign _04640_ = _02531_ | _02532_;
  assign _04641_ = _02534_ | _02535_;
  assign _04642_ = _02537_ | _02538_;
  assign _04645_ = _02540_ | _02541_;
  assign _04646_ = _02543_ | _02544_;
  assign _04647_ = _02546_ | _02547_;
  assign _04648_ = _02549_ | _02550_;
  assign _04649_ = _02552_ | _02553_;
  assign _04650_ = _02555_ | _02556_;
  assign _04651_ = _02558_ | _02559_;
  assign _04652_ = _02561_ | _02562_;
  assign _04653_ = _02564_ | _02565_;
  assign _04654_ = _02567_ | _02568_;
  assign _04655_ = _02570_ | _02571_;
  assign _04656_ = _02573_ | _02574_;
  assign _04657_ = _02576_ | _02577_;
  assign _04658_ = _02579_ | _02580_;
  assign _04659_ = _02582_ | _02583_;
  assign _04660_ = _02585_ | _02586_;
  assign _04663_ = _02588_ | _02589_;
  assign _04666_ = _02591_ | _02592_;
  assign _04667_ = _02594_ | _02595_;
  assign _04670_ = _02597_ | _02598_;
  assign _04671_ = _02600_ | _02601_;
  assign _04672_ = _02603_ | _02604_;
  assign _04673_ = _02606_ | _02607_;
  assign _04676_ = _02609_ | _02610_;
  assign _04677_ = _02612_ | _02613_;
  assign _04678_ = _02615_ | _02616_;
  assign _04679_ = _02618_ | _02619_;
  assign _04680_ = _02621_ | _02622_;
  assign _04681_ = _02624_ | _02625_;
  assign _04682_ = _02627_ | _02628_;
  assign _04683_ = _02630_ | _02631_;
  assign _04686_ = _02633_ | _02634_;
  assign _04687_ = _02636_ | _02637_;
  assign _04688_ = _02639_ | _02640_;
  assign _04689_ = _02642_ | _02643_;
  assign _04690_ = _02645_ | _02646_;
  assign _04691_ = _02648_ | _02649_;
  assign _04692_ = _02651_ | _02652_;
  assign _04693_ = _02654_ | _02655_;
  assign _04694_ = _02657_ | _02658_;
  assign _04695_ = _02660_ | _02661_;
  assign _04696_ = _02663_ | _02664_;
  assign _04697_ = _02666_ | _02667_;
  assign _04698_ = _02669_ | _02670_;
  assign _04699_ = _02672_ | _02673_;
  assign _04700_ = _02675_ | _02676_;
  assign _04701_ = _02678_ | _02679_;
  assign _04750_ = _02796_ | _02797_;
  assign _04753_ = _02801_ | _02802_;
  assign _04754_ = _02806_ | _02807_;
  assign _00013_ = _02809_ | _02810_;
  assign _04763_ = _02811_ | _02812_;
  assign _04765_ = _02815_ | _02795_;
  assign _04770_ = _02820_ | _02821_;
  assign _04774_ = _02825_ | _02826_;
  assign _04783_ = _02840_ | _02841_;
  assign _04788_ = _02847_ | _02848_;
  assign _04792_ = _02850_ | _02851_;
  assign _00010_ = _02853_ | _02854_;
  assign _04795_ = _02855_ | _02856_;
  assign _04796_ = _02858_ | _02859_;
  assign _00007_ = _02861_ | _02862_;
  assign _04798_ = _02865_ | _02817_;
  assign _04807_ = _02869_ | _02870_;
  assign _04808_ = _02872_ | _02873_;
  assign _04811_ = _02875_ | _02876_;
  assign _04823_ = _02890_ | _02891_;
  assign _04826_ = _02893_ | _02894_;
  assign _04832_ = _02900_ | _02901_;
  assign _04835_ = _02903_ | _02904_;
  assign _04843_ = _02912_ | _02913_;
  assign _04844_ = _02915_ | _02916_;
  assign _04845_ = _02918_ | _02919_;
  assign _04846_ = _02921_ | _02922_;
  assign _04849_ = _02924_ | _02925_;
  assign _04850_ = _02927_ | _02928_;
  assign _04853_ = _02930_ | _02931_;
  assign _04856_ = _02933_ | _02934_;
  assign _04857_ = _02936_ | _02937_;
  assign _04858_ = _02939_ | _02940_;
  assign _04863_ = _02946_ | _02947_;
  assign _04866_ = _02949_ | _02950_;
  assign _04871_ = _02956_ | _02957_;
  assign _04874_ = _02959_ | _02960_;
  assign _04879_ = _02966_ | _02967_;
  assign _04880_ = _02973_ | _02974_;
  assign _04881_ = _02973_ | _02978_;
  assign _04882_ = _02980_ | _02981_;
  assign _04883_ = _02985_ | _02986_;
  assign _04884_ = _02994_ | _02995_;
  assign _04885_ = _02985_ | _02997_;
  assign _04886_ = _02999_ | _03000_;
  assign _04887_ = _03004_ | _03005_;
  assign _04888_ = _03007_ | _03008_;
  assign _04889_ = _03010_ | _03011_;
  assign _04891_ = _03015_ | _03016_;
  assign _04895_ = _03020_ | _03021_;
  assign _04896_ = _03024_ | _03025_;
  assign _04900_ = _03029_ | _03030_;
  assign _04905_ = _03036_ | _03037_;
  assign _04908_ = _03044_ | _03045_;
  assign _04911_ = _03047_ | _03048_;
  assign _04913_ = _03054_ | _03055_;
  assign _04917_ = _03063_ | _03064_;
  assign _04918_ = _03066_ | _03067_;
  assign _04920_ = _03073_ | _03074_;
  assign _04921_ = _03080_ | _03081_;
  assign _04922_ = _03083_ | _03084_;
  assign _04923_ = _03086_ | _03087_;
  assign _04925_ = _03091_ | _03092_;
  assign _04926_ = _03094_ | _03095_;
  assign _04927_ = _03099_ | _03100_;
  assign _04928_ = _03102_ | _03103_;
  assign _04929_ = _03105_ | _03106_;
  assign _04930_ = _03108_ | _03109_;
  assign _04933_ = _03111_ | _03112_;
  assign _04934_ = _03114_ | _03115_;
  assign _04937_ = _03117_ | _03118_;
  assign _04940_ = _03120_ | _03121_;
  assign _04941_ = _03123_ | _03124_;
  assign _04944_ = _03126_ | _03127_;
  assign _04947_ = _03129_ | _03130_;
  assign _04953_ = _03132_ | _03133_;
  assign _04959_ = _03138_ | _03139_;
  assign _04963_ = _03143_ | _03144_;
  assign _04968_ = _03150_ | _03151_;
  assign _04972_ = _03165_ | _03166_;
  assign _04975_ = _03172_ | _03173_;
  assign _04976_ = _03175_ | _03176_;
  assign _04977_ = _03180_ | _03181_;
  assign _04978_ = _03183_ | _03184_;
  assign _04981_ = _03186_ | _03187_;
  assign _04983_ = _03193_ | _03194_;
  assign _04986_ = _03196_ | _03197_;
  assign _04989_ = _03199_ | _03200_;
  assign _04990_ = _03202_ | _03203_;
  assign _04991_ = _03205_ | _03206_;
  assign _04994_ = _03208_ | _03209_;
  assign _04997_ = _03211_ | _03212_;
  assign _04998_ = _03214_ | _03215_;
  assign _05001_ = _03217_ | _03218_;
  assign _05015_ = _03242_ | _03243_;
  assign _05019_ = _03247_ | _03248_;
  assign _05022_ = _03250_ | _03251_;
  assign _05023_ = _03253_ | _03254_;
  assign _05024_ = _03256_ | _03257_;
  assign _05025_ = _03253_ | _03259_;
  assign _05028_ = _03261_ | _03262_;
  assign _05031_ = _03264_ | _03265_;
  assign _05040_ = _03279_ | _03280_;
  assign _05043_ = _03282_ | _03283_;
  assign _05046_ = _03285_ | _03286_;
  assign _05049_ = _03288_ | _03289_;
  assign _05052_ = _03292_ | _03293_;
  assign _05055_ = _03295_ | _03296_;
  assign _05059_ = _03302_ | _03303_;
  assign _05071_ = _03325_ | _03326_;
  assign _05074_ = _03328_ | _03329_;
  assign _05079_ = _03335_ | _03336_;
  assign _05082_ = _03338_ | _03339_;
  assign _05087_ = _03345_ | _03346_;
  assign _05090_ = _03348_ | _03349_;
  assign _05093_ = _03351_ | _03352_;
  assign _05096_ = _03354_ | _03355_;
  assign _05099_ = _03357_ | _03358_;
  assign _05509_ = decoded_rs1 ^ { _07274_, _07312_ };
  assign _05510_ = _05738_ ^ _07126_;
  assign _05511_ = _06106_ ^ _07122_;
  assign _05512_ = mem_rdata_word ^ { mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15:0] };
  assign _05513_ = _06110_ ^ { mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7:0] };
  assign _05514_ = _07132_ ^ _07130_;
  assign _05515_ = _06122_ ^ _07136_;
  assign _05516_ = _06116_ ^ _00096_;
  assign _05517_ = _06118_ ^ _06114_;
  assign _05518_ = _07134_ ^ _06128_;
  assign _05519_ = count_instr[31:0] ^ count_instr[63:32];
  assign _05520_ = count_cycle[31:0] ^ count_cycle[63:32];
  assign _05521_ = _06126_ ^ _06124_;
  assign _05522_ = _06136_ ^ cpuregs_rs2[4:0];
  assign _05523_ = _06130_ ^ _07140_;
  assign _05524_ = cpuregs_rs2[4:0] ^ decoded_rs2;
  assign _05525_ = decoded_rd ^ _07144_;
  assign _05528_ = _07153_ ^ _07151_;
  assign _05531_ = _06150_ ^ _07159_;
  assign _05532_ = _06152_ ^ _06148_;
  assign _05533_ = _07169_ ^ _07165_;
  assign _05534_ = _06157_ ^ _07163_;
  assign _05535_ = _06184_ ^ _06172_;
  assign _05536_ = cpu_state ^ _07177_;
  assign _05537_ = _06163_ ^ _06161_;
  assign _05538_ = _06165_ ^ _06159_;
  assign _05540_ = _06170_ ^ _06169_;
  assign _05543_ = _06175_ ^ { _05539_[7:4], _07173_[3], _05539_[2:0] };
  assign _05545_ = _06182_ ^ _06178_;
  assign _05546_ = _07192_ ^ _07194_;
  assign _05547_ = _06188_ ^ cpuregs_rs2;
  assign _05548_ = _06201_ ^ _07202_;
  assign _05549_ = _07206_ ^ _06213_;
  assign _05550_ = _06194_ ^ _06192_;
  assign _05551_ = mem_do_prefetch ^ _07204_;
  assign _05552_ = _06199_ ^ _06198_;
  assign _05553_ = _06205_ ^ _07204_;
  assign _05554_ = _06211_ ^ _06207_;
  assign _05557_ = _06218_ ^ _07213_;
  assign _05559_ = _06228_ ^ cpuregs_rs2;
  assign _05560_ = _06226_ ^ decoded_imm;
  assign _05561_ = _07224_ ^ _07220_;
  assign _05562_ = _06246_ ^ _07228_;
  assign _05563_ = _06232_ ^ _06230_;
  assign _05564_ = { pcpi_rs1[30:0], 1'h0 } ^ { 1'h0, pcpi_rs1[31:1] };
  assign _05565_ = _06236_ ^ { 1'hx, pcpi_rs1[31:1] };
  assign _05566_ = { pcpi_rs1[27:0], 4'h0 } ^ { 4'h0, pcpi_rs1[31:4] };
  assign _05567_ = _06240_ ^ { 1'hx, pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31:4] };
  assign _05568_ = _06244_ ^ _07597_;
  assign _05569_ = _00086_ ^ { _00110_[31:1], _07592_[0] };
  assign _05570_ = _07094_ ^ _00108_;
  assign _05571_ = alu_add_sub ^ { 31'h00000000, alu_out_0 };
  assign _05572_ = _06250_ ^ _07609_;
  assign _05573_ = _06252_ ^ _06248_;
  assign _05574_ = _06826_ ^ alu_lts;
  assign _05575_ = _06254_ ^ alu_ltu;
  assign _05576_ = alu_eq ^ _06824_;
  assign _05577_ = _06258_ ^ _06825_;
  assign _05578_ = _06260_ ^ _06256_;
  assign _05580_ = _06262_ ^ _07245_;
  assign _05581_ = _06278_ ^ _06264_;
  assign _05583_ = _06268_ ^ _06266_;
  assign _05584_ = _07260_ ^ _00106_[4];
  assign _05585_ = _06274_ ^ _07263_;
  assign _05586_ = _06276_ ^ _06272_;
  assign _05589_ = _06282_ ^ _07301_;
  assign _05590_ = _06284_ ^ _06280_;
  assign _05591_ = _06300_ ^ _06286_;
  assign _05593_ = _06290_ ^ _06288_;
  assign _05594_ = _07307_ ^ _00106_[3:0];
  assign _05595_ = _06296_ ^ _07310_;
  assign _05596_ = _06298_ ^ _06294_;
  assign _05597_ = _06302_ ^ _00106_[3:0];
  assign _05598_ = _06557_ ^ _07322_;
  assign _05599_ = _06305_ ^ _07318_;
  assign _05600_ = _06319_ ^ _07328_;
  assign _05601_ = _06555_ ^ _07338_;
  assign _05602_ = _06311_ ^ _06309_;
  assign _05603_ = _07336_ ^ _07332_;
  assign _05604_ = _06317_ ^ _06315_;
  assign _05605_ = _06551_ ^ _07358_;
  assign _05606_ = _06321_ ^ _07356_;
  assign _05607_ = { mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31:20] } ^ { mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[7], mem_rdata_q[30:25], mem_rdata_q[11:8], 1'h0 };
  assign _05608_ = _06325_ ^ { mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31:25], mem_rdata_q[11:7] };
  assign _05609_ = _06329_ ^ { mem_rdata_q[31:12], 12'h000 };
  assign _05610_ = _06331_ ^ _06327_;
  assign _05611_ = _07367_ ^ mem_rdata_latched[6:2];
  assign _05613_ = _06337_ ^ _06335_;
  assign _05614_ = _07373_ ^ _06339_;
  assign _05616_ = _06343_ ^ _06341_;
  assign _05617_ = _07386_ ^ _07384_;
  assign _05619_ = _06349_ ^ _06347_;
  assign _05620_ = _06365_ ^ _06351_;
  assign _05622_ = _06355_ ^ _06353_;
  assign _05623_ = _07395_ ^ _07393_;
  assign _05624_ = _06361_ ^ mem_rdata_latched[11:7];
  assign _05625_ = _06363_ ^ _06359_;
  assign _05626_ = _07444_ ^ _07443_;
  assign _05627_ = _07450_ ^ _07447_;
  assign _05628_ = _06369_ ^ _06367_;
  assign _05629_ = _07465_ ^ _07461_;
  assign _05630_ = _06373_ ^ _07460_;
  assign _05631_ = _05831_ ^ _07472_;
  assign _05633_ = _06388_ ^ _06378_;
  assign _05634_ = _05831_ ^ _07481_;
  assign _05635_ = _06382_ ^ _06380_;
  assign _05636_ = _05831_ ^ _07479_;
  assign _05637_ = _06386_ ^ mem_rdata_latched[12];
  assign _05638_ = _05840_ ^ _07486_;
  assign _05639_ = _06390_ ^ _07484_;
  assign _05640_ = _05844_ ^ { mem_rdata_latched[6:4], 2'h0 };
  assign _05641_ = _06394_ ^ _07490_;
  assign _05642_ = _06408_ ^ _06396_;
  assign _05643_ = _05844_ ^ _06412_;
  assign _05644_ = _06400_ ^ _06398_;
  assign _05645_ = _07494_ ^ _07492_;
  assign _05646_ = _05844_ ^ mem_rdata_latched[6:2];
  assign _05647_ = _06406_ ^ _06404_;
  assign _05648_ = _05844_ ^ { mem_rdata_latched[11], mem_rdata_latched[5], mem_rdata_latched[6], 2'h0 };
  assign _05649_ = _06410_ ^ { mem_rdata_latched[11:10], mem_rdata_latched[6], 2'h0 };
  assign _05652_ = _06416_ ^ _06414_;
  assign _05653_ = _06432_ ^ _06418_;
  assign _05654_ = { _05651_[2:1], _05659_[0] } ^ _06436_;
  assign _05655_ = _06422_ ^ _06420_;
  assign _05656_ = { _05651_[2:1], _05659_[0] } ^ _07525_;
  assign _05657_ = _06428_ ^ _07523_;
  assign _05658_ = _06430_ ^ _06426_;
  assign _05661_ = _07531_ ^ _07529_;
  assign _05662_ = _07527_ ^ _07533_;
  assign _05663_ = _06440_ ^ _06438_;
  assign _05664_ = _07539_ ^ { 3'h0, mem_rdata_latched[8:7], mem_rdata_latched[12] };
  assign _05666_ = _06446_ ^ { 3'h0, mem_rdata_latched[3:2], mem_rdata_latched[12] };
  assign _05667_ = _06448_ ^ _06444_;
  assign _05668_ = _06464_ ^ _06450_;
  assign _05669_ = _05665_ ^ _06468_;
  assign _05670_ = _06454_ ^ _06452_;
  assign _05671_ = _07547_ ^ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[6:5], mem_rdata_latched[2] };
  assign _05672_ = _05665_ ^ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] };
  assign _05673_ = _06460_ ^ _07549_;
  assign _05674_ = _06462_ ^ _06458_;
  assign _05675_ = _05665_ ^ { 1'h0, mem_rdata_latched[10:7], mem_rdata_latched[12] };
  assign _05676_ = _06466_ ^ { 4'h0, mem_rdata_latched[5], mem_rdata_latched[12] };
  assign _05677_ = { 24'h000000, mem_rdata[23:16] } ^ { 24'h000000, mem_rdata[31:24] };
  assign _05678_ = { 24'h000000, mem_rdata[7:0] } ^ { 24'h000000, mem_rdata[15:8] };
  assign _05679_ = _06472_ ^ _06470_;
  assign _05680_ = { 16'h0000, mem_rdata[15:0] } ^ { 16'h0000, mem_rdata[31:16] };
  assign _05681_ = mem_rdata ^ _00047_;
  assign _05682_ = _06474_ ^ _00064_;
  assign _05683_ = _06476_ ^ _07581_;
  assign _05684_ = pcpi_rs2 ^ { pcpi_rs2[15:0], pcpi_rs2[15:0] };
  assign _05685_ = _06478_ ^ { pcpi_rs2[7:0], pcpi_rs2[7:0], pcpi_rs2[7:0], pcpi_rs2[7:0] };
  assign _05686_ = pcpi_mul_rd ^ pcpi_div_rd;
  assign _05687_ = _06480_ ^ pcpi_div_wr;
  assign _05688_ = _06901_ ^ _06903_;
  assign _05689_ = _06905_ ^ _06907_;
  assign _05690_ = _06909_ ^ _06911_;
  assign _05691_ = _06913_ ^ _06915_;
  assign _05692_ = _06917_ ^ _06919_;
  assign _05693_ = _06921_ ^ _06923_;
  assign _05694_ = _06925_ ^ _06927_;
  assign _05695_ = _06929_ ^ _06931_;
  assign _05696_ = _06933_ ^ _06935_;
  assign _05697_ = _06937_ ^ _06939_;
  assign _05698_ = _06941_ ^ _06943_;
  assign _05699_ = _06945_ ^ _06947_;
  assign _05700_ = _06949_ ^ _06951_;
  assign _05701_ = _06953_ ^ _06955_;
  assign _05702_ = _06957_ ^ _06959_;
  assign _05703_ = \cpuregs[0]  ^ \cpuregs[1] ;
  assign _05704_ = \cpuregs[20]  ^ \cpuregs[21] ;
  assign _05705_ = \cpuregs[22]  ^ \cpuregs[23] ;
  assign _05706_ = \cpuregs[24]  ^ \cpuregs[25] ;
  assign _05707_ = \cpuregs[26]  ^ \cpuregs[27] ;
  assign _05708_ = \cpuregs[28]  ^ \cpuregs[29] ;
  assign _05709_ = \cpuregs[30]  ^ \cpuregs[31] ;
  assign _05710_ = \cpuregs[2]  ^ \cpuregs[3] ;
  assign _05711_ = \cpuregs[4]  ^ \cpuregs[5] ;
  assign _05712_ = \cpuregs[6]  ^ \cpuregs[7] ;
  assign _05713_ = \cpuregs[8]  ^ \cpuregs[9] ;
  assign _05714_ = \cpuregs[10]  ^ \cpuregs[11] ;
  assign _05715_ = \cpuregs[12]  ^ \cpuregs[13] ;
  assign _05716_ = \cpuregs[14]  ^ \cpuregs[15] ;
  assign _05717_ = \cpuregs[16]  ^ \cpuregs[17] ;
  assign _05718_ = \cpuregs[18]  ^ \cpuregs[19] ;
  assign _05719_ = _06961_ ^ _06963_;
  assign _05720_ = _06965_ ^ _06967_;
  assign _05721_ = _06969_ ^ _06971_;
  assign _05722_ = _06973_ ^ _06975_;
  assign _05723_ = _06977_ ^ _06979_;
  assign _05724_ = _06981_ ^ _06983_;
  assign _05725_ = _06985_ ^ _06987_;
  assign _05726_ = _06989_ ^ _06991_;
  assign _05727_ = _06993_ ^ _06995_;
  assign _05728_ = _06997_ ^ _06999_;
  assign _05729_ = _07001_ ^ _07003_;
  assign _05730_ = _07005_ ^ _07007_;
  assign _05731_ = _07009_ ^ _07011_;
  assign _05732_ = _07013_ ^ _07015_;
  assign _05733_ = _07017_ ^ _07019_;
  assign _05734_ = _07108_ ^ _07599_;
  assign _05735_ = _07112_ ^ latched_rd;
  assign _05736_ = reg_next_pc ^ _07594_;
  assign _05737_ = _05738_ ^ _07120_;
  assign _05739_ = _05738_ ^ _07124_;
  assign _05740_ = _07589_[4:0] ^ _07587_[4:0];
  assign _05741_ = instr_jalr ^ alu_out_0;
  assign _05743_ = latched_store ^ pcpi_int_wr;
  assign _05744_ = cpu_state ^ _07161_;
  assign _05747_ = cpu_state ^ _07175_;
  assign _05751_ = { _07179_[7], _05749_[6:0] } ^ _07183_;
  assign _05752_ = cpuregs_rs2 ^ _07192_;
  assign _05753_ = cpuregs_rs1 ^ _07196_;
  assign _05754_ = _07196_ ^ _07198_;
  assign _05755_ = _06609_ ^ _05742_;
  assign _05757_ = _06238_ ^ _06242_;
  assign _05758_ = _00090_ ^ _00094_;
  assign _05759_ = _00060_ ^ _07230_;
  assign _05762_ = _07241_ ^ mem_rdata_latched[11];
  assign _05763_ = _07243_ ^ mem_rdata_latched[11];
  assign _05764_ = _07256_ ^ _00106_[4];
  assign _05765_ = _07258_ ^ _00106_[4];
  assign _05767_ = mem_rdata_latched[19] ^ _06270_;
  assign _05768_ = mem_rdata_latched[30] ^ mem_rdata_latched[8];
  assign _05769_ = mem_rdata_latched[27] ^ mem_rdata_latched[6];
  assign _05770_ = mem_rdata_latched[26] ^ mem_rdata_latched[7];
  assign _05771_ = mem_rdata_latched[23:21] ^ mem_rdata_latched[5:3];
  assign _05772_ = mem_rdata_latched[25] ^ mem_rdata_latched[2];
  assign _05773_ = mem_rdata_latched[29:28] ^ mem_rdata_latched[10:9];
  assign _05774_ = { mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31] } ^ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] };
  assign _05775_ = mem_rdata_latched[24] ^ mem_rdata_latched[11];
  assign _05776_ = mem_rdata_latched[20] ^ mem_rdata_latched[12];
  assign _05778_ = _07295_ ^ mem_rdata_latched[10:7];
  assign _05779_ = _07297_ ^ mem_rdata_latched[10:7];
  assign _05780_ = _07303_ ^ _00106_[3:0];
  assign _05781_ = _07305_ ^ _00106_[3:0];
  assign _05783_ = mem_rdata_latched[18:15] ^ _06292_;
  assign _05784_ = _06557_ ^ _07316_;
  assign _05785_ = _06557_ ^ _07320_;
  assign _05786_ = _06557_ ^ _06307_;
  assign _05787_ = _06555_ ^ _07326_;
  assign _05788_ = _06555_ ^ _07334_;
  assign _05789_ = _06555_ ^ _07575_;
  assign _05790_ = _06555_ ^ _06313_;
  assign _05791_ = _06549_ ^ _07342_;
  assign _05792_ = _06549_ ^ _07344_;
  assign _05793_ = _06553_ ^ _07348_;
  assign _05794_ = _06553_ ^ _07350_;
  assign _05795_ = _06551_ ^ _07354_;
  assign _05796_ = _06551_ ^ _06323_;
  assign _05797_ = _07365_ ^ mem_rdata_latched[6:2];
  assign _05798_ = _07370_ ^ _00104_[4:0];
  assign _05800_ = mem_rdata_latched[24:20] ^ _06345_;
  assign _05801_ = mem_rdata_latched[19:12] ^ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] };
  assign _05803_ = _07382_ ^ mem_rdata_latched[11:7];
  assign _05804_ = _07389_ ^ _00106_[4:0];
  assign _05805_ = _07391_ ^ _00106_[4:0];
  assign _05806_ = mem_rdata_latched[11:7] ^ _06357_;
  assign _05807_ = _06675_ ^ _07403_;
  assign _05808_ = _06675_ ^ _07405_;
  assign _05809_ = _06675_ ^ _07407_;
  assign _05810_ = _06543_ ^ _07411_;
  assign _05811_ = _06543_ ^ _07415_;
  assign _05812_ = _06539_ ^ _07419_;
  assign _05813_ = _06539_ ^ _07421_;
  assign _05814_ = _06539_ ^ _07423_;
  assign _05815_ = _06539_ ^ _07425_;
  assign _05819_ = q_insn_rs2 ^ _00045_;
  assign _05820_ = q_insn_rs1 ^ _00043_;
  assign _05821_ = { rvfi_insn[31:25], 5'hxx, rvfi_insn[19:15], 3'hx, rvfi_insn[11:0] } ^ _00041_;
  assign _05822_ = { 16'h0000, next_insn_opcode[15:0] } ^ next_insn_opcode;
  assign _05823_ = _07433_ ^ _07435_;
  assign _05825_ = _06371_ ^ _07452_;
  assign _05826_ = mem_wstrb ^ _00112_;
  assign _05828_ = _05827_ ^ _07454_;
  assign _05829_ = _06375_ ^ _07467_;
  assign _05830_ = mem_rdata_q[31] ^ mem_rdata_latched[31];
  assign _05836_ = _07475_ ^ mem_rdata_latched[12];
  assign _05837_ = _07477_ ^ _07607_[6];
  assign _05838_ = _05831_ ^ _06384_;
  assign _05839_ = mem_rdata_q[7] ^ mem_rdata_latched[7];
  assign _05841_ = _05840_ ^ mem_rdata_latched[12];
  assign _05842_ = _05840_ ^ _06392_;
  assign _05843_ = mem_rdata_q[24:20] ^ mem_rdata_latched[24:20];
  assign _05846_ = { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] } ^ { mem_rdata_latched[6], 4'h0 };
  assign _05847_ = _05844_ ^ _06402_;
  assign _05848_ = mem_rdata_q[19:15] ^ mem_rdata_latched[19:15];
  assign _05849_ = { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[6:5] } ^ _07496_;
  assign _05850_ = _07496_ ^ _07498_;
  assign _05851_ = _07496_ ^ _07500_;
  assign _05852_ = _07496_ ^ _07502_;
  assign _05853_ = mem_rdata_q[14:12] ^ mem_rdata_latched[14:12];
  assign _05861_ = _05858_ ^ _07521_;
  assign _05862_ = { _05651_[2:1], _05659_[0] } ^ _06424_;
  assign _05863_ = mem_rdata_q[11:8] ^ mem_rdata_latched[11:8];
  assign _05864_ = _07527_ ^ { mem_rdata_latched[11:9], 1'h0 };
  assign _05865_ = _07527_ ^ { mem_rdata_latched[11:10], mem_rdata_latched[4:3] };
  assign _05866_ = _07527_ ^ { mem_rdata_latched[11:10], mem_rdata_latched[6], 1'h0 };
  assign _05867_ = _07527_ ^ _06442_;
  assign _05868_ = mem_rdata_q[30:25] ^ mem_rdata_latched[30:25];
  assign _05873_ = _07543_ ^ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] };
  assign _05874_ = _07545_ ^ _07607_[5:0];
  assign _05875_ = { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] } ^ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[4:3], mem_rdata_latched[5], mem_rdata_latched[2] };
  assign _05876_ = _05665_ ^ _06456_;
  assign _05877_ = mem_la_firstword ^ mem_la_firstword_reg;
  assign _05878_ = _00053_ ^ { rvfi_rd_wdata, 32'h00000000 };
  assign _05879_ = _00049_ ^ { rvfi_rd_wdata, 32'h00000000 };
  assign _05884_ = reg_next_pc ^ { reg_out[31:1], 1'h0 };
  assign _05885_ = _00084_ ^ _07583_;
  assign _05888_ = reg_next_pc ^ { _00110_[31:1], 1'h0 };
  assign _05889_ = reg_out ^ alu_out_q;
  assign _05890_ = { pcpi_rs1[31:2], 2'h0 } ^ { _00102_, 2'h0 };
  assign _05891_ = mem_rdata_q ^ mem_rdata;
  assign _05892_ = _07604_ ^ { 16'hxxxx, mem_16bit_buffer };
  assign _05893_ = mem_rdata_latched_noshuffle ^ { 16'hxxxx, mem_rdata_latched_noshuffle[31:16] };
  assign _05894_ = _07602_ ^ { mem_rdata_latched_noshuffle[15:0], mem_16bit_buffer };
  assign _01329_ = { _06608_, _06608_, _06608_, _06608_, _06608_ } & _05508_;
  assign _01332_ = { _06608_, _06608_, _06608_, _06608_, _06608_ } & _05509_;
  assign _01573_ = _06492_ & _05510_;
  assign _01576_ = _01098_ & _05511_;
  assign _01579_ = { latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0, latched_is_lh_t0 } & _05512_;
  assign _01582_ = { latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0, latched_is_lb_t0 } & _05513_;
  assign _01585_ = { _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_ } & _05514_;
  assign _01588_ = { _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_ } & _05515_;
  assign _01591_ = { _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_, _06492_ } & _05516_;
  assign _01594_ = { _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_, _05101_ } & _05517_;
  assign _01597_ = { is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0 } & _05518_;
  assign _01600_ = { instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0, instr_rdinstrh_t0 } & _05519_;
  assign _01603_ = { instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0, instr_rdcycleh_t0 } & _05520_;
  assign _01606_ = { _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_, _05103_ } & _05521_;
  assign _01609_ = { _06490_, _06490_, _06490_, _06490_, _06490_ } & _05522_;
  assign _01612_ = { _06494_, _06494_, _06494_, _06494_, _06494_ } & _05523_;
  assign _01615_ = { is_slli_srli_srai_t0, is_slli_srli_srai_t0, is_slli_srli_srai_t0, is_slli_srli_srai_t0, is_slli_srli_srai_t0 } & _05524_;
  assign _01617_ = { _06492_, _06492_, _06492_, _06492_, _06492_ } & _05525_;
  assign _01619_ = _06498_ & _05526_;
  assign _01621_ = _06498_ & _05527_;
  assign _01624_ = _06492_ & _05528_;
  assign _06147_ = _06492_ & _05529_;
  assign _01626_ = _01083_ & _00814_;
  assign _01628_ = _06488_ & _05530_;
  assign _01631_ = _06490_ & _05531_;
  assign _01634_ = _05105_ & _05532_;
  assign _01636_ = is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0 & _00813_;
  assign _01639_ = { _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_ } & _05533_;
  assign _01642_ = { _01098_, _01098_, _01098_, _01098_, _01098_, _01098_, _01098_, _01098_ } & _05534_;
  assign _01645_ = { _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_ } & _05535_;
  assign _01648_ = { _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_ } & _05536_;
  assign _01651_ = { _05107_, _05107_, _05107_, _05107_, _05107_, _05107_, _05107_, _05107_ } & _05537_;
  assign _01654_ = { _00868_, _00868_, _00868_, _00868_, _00868_, _00868_, _00868_, _00868_ } & _05538_;
  assign _01656_ = { instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0 } & { _05539_[7:4], _00827_, _05539_[2:0] };
  assign _01659_ = { _05109_, _05109_, _05109_, _05109_, _05109_, _05109_, _05109_, _05109_ } & _05540_;
  assign _01661_ = { is_sll_srl_sra_t0, is_sll_srl_sra_t0, is_sll_srl_sra_t0, is_sll_srl_sra_t0, is_sll_srl_sra_t0, is_sll_srl_sra_t0, is_sll_srl_sra_t0, is_sll_srl_sra_t0 } & { _05541_[7:3], _00822_, _05541_[1:0] };
  assign _01663_ = { _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_ } & { _05542_[7:4], _00826_, _05542_[2:0] };
  assign _01665_ = { instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0, instr_trap_t0 } & _05543_;
  assign _01667_ = { is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0, is_rdcycle_rdcycleh_rdinstr_rdinstrh_t0 } & { _05544_[7], _00825_, _05544_[5:0] };
  assign _01670_ = { _00870_, _00870_, _00870_, _00870_, _00870_, _00870_, _00870_, _00870_ } & _05545_;
  assign _01673_ = { _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_ } & _05546_;
  assign _01676_ = { _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_ } & _05547_;
  assign _01679_ = _06494_ & _05548_;
  assign _01682_ = _06488_ & _05549_;
  assign _01685_ = _05111_ & _05550_;
  assign _01688_ = instr_trap_t0 & _05551_;
  assign _01690_ = _05109_ & _05552_;
  assign _01692_ = is_sb_sh_sw_t0 & _00474_;
  assign _01694_ = instr_trap_t0 & _05553_;
  assign _01696_ = _06614_ & _00815_;
  assign _01699_ = _05113_ & _05554_;
  assign _01701_ = { instr_lw_t0, instr_lw_t0 } & _05555_;
  assign _01703_ = { _06496_, _06496_ } & _05556_;
  assign _01706_ = { _06498_, _06498_ } & _05557_;
  assign _01708_ = { instr_sw_t0, instr_sw_t0 } & _05558_;
  assign _01710_ = { _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_, _06490_ } & _05559_;
  assign _01713_ = { _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_, _01081_ } & _05560_;
  assign _01716_ = { _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_, _06498_ } & _05561_;
  assign _01719_ = { _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_, _06494_ } & _05562_;
  assign _01722_ = { _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_, _05115_ } & _05563_;
  assign _01725_ = { _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_ } & _05564_;
  assign _01728_ = { _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_ } & _05565_;
  assign _01731_ = { _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_, _06860_ } & _05566_;
  assign _01734_ = { _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_, _06850_ } & _05567_;
  assign _01737_ = { is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0, is_lui_auipc_jal_t0 } & _05568_;
  assign _01740_ = { _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_, _06602_ } & _05569_;
  assign _01743_ = { _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_, _06856_ } & _05570_;
  assign _01746_ = { is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0, is_compare_t0 } & _05571_;
  assign _01749_ = { _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_, _06852_ } & _05572_;
  assign _01752_ = { _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_, _05117_ } & _05573_;
  assign _01755_ = is_slti_blt_slt_t0 & _05574_;
  assign _01758_ = is_sltiu_bltu_sltu_t0 & _05575_;
  assign _01761_ = instr_bne_t0 & _05576_;
  assign _01764_ = instr_bge_t0 & _05577_;
  assign _01767_ = _00872_ & _05578_;
  assign _01769_ = _06303_[1] & _05579_;
  assign _01772_ = _07248_ & _05580_;
  assign _01775_ = _07252_ & _05581_;
  assign _01777_ = _07273_ & _05582_;
  assign _01780_ = _05119_ & _05583_;
  assign _01783_ = _01079_ & _05584_;
  assign _01785_ = _06303_[1] & mem_rdata_latched[11];
  assign _01788_ = _07266_ & _05585_;
  assign _01791_ = _05121_ & _05586_;
  assign _01793_ = { _07255_, _07255_, _07255_, _07255_ } & { _05587_[3:2], _00818_, _05587_[0] };
  assign _01795_ = { _06303_[1], _06303_[1], _06303_[1], _06303_[1] } & _05588_;
  assign _01798_ = { _07271_, _07271_, _07271_, _07271_ } & _05589_;
  assign _01801_ = { _05123_, _05123_, _05123_, _05123_ } & _05590_;
  assign _01804_ = { _07252_, _07252_, _07252_, _07252_ } & _05591_;
  assign _01806_ = { _07273_, _07273_, _07273_, _07273_ } & _05592_;
  assign _01809_ = { _05119_, _05119_, _05119_, _05119_ } & _05593_;
  assign _01812_ = { _01079_, _01079_, _01079_, _01079_ } & _05594_;
  assign _01814_ = { _06303_[1], _06303_[1], _06303_[1], _06303_[1] } & mem_rdata_latched[10:7];
  assign _01817_ = { _07266_, _07266_, _07266_, _07266_ } & _05595_;
  assign _01820_ = { _05121_, _05121_, _05121_, _05121_ } & _05596_;
  assign _01823_ = { _01077_, _01077_, _01077_, _01077_ } & _05597_;
  assign _01826_ = _07268_ & _05598_;
  assign _01829_ = _07252_ & _05599_;
  assign _01832_ = _07252_ & _05600_;
  assign _01835_ = _07273_ & _05601_;
  assign _01838_ = _05119_ & _05602_;
  assign _01841_ = _07248_ & _05603_;
  assign _01843_ = _00866_ & _00802_;
  assign _01846_ = _05125_ & _05604_;
  assign _01849_ = _07273_ & _05605_;
  assign _01852_ = _07252_ & _05606_;
  assign _01855_ = { is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0 } & _05607_;
  assign _01858_ = { is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0, is_sb_sh_sw_t0 } & _05608_;
  assign _01860_ = { instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0 } & { decoded_imm_j[31:1], 1'hx };
  assign _01863_ = { _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_, _07364_ } & _05609_;
  assign _01866_ = { _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_, _00874_ } & _05610_;
  assign _01869_ = { _07255_, _07255_, _07255_, _07255_, _07255_ } & _05611_;
  assign _01871_ = { _06303_[1], _06303_[1], _06303_[1], _06303_[1], _06303_[1] } & _05612_;
  assign _01874_ = { _05123_, _05123_, _05123_, _05123_, _05123_ } & _05613_;
  assign _01877_ = { _07252_, _07252_, _07252_, _07252_, _07252_ } & _05614_;
  assign _01879_ = { _07273_, _07273_, _07273_, _07273_, _07273_ } & _05615_;
  assign _01882_ = { _05119_, _05119_, _05119_, _05119_, _05119_ } & _05616_;
  assign _01885_ = { _07248_, _07248_, _07248_, _07248_, _07248_ } & _05617_;
  assign _01887_ = { _06303_[1], _06303_[1], _06303_[1], _06303_[1], _06303_[1] } & _05618_;
  assign _01890_ = { _05127_, _05127_, _05127_, _05127_, _05127_ } & _05619_;
  assign _01893_ = { _07252_, _07252_, _07252_, _07252_, _07252_ } & _05620_;
  assign _01895_ = { _07273_, _07273_, _07273_, _07273_, _07273_ } & _05621_;
  assign _01898_ = { _05119_, _05119_, _05119_, _05119_, _05119_ } & _05622_;
  assign _01901_ = { _07248_, _07248_, _07248_, _07248_, _07248_ } & _05623_;
  assign _01904_ = { _00866_, _00866_, _00866_, _00866_, _00866_ } & _05624_;
  assign _01907_ = { _05125_, _05125_, _05125_, _05125_, _05125_ } & _05625_;
  assign _06368_ = { _06538_, _06538_ } & _05626_;
  assign _01910_ = { _07440_, _07440_ } & _05627_;
  assign _01913_ = { _05129_, _05129_ } & _05628_;
  assign _01916_ = _07440_ & _05629_;
  assign _01918_ = _06536_ & _05630_;
  assign _01921_ = _07248_ & _05631_;
  assign _01923_ = _00862_ & _05632_;
  assign _01926_ = _07252_ & _05633_;
  assign _01929_ = _07273_ & _05634_;
  assign _01932_ = _05119_ & _05635_;
  assign _01934_ = _07248_ & _05636_;
  assign _01937_ = _01091_ & _05637_;
  assign _01940_ = _07268_ & _05638_;
  assign _01943_ = _00864_ & _05639_;
  assign _01946_ = { _07271_, _07271_, _07271_, _07271_, _07271_ } & _05640_;
  assign _01949_ = { _07248_, _07248_, _07248_, _07248_, _07248_ } & _05641_;
  assign _01952_ = { _07252_, _07252_, _07252_, _07252_, _07252_ } & _05642_;
  assign _01955_ = { _07273_, _07273_, _07273_, _07273_, _07273_ } & _05643_;
  assign _01958_ = { _05119_, _05119_, _05119_, _05119_, _05119_ } & _05644_;
  assign _01961_ = { _07248_, _07248_, _07248_, _07248_, _07248_ } & _05645_;
  assign _01964_ = { _00866_, _00866_, _00866_, _00866_, _00866_ } & _05646_;
  assign _01967_ = { _05125_, _05125_, _05125_, _05125_, _05125_ } & _05647_;
  assign _01970_ = { _06303_[1], _06303_[1], _06303_[1], _06303_[1], _06303_[1] } & _05648_;
  assign _01973_ = { _07271_, _07271_, _07271_, _07271_, _07271_ } & _05649_;
  assign _01975_ = { _01077_, _01077_, _01077_ } & { _05650_[2], _00829_, _05650_[0] };
  assign _01977_ = { _06303_[1], _06303_[1], _06303_[1] } & { _05651_[2:1], _00830_ };
  assign _01980_ = { _05131_, _05131_, _05131_ } & _05652_;
  assign _01983_ = { _07252_, _07252_, _07252_ } & _05653_;
  assign _01986_ = { _07273_, _07273_, _07273_ } & _05654_;
  assign _01989_ = { _05119_, _05119_, _05119_ } & _05655_;
  assign _01992_ = { _07266_, _07266_, _07266_ } & _05656_;
  assign _01995_ = { _07248_, _07248_, _07248_ } & _05657_;
  assign _01998_ = { _05133_, _05133_, _05133_ } & _05658_;
  assign _01999_ = { _06303_[1], _06303_[1], _06303_[1] } & { _05651_[2:1], _05659_[0] };
  assign _02001_ = { _01077_, _01077_, _01077_ } & { _05660_[2], _00837_, _05660_[0] };
  assign _02004_ = { _07252_, _07252_, _07252_, _07252_ } & _05661_;
  assign _02007_ = { _07273_, _07273_, _07273_, _07273_ } & _05662_;
  assign _02010_ = { _05119_, _05119_, _05119_, _05119_ } & _05663_;
  assign _02013_ = { _07255_, _07255_, _07255_, _07255_, _07255_, _07255_ } & _05664_;
  assign _02015_ = { _06303_[1], _06303_[1], _06303_[1], _06303_[1], _06303_[1], _06303_[1] } & _05665_;
  assign _02018_ = { _07271_, _07271_, _07271_, _07271_, _07271_, _07271_ } & _05666_;
  assign _02021_ = { _05123_, _05123_, _05123_, _05123_, _05123_, _05123_ } & _05667_;
  assign _02024_ = { _07252_, _07252_, _07252_, _07252_, _07252_, _07252_ } & _05668_;
  assign _02027_ = { _07273_, _07273_, _07273_, _07273_, _07273_, _07273_ } & _05669_;
  assign _02030_ = { _05119_, _05119_, _05119_, _05119_, _05119_, _05119_ } & _05670_;
  assign _02033_ = { _01079_, _01079_, _01079_, _01079_, _01079_, _01079_ } & _05671_;
  assign _02036_ = { _00866_, _00866_, _00866_, _00866_, _00866_, _00866_ } & _05672_;
  assign _02039_ = { _07266_, _07266_, _07266_, _07266_, _07266_, _07266_ } & _05673_;
  assign _02042_ = { _05121_, _05121_, _05121_, _05121_, _05121_, _05121_ } & _05674_;
  assign _02044_ = { _06303_[1], _06303_[1], _06303_[1], _06303_[1], _06303_[1], _06303_[1] } & _05675_;
  assign _02047_ = { _01077_, _01077_, _01077_, _01077_, _01077_, _01077_ } & _05676_;
  assign _02050_ = { _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_, _07552_ } & _05677_;
  assign _02053_ = { _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_, _07556_ } & _05678_;
  assign _02056_ = { _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_, _05135_ } & _05679_;
  assign _02059_ = { pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1], pcpi_rs1_t0[1] } & _05680_;
  assign _02062_ = { _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_ } & _05681_;
  assign _02065_ = { _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_ } & _05682_;
  assign _02067_ = { _06504_, _06504_, _06504_, _06504_ } & _00816_;
  assign _02070_ = { _07558_, _07558_, _07558_, _07558_ } & _05683_;
  assign _02073_ = { _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_, _06504_ } & _05684_;
  assign _02076_ = { _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_, _07558_ } & _05685_;
  assign _02079_ = { pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0, pcpi_div_ready_t0 } & _05686_;
  assign _02081_ = pcpi_mul_ready_t0 & pcpi_mul_wr;
  assign _02084_ = pcpi_div_ready_t0 & _05687_;
  assign _02497_ = { _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4], _00081_[4] } & _05688_;
  assign _02500_ = { _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3] } & _05689_;
  assign _02503_ = { _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3], _00081_[3] } & _05690_;
  assign _02506_ = { _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2] } & _05691_;
  assign _02509_ = { _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2] } & _05692_;
  assign _02512_ = { _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2] } & _05693_;
  assign _02515_ = { _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2], _00081_[2] } & _05694_;
  assign _02518_ = { _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1] } & _05695_;
  assign _02521_ = { _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1] } & _05696_;
  assign _02524_ = { _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1] } & _05697_;
  assign _02527_ = { _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1] } & _05698_;
  assign _02530_ = { _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1] } & _05699_;
  assign _02533_ = { _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1] } & _05700_;
  assign _02536_ = { _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1] } & _05701_;
  assign _02539_ = { _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1], _00081_[1] } & _05702_;
  assign _02542_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } & _05703_;
  assign _02545_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } & _05704_;
  assign _02548_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } & _05705_;
  assign _02551_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } & _05706_;
  assign _02554_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } & _05707_;
  assign _02557_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } & _05708_;
  assign _02560_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } & _05709_;
  assign _02563_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } & _05710_;
  assign _02566_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } & _05711_;
  assign _02569_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } & _05712_;
  assign _02572_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } & _05713_;
  assign _02575_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } & _05714_;
  assign _02578_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } & _05715_;
  assign _02581_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } & _05716_;
  assign _02584_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } & _05717_;
  assign _02587_ = { _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0], _00081_[0] } & _05718_;
  assign _02590_ = { _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4], _00083_[4] } & _05719_;
  assign _02593_ = { _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3] } & _05720_;
  assign _02596_ = { _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3], _00083_[3] } & _05721_;
  assign _02599_ = { _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2] } & _05722_;
  assign _02602_ = { _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2] } & _05723_;
  assign _02605_ = { _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2] } & _05724_;
  assign _02608_ = { _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2], _00083_[2] } & _05725_;
  assign _02611_ = { _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1] } & _05726_;
  assign _02614_ = { _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1] } & _05727_;
  assign _02617_ = { _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1] } & _05728_;
  assign _02620_ = { _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1] } & _05729_;
  assign _02623_ = { _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1] } & _05730_;
  assign _02626_ = { _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1] } & _05731_;
  assign _02629_ = { _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1] } & _05732_;
  assign _02632_ = { _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1], _00083_[1] } & _05733_;
  assign _02635_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } & _05703_;
  assign _02638_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } & _05704_;
  assign _02641_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } & _05705_;
  assign _02644_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } & _05706_;
  assign _02647_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } & _05707_;
  assign _02650_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } & _05708_;
  assign _02653_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } & _05709_;
  assign _02656_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } & _05710_;
  assign _02659_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } & _05711_;
  assign _02662_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } & _05712_;
  assign _02665_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } & _05713_;
  assign _02668_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } & _05714_;
  assign _02671_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } & _05715_;
  assign _02674_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } & _05716_;
  assign _02677_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } & _05717_;
  assign _02680_ = { _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0], _00083_[0] } & _05718_;
  assign _02784_ = { _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_ } & _00070_;
  assign _02786_ = { _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_ } & _00072_;
  assign _02788_ = { _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_ } & _00066_;
  assign _02790_ = { _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_, _06632_ } & _00068_;
  assign _02792_ = { cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0 } & _05734_;
  assign _02794_ = { cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0, cpuregs_write_t0 } & _05735_;
  assign _02798_ = { latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0, latched_branch_t0 } & _05736_;
  assign _02800_ = _06616_ & _00131_;
  assign _02803_ = _06866_ & _05737_;
  assign _02805_ = alu_out_0_t0 & _05738_;
  assign _02808_ = is_beq_bne_blt_bge_bltu_bgeu_t0 & _05739_;
  assign _02813_ = { _06598_, _06598_, _06598_, _06598_, _06598_ } & _05740_;
  assign _02816_ = is_beq_bne_blt_bge_bltu_bgeu_t0 & _05741_;
  assign _02818_ = decoder_trigger_t0 & _05742_;
  assign _02819_ = is_beq_bne_blt_bge_bltu_bgeu_t0 & _00667_;
  assign _02822_ = pcpi_int_ready_t0 & _05743_;
  assign _02824_ = { _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_, _06616_ } & { cpu_state[7], _00820_, cpu_state[5:0] };
  assign _02827_ = { _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_, _06866_ } & _05744_;
  assign _02829_ = { _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_, _06500_ } & { cpu_state[7], _00820_, cpu_state[5:0] };
  assign _02831_ = { mem_done_t0, mem_done_t0, mem_done_t0, mem_done_t0, mem_done_t0, mem_done_t0, mem_done_t0, mem_done_t0 } & { cpu_state[7], _00820_, cpu_state[5:0] };
  assign _02833_ = { is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0, is_beq_bne_blt_bge_bltu_bgeu_t0 } & { _05745_[7], _00821_, _05745_[5:0] };
  assign _02835_ = { _06612_, _06612_, _06612_, _06612_, _06612_, _06612_, _06612_, _06612_ } & { _00823_, cpu_state[6:0] };
  assign _02837_ = { pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0, pcpi_int_ready_t0 } & { _05746_[7], _00824_, _05746_[5:0] };
  assign _02839_ = { instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0 } & { cpu_state[7:6], _00828_, cpu_state[4:0] };
  assign _02842_ = { decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0 } & _05747_;
  assign _02844_ = { _06620_, _06620_, _06620_, _06620_, _06620_, _06620_, _06620_, _06620_ } & { _00841_, _05749_[6:0] };
  assign _02846_ = { _06622_, _06622_, _06622_, _06622_, _06622_, _06622_, _06622_, _06622_ } & { _00842_, _05750_[6:0] };
  assign _02849_ = { _06618_, _06618_, _06618_, _06618_, _06618_, _06618_, _06618_, _06618_ } & _05751_;
  assign _02852_ = { _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_, _00856_ } & _05752_;
  assign _02857_ = { _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_, _00860_ } & _05753_;
  assign _02860_ = { _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_, _06488_ } & _05754_;
  assign _02864_ = pcpi_int_ready_t0 & _00476_;
  assign _02866_ = decoder_trigger_t0 & _05755_;
  assign _02868_ = _06873_ & _05756_;
  assign _02871_ = { _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_, _06598_ } & _05757_;
  assign _02874_ = { instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0, instr_jal_t0 } & _05758_;
  assign _02877_ = { decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0, decoder_trigger_t0 } & _05759_;
  assign _02879_ = pcpi_int_ready_t0 & _05760_;
  assign _02881_ = _06486_ & _00039_;
  assign _02883_ = _06864_ & _00799_;
  assign _02885_ = prefetched_high_word_t0 & clear_prefetched_high_word_q;
  assign _02887_ = _06684_ & mem_rdata_latched[11];
  assign _02889_ = _06668_ & _05761_;
  assign _02892_ = _06672_ & _05762_;
  assign _02895_ = _06674_ & _05763_;
  assign _02897_ = mem_rdata_latched_t0[12] & mem_rdata_latched[11];
  assign _02899_ = _06680_ & _00106_[4];
  assign _02902_ = _06522_ & _05764_;
  assign _02905_ = _06524_ & _05765_;
  assign _02907_ = _06516_ & mem_rdata_latched[11];
  assign _02909_ = _06896_ & _05766_;
  assign _02911_ = _01077_ & _00106_[4];
  assign _02914_ = _06678_ & _05767_;
  assign _02917_ = _06678_ & _05768_;
  assign _02920_ = _06678_ & _05769_;
  assign _02923_ = _06678_ & _05770_;
  assign _02926_ = { _06678_, _06678_, _06678_ } & _05771_;
  assign _02929_ = _06678_ & _05772_;
  assign _02932_ = { _06678_, _06678_ } & _05773_;
  assign _02935_ = { _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_ } & _05774_;
  assign _02938_ = _06678_ & _05775_;
  assign _02941_ = _06678_ & _05776_;
  assign _02943_ = { _06684_, _06684_, _06684_, _06684_ } & mem_rdata_latched[10:7];
  assign _02945_ = { _06668_, _06668_, _06668_, _06668_ } & _05777_;
  assign _02948_ = { _06672_, _06672_, _06672_, _06672_ } & _05778_;
  assign _02951_ = { _06674_, _06674_, _06674_, _06674_ } & _05779_;
  assign _02953_ = { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] } & mem_rdata_latched[10:7];
  assign _02955_ = { _06680_, _06680_, _06680_, _06680_ } & _00106_[3:0];
  assign _02958_ = { _06522_, _06522_, _06522_, _06522_ } & _05780_;
  assign _02961_ = { _06524_, _06524_, _06524_, _06524_ } & _05781_;
  assign _02963_ = { _06516_, _06516_, _06516_, _06516_ } & mem_rdata_latched[10:7];
  assign _02965_ = { _06896_, _06896_, _06896_, _06896_ } & _05782_;
  assign _02968_ = { _06678_, _06678_, _06678_, _06678_ } & _05783_;
  assign _02970_ = _06668_ & _00800_;
  assign _02972_ = _06674_ & _00801_;
  assign _02975_ = _07248_ & _05784_;
  assign _02977_ = _06524_ & _00800_;
  assign _02979_ = _07248_ & _05785_;
  assign _02982_ = _06678_ & _05786_;
  assign _02984_ = mem_rdata_latched_t0[12] & _00802_;
  assign _02987_ = _06303_[1] & _05787_;
  assign _02989_ = _06680_ & _00802_;
  assign _02991_ = _06522_ & _00803_;
  assign _02993_ = _06516_ & _00802_;
  assign _02996_ = _06896_ & _05788_;
  assign _02998_ = _06303_[1] & _05789_;
  assign _03001_ = _06678_ & _05790_;
  assign _03003_ = _01079_ & _00807_;
  assign _03006_ = _07268_ & _05791_;
  assign _03009_ = _06678_ & _05792_;
  assign _03012_ = _00864_ & _05793_;
  assign _03014_ = _07255_ & _00806_;
  assign _03017_ = _06678_ & _05794_;
  assign _03019_ = _07091_ & _00804_;
  assign _03022_ = _07271_ & _05795_;
  assign _03023_ = _07271_ & _00804_;
  assign _03026_ = _06678_ & _05796_;
  assign _03028_ = { _06668_, _06668_, _06668_, _06668_, _06668_ } & mem_rdata_latched[6:2];
  assign _03031_ = { _06674_, _06674_, _06674_, _06674_, _06674_ } & _05797_;
  assign _03033_ = { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] } & mem_rdata_latched[6:2];
  assign _03035_ = { _06680_, _06680_, _06680_, _06680_, _06680_ } & mem_rdata_latched[6:2];
  assign _03038_ = { _06524_, _06524_, _06524_, _06524_, _06524_ } & _05798_;
  assign _03040_ = { _07248_, _07248_, _07248_, _07248_, _07248_ } & _05799_;
  assign _03042_ = { _07255_, _07255_, _07255_, _07255_, _07255_ } & _00104_[4:0];
  assign _03046_ = { _06678_, _06678_, _06678_, _06678_, _06678_ } & _05800_;
  assign _03049_ = { _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_, _06678_ } & _05801_;
  assign _03051_ = { _06668_, _06668_, _06668_, _06668_, _06668_ } & mem_rdata_latched[11:7];
  assign _03053_ = { _06672_, _06672_, _06672_, _06672_, _06672_ } & { _05802_[4:1], _00819_ };
  assign _03056_ = { _06674_, _06674_, _06674_, _06674_, _06674_ } & _05803_;
  assign _03058_ = { _07091_, _07091_, _07091_, _07091_, _07091_ } & mem_rdata_latched[11:7];
  assign _03060_ = { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] } & mem_rdata_latched[11:7];
  assign _03062_ = { _06680_, _06680_, _06680_, _06680_, _06680_ } & _00106_[4:0];
  assign _03065_ = { _06522_, _06522_, _06522_, _06522_, _06522_ } & _05804_;
  assign _03068_ = { _06524_, _06524_, _06524_, _06524_, _06524_ } & _05805_;
  assign _03070_ = { _06896_, _06896_, _06896_, _06896_, _06896_ } & mem_rdata_latched[11:7];
  assign _03072_ = { _00866_, _00866_, _00866_, _00866_, _00866_ } & _00104_[4:0];
  assign _03075_ = { _06678_, _06678_, _06678_, _06678_, _06678_ } & _05806_;
  assign _03077_ = _06684_ & _00809_;
  assign _03079_ = _06672_ & _00810_;
  assign _03082_ = _07248_ & _05807_;
  assign _03085_ = _07252_ & _05808_;
  assign _03088_ = _06678_ & _05809_;
  assign _03090_ = _01089_ & _00811_;
  assign _03093_ = _07268_ & _05810_;
  assign _03096_ = _06678_ & _05811_;
  assign _03098_ = _06516_ & _00812_;
  assign _03101_ = _06896_ & _05812_;
  assign _03104_ = _07266_ & _05813_;
  assign _03107_ = _07268_ & _05814_;
  assign _03110_ = _06678_ & _05815_;
  assign _03113_ = { decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0 } & _05816_;
  assign _03116_ = { decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0 } & _05817_;
  assign _03119_ = { decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0, decoder_pseudo_trigger_q_t0 } & _05818_;
  assign _03122_ = { dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0 } & _05819_;
  assign _03125_ = { dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0 } & _05820_;
  assign _03128_ = { dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0, dbg_next_t0 } & _05821_;
  assign _03131_ = { _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_, _07430_ } & _05822_;
  assign _03134_ = { mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0, mem_la_read_t0 } & _05823_;
  assign _07451_ = { mem_do_wdata_t0, mem_do_wdata_t0 } & { _00817_, _05824_[0] };
  assign _03137_ = { _00797_, _00797_ } & _05825_;
  assign _03140_ = { _06892_, _06892_, _06892_, _06892_ } & _05826_;
  assign _03142_ = { _06885_, _06885_, _06885_, _06885_ } & _05827_;
  assign _03145_ = { _06837_, _06837_, _06837_, _06837_ } & _05828_;
  assign _03147_ = mem_do_wdata_t0 & _00808_;
  assign _03149_ = _00797_ & _05829_;
  assign _03152_ = mem_xfer_t0 & _05830_;
  assign _03154_ = _06666_ & _05831_;
  assign _03156_ = _06668_ & _05832_;
  assign _03158_ = _06672_ & _05833_;
  assign _03160_ = _06674_ & _05834_;
  assign _03162_ = _06518_ & _05831_;
  assign _03164_ = _06520_ & _05835_;
  assign _03167_ = _06522_ & _05836_;
  assign _03169_ = _06524_ & _05837_;
  assign _03171_ = _00862_ & _05831_;
  assign _03174_ = _06664_ & _05838_;
  assign _03177_ = mem_xfer_t0 & _05839_;
  assign _03179_ = _07255_ & _05840_;
  assign _03182_ = _01079_ & _05841_;
  assign _03185_ = _06664_ & _05842_;
  assign _03188_ = { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 } & _05843_;
  assign _03190_ = { _06666_, _06666_, _06666_, _06666_, _06666_ } & _05844_;
  assign _03192_ = { _06672_, _06672_, _06672_, _06672_, _06672_ } & _05845_;
  assign _03195_ = { _06522_, _06522_, _06522_, _06522_, _06522_ } & _05646_;
  assign _03198_ = { _06516_, _06516_, _06516_, _06516_, _06516_ } & _05846_;
  assign _03201_ = { _06664_, _06664_, _06664_, _06664_, _06664_ } & _05847_;
  assign _03204_ = { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 } & _05848_;
  assign _03207_ = { _06516_, _06516_, _06516_, _06516_, _06516_ } & _05849_;
  assign _03210_ = { _07266_, _07266_, _07266_, _07266_, _07266_ } & _05850_;
  assign _03213_ = { _07268_, _07268_, _07268_, _07268_, _07268_ } & _05851_;
  assign _03216_ = { _06664_, _06664_, _06664_, _06664_, _06664_ } & _05852_;
  assign _03219_ = { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 } & _05853_;
  assign _03221_ = { _06666_, _06666_, _06666_ } & { _05651_[2:1], _05659_[0] };
  assign _03223_ = { _06668_, _06668_, _06668_ } & _05854_;
  assign _03225_ = { _06672_, _06672_, _06672_ } & _05855_;
  assign _03227_ = { _06674_, _06674_, _06674_ } & _05856_;
  assign _03229_ = { _06518_, _06518_, _06518_ } & { _00831_[1], _05651_[1], _00831_[0] };
  assign _03231_ = { _06520_, _06520_, _06520_ } & { _00832_[1], _05857_[1], _00832_[0] };
  assign _03233_ = { _06522_, _06522_, _06522_ } & _00833_;
  assign _03235_ = { _06526_, _06526_, _06526_ } & _05858_;
  assign _03237_ = { _06528_, _06528_, _06528_ } & { _00834_, _05859_[1:0] };
  assign _03239_ = { _06530_, _06530_, _06530_ } & { _00835_, _05860_[0] };
  assign _03241_ = { _06532_, _06532_, _06532_ } & _00836_;
  assign _03244_ = { _06524_, _06524_, _06524_ } & _05861_;
  assign _03246_ = { _06516_, _06516_, _06516_ } & mem_rdata_latched[4:2];
  assign _03249_ = { _06664_, _06664_, _06664_ } & _05862_;
  assign _03252_ = { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 } & _05863_;
  assign _03255_ = { _07255_, _07255_, _07255_, _07255_ } & _05864_;
  assign _03258_ = { _01079_, _01079_, _01079_, _01079_ } & _05865_;
  assign _03260_ = { _07255_, _07255_, _07255_, _07255_ } & _05866_;
  assign _03263_ = { _06664_, _06664_, _06664_, _06664_ } & _05867_;
  assign _03266_ = { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 } & _05868_;
  assign _03268_ = { _06666_, _06666_, _06666_, _06666_, _06666_, _06666_ } & _05665_;
  assign _03270_ = { _06668_, _06668_, _06668_, _06668_, _06668_, _06668_ } & _05869_;
  assign _03272_ = { _06672_, _06672_, _06672_, _06672_, _06672_, _06672_ } & _05870_;
  assign _03274_ = { _06674_, _06674_, _06674_, _06674_, _06674_, _06674_ } & _05871_;
  assign _03276_ = { _06518_, _06518_, _06518_, _06518_, _06518_, _06518_ } & _05665_;
  assign _03278_ = { _06520_, _06520_, _06520_, _06520_, _06520_, _06520_ } & { _00838_, _05872_[4:0] };
  assign _03281_ = { _06522_, _06522_, _06522_, _06522_, _06522_, _06522_ } & _05873_;
  assign _03284_ = { _06524_, _06524_, _06524_, _06524_, _06524_, _06524_ } & _05874_;
  assign _03287_ = { _06516_, _06516_, _06516_, _06516_, _06516_, _06516_ } & _05875_;
  assign _03290_ = { _06664_, _06664_, _06664_, _06664_, _06664_, _06664_ } & _05876_;
  assign _03294_ = last_mem_valid_t0 & _05877_;
  assign _03297_ = { _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_ } & _05878_;
  assign _03299_ = { _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_, _06514_ } & { _00839_, _00055_[31:0] };
  assign _03301_ = { _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31] } & { 32'h00000000, rvfi_rd_wdata };
  assign _03304_ = { _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_ } & _05879_;
  assign _03306_ = { _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_, _06511_ } & { _00840_, _00051_[31:0] };
  assign _03308_ = { _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31] } & { 32'h00000000, rvfi_rd_wdata };
  assign _03327_ = { _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_, _06600_ } & _05884_;
  assign _03330_ = { instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0, instr_sub_t0 } & _05885_;
  assign _03332_ = { _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_, _07565_ } & _05886_;
  assign _03334_ = { _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_, _07567_ } & _05887_;
  assign _03337_ = { latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0, latched_store_t0 } & _05888_;
  assign _03340_ = { latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0, latched_stalu_t0 } & _05889_;
  assign _03342_ = { instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0, instr_lui_t0 } & reg_pc;
  assign _03344_ = { _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_, _07569_ } & cpuregs_wrdata;
  assign _03347_ = { _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_, _06634_ } & _05890_;
  assign _03350_ = { mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0, mem_xfer_t0 } & _05891_;
  assign _03353_ = { mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0, mem_la_use_prefetched_high_word_t0 } & _05892_;
  assign _03356_ = { mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0, mem_la_firstword_t0 } & _05893_;
  assign _03359_ = { mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0, mem_la_secondword_t0 } & _05894_;
  assign _06103_ = _01329_ | _03983_;
  assign _06105_ = _01332_ | _03984_;
  assign _06107_ = _01573_ | _04075_;
  assign _06109_ = _01576_ | _04078_;
  assign _06111_ = _01579_ | _04081_;
  assign _06113_ = _01582_ | _04084_;
  assign _06115_ = _01585_ | _04087_;
  assign _06117_ = _01588_ | _04090_;
  assign _06119_ = _01591_ | _04093_;
  assign _06121_ = _01594_ | _04096_;
  assign _06123_ = _01597_ | _04099_;
  assign _06125_ = _01600_ | _04102_;
  assign _06127_ = _01603_ | _04105_;
  assign _06129_ = _01606_ | _04108_;
  assign _06131_ = _01609_ | _04111_;
  assign _06133_ = _01612_ | _04114_;
  assign _06135_ = _01615_ | _04117_;
  assign _06139_ = _01617_ | _01616_;
  assign _06141_ = _01619_ | _01618_;
  assign _06143_ = _01621_ | _01620_;
  assign _06145_ = _01624_ | _04120_;
  assign _06149_ = _01626_ | _01625_;
  assign _06151_ = _01628_ | _01627_;
  assign _06153_ = _01631_ | _04126_;
  assign _06155_ = _01634_ | _04129_;
  assign _06156_ = _01636_ | _01635_;
  assign _06158_ = _01639_ | _04133_;
  assign _06160_ = _01642_ | _04136_;
  assign _06162_ = _01645_ | _04139_;
  assign _06164_ = _01648_ | _04142_;
  assign _06166_ = _01651_ | _04145_;
  assign _06168_ = _01654_ | _04148_;
  assign _06171_ = _01656_ | _01655_;
  assign _06173_ = _01659_ | _04154_;
  assign _06176_ = _01661_ | _01660_;
  assign _06179_ = _01663_ | _01662_;
  assign _06181_ = _01665_ | _04156_;
  assign _06183_ = _01667_ | _01666_;
  assign _06185_ = _01670_ | _04160_;
  assign _06189_ = _01673_ | _04163_;
  assign _06191_ = _01676_ | _04164_;
  assign _06193_ = _01679_ | _04167_;
  assign _06195_ = _01682_ | _04168_;
  assign _06197_ = _01685_ | _04171_;
  assign _06200_ = _01688_ | _04175_;
  assign _06202_ = _01690_ | _01689_;
  assign _06204_ = _01692_ | _01691_;
  assign _06210_ = _01694_ | _04179_;
  assign _06212_ = _01696_ | _01695_;
  assign _06214_ = _01699_ | _04183_;
  assign _06217_ = _01701_ | _01700_;
  assign _06219_ = _01703_ | _01702_;
  assign _06221_ = _01706_ | _04188_;
  assign _06223_ = _01708_ | _01707_;
  assign _06225_ = _01710_ | _04190_;
  assign _06229_ = _01713_ | _04194_;
  assign _06231_ = _01716_ | _04195_;
  assign _06233_ = _01719_ | _04198_;
  assign _06235_ = _01722_ | _04201_;
  assign _06237_ = _01725_ | _04204_;
  assign _06239_ = _01728_ | _04207_;
  assign _06241_ = _01731_ | _04208_;
  assign _06243_ = _01734_ | _04209_;
  assign _06247_ = _01737_ | _04212_;
  assign _00038_ = _01740_ | _04215_;
  assign _06249_ = _01743_ | _04218_;
  assign _06251_ = _01746_ | _04221_;
  assign _06253_ = _01749_ | _04224_;
  assign alu_out_t0 = _01752_ | _04227_;
  assign _06255_ = _01755_ | _04230_;
  assign _06257_ = _01758_ | _04233_;
  assign _06259_ = _01761_ | _04236_;
  assign _06261_ = _01764_ | _04239_;
  assign alu_out_0_t0 = _01767_ | _04242_;
  assign _06263_ = _01769_ | _01768_;
  assign _06265_ = _01772_ | _04247_;
  assign _06267_ = _01775_ | _04250_;
  assign _06269_ = _01777_ | _01776_;
  assign _06271_ = _01780_ | _04255_;
  assign _06273_ = _01783_ | _04258_;
  assign _06275_ = _01785_ | _01784_;
  assign _06277_ = _01788_ | _04261_;
  assign _06279_ = _01791_ | _04264_;
  assign _06281_ = _01793_ | _01792_;
  assign _06283_ = _01795_ | _01794_;
  assign _06285_ = _01798_ | _04270_;
  assign _06287_ = _01801_ | _04273_;
  assign _06289_ = _01804_ | _04276_;
  assign _06291_ = _01806_ | _01805_;
  assign _06293_ = _01809_ | _04281_;
  assign _06295_ = _01812_ | _04284_;
  assign _06297_ = _01814_ | _01813_;
  assign _06299_ = _01817_ | _04287_;
  assign _06301_ = _01820_ | _04290_;
  assign _06304_ = _01823_ | _04293_;
  assign _06306_ = _01826_ | _04296_;
  assign _06308_ = _01829_ | _04297_;
  assign _06310_ = _01832_ | _04298_;
  assign _06312_ = _01835_ | _04299_;
  assign _06314_ = _01838_ | _04300_;
  assign _06316_ = _01841_ | _04301_;
  assign _06318_ = _01843_ | _01842_;
  assign _06320_ = _01846_ | _04305_;
  assign _06322_ = _01849_ | _04306_;
  assign _06324_ = _01852_ | _04307_;
  assign _06326_ = _01855_ | _04310_;
  assign _06328_ = _01858_ | _04313_;
  assign _06330_ = _01860_ | _01859_;
  assign _06332_ = _01863_ | _04318_;
  assign _06334_ = _01866_ | _04321_;
  assign _06336_ = _01869_ | _04324_;
  assign _06338_ = _01871_ | _01870_;
  assign _06340_ = _01874_ | _04329_;
  assign _06342_ = _01877_ | _04332_;
  assign _06344_ = _01879_ | _01878_;
  assign _06346_ = _01882_ | _04337_;
  assign _06348_ = _01885_ | _04340_;
  assign _06350_ = _01887_ | _01886_;
  assign _06352_ = _01890_ | _04343_;
  assign _06354_ = _01893_ | _04344_;
  assign _06356_ = _01895_ | _01894_;
  assign _06358_ = _01898_ | _04345_;
  assign _06360_ = _01901_ | _04346_;
  assign _06364_ = _01904_ | _04349_;
  assign _06366_ = _01907_ | _04352_;
  assign _06370_ = _01910_ | _04355_;
  assign _06372_ = _01913_ | _04358_;
  assign _06374_ = _01916_ | _04361_;
  assign _06376_ = _01918_ | _01917_;
  assign _06377_ = _01921_ | _04363_;
  assign _06379_ = _01923_ | _01922_;
  assign _06381_ = _01926_ | _04365_;
  assign _06383_ = _01929_ | _04366_;
  assign _06385_ = _01932_ | _04367_;
  assign _06387_ = _01934_ | _04368_;
  assign _06389_ = _01937_ | _04371_;
  assign _06391_ = _01940_ | _04372_;
  assign _06393_ = _01943_ | _04375_;
  assign _06395_ = _01946_ | _04378_;
  assign _06397_ = _01949_ | _04379_;
  assign _06399_ = _01952_ | _04380_;
  assign _06401_ = _01955_ | _04381_;
  assign _06403_ = _01958_ | _04382_;
  assign _06405_ = _01961_ | _04383_;
  assign _06407_ = _01964_ | _04384_;
  assign _06409_ = _01967_ | _04385_;
  assign _06411_ = _01970_ | _04386_;
  assign _06413_ = _01973_ | _04387_;
  assign _06415_ = _01975_ | _01974_;
  assign _06417_ = _01977_ | _01976_;
  assign _06419_ = _01980_ | _04392_;
  assign _06421_ = _01983_ | _04395_;
  assign _06423_ = _01986_ | _04398_;
  assign _06425_ = _01989_ | _04401_;
  assign _06429_ = _01992_ | _04404_;
  assign _06431_ = _01995_ | _04407_;
  assign _06433_ = _01998_ | _04410_;
  assign _06435_ = _01999_ | _01976_;
  assign _06437_ = _02001_ | _02000_;
  assign _06439_ = _02004_ | _04411_;
  assign _06441_ = _02007_ | _04412_;
  assign _06443_ = _02010_ | _04413_;
  assign _06445_ = _02013_ | _04416_;
  assign _06447_ = _02015_ | _02014_;
  assign _06449_ = _02018_ | _04421_;
  assign _06451_ = _02021_ | _04424_;
  assign _06453_ = _02024_ | _04427_;
  assign _06455_ = _02027_ | _04430_;
  assign _06457_ = _02030_ | _04433_;
  assign _06459_ = _02033_ | _04436_;
  assign _06461_ = _02036_ | _04439_;
  assign _06463_ = _02039_ | _04442_;
  assign _06465_ = _02042_ | _04445_;
  assign _06467_ = _02044_ | _04446_;
  assign _06469_ = _02047_ | _04449_;
  assign _06471_ = _02050_ | _04452_;
  assign _06473_ = _02053_ | _04455_;
  assign _00065_ = _02056_ | _04458_;
  assign _00048_ = _02059_ | _04461_;
  assign _06475_ = _02062_ | _04464_;
  assign mem_rdata_word_t0 = _02065_ | _04467_;
  assign _06477_ = _02067_ | _02066_;
  assign mem_la_wstrb_t0 = _02070_ | _04471_;
  assign _06479_ = _02073_ | _04472_;
  assign mem_la_wdata_t0 = _02076_ | _04473_;
  assign pcpi_int_rd_t0 = _02079_ | _04476_;
  assign _06481_ = _02081_ | _02080_;
  assign pcpi_int_wr_t0 = _02084_ | _04480_;
  assign _07086_ = _02497_ | _04622_;
  assign _06902_ = _02500_ | _04625_;
  assign _06904_ = _02503_ | _04626_;
  assign _06906_ = _02506_ | _04629_;
  assign _06908_ = _02509_ | _04630_;
  assign _06910_ = _02512_ | _04631_;
  assign _06912_ = _02515_ | _04632_;
  assign _06914_ = _02518_ | _04635_;
  assign _06916_ = _02521_ | _04636_;
  assign _06918_ = _02524_ | _04637_;
  assign _06920_ = _02527_ | _04638_;
  assign _06922_ = _02530_ | _04639_;
  assign _06924_ = _02533_ | _04640_;
  assign _06926_ = _02536_ | _04641_;
  assign _06928_ = _02539_ | _04642_;
  assign _06930_ = _02542_ | _04645_;
  assign _06950_ = _02545_ | _04646_;
  assign _06952_ = _02548_ | _04647_;
  assign _06954_ = _02551_ | _04648_;
  assign _06956_ = _02554_ | _04649_;
  assign _06958_ = _02557_ | _04650_;
  assign _06960_ = _02560_ | _04651_;
  assign _06932_ = _02563_ | _04652_;
  assign _06934_ = _02566_ | _04653_;
  assign _06936_ = _02569_ | _04654_;
  assign _06938_ = _02572_ | _04655_;
  assign _06940_ = _02575_ | _04656_;
  assign _06942_ = _02578_ | _04657_;
  assign _06944_ = _02581_ | _04658_;
  assign _06946_ = _02584_ | _04659_;
  assign _06948_ = _02587_ | _04660_;
  assign _07085_ = _02590_ | _04663_;
  assign _06962_ = _02593_ | _04666_;
  assign _06964_ = _02596_ | _04667_;
  assign _06966_ = _02599_ | _04670_;
  assign _06968_ = _02602_ | _04671_;
  assign _06970_ = _02605_ | _04672_;
  assign _06972_ = _02608_ | _04673_;
  assign _06974_ = _02611_ | _04676_;
  assign _06976_ = _02614_ | _04677_;
  assign _06978_ = _02617_ | _04678_;
  assign _06980_ = _02620_ | _04679_;
  assign _06982_ = _02623_ | _04680_;
  assign _06984_ = _02626_ | _04681_;
  assign _06986_ = _02629_ | _04682_;
  assign _06988_ = _02632_ | _04683_;
  assign _06990_ = _02635_ | _04686_;
  assign _07010_ = _02638_ | _04687_;
  assign _07012_ = _02641_ | _04688_;
  assign _07014_ = _02644_ | _04689_;
  assign _07016_ = _02647_ | _04690_;
  assign _07018_ = _02650_ | _04691_;
  assign _07020_ = _02653_ | _04692_;
  assign _06992_ = _02656_ | _04693_;
  assign _06994_ = _02659_ | _04694_;
  assign _06996_ = _02662_ | _04695_;
  assign _06998_ = _02665_ | _04696_;
  assign _07000_ = _02668_ | _04697_;
  assign _07002_ = _02671_ | _04698_;
  assign _07004_ = _02674_ | _04699_;
  assign _07006_ = _02677_ | _04700_;
  assign _07008_ = _02680_ | _04701_;
  assign rvfi_csr_minstret_rdata_t0 = _02784_ | _02783_;
  assign rvfi_csr_minstret_rmask_t0 = _02786_ | _02785_;
  assign rvfi_csr_mcycle_rdata_t0 = _02788_ | _02787_;
  assign rvfi_csr_mcycle_rmask_t0 = _02790_ | _02789_;
  assign _07110_ = _02792_ | _02791_;
  assign _07114_ = _02794_ | _02793_;
  assign _07116_ = _02798_ | _04750_;
  assign _07121_ = _02800_ | _02799_;
  assign _07123_ = _02803_ | _04753_;
  assign _07125_ = _02805_ | _02804_;
  assign _07127_ = _02808_ | _04754_;
  assign _07139_ = _02813_ | _04763_;
  assign _07152_ = _02816_ | _04765_;
  assign _07154_ = _02818_ | _02817_;
  assign _07156_ = _02819_ | _02795_;
  assign _07158_ = _02822_ | _04770_;
  assign _07162_ = _02824_ | _02823_;
  assign _07164_ = _02827_ | _04774_;
  assign _07166_ = _02829_ | _02828_;
  assign _07168_ = _02831_ | _02830_;
  assign _07170_ = _02833_ | _02832_;
  assign _07172_ = _02835_ | _02834_;
  assign _07174_ = _02837_ | _02836_;
  assign _07176_ = _02839_ | _02838_;
  assign _07178_ = _02842_ | _04783_;
  assign _07182_ = _02844_ | _02843_;
  assign _07184_ = _02846_ | _02845_;
  assign _07186_ = _02849_ | _04788_;
  assign _07195_ = _02852_ | _04792_;
  assign _07199_ = _02857_ | _04795_;
  assign _07201_ = _02860_ | _04796_;
  assign _07205_ = _02864_ | _02863_;
  assign _07207_ = _02866_ | _04798_;
  assign _07210_ = _02868_ | _02867_;
  assign _07227_ = _02871_ | _04807_;
  assign _07231_ = _02874_ | _04808_;
  assign _07233_ = _02877_ | _04811_;
  assign _07235_ = _02879_ | _02878_;
  assign cpuregs_write_t0 = _02881_ | _02880_;
  assign clear_prefetched_high_word_t0 = _02883_ | _02882_;
  assign _00036_ = _02885_ | _02884_;
  assign _07240_ = _02887_ | _02886_;
  assign _07242_ = _02889_ | _02888_;
  assign _07244_ = _02892_ | _04823_;
  assign _07246_ = _02895_ | _04826_;
  assign _07249_ = _02897_ | _02896_;
  assign _07257_ = _02899_ | _02898_;
  assign _07259_ = _02902_ | _04832_;
  assign _07261_ = _02905_ | _04835_;
  assign _07262_ = _02907_ | _02906_;
  assign _07264_ = _02909_ | _02908_;
  assign _07269_ = _02911_ | _02910_;
  assign _07275_ = _02914_ | _04843_;
  assign _07277_ = _02917_ | _04844_;
  assign _07279_ = _02920_ | _04845_;
  assign _07281_ = _02923_ | _04846_;
  assign _07283_ = _02926_ | _04849_;
  assign _07285_ = _02929_ | _04850_;
  assign _07287_ = _02932_ | _04853_;
  assign _07289_ = _02935_ | _04856_;
  assign _07291_ = _02938_ | _04857_;
  assign _07293_ = _02941_ | _04858_;
  assign _07294_ = _02943_ | _02942_;
  assign _07296_ = _02945_ | _02944_;
  assign _07298_ = _02948_ | _04863_;
  assign _07300_ = _02951_ | _04866_;
  assign _07302_ = _02953_ | _02952_;
  assign _07304_ = _02955_ | _02954_;
  assign _07306_ = _02958_ | _04871_;
  assign _07308_ = _02961_ | _04874_;
  assign _07309_ = _02963_ | _02962_;
  assign _07311_ = _02965_ | _02964_;
  assign _07313_ = _02968_ | _04879_;
  assign _07315_ = _02970_ | _02969_;
  assign _07317_ = _02972_ | _02971_;
  assign _07319_ = _02975_ | _04880_;
  assign _07321_ = _02977_ | _02976_;
  assign _07323_ = _02979_ | _04881_;
  assign _07325_ = _02982_ | _04882_;
  assign _07327_ = _02984_ | _02983_;
  assign _07329_ = _02987_ | _04883_;
  assign _07331_ = _02989_ | _02988_;
  assign _07333_ = _02991_ | _02990_;
  assign _07335_ = _02993_ | _02992_;
  assign _07337_ = _02996_ | _04884_;
  assign _07339_ = _02998_ | _04885_;
  assign _07341_ = _03001_ | _04886_;
  assign _07343_ = _03003_ | _03002_;
  assign _07345_ = _03006_ | _04887_;
  assign _07347_ = _03009_ | _04888_;
  assign _07351_ = _03012_ | _04889_;
  assign _07349_ = _03014_ | _03013_;
  assign _07353_ = _03017_ | _04891_;
  assign _07355_ = _03019_ | _03018_;
  assign _07357_ = _03022_ | _04895_;
  assign _07359_ = _03023_ | _03020_;
  assign _07361_ = _03026_ | _04896_;
  assign _07366_ = _03028_ | _03027_;
  assign _07368_ = _03031_ | _04900_;
  assign _07369_ = _03033_ | _03032_;
  assign _07371_ = _03035_ | _03034_;
  assign _07372_ = _03038_ | _04905_;
  assign _07374_ = _03040_ | _03039_;
  assign _07375_ = _03042_ | _03041_;
  assign _07377_ = _03046_ | _04908_;
  assign _07379_ = _03049_ | _04911_;
  assign _07381_ = _03051_ | _03050_;
  assign _07383_ = _03053_ | _03052_;
  assign _07385_ = _03056_ | _04913_;
  assign _07387_ = _03058_ | _03057_;
  assign _07388_ = _03060_ | _03059_;
  assign _07390_ = _03062_ | _03061_;
  assign _07392_ = _03065_ | _04917_;
  assign _07394_ = _03068_ | _04918_;
  assign _07396_ = _03070_ | _03069_;
  assign _07398_ = _03072_ | _03071_;
  assign _07400_ = _03075_ | _04920_;
  assign _07402_ = _03077_ | _03076_;
  assign _07404_ = _03079_ | _03078_;
  assign _07406_ = _03082_ | _04921_;
  assign _07408_ = _03085_ | _04922_;
  assign _07410_ = _03088_ | _04923_;
  assign _07412_ = _03090_ | _03089_;
  assign _07416_ = _03093_ | _04925_;
  assign _07418_ = _03096_ | _04926_;
  assign _07420_ = _03098_ | _03097_;
  assign _07422_ = _03101_ | _04927_;
  assign _07424_ = _03104_ | _04928_;
  assign _07426_ = _03107_ | _04929_;
  assign _07428_ = _03110_ | _04930_;
  assign _00046_ = _03113_ | _04933_;
  assign _00044_ = _03116_ | _04934_;
  assign _00042_ = _03119_ | _04937_;
  assign dbg_insn_rs2_t0 = _03122_ | _04940_;
  assign dbg_insn_rs1_t0 = _03125_ | _04941_;
  assign dbg_insn_opcode_t0 = _03128_ | _04944_;
  assign _00063_ = _03131_ | _04947_;
  assign _07438_ = _03134_ | _04953_;
  assign _00023_ = _03137_ | _03136_;
  assign _07453_ = _03140_ | _04959_;
  assign _07455_ = _03142_ | _03141_;
  assign _07457_ = _03145_ | _04963_;
  assign _07466_ = _03147_ | _03146_;
  assign _00025_ = _03149_ | _03148_;
  assign _07468_ = _03152_ | _04968_;
  assign _07469_ = _03154_ | _03153_;
  assign _07470_ = _03156_ | _03155_;
  assign _07471_ = _03158_ | _03157_;
  assign _07473_ = _03160_ | _03159_;
  assign _07474_ = _03162_ | _03161_;
  assign _07476_ = _03164_ | _03163_;
  assign _07478_ = _03167_ | _04972_;
  assign _07480_ = _03169_ | _03168_;
  assign _07482_ = _03171_ | _03170_;
  assign _00021_[31] = _03174_ | _04975_;
  assign _07483_ = _03177_ | _04976_;
  assign _07485_ = _03179_ | _03178_;
  assign _07487_ = _03182_ | _04977_;
  assign _00021_[7] = _03185_ | _04978_;
  assign _07488_ = _03188_ | _04981_;
  assign _07489_ = _03190_ | _03189_;
  assign _07491_ = _03192_ | _03191_;
  assign _07493_ = _03195_ | _04983_;
  assign _07495_ = _03198_ | _04986_;
  assign _00021_[24:20] = _03201_ | _04989_;
  assign _07497_ = _03204_ | _04990_;
  assign _07499_ = _03207_ | _04991_;
  assign _07501_ = _03210_ | _04994_;
  assign _07503_ = _03213_ | _04997_;
  assign _00021_[19:15] = _03216_ | _04998_;
  assign _07504_ = _03219_ | _05001_;
  assign _07505_ = _03221_ | _03220_;
  assign _07506_ = _03223_ | _03222_;
  assign _07507_ = _03225_ | _03224_;
  assign _07509_ = _03227_ | _03226_;
  assign _07511_ = _03229_ | _03228_;
  assign _07513_ = _03231_ | _03230_;
  assign _07514_ = _03233_ | _03232_;
  assign _07516_ = _03235_ | _03234_;
  assign _07518_ = _03237_ | _03236_;
  assign _07520_ = _03239_ | _03238_;
  assign _07522_ = _03241_ | _03240_;
  assign _07524_ = _03244_ | _05015_;
  assign _07526_ = _03246_ | _03245_;
  assign _00021_[14:12] = _03249_ | _05019_;
  assign _07528_ = _03252_ | _05022_;
  assign _07530_ = _03255_ | _05023_;
  assign _07532_ = _03258_ | _05024_;
  assign _07534_ = _03260_ | _05025_;
  assign _00021_[11:8] = _03263_ | _05028_;
  assign _07535_ = _03266_ | _05031_;
  assign _07536_ = _03268_ | _03267_;
  assign _07537_ = _03270_ | _03269_;
  assign _07538_ = _03272_ | _03271_;
  assign _07540_ = _03274_ | _03273_;
  assign _07542_ = _03276_ | _03275_;
  assign _07544_ = _03278_ | _03277_;
  assign _07546_ = _03281_ | _05040_;
  assign _07548_ = _03284_ | _05043_;
  assign _07550_ = _03287_ | _05046_;
  assign _00021_[30:25] = _03290_ | _05049_;
  assign _07560_ = _03294_ | _05052_;
  assign _00071_ = _03297_ | _05055_;
  assign _00073_ = _03299_ | _03298_;
  assign _00054_ = _03301_ | _03300_;
  assign _00067_ = _03304_ | _05059_;
  assign _00069_ = _03306_ | _03305_;
  assign _00050_ = _03308_ | _03307_;
  assign next_pc_t0 = _03327_ | _05071_;
  assign alu_add_sub_t0 = _03330_ | _05074_;
  assign cpuregs_rs1_t0 = _03332_ | _03331_;
  assign cpuregs_rs2_t0 = _03334_ | _03333_;
  assign _07595_ = _03337_ | _05079_;
  assign { _00111_[31:1], _07593_[0] } = _03340_ | _05082_;
  assign _07598_ = _03342_ | _03341_;
  assign _07600_ = _03344_ | _03343_;
  assign mem_la_addr_t0 = _03347_ | _05087_;
  assign mem_rdata_latched_noshuffle_t0 = _03350_ | _05090_;
  assign mem_rdata_latched_t0 = _03353_ | _05093_;
  assign _07603_ = _03356_ | _05096_;
  assign _07605_ = _03359_ | _05099_;
  assign _00943_ = | { _06893_, mem_la_read, mem_do_rdata };
  assign _00945_ = { mem_la_read, mem_do_rdata } != 2'h1;
  assign _00947_ = { mem_la_read, mem_la_use_prefetched_high_word } != 2'h3;
  assign _00949_ = { _06888_, resetn } != 2'h3;
  assign _00951_ = { _06537_, _06888_, mem_do_rinst } != 3'h4;
  assign _00953_ = { _06836_, _06888_, _06884_, mem_do_wdata } != 4'h8;
  assign _00955_ = { _07439_, _06888_, mem_xfer } != 3'h4;
  assign _00957_ = { _06535_, _06888_, mem_xfer } != 3'h4;
  assign _00959_ = { _07439_, _06888_, mem_la_read, mem_xfer } != 4'hb;
  assign _00961_ = | { _06836_, _06535_, _06537_, _07439_, _06888_ };
  assign _00963_ = | { _06884_, mem_do_wdata };
  assign _00965_ = { _06888_, _06889_ } != 2'h2;
  assign _00967_ = | { _06836_, _06535_, _07439_, _06888_ };
  assign _00969_ = | { _06487_, _06489_ };
  assign _00971_ = | { _06627_, mem_instr };
  assign _00973_ = { _06491_, is_beq_bne_blt_bge_bltu_bgeu } != 2'h2;
  assign _00975_ = | { _06485_, _06491_ };
  assign _00977_ = { _06497_, _06865_, mem_do_rdata } != 3'h7;
  assign _00979_ = { _06497_, _06865_ } != 2'h2;
  assign _00981_ = | { _06485_, _06497_ };
  assign _00983_ = { _06491_, is_beq_bne_blt_bge_bltu_bgeu } != 2'h3;
  assign _00985_ = { _06487_, is_rdcycle_rdcycleh_rdinstr_rdinstrh, instr_trap } != 3'h4;
  assign _00987_ = { _06489_, instr_trap } != 2'h2;
  assign _00989_ = | { _06487_, _06489_, _06485_, _06491_, _01082_ };
  assign _00991_ = | { _06872_, resetn };
  assign _00993_ = { _01080_, _06487_, _01092_, _06872_, _06613_, instr_trap, is_sll_srl_sra, resetn } != 8'h43;
  assign _00995_ = { _06489_, _06872_, is_sll_srl_sra, resetn } != 4'hb;
  assign _00997_ = { _06493_, _06872_, _06499_, resetn } != 4'h9;
  assign _00999_ = { _06487_, _01092_, _06872_, resetn } != 4'hd;
  assign _01001_ = { _06487_, _06489_, _06485_, _06493_, _06872_, resetn } != 6'h01;
  assign _01003_ = { _06495_, _06865_, mem_do_wdata } != 3'h7;
  assign _01005_ = { _06493_, _06849_, _06859_, _06857_, _06597_, _06499_ } != 6'h20;
  assign _01007_ = { _06493_, _06849_, _06597_, _06499_ } != 4'hc;
  assign _01009_ = { _06493_, _06849_, _06859_, _06857_, _06597_, _06499_ } != 6'h22;
  assign _01011_ = { _06493_, _06849_, _06597_, _06499_ } != 4'he;
  assign _01013_ = { _06493_, _06499_ } != 2'h3;
  assign _01015_ = { _06495_, _06865_ } != 2'h2;
  assign _01017_ = | { _06487_, _06493_, _06495_, _06497_ };
  assign _01019_ = { _06497_, _06869_, _06867_, _06865_, instr_lw, mem_do_rdata } != 6'h24;
  assign _01021_ = { _06495_, _06865_, instr_sw, instr_sh, instr_sb, mem_do_wdata } != 6'h30;
  assign _01023_ = | { _06485_, _06495_, _06497_ };
  assign _01025_ = | { cpuregs_write, rvfi_valid };
  assign _01027_ = { _00857_, instr_trap } != 2'h2;
  assign _01029_ = & { _00175_, _07439_, _00945_, _00943_, _00947_, mem_xfer };
  assign _01031_ = & { _00472_, _00467_, _07439_, mem_xfer };
  assign _01033_ = & { _07439_, mem_xfer };
  assign _01035_ = & { _00951_, _00949_, _00959_, _00961_, _00953_, _00955_, _00957_ };
  assign _01037_ = & { _00175_, _00963_, _06836_ };
  assign _01039_ = & { _00175_, _06891_ };
  assign _01041_ = & { _00953_, _00955_, _00957_, _00967_, _00965_ };
  assign _01043_ = & { _00175_, mem_la_write };
  assign _01045_ = & { _00975_, _00973_, resetn };
  assign _01047_ = & { _00981_, _00979_, _00977_ };
  assign _01049_ = & { _06485_, resetn };
  assign _01051_ = & { _00983_, _00975_ };
  assign _01053_ = & { _00989_, _00987_, _00985_ };
  assign _01055_ = & { _01001_, _00999_, _00997_, _00995_, _00993_, _00991_ };
  assign _01057_ = & { _00969_, resetn };
  assign _01059_ = & { _01017_, _01015_, _01013_, _01011_, _01009_, _01007_, _01005_, _01003_, _00979_, _00977_, resetn };
  assign _01061_ = & { _01017_, _01015_, _01013_, _01009_, _01005_, _01003_, _00979_, _00977_, resetn };
  assign _01063_ = & { _01023_, _01021_, _01019_, _01015_, _01003_, _00979_, _00977_, resetn };
  assign _01065_ = & { _00675_, _06485_, decoder_trigger, resetn };
  assign _01067_ = & { _06485_, decoder_trigger };
  assign _01069_ = & { _01027_, _00969_ };
  assign _00798_ = ~ dbg_rs1val_valid;
  assign _01071_ = | { _06888_, clear_prefetched_high_word };
  assign _01072_ = | { _00670_, _06685_ };
  assign _01073_ = | { _00670_, _07111_ };
  assign _01074_ = | { _00798_, _07097_, _07096_ };
  assign _01075_ = & { _06865_, _01097_, resetn };
  assign _00799_ = ~ _00035_;
  assign _00800_ = ~ _06557_;
  assign _00801_ = ~ _07314_;
  assign _00802_ = ~ _06555_;
  assign _00803_ = ~ _07330_;
  assign _00804_ = ~ _06551_;
  assign _00805_ = ~ dbg_valid_insn;
  assign _00806_ = ~ _06553_;
  assign _00807_ = ~ _06549_;
  assign _00808_ = ~ _07463_;
  assign _00809_ = ~ _06675_;
  assign _00810_ = ~ _07401_;
  assign _00811_ = ~ _06543_;
  assign _00812_ = ~ _06539_;
  assign _00813_ = ~ _07157_;
  assign _00814_ = ~ _07155_;
  assign _00815_ = ~ _06209_;
  assign _00816_ = ~ _07606_;
  assign _00817_ = ~ _07449_[1];
  assign _00818_ = ~ _07299_[1];
  assign _00819_ = ~ _07380_[0];
  assign _00821_ = ~ _07167_[6];
  assign _00820_ = ~ cpu_state[6];
  assign _00822_ = ~ _06174_[2];
  assign _00823_ = ~ cpu_state[7];
  assign _00824_ = ~ _07171_[6];
  assign _00825_ = ~ _06180_[6];
  assign _00826_ = ~ _06177_[3];
  assign _00827_ = ~ _07173_[3];
  assign _00828_ = ~ cpu_state[5];
  assign _00829_ = ~ _07508_[1];
  assign _00830_ = ~ _05659_[0];
  assign _00831_ = ~ { _05651_[2], _05659_[0] };
  assign _00832_ = ~ { _07510_[2], _07510_[0] };
  assign _00833_ = ~ _07512_;
  assign _00834_ = ~ _07515_[2];
  assign _00835_ = ~ _07517_[2:1];
  assign _00836_ = ~ _07519_;
  assign _00837_ = ~ _06434_[1];
  assign _00838_ = ~ _07541_[5];
  assign _00839_ = ~ _00055_[63:32];
  assign _00840_ = ~ _00051_[63:32];
  assign _00841_ = ~ _07179_[7];
  assign _00842_ = ~ _07181_[7];
  assign _01080_ = | { is_jalr_addi_slti_sltiu_xori_ori_andi, is_lui_auipc_jal };
  assign _01082_ = | { _06497_, _06493_ };
  assign _01084_ = | { _06613_, is_jalr_addi_slti_sltiu_xori_ori_andi, is_lui_auipc_jal, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle };
  assign _01086_ = | { _06497_, _06495_, _06493_, _06489_, _06487_, _06485_, _06483_ };
  assign _01087_ = | { _06497_, _06493_, _06491_, _06489_, _06487_, _06485_, _06483_ };
  assign _01088_ = | { _07413_, _07397_ };
  assign _01076_ = | { _07270_, _07254_ };
  assign _01078_ = | { _07254_, _07253_ };
  assign _01090_ = | { _07270_, _07265_, _07254_, _07253_, _07250_ };
  assign _01092_ = | { is_slli_srli_srai, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle };
  assign _01094_ = | { _06601_, latched_branch };
  assign _01095_ = | { _06613_, is_slli_srli_srai, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle };
  assign _01097_ = | { _06497_, _06495_ };
  assign _00843_ = ~ instr_rdinstr;
  assign _00844_ = ~ _01092_;
  assign _00845_ = ~ _06495_;
  assign _00846_ = ~ _06853_;
  assign _00847_ = ~ _07553_;
  assign _00848_ = ~ pcpi_rs1;
  assign _00849_ = ~ instr_rdinstrh;
  assign _00850_ = ~ _06855_;
  assign _00851_ = ~ _06537_;
  assign _00852_ = ~ _07253_;
  assign _00853_ = ~ _07551_;
  assign _00854_ = ~ pcpi_rs2;
  assign _01513_ = _06494_ & _00516_;
  assign _01516_ = instr_rdinstr_t0 & _00849_;
  assign _01519_ = _06492_ & _00534_;
  assign _01522_ = _06488_ & _00536_;
  assign _01525_ = _06490_ & _00552_;
  assign _01528_ = is_sb_sh_sw_t0 & _00554_;
  assign _01531_ = _01093_ & _00558_;
  assign _01534_ = _06496_ & _00516_;
  assign _01537_ = _06854_ & _00850_;
  assign _01540_ = _07271_ & _00582_;
  assign _01543_ = _06536_ & _00851_;
  assign _01546_ = _07266_ & _00582_;
  assign _01549_ = _07248_ & _00710_;
  assign _01552_ = _00862_ & _00852_;
  assign _01555_ = _07248_ & _00722_;
  assign _01558_ = _07268_ & _00583_;
  assign _01561_ = _07248_ & _00586_;
  assign _01564_ = _07554_ & _00853_;
  assign _02780_ = pcpi_rs1_t0 & _00854_;
  assign _01514_ = _06498_ & _00552_;
  assign _01517_ = instr_rdinstrh_t0 & _00843_;
  assign _01520_ = _01083_ & _00517_;
  assign _01523_ = _06490_ & _00535_;
  assign _01526_ = _06494_ & _00536_;
  assign _01529_ = is_sll_srl_sra_t0 & _00557_;
  assign _01532_ = _01081_ & _00844_;
  assign _01535_ = _06498_ & _00845_;
  assign _01538_ = _06856_ & _00846_;
  assign _01541_ = _07248_ & _00724_;
  assign _01544_ = _06538_ & _00620_;
  assign _01547_ = _07248_ & _00587_;
  assign _01550_ = _01077_ & _00582_;
  assign _01553_ = _06427_[0] & _00621_;
  assign _01556_ = _07255_ & _00582_;
  assign _01559_ = _07252_ & _00599_;
  assign _01562_ = _01079_ & _00582_;
  assign _01565_ = _07552_ & _00847_;
  assign _02781_ = pcpi_rs2_t0 & _00848_;
  assign _01515_ = _06494_ & _06498_;
  assign _01518_ = instr_rdinstr_t0 & instr_rdinstrh_t0;
  assign _01521_ = _06492_ & _01083_;
  assign _01524_ = _06488_ & _06490_;
  assign _01527_ = _06490_ & _06494_;
  assign _01530_ = is_sb_sh_sw_t0 & is_sll_srl_sra_t0;
  assign _01533_ = _01093_ & _01081_;
  assign _01536_ = _06496_ & _06498_;
  assign _01539_ = _06854_ & _06856_;
  assign _01542_ = _07271_ & _07248_;
  assign _01545_ = _06536_ & _06538_;
  assign _01548_ = _07266_ & _07248_;
  assign _01551_ = _07248_ & _01077_;
  assign _01554_ = _00862_ & _06427_[0];
  assign _01557_ = _07248_ & _07255_;
  assign _01560_ = _07268_ & _07252_;
  assign _01563_ = _07248_ & _01079_;
  assign _01566_ = _07554_ & _07552_;
  assign _04054_ = _01513_ | _01514_;
  assign _04055_ = _01516_ | _01517_;
  assign _04056_ = _01519_ | _01520_;
  assign _04057_ = _01522_ | _01523_;
  assign _04058_ = _01525_ | _01526_;
  assign _04059_ = _01528_ | _01529_;
  assign _04060_ = _01531_ | _01532_;
  assign _04061_ = _01534_ | _01535_;
  assign _04062_ = _01537_ | _01538_;
  assign _04063_ = _01540_ | _01541_;
  assign _04064_ = _01543_ | _01544_;
  assign _04065_ = _01546_ | _01547_;
  assign _04066_ = _01549_ | _01550_;
  assign _04067_ = _01552_ | _01553_;
  assign _04068_ = _01555_ | _01556_;
  assign _04069_ = _01558_ | _01559_;
  assign _04070_ = _01561_ | _01562_;
  assign _04071_ = _01564_ | _01565_;
  assign _04734_ = _02780_ | _02781_;
  assign _05101_ = _04054_ | _01515_;
  assign _05103_ = _04055_ | _01518_;
  assign _05105_ = _04056_ | _01521_;
  assign _05107_ = _04057_ | _01524_;
  assign _05111_ = _04058_ | _01527_;
  assign _05109_ = _04059_ | _01530_;
  assign _05113_ = _04060_ | _01533_;
  assign _05115_ = _04061_ | _01536_;
  assign _05117_ = _04062_ | _01539_;
  assign _05127_ = _04063_ | _01542_;
  assign _05129_ = _04064_ | _01545_;
  assign _05125_ = _04065_ | _01548_;
  assign _05131_ = _04066_ | _01551_;
  assign _05133_ = _04067_ | _01554_;
  assign _05123_ = _04068_ | _01557_;
  assign _05119_ = _04069_ | _01560_;
  assign _05121_ = _04070_ | _01563_;
  assign _05135_ = _04071_ | _01566_;
  assign _07095_ = _04734_ | _02782_;
  assign _00857_ = | { _06489_, _06487_ };
  assign _00855_ = | { _06613_, is_jalr_addi_slti_sltiu_xori_ori_andi, is_slli_srli_srai, is_lui_auipc_jal, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle };
  assign _00859_ = | { is_lui_auipc_jal, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle };
  assign _00863_ = | { _07272_, _07251_ };
  assign _00865_ = | { _07270_, _07250_ };
  assign _00861_ = | { _07270_, _07254_, _07250_ };
  assign pcpi_int_ready = | { pcpi_div_ready, pcpi_mul_ready };
  assign _05100_ = _06493_ | _06497_;
  assign _05102_ = instr_rdinstr | instr_rdinstrh;
  assign _05104_ = _06491_ | _01082_;
  assign _05106_ = _06487_ | _06489_;
  assign _05110_ = _06489_ | _06493_;
  assign _05108_ = is_sb_sh_sw | is_sll_srl_sra;
  assign _05112_ = _01092_ | _01080_;
  assign _05114_ = _06495_ | _06497_;
  assign _05116_ = _06853_ | _06855_;
  assign _05126_ = _07270_ | _07247_;
  assign _05128_ = _06535_ | _06537_;
  assign _05124_ = _07265_ | _07247_;
  assign _05130_ = _07247_ | _01076_;
  assign _05132_ = _00861_ | _07253_;
  assign _05122_ = _07247_ | _07254_;
  assign _05118_ = _07267_ | _07251_;
  assign _05120_ = _07247_ | _01078_;
  assign _05134_ = _07553_ | _07551_;
  assign _00867_ = | { _06497_, _06495_, _06493_, _06491_ };
  assign _00869_ = | { _06613_, is_jalr_addi_slti_sltiu_xori_ori_andi, is_slli_srli_srai, is_lui_auipc_jal };
  assign _00871_ = | { is_sltiu_bltu_sltu, is_slti_blt_slt, instr_bgeu };
  assign _00873_ = | { is_alu_reg_imm, is_beq_bne_blt_bge_bltu_bgeu, is_sb_sh_sw, is_lb_lh_lw_lbu_lhu, instr_jalr };
  assign _00059_ = _01087_ ? 1'h0 : _00076_;
  assign _00057_ = _06497_ ? _00074_ : 1'h0;
  assign _00058_ = _01086_ ? 1'h0 : _00075_;
  assign _06106_ = _06491_ ? _07126_ : _05738_;
  assign _06108_ = _01097_ ? _07122_ : _06106_;
  assign _06110_ = latched_is_lh ? { mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15:0] } : mem_rdata_word;
  assign _06112_ = latched_is_lb ? { mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7:0] } : _06110_;
  assign _06114_ = _06497_ ? _07130_ : _07132_;
  assign _06116_ = _06489_ ? _07136_ : _06122_;
  assign _06118_ = _06491_ ? _00096_ : _06116_;
  assign _06120_ = _05100_ ? _06114_ : _06118_;
  assign _06122_ = is_rdcycle_rdcycleh_rdinstr_rdinstrh ? _06128_ : _07134_;
  assign _06124_ = instr_rdinstrh ? count_instr[63:32] : count_instr[31:0];
  assign _06126_ = instr_rdcycleh ? count_cycle[63:32] : count_cycle[31:0];
  assign _06128_ = _05102_ ? _06124_ : _06126_;
  assign _06130_ = _06489_ ? cpuregs_rs2[4:0] : _06136_;
  assign _06132_ = _06493_ ? _07140_ : _06130_;
  assign _06134_ = is_slli_srli_srai ? decoded_rs2 : cpuregs_rs2[4:0];
  assign _06136_ = _01084_ ? 5'hxx : _06134_;
  assign _06138_ = _06491_ ? _07144_ : decoded_rd;
  assign _06140_ = _06497_ ? _05526_ : 1'h0;
  assign _06142_ = _06497_ ? _05527_ : 1'h0;
  assign _06144_ = _06491_ ? _07151_ : _07153_;
  assign _06146_ = _06491_ ? _05529_ : 1'h0;
  assign _06148_ = _01082_ ? 1'h1 : _07155_;
  assign _06150_ = _06487_ ? _05530_ : 1'h0;
  assign _06152_ = _06489_ ? _07159_ : _06150_;
  assign _06154_ = _05104_ ? _06148_ : _06152_;
  assign _05530_ = is_rdcycle_rdcycleh_rdinstr_rdinstrh ? 1'h1 : _07157_;
  assign _06157_ = _06493_ ? _07165_ : _07169_;
  assign _06159_ = _01097_ ? _07163_ : _06157_;
  assign _06161_ = _06489_ ? _06172_ : _06184_;
  assign _06163_ = _06485_ ? _07177_ : cpu_state;
  assign _06165_ = _05106_ ? _06161_ : _06163_;
  assign { _05748_[7], _06167_[6], _05748_[5:0] } = _00867_ ? _06159_ : _06165_;
  assign _06169_ = is_sll_srl_sra ? 8'h04 : 8'h02;
  assign _06170_ = instr_trap ? { _05539_[7:4], _07173_[3], _05539_[2:0] } : 8'h08;
  assign _06172_ = _05108_ ? _06169_ : _06170_;
  assign { _05541_[7:3], _06174_[2], _05541_[1:0] } = is_sb_sh_sw ? 8'h02 : 8'h08;
  assign _06175_ = is_sll_srl_sra ? 8'h04 : { _05541_[7:3], _06174_[2], _05541_[1:0] };
  assign { _05542_[7:4], _06177_[3], _05542_[2:0] } = is_slli_srli_srai ? 8'h04 : 8'h01;
  assign _06178_ = _01080_ ? 8'h08 : { _05542_[7:4], _06177_[3], _05542_[2:0] };
  assign { _05544_[7], _06180_[6], _05544_[5:0] } = instr_trap ? { _05539_[7:4], _07173_[3], _05539_[2:0] } : _06175_;
  assign _06182_ = is_rdcycle_rdcycleh_rdinstr_rdinstrh ? 8'h40 : { _05544_[7], _06180_[6], _05544_[5:0] };
  assign _06184_ = _00869_ ? _06178_ : _06182_;
  assign _06186_ = _06487_ ? _07188_ : _07187_;
  assign _06187_ = _06489_ ? 1'h1 : _06186_;
  assign _06188_ = _06487_ ? _07194_ : _07192_;
  assign _06190_ = _06489_ ? cpuregs_rs2 : _06188_;
  assign _06192_ = _06493_ ? _07202_ : _06201_;
  assign _06194_ = _06487_ ? _06213_ : _07206_;
  assign _06196_ = _05110_ ? _06192_ : _06194_;
  assign _06198_ = is_sll_srl_sra ? 1'hx : 1'h1;
  assign _06199_ = instr_trap ? _07204_ : mem_do_prefetch;
  assign _06201_ = _05108_ ? _06198_ : _06199_;
  assign _06203_ = is_sb_sh_sw ? 1'h1 : mem_do_prefetch;
  assign _06205_ = is_sll_srl_sra ? 1'hx : _06203_;
  assign _06207_ = _01080_ ? mem_do_prefetch : 1'hx;
  assign _06209_ = instr_trap ? _07204_ : _06205_;
  assign _06211_ = _06613_ ? 1'h1 : _06209_;
  assign _06213_ = _05112_ ? _06207_ : _06211_;
  assign _05555_ = _06869_ ? 2'h1 : 2'h2;
  assign _06216_ = instr_lw ? 2'h0 : _05555_;
  assign _06218_ = _06495_ ? _05556_ : 2'h0;
  assign _06220_ = _06497_ ? _07213_ : _06218_;
  assign _05558_ = instr_sh ? 2'h1 : 2'h2;
  assign _06222_ = instr_sw ? 2'h0 : _05558_;
  assign _06224_ = _06489_ ? cpuregs_rs2 : _06228_;
  assign _06226_ = _01095_ ? 32'hxxxxxxxx : cpuregs_rs2;
  assign _06228_ = _01080_ ? decoded_imm : _06226_;
  assign _06230_ = _06497_ ? _07220_ : _07224_;
  assign _06232_ = _06493_ ? _07228_ : _06246_;
  assign _06234_ = _05114_ ? _06230_ : _06232_;
  assign _06236_ = _06859_ ? { 1'h0, pcpi_rs1[31:1] } : { pcpi_rs1[30:0], 1'h0 };
  assign _06238_ = _06849_ ? { 1'hx, pcpi_rs1[31:1] } : _06236_;
  assign _06240_ = _06859_ ? { 4'h0, pcpi_rs1[31:4] } : { pcpi_rs1[27:0], 4'h0 };
  assign _06242_ = _06849_ ? { 1'hx, pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31:4] } : _06240_;
  assign _06244_ = is_rdcycle_rdcycleh_rdinstr_rdinstrh ? 32'hxxxxxxxx : cpuregs_rs1;
  assign _06246_ = is_lui_auipc_jal ? _07597_ : _06244_;
  assign _00037_ = _06601_ ? { _00110_[31:1], _07592_[0] } : _00086_;
  assign _06248_ = _06855_ ? _00108_ : _07094_;
  assign _06250_ = is_compare ? { 31'h00000000, alu_out_0 } : alu_add_sub;
  assign _06252_ = _06851_ ? _07609_ : _06250_;
  assign alu_out = _05116_ ? _06248_ : _06252_;
  assign _06254_ = is_slti_blt_slt ? alu_lts : _06826_;
  assign _06256_ = is_sltiu_bltu_sltu ? alu_ltu : _06254_;
  assign _06258_ = instr_bne ? _06824_ : alu_eq;
  assign _06260_ = instr_bge ? _06825_ : _06258_;
  assign alu_out_0 = _00871_ ? _06256_ : _06260_;
  assign _06262_ = _07250_ ? _05579_ : 1'h0;
  assign _06264_ = _07247_ ? _07245_ : _06262_;
  assign _06266_ = _07251_ ? _06264_ : _06278_;
  assign _06268_ = _07272_ ? _05582_ : 1'h0;
  assign _06270_ = _05118_ ? _06266_ : _06268_;
  assign _06272_ = _01078_ ? _00106_[4] : _07260_;
  assign _06274_ = _07250_ ? mem_rdata_latched[11] : 1'h0;
  assign _06276_ = _07265_ ? _07263_ : _06274_;
  assign _06278_ = _05120_ ? _06272_ : _06276_;
  assign _06280_ = _07254_ ? 4'h2 : { _05587_[3:2], _07299_[1], _05587_[0] };
  assign _06282_ = _07250_ ? _05588_ : 4'h0;
  assign _06284_ = _07270_ ? _07301_ : _06282_;
  assign _06286_ = _05122_ ? _06280_ : _06284_;
  assign _06288_ = _07251_ ? _06286_ : _06300_;
  assign _06290_ = _07272_ ? _05592_ : 4'h0;
  assign _06292_ = _05118_ ? _06288_ : _06290_;
  assign _06294_ = _01078_ ? _00106_[3:0] : _07307_;
  assign _06296_ = _07250_ ? mem_rdata_latched[10:7] : 4'h0;
  assign _06298_ = _07265_ ? _07310_ : _06296_;
  assign _06300_ = _05120_ ? _06294_ : _06298_;
  assign _06302_ = _07250_ ? 4'h2 : 4'h0;
  assign _05592_ = _01076_ ? _00106_[3:0] : _06302_;
  assign _06305_ = _07267_ ? _07322_ : _06557_;
  assign _06307_ = _07251_ ? _07318_ : _06305_;
  assign _06309_ = _07251_ ? _07328_ : _06319_;
  assign _06311_ = _07272_ ? _07338_ : _06555_;
  assign _06313_ = _05118_ ? _06309_ : _06311_;
  assign _06315_ = _07247_ ? _07332_ : _07336_;
  assign _06317_ = _00865_ ? 1'h1 : _06555_;
  assign _06319_ = _05124_ ? _06315_ : _06317_;
  assign _06321_ = _07272_ ? _07358_ : _06551_;
  assign _06323_ = _07251_ ? _07356_ : _06321_;
  assign _06325_ = is_beq_bne_blt_bge_bltu_bgeu ? { mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[7], mem_rdata_q[30:25], mem_rdata_q[11:8], 1'h0 } : { mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31:20] };
  assign _06327_ = is_sb_sh_sw ? { mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31:25], mem_rdata_q[11:7] } : _06325_;
  assign _06329_ = instr_jal ? { decoded_imm_j[31:1], 1'h0 } : 32'b0000000000000000000000000000000x;
  assign _06331_ = _07363_ ? { mem_rdata_q[31:12], 12'h000 } : _06329_;
  assign _06333_ = _00873_ ? _06327_ : _06331_;
  assign _06335_ = _07254_ ? mem_rdata_latched[6:2] : _07367_;
  assign _06337_ = _07250_ ? _05612_ : 5'h00;
  assign _06339_ = _05122_ ? _06335_ : _06337_;
  assign _06341_ = _07251_ ? _06339_ : _07373_;
  assign _06343_ = _07272_ ? _05615_ : 5'h00;
  assign _06345_ = _05118_ ? _06341_ : _06343_;
  assign _06347_ = _07247_ ? _07384_ : _07386_;
  assign _06349_ = _07250_ ? _05618_ : 5'h00;
  assign _06351_ = _05126_ ? _06347_ : _06349_;
  assign _06353_ = _07251_ ? _06351_ : _06365_;
  assign _06355_ = _07272_ ? _05621_ : 5'h00;
  assign _06357_ = _05118_ ? _06353_ : _06355_;
  assign _06359_ = _07247_ ? _07393_ : _07395_;
  assign _06361_ = _07397_ ? 5'h01 : 5'h00;
  assign _06363_ = _00865_ ? mem_rdata_latched[11:7] : _06361_;
  assign _06365_ = _05124_ ? _06359_ : _06363_;
  assign _06367_ = _06537_ ? _07443_ : _07444_;
  assign _06369_ = _07439_ ? _07447_ : _07450_;
  assign _06371_ = _05128_ ? _06367_ : _06369_;
  assign _06373_ = _07439_ ? _07461_ : _07465_;
  assign _06375_ = _06535_ ? _07460_ : _06373_;
  assign _05632_ = _07247_ ? _07472_ : _05831_;
  assign _06378_ = _00861_ ? 1'h0 : _05632_;
  assign _06380_ = _07251_ ? _06378_ : _06388_;
  assign _06382_ = _07272_ ? _07481_ : _05831_;
  assign _06384_ = _05118_ ? _06380_ : _06382_;
  assign _06386_ = _07247_ ? _07479_ : _05831_;
  assign _06388_ = _01090_ ? mem_rdata_latched[12] : _06386_;
  assign _06390_ = _07267_ ? _07486_ : _05840_;
  assign _06392_ = _00863_ ? _07484_ : _06390_;
  assign _06394_ = _07270_ ? { mem_rdata_latched[6:4], 2'h0 } : _05844_;
  assign _06396_ = _07247_ ? _07490_ : _06394_;
  assign _06398_ = _07251_ ? _06396_ : _06408_;
  assign _06400_ = _07272_ ? _06412_ : _05844_;
  assign _06402_ = _05118_ ? _06398_ : _06400_;
  assign _06404_ = _07247_ ? _07492_ : _07494_;
  assign _06406_ = _00865_ ? mem_rdata_latched[6:2] : _05844_;
  assign _06408_ = _05124_ ? _06404_ : _06406_;
  assign _06410_ = _07250_ ? { mem_rdata_latched[11], mem_rdata_latched[5], mem_rdata_latched[6], 2'h0 } : _05844_;
  assign _06412_ = _07270_ ? { mem_rdata_latched[11:10], mem_rdata_latched[6], 2'h0 } : _06410_;
  assign _06414_ = _01076_ ? 3'h2 : { _05650_[2], _07508_[1], _05650_[0] };
  assign _06416_ = _07250_ ? 3'h1 : { _05651_[2:1], _05659_[0] };
  assign _06418_ = _05130_ ? _06414_ : _06416_;
  assign _06420_ = _07251_ ? _06418_ : _06432_;
  assign _06422_ = _07272_ ? _06436_ : { _05651_[2:1], _05659_[0] };
  assign _06424_ = _05118_ ? _06420_ : _06422_;
  assign _06426_ = _07253_ ? 3'h1 : 3'h0;
  assign _06428_ = _07265_ ? _07525_ : { _05651_[2:1], _05659_[0] };
  assign _06430_ = _07247_ ? _07523_ : _06428_;
  assign _06432_ = _05132_ ? _06426_ : _06430_;
  assign { _05660_[2], _06434_[1], _05660_[0] } = _07250_ ? 3'h0 : { _05651_[2:1], _05659_[0] };
  assign _06436_ = _01076_ ? 3'h2 : { _05660_[2], _06434_[1], _05660_[0] };
  assign _06438_ = _07251_ ? _07529_ : _07531_;
  assign _06440_ = _07272_ ? _07533_ : _07527_;
  assign _06442_ = _05118_ ? _06438_ : _06440_;
  assign _06444_ = _07254_ ? { 3'h0, mem_rdata_latched[8:7], mem_rdata_latched[12] } : _07539_;
  assign _06446_ = _07250_ ? 6'h00 : _05665_;
  assign _06448_ = _07270_ ? { 3'h0, mem_rdata_latched[3:2], mem_rdata_latched[12] } : _06446_;
  assign _06450_ = _05122_ ? _06444_ : _06448_;
  assign _06452_ = _07251_ ? _06450_ : _06464_;
  assign _06454_ = _07272_ ? _06468_ : _05665_;
  assign _06456_ = _05118_ ? _06452_ : _06454_;
  assign _06458_ = _01078_ ? { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[6:5], mem_rdata_latched[2] } : _07547_;
  assign _06460_ = _00865_ ? { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] } : _05665_;
  assign _06462_ = _07265_ ? _07549_ : _06460_;
  assign _06464_ = _05120_ ? _06458_ : _06462_;
  assign _06466_ = _07250_ ? { 1'h0, mem_rdata_latched[10:7], mem_rdata_latched[12] } : _05665_;
  assign _06468_ = _01076_ ? { 4'h0, mem_rdata_latched[5], mem_rdata_latched[12] } : _06466_;
  assign _06470_ = _07551_ ? { 24'h000000, mem_rdata[31:24] } : { 24'h000000, mem_rdata[23:16] };
  assign _06472_ = _07555_ ? { 24'h000000, mem_rdata[15:8] } : { 24'h000000, mem_rdata[7:0] };
  assign _00064_ = _05134_ ? _06470_ : _06472_;
  assign _00047_ = pcpi_rs1[1] ? { 16'h0000, mem_rdata[31:16] } : { 16'h0000, mem_rdata[15:0] };
  assign _06474_ = _06503_ ? _00047_ : mem_rdata;
  assign mem_rdata_word = _07557_ ? _00064_ : _06474_;
  assign _06476_ = _06503_ ? _07606_ : 4'hf;
  assign mem_la_wstrb = _07557_ ? _07581_ : _06476_;
  assign _06478_ = _06503_ ? { pcpi_rs2[15:0], pcpi_rs2[15:0] } : pcpi_rs2;
  assign mem_la_wdata = _07557_ ? { pcpi_rs2[7:0], pcpi_rs2[7:0], pcpi_rs2[7:0], pcpi_rs2[7:0] } : _06478_;
  assign pcpi_int_rd = pcpi_div_ready ? pcpi_div_rd : pcpi_mul_rd;
  assign _06480_ = pcpi_mul_ready ? pcpi_mul_wr : 1'h0;
  assign pcpi_int_wr = pcpi_div_ready ? pcpi_div_wr : _06480_;
  assign _00875_ = | { _00797_, _07440_, _00948_, _00946_, _00944_, mem_xfer_t0 };
  assign _00876_ = | { _07440_, mem_do_rdata_t0, mem_la_read_t0, mem_xfer_t0 };
  assign _00877_ = | { _07440_, mem_xfer_t0 };
  assign _00878_ = | { _00962_, _00960_, _00958_, _00956_, _00954_, _00952_, _00950_ };
  assign _00879_ = | { _00797_, _00964_, _06837_ };
  assign _00880_ = | { _06892_, _00797_ };
  assign _00881_ = | { _00968_, _00966_, _00958_, _00956_, _00954_ };
  assign _00882_ = | { _00797_, mem_la_write_t0 };
  assign _00883_ = | { _00974_, _00976_ };
  assign _00884_ = | { _00982_, _00980_, _00978_ };
  assign _00885_ = | { _00984_, _00976_ };
  assign _00886_ = | { _00990_, _00988_, _00986_ };
  assign _00887_ = | { _01002_, _01000_, _00998_, _00996_, _00994_, _00992_ };
  assign _00888_ = | { _01018_, _01016_, _01014_, _01012_, _01010_, _01008_, _01006_, _01004_, _00980_, _00978_ };
  assign _00889_ = | { _01018_, _01016_, _01014_, _01010_, _01006_, _01004_, _00980_, _00978_ };
  assign _00890_ = | { _01024_, _01022_, _01020_, _01016_, _01004_, _00980_, _00978_ };
  assign _00891_ = | { decoder_trigger_t0, _06486_, instr_jal_t0 };
  assign _00892_ = | { decoder_trigger_t0, _06486_ };
  assign _00893_ = | { _01028_, _00970_ };
  assign _00894_ = | mem_rdata_t0[1:0];
  assign _00895_ = | next_insn_opcode_t0[1:0];
  assign _04033_ = { _07439_, _00945_, _00943_, _00947_, _00175_, mem_xfer } | { _07440_, _00946_, _00944_, _00948_, _00797_, mem_xfer_t0 };
  assign _04034_ = { _00472_, _07439_, _00467_, mem_xfer } | { mem_la_read_t0, _07440_, mem_do_rdata_t0, mem_xfer_t0 };
  assign _04035_ = { _07439_, mem_xfer } | { _07440_, mem_xfer_t0 };
  assign _04036_ = { _00951_, _00949_, _00959_, _00961_, _00953_, _00955_, _00957_ } | { _00952_, _00950_, _00960_, _00962_, _00954_, _00956_, _00958_ };
  assign _04037_ = { _00963_, _00175_, _06836_ } | { _00964_, _00797_, _06837_ };
  assign _04038_ = { _00175_, _06891_ } | { _00797_, _06892_ };
  assign _04039_ = { _00953_, _00955_, _00957_, _00967_, _00965_ } | { _00954_, _00956_, _00958_, _00968_, _00966_ };
  assign _04040_ = { _00175_, mem_la_write } | { _00797_, mem_la_write_t0 };
  assign _04041_ = { _00975_, _00973_, resetn } | { _00976_, _00974_, 1'h0 };
  assign _04042_ = { _00981_, _00979_, _00977_ } | { _00982_, _00980_, _00978_ };
  assign _04043_ = { _06485_, resetn } | { _06486_, 1'h0 };
  assign _04044_ = { _00983_, _00975_ } | { _00984_, _00976_ };
  assign _04045_ = { _00989_, _00987_, _00985_ } | { _00990_, _00988_, _00986_ };
  assign _04046_ = { _01001_, _00999_, _00997_, _00995_, _00993_, _00991_ } | { _01002_, _01000_, _00998_, _00996_, _00994_, _00992_ };
  assign _04047_ = { _00969_, resetn } | { _00970_, 1'h0 };
  assign _04048_ = { _01017_, _01015_, _01013_, _01011_, _01009_, _01007_, _01005_, _01003_, _00979_, _00977_, resetn } | { _01018_, _01016_, _01014_, _01012_, _01010_, _01008_, _01006_, _01004_, _00980_, _00978_, 1'h0 };
  assign _04049_ = { _01017_, _01015_, _01013_, _01009_, _01005_, _01003_, _00979_, _00977_, resetn } | { _01018_, _01016_, _01014_, _01010_, _01006_, _01004_, _00980_, _00978_, 1'h0 };
  assign _04050_ = { _01023_, _01021_, _01019_, _01015_, _01003_, _00979_, _00977_, resetn } | { _01024_, _01022_, _01020_, _01016_, _01004_, _00980_, _00978_, 1'h0 };
  assign _04051_ = { _00675_, _06485_, decoder_trigger, resetn } | { instr_jal_t0, _06486_, decoder_trigger_t0, 1'h0 };
  assign _04052_ = { _06485_, decoder_trigger } | { _06486_, decoder_trigger_t0 };
  assign _04053_ = { _01027_, _00969_ } | { _01028_, _00970_ };
  assign _05060_ = mem_state | mem_state_t0;
  assign _05061_ = mem_rdata_latched[1:0] | mem_rdata_latched_t0[1:0];
  assign _05062_ = mem_rdata[1:0] | mem_rdata_t0[1:0];
  assign _05063_ = next_insn_opcode[1:0] | next_insn_opcode_t0[1:0];
  assign _00896_ = & _04033_;
  assign _00897_ = & _04034_;
  assign _00898_ = & _04035_;
  assign _00899_ = & _04036_;
  assign _00900_ = & _04037_;
  assign _00901_ = & _04038_;
  assign _00902_ = & _04039_;
  assign _00903_ = & _04040_;
  assign _00904_ = & _04041_;
  assign _00905_ = & _04042_;
  assign _00906_ = & _04043_;
  assign _00907_ = & _04044_;
  assign _00908_ = & _04045_;
  assign _00909_ = & _04046_;
  assign _00910_ = & _04047_;
  assign _00911_ = & _04048_;
  assign _00912_ = & _04049_;
  assign _00913_ = & _04050_;
  assign _00914_ = & _04051_;
  assign _00915_ = & _04052_;
  assign _00916_ = & _04053_;
  assign _00917_ = & _05060_;
  assign _00918_ = & _05061_;
  assign _00919_ = & _05062_;
  assign _00920_ = & _05063_;
  assign _01030_ = _00875_ & _00896_;
  assign _01032_ = _00876_ & _00897_;
  assign _01034_ = _00877_ & _00898_;
  assign _01036_ = _00878_ & _00899_;
  assign _01038_ = _00879_ & _00900_;
  assign _01040_ = _00880_ & _00901_;
  assign _01042_ = _00881_ & _00902_;
  assign _01044_ = _00882_ & _00903_;
  assign _01046_ = _00883_ & _00904_;
  assign _01048_ = _00884_ & _00905_;
  assign _01050_ = _06486_ & _00906_;
  assign _01052_ = _00885_ & _00907_;
  assign _01054_ = _00886_ & _00908_;
  assign _01056_ = _00887_ & _00909_;
  assign _01058_ = _00970_ & _00910_;
  assign _01060_ = _00888_ & _00911_;
  assign _01062_ = _00889_ & _00912_;
  assign _01064_ = _00890_ & _00913_;
  assign _01066_ = _00891_ & _00914_;
  assign _01068_ = _00892_ & _00915_;
  assign _01070_ = _00893_ & _00916_;
  assign _07562_ = _00223_ & _00917_;
  assign _06822_ = _00220_ & _00918_;
  assign _06820_ = _00894_ & _00919_;
  assign _07430_ = _00895_ & _00920_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_timeout_t0 */
  always_ff @(posedge clk)
    if (!resetn) pcpi_timeout_t0 <= 1'h0;
    else pcpi_timeout_t0 <= _06830_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME count_cycle_t0 */
  always_ff @(posedge clk)
    if (!resetn) count_cycle_t0 <= 64'h0000000000000000;
    else count_cycle_t0 <= _00089_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rs2_rdata_t0 */
  always_ff @(posedge clk)
    if (!dbg_rs2val_valid) rvfi_rs2_rdata_t0 <= 32'd0;
    else rvfi_rs2_rdata_t0 <= dbg_rs2val_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rs1_rdata_t0 */
  always_ff @(posedge clk)
    if (_01074_) rvfi_rs1_rdata_t0 <= 32'd0;
    else rvfi_rs1_rdata_t0 <= dbg_rs1val_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rs2_addr_t0 */
  always_ff @(posedge clk)
    if (!dbg_rs2val_valid) rvfi_rs2_addr_t0 <= 5'h00;
    else rvfi_rs2_addr_t0 <= dbg_insn_rs2_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rs1_addr_t0 */
  always_ff @(posedge clk)
    if (_01074_) rvfi_rs1_addr_t0 <= 5'h00;
    else rvfi_rs1_addr_t0 <= dbg_insn_rs1_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_order_t0 */
  always_ff @(posedge clk)
    if (!resetn) rvfi_order_t0 <= 64'h0000000000000000;
    else rvfi_order_t0 <= _00101_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME cpu_state_t0 */
  always_ff @(posedge clk)
    if (_06624_) cpu_state_t0 <= 8'h00;
    else cpu_state_t0 <= _07186_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoder_pseudo_trigger_t0 */
  always_ff @(posedge clk)
    if (!_01075_) decoder_pseudo_trigger_t0 <= 1'h0;
    else decoder_pseudo_trigger_t0 <= _06616_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME last_mem_valid_t0 */
  always_ff @(posedge clk)
    if (!resetn) last_mem_valid_t0 <= 1'h0;
    else last_mem_valid_t0 <= _06662_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_la_firstword_reg_t0 */
  always_ff @(posedge clk)
    if (!resetn) mem_la_firstword_reg_t0 <= 1'h0;
    else mem_la_firstword_reg_t0 <= _07560_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_compare_t0 */
  always_ff @(posedge clk)
    if (_01072_) is_compare_t0 <= 1'h0;
    else is_compare_t0 <= _07574_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME trap_t0 */
  always_ff @(posedge clk)
    if (!resetn) trap_t0 <= 1'h0;
    else trap_t0 <= _06484_;
  assign _00921_ = ~ _00971_;
  assign _00922_ = ~ _01037_;
  assign _05458_ = _07102_ ^ rvfi_mem_wmask;
  assign _05459_ = _07104_ ^ rvfi_mem_rmask;
  assign _05464_ = _07100_ ^ rvfi_mem_rdata;
  assign _05467_ = _07106_ ^ rvfi_mem_addr;
  assign _05474_ = reg_next_pc[0] ^ rvfi_pc_wdata[0];
  assign _05912_ = _07458_ ^ mem_instr;
  assign _05937_ = _07098_ ^ rvfi_mem_wdata;
  assign _03777_ = _07103_ | rvfi_mem_wmask_t0;
  assign _03781_ = _07105_ | rvfi_mem_rmask_t0;
  assign _03805_ = _07101_ | rvfi_mem_rdata_t0;
  assign _03817_ = _07107_ | rvfi_mem_addr_t0;
  assign _03845_ = reg_next_pc_t0[0] | rvfi_pc_wdata_t0[0];
  assign _05190_ = _07459_ | mem_instr_t0;
  assign _05308_ = _07099_ | rvfi_mem_wdata_t0;
  assign _03778_ = _05458_ | _03777_;
  assign _03782_ = _05459_ | _03781_;
  assign _03806_ = _05464_ | _03805_;
  assign _03818_ = _05467_ | _03817_;
  assign _03846_ = _05474_ | _03845_;
  assign _05191_ = _05912_ | _05190_;
  assign _05309_ = _05937_ | _05308_;
  assign _01173_ = { _00971_, _00971_, _00971_, _00971_ } & _07103_;
  assign _01176_ = { _00971_, _00971_, _00971_, _00971_ } & _07105_;
  assign _01195_ = { _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_ } & _07101_;
  assign _01204_ = { _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_ } & _07107_;
  assign _01225_ = launch_next_insn & reg_next_pc_t0[0];
  assign _03496_ = _01037_ & _07459_;
  assign _03585_ = { _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_, _00971_ } & _07099_;
  assign _01174_ = { _00921_, _00921_, _00921_, _00921_ } & rvfi_mem_wmask_t0;
  assign _01177_ = { _00921_, _00921_, _00921_, _00921_ } & rvfi_mem_rmask_t0;
  assign _01196_ = { _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_ } & rvfi_mem_rdata_t0;
  assign _01205_ = { _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_ } & rvfi_mem_addr_t0;
  assign _01226_ = _00139_ & rvfi_pc_wdata_t0[0];
  assign _03497_ = _00922_ & mem_instr_t0;
  assign _03586_ = { _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_, _00921_ } & rvfi_mem_wdata_t0;
  assign _01175_ = _03778_ & { _00972_, _00972_, _00972_, _00972_ };
  assign _01178_ = _03782_ & { _00972_, _00972_, _00972_, _00972_ };
  assign _01197_ = _03806_ & { _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_ };
  assign _01206_ = _03818_ & { _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_ };
  assign _01227_ = _03846_ & launch_next_insn_t0;
  assign _03498_ = _05191_ & _01038_;
  assign _03587_ = _05309_ & { _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_, _00972_ };
  assign _03779_ = _01173_ | _01174_;
  assign _03783_ = _01176_ | _01177_;
  assign _03807_ = _01195_ | _01196_;
  assign _03819_ = _01204_ | _01205_;
  assign _03847_ = _01225_ | _01226_;
  assign _05192_ = _03496_ | _03497_;
  assign _05310_ = _03585_ | _03586_;
  assign _03780_ = _03779_ | _01175_;
  assign _03784_ = _03783_ | _01178_;
  assign _03808_ = _03807_ | _01197_;
  assign _03820_ = _03819_ | _01206_;
  assign _03848_ = _03847_ | _01227_;
  assign _05193_ = _05192_ | _03498_;
  assign _05311_ = _05310_ | _03587_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_wmask_t0 */
  always_ff @(posedge clk)
    if (mem_instr) rvfi_mem_wmask_t0 <= 4'h0;
    else rvfi_mem_wmask_t0 <= _03780_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_rmask_t0 */
  always_ff @(posedge clk)
    if (mem_instr) rvfi_mem_rmask_t0 <= 4'h0;
    else rvfi_mem_rmask_t0 <= _03784_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_rdata_t0 */
  always_ff @(posedge clk)
    if (mem_instr) rvfi_mem_rdata_t0 <= 32'd0;
    else rvfi_mem_rdata_t0 <= _03808_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_addr_t0 */
  always_ff @(posedge clk)
    if (mem_instr) rvfi_mem_addr_t0 <= 32'd0;
    else rvfi_mem_addr_t0 <= _03820_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_pc_wdata_t0[0] */
  always_ff @(posedge clk)
    if (_06599_) rvfi_pc_wdata_t0[0] <= 1'h0;
    else rvfi_pc_wdata_t0[0] <= _03848_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_instr_t0 */
  always_ff @(posedge clk)
    if (mem_do_wdata) mem_instr_t0 <= 1'h0;
    else mem_instr_t0 <= _05193_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_wdata_t0 */
  always_ff @(posedge clk)
    if (mem_instr) rvfi_mem_wdata_t0 <= 32'd0;
    else rvfi_mem_wdata_t0 <= _05311_;
  assign _00923_ = ~ _07143_;
  assign _00924_ = ~ _01047_;
  assign _00925_ = ~ _00975_;
  assign _00926_ = ~ _01051_;
  assign _00927_ = ~ _01053_;
  assign _00928_ = ~ _01055_;
  assign _00929_ = ~ _01025_;
  assign _00930_ = ~ _01065_;
  assign _00931_ = ~ _01067_;
  assign _00932_ = ~ _01069_;
  assign _00933_ = ~ _01031_;
  assign _00934_ = ~ _01033_;
  assign _05437_ = _06697_ ^ instr_bgeu;
  assign _05438_ = _06695_ ^ instr_bltu;
  assign _05439_ = _06693_ ^ instr_bge;
  assign _05440_ = _06691_ ^ instr_blt;
  assign _05441_ = _06689_ ^ instr_bne;
  assign _05442_ = _06687_ ^ instr_beq;
  assign _05448_ = _07585_[3:0] ^ pcpi_timeout_counter;
  assign _05450_ = _06140_ ^ latched_is_lb;
  assign _05451_ = _06142_ ^ latched_is_lh;
  assign _05453_ = _06144_ ^ latched_branch;
  assign _05454_ = _06146_ ^ latched_stalu;
  assign _05455_ = _06154_ ^ latched_store;
  assign _05456_ = _00060_ ^ reg_pc;
  assign _05457_ = _07232_ ^ reg_next_pc;
  assign _05460_ = _07209_ ^ mem_do_rinst;
  assign _05466_ = _06745_ ^ instr_sll;
  assign _05468_ = _07109_ ^ rvfi_rd_wdata;
  assign _05469_ = _07113_ ^ rvfi_rd_addr;
  assign _05471_ = _06610_ ^ mem_do_prefetch;
  assign _05472_ = _00092_ ^ count_instr;
  assign _05473_ = _07238_ ^ pcpi_valid;
  assign _05908_ = _07441_ ^ prefetched_high_word;
  assign _05909_ = _07442_ ^ mem_la_secondword;
  assign _05917_ = _06805_ ^ instr_fence;
  assign _05919_ = _07346_ ^ is_beq_bne_blt_bge_bltu_bgeu;
  assign _05946_ = _06771_ ^ instr_and;
  assign _05947_ = _06767_ ^ instr_or;
  assign _05948_ = _06763_ ^ instr_sra;
  assign _05949_ = _06761_ ^ instr_srl;
  assign _05950_ = _06757_ ^ instr_xor;
  assign _05951_ = _06753_ ^ instr_sltu;
  assign _05952_ = _06749_ ^ instr_slt;
  assign _05953_ = _06741_ ^ instr_sub;
  assign _05954_ = _06739_ ^ instr_add;
  assign _05958_ = _06725_ ^ instr_andi;
  assign _05959_ = _06723_ ^ instr_ori;
  assign _05960_ = _06721_ ^ instr_xori;
  assign _05961_ = _06719_ ^ instr_sltiu;
  assign _05962_ = _06717_ ^ instr_slti;
  assign _05963_ = _06715_ ^ instr_addi;
  assign _03693_ = _06698_ | instr_bgeu_t0;
  assign _03697_ = _06696_ | instr_bltu_t0;
  assign _03701_ = _06694_ | instr_bge_t0;
  assign _03705_ = _06692_ | instr_blt_t0;
  assign _03709_ = _06690_ | instr_bne_t0;
  assign _03713_ = _06688_ | instr_beq_t0;
  assign _03737_ = _07586_[3:0] | pcpi_timeout_counter_t0;
  assign _03745_ = _06141_ | latched_is_lb_t0;
  assign _03749_ = _06143_ | latched_is_lh_t0;
  assign _03757_ = _06145_ | latched_branch_t0;
  assign _03761_ = _06147_ | latched_stalu_t0;
  assign _03765_ = _06155_ | latched_store_t0;
  assign _03769_ = _00061_ | reg_pc_t0;
  assign _03773_ = _07233_ | reg_next_pc_t0;
  assign _03789_ = _07210_ | mem_do_rinst_t0;
  assign _03813_ = _06746_ | instr_sll_t0;
  assign _03821_ = _07110_ | rvfi_rd_wdata_t0;
  assign _03825_ = _07114_ | rvfi_rd_addr_t0;
  assign _03833_ = instr_jalr_t0 | mem_do_prefetch_t0;
  assign _03837_ = _00093_ | count_instr_t0;
  assign _03841_ = _07239_ | pcpi_valid_t0;
  assign _05174_ = _06894_ | prefetched_high_word_t0;
  assign _05178_ = mem_la_read_t0 | mem_la_secondword_t0;
  assign _05224_ = _06806_ | instr_fence_t0;
  assign _05232_ = _07347_ | is_beq_bne_blt_bge_bltu_bgeu_t0;
  assign _05344_ = _06772_ | instr_and_t0;
  assign _05348_ = _06768_ | instr_or_t0;
  assign _05352_ = _06764_ | instr_sra_t0;
  assign _05356_ = _06762_ | instr_srl_t0;
  assign _05360_ = _06758_ | instr_xor_t0;
  assign _05364_ = _06754_ | instr_sltu_t0;
  assign _05368_ = _06750_ | instr_slt_t0;
  assign _05372_ = _06742_ | instr_sub_t0;
  assign _05376_ = _06740_ | instr_add_t0;
  assign _05392_ = _06726_ | instr_andi_t0;
  assign _05396_ = _06724_ | instr_ori_t0;
  assign _05400_ = _06722_ | instr_xori_t0;
  assign _05404_ = _06720_ | instr_sltiu_t0;
  assign _05408_ = _06718_ | instr_slti_t0;
  assign _05412_ = _06716_ | instr_addi_t0;
  assign _03694_ = _05437_ | _03693_;
  assign _03698_ = _05438_ | _03697_;
  assign _03702_ = _05439_ | _03701_;
  assign _03706_ = _05440_ | _03705_;
  assign _03710_ = _05441_ | _03709_;
  assign _03714_ = _05442_ | _03713_;
  assign _03738_ = _05448_ | _03737_;
  assign _03746_ = _05450_ | _03745_;
  assign _03750_ = _05451_ | _03749_;
  assign _03758_ = _05453_ | _03757_;
  assign _03762_ = _05454_ | _03761_;
  assign _03766_ = _05455_ | _03765_;
  assign _03770_ = _05456_ | _03769_;
  assign _03774_ = _05457_ | _03773_;
  assign _03790_ = _05460_ | _03789_;
  assign _03814_ = _05466_ | _03813_;
  assign _03822_ = _05468_ | _03821_;
  assign _03826_ = _05469_ | _03825_;
  assign _03834_ = _05471_ | _03833_;
  assign _03838_ = _05472_ | _03837_;
  assign _03842_ = _05473_ | _03841_;
  assign _05175_ = _05908_ | _05174_;
  assign _05179_ = _05909_ | _05178_;
  assign _05214_ = _00805_ | dbg_valid_insn_t0;
  assign _05225_ = _05917_ | _05224_;
  assign _05233_ = _05919_ | _05232_;
  assign _05345_ = _05946_ | _05344_;
  assign _05349_ = _05947_ | _05348_;
  assign _05353_ = _05948_ | _05352_;
  assign _05357_ = _05949_ | _05356_;
  assign _05361_ = _05950_ | _05360_;
  assign _05365_ = _05951_ | _05364_;
  assign _05369_ = _05952_ | _05368_;
  assign _05373_ = _05953_ | _05372_;
  assign _05377_ = _05954_ | _05376_;
  assign _05393_ = _05958_ | _05392_;
  assign _05397_ = _05959_ | _05396_;
  assign _05401_ = _05960_ | _05400_;
  assign _05405_ = _05961_ | _05404_;
  assign _05409_ = _05962_ | _05408_;
  assign _05413_ = _05963_ | _05412_;
  assign _01110_ = _06685_ & _06698_;
  assign _01113_ = _06685_ & _06696_;
  assign _01116_ = _06685_ & _06694_;
  assign _01119_ = _06685_ & _06692_;
  assign _01122_ = _06685_ & _06690_;
  assign _01125_ = _06685_ & _06688_;
  assign _01143_ = { _07143_, _07143_, _07143_, _07143_ } & _07586_[3:0];
  assign _01149_ = _01047_ & _06141_;
  assign _01152_ = _01047_ & _06143_;
  assign _01158_ = _00975_ & _06145_;
  assign _01161_ = _01051_ & _06147_;
  assign _01164_ = _01053_ & _06155_;
  assign _01167_ = { _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_ } & _00061_;
  assign _01170_ = { _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_, _06485_ } & _07233_;
  assign _01183_ = _01055_ & _07210_;
  assign _01201_ = _06685_ & _06746_;
  assign _01207_ = { _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_, _01025_ } & _07110_;
  assign _01210_ = { _01025_, _01025_, _01025_, _01025_, _01025_ } & _07114_;
  assign _01216_ = _01065_ & instr_jalr_t0;
  assign _01219_ = { _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_, _01067_ } & _00093_;
  assign _01222_ = _01069_ & _07239_;
  assign _03484_ = _01031_ & _06894_;
  assign _03487_ = _01033_ & mem_la_read_t0;
  assign _03522_ = _06685_ & _06806_;
  assign _03528_ = _05738_ & _07347_;
  assign _03612_ = _06685_ & _06772_;
  assign _03615_ = _06685_ & _06768_;
  assign _03618_ = _06685_ & _06764_;
  assign _03621_ = _06685_ & _06762_;
  assign _03624_ = _06685_ & _06758_;
  assign _03627_ = _06685_ & _06754_;
  assign _03630_ = _06685_ & _06750_;
  assign _03633_ = _06685_ & _06742_;
  assign _03636_ = _06685_ & _06740_;
  assign _03648_ = _06685_ & _06726_;
  assign _03651_ = _06685_ & _06724_;
  assign _03654_ = _06685_ & _06722_;
  assign _03657_ = _06685_ & _06720_;
  assign _03660_ = _06685_ & _06718_;
  assign _03663_ = _06685_ & _06716_;
  assign _01111_ = _00130_ & instr_bgeu_t0;
  assign _01114_ = _00130_ & instr_bltu_t0;
  assign _01117_ = _00130_ & instr_bge_t0;
  assign _01120_ = _00130_ & instr_blt_t0;
  assign _01123_ = _00130_ & instr_bne_t0;
  assign _01126_ = _00130_ & instr_beq_t0;
  assign _01144_ = { _00923_, _00923_, _00923_, _00923_ } & pcpi_timeout_counter_t0;
  assign _01150_ = _00924_ & latched_is_lb_t0;
  assign _01153_ = _00924_ & latched_is_lh_t0;
  assign _01159_ = _00925_ & latched_branch_t0;
  assign _01162_ = _00926_ & latched_stalu_t0;
  assign _01165_ = _00927_ & latched_store_t0;
  assign _01168_ = { _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_ } & reg_pc_t0;
  assign _01171_ = { _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_, _00698_ } & reg_next_pc_t0;
  assign _01179_ = _00691_ & mem_do_wdata_t0;
  assign _01181_ = _00691_ & mem_do_rdata_t0;
  assign _01184_ = _00928_ & mem_do_rinst_t0;
  assign _01202_ = _00130_ & instr_sll_t0;
  assign _01208_ = { _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_, _00929_ } & rvfi_rd_wdata_t0;
  assign _01211_ = { _00929_, _00929_, _00929_, _00929_, _00929_ } & rvfi_rd_addr_t0;
  assign _01217_ = _00930_ & mem_do_prefetch_t0;
  assign _01220_ = { _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_, _00931_ } & count_instr_t0;
  assign _01223_ = _00932_ & pcpi_valid_t0;
  assign _03485_ = _00933_ & prefetched_high_word_t0;
  assign _03488_ = _00934_ & mem_la_secondword_t0;
  assign _03514_ = _00139_ & dbg_valid_insn_t0;
  assign _03523_ = _00130_ & instr_fence_t0;
  assign _03529_ = _00131_ & is_beq_bne_blt_bge_bltu_bgeu_t0;
  assign _03613_ = _00130_ & instr_and_t0;
  assign _03616_ = _00130_ & instr_or_t0;
  assign _03619_ = _00130_ & instr_sra_t0;
  assign _03622_ = _00130_ & instr_srl_t0;
  assign _03625_ = _00130_ & instr_xor_t0;
  assign _03628_ = _00130_ & instr_sltu_t0;
  assign _03631_ = _00130_ & instr_slt_t0;
  assign _03634_ = _00130_ & instr_sub_t0;
  assign _03637_ = _00130_ & instr_add_t0;
  assign _03649_ = _00130_ & instr_andi_t0;
  assign _03652_ = _00130_ & instr_ori_t0;
  assign _03655_ = _00130_ & instr_xori_t0;
  assign _03658_ = _00130_ & instr_sltiu_t0;
  assign _03661_ = _00130_ & instr_slti_t0;
  assign _03664_ = _00130_ & instr_addi_t0;
  assign _01112_ = _03694_ & _06686_;
  assign _01115_ = _03698_ & _06686_;
  assign _01118_ = _03702_ & _06686_;
  assign _01121_ = _03706_ & _06686_;
  assign _01124_ = _03710_ & _06686_;
  assign _01127_ = _03714_ & _06686_;
  assign _01145_ = _03738_ & { _06830_, _06830_, _06830_, _06830_ };
  assign _01151_ = _03746_ & _01048_;
  assign _01154_ = _03750_ & _01048_;
  assign _01160_ = _03758_ & _00976_;
  assign _01163_ = _03762_ & _01052_;
  assign _01166_ = _03766_ & _01054_;
  assign _01169_ = _03770_ & { _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_ };
  assign _01172_ = _03774_ & { _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_, _06486_ };
  assign _01180_ = _03785_ & _06873_;
  assign _01182_ = _03787_ & _06873_;
  assign _01185_ = _03790_ & _01056_;
  assign _01203_ = _03814_ & _06686_;
  assign _01209_ = _03822_ & { _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_, _01026_ };
  assign _01212_ = _03826_ & { _01026_, _01026_, _01026_, _01026_, _01026_ };
  assign _01218_ = _03834_ & _01066_;
  assign _01221_ = _03838_ & { _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_, _01068_ };
  assign _01224_ = _03842_ & _01070_;
  assign _03486_ = _05175_ & _01032_;
  assign _03489_ = _05179_ & _01034_;
  assign _03515_ = _05214_ & launch_next_insn_t0;
  assign _03524_ = _05225_ & _06686_;
  assign _03530_ = _05233_ & _06608_;
  assign _03614_ = _05345_ & _06686_;
  assign _03617_ = _05349_ & _06686_;
  assign _03620_ = _05353_ & _06686_;
  assign _03623_ = _05357_ & _06686_;
  assign _03626_ = _05361_ & _06686_;
  assign _03629_ = _05365_ & _06686_;
  assign _03632_ = _05369_ & _06686_;
  assign _03635_ = _05373_ & _06686_;
  assign _03638_ = _05377_ & _06686_;
  assign _03650_ = _05393_ & _06686_;
  assign _03653_ = _05397_ & _06686_;
  assign _03656_ = _05401_ & _06686_;
  assign _03659_ = _05405_ & _06686_;
  assign _03662_ = _05409_ & _06686_;
  assign _03665_ = _05413_ & _06686_;
  assign _03695_ = _01110_ | _01111_;
  assign _03699_ = _01113_ | _01114_;
  assign _03703_ = _01116_ | _01117_;
  assign _03707_ = _01119_ | _01120_;
  assign _03711_ = _01122_ | _01123_;
  assign _03715_ = _01125_ | _01126_;
  assign _03739_ = _01143_ | _01144_;
  assign _03747_ = _01149_ | _01150_;
  assign _03751_ = _01152_ | _01153_;
  assign _03759_ = _01158_ | _01159_;
  assign _03763_ = _01161_ | _01162_;
  assign _03767_ = _01164_ | _01165_;
  assign _03771_ = _01167_ | _01168_;
  assign _03775_ = _01170_ | _01171_;
  assign _03791_ = _01183_ | _01184_;
  assign _03815_ = _01201_ | _01202_;
  assign _03823_ = _01207_ | _01208_;
  assign _03827_ = _01210_ | _01211_;
  assign _03835_ = _01216_ | _01217_;
  assign _03839_ = _01219_ | _01220_;
  assign _03843_ = _01222_ | _01223_;
  assign _05176_ = _03484_ | _03485_;
  assign _05180_ = _03487_ | _03488_;
  assign _05226_ = _03522_ | _03523_;
  assign _05234_ = _03528_ | _03529_;
  assign _05346_ = _03612_ | _03613_;
  assign _05350_ = _03615_ | _03616_;
  assign _05354_ = _03618_ | _03619_;
  assign _05358_ = _03621_ | _03622_;
  assign _05362_ = _03624_ | _03625_;
  assign _05366_ = _03627_ | _03628_;
  assign _05370_ = _03630_ | _03631_;
  assign _05374_ = _03633_ | _03634_;
  assign _05378_ = _03636_ | _03637_;
  assign _05394_ = _03648_ | _03649_;
  assign _05398_ = _03651_ | _03652_;
  assign _05402_ = _03654_ | _03655_;
  assign _05406_ = _03657_ | _03658_;
  assign _05410_ = _03660_ | _03661_;
  assign _05414_ = _03663_ | _03664_;
  assign _03696_ = _03695_ | _01112_;
  assign _03700_ = _03699_ | _01115_;
  assign _03704_ = _03703_ | _01118_;
  assign _03708_ = _03707_ | _01121_;
  assign _03712_ = _03711_ | _01124_;
  assign _03716_ = _03715_ | _01127_;
  assign _03740_ = _03739_ | _01145_;
  assign _03748_ = _03747_ | _01151_;
  assign _03752_ = _03751_ | _01154_;
  assign _03760_ = _03759_ | _01160_;
  assign _03764_ = _03763_ | _01163_;
  assign _03768_ = _03767_ | _01166_;
  assign _03772_ = _03771_ | _01169_;
  assign _03776_ = _03775_ | _01172_;
  assign _03786_ = _01179_ | _01180_;
  assign _03788_ = _01181_ | _01182_;
  assign _03792_ = _03791_ | _01185_;
  assign _03816_ = _03815_ | _01203_;
  assign _03824_ = _03823_ | _01209_;
  assign _03828_ = _03827_ | _01212_;
  assign _03836_ = _03835_ | _01218_;
  assign _03840_ = _03839_ | _01221_;
  assign _03844_ = _03843_ | _01224_;
  assign _05177_ = _05176_ | _03486_;
  assign _05181_ = _05180_ | _03489_;
  assign _05215_ = _03514_ | _03515_;
  assign _05227_ = _05226_ | _03524_;
  assign _05235_ = _05234_ | _03530_;
  assign _05347_ = _05346_ | _03614_;
  assign _05351_ = _05350_ | _03617_;
  assign _05355_ = _05354_ | _03620_;
  assign _05359_ = _05358_ | _03623_;
  assign _05363_ = _05362_ | _03626_;
  assign _05367_ = _05366_ | _03629_;
  assign _05371_ = _05370_ | _03632_;
  assign _05375_ = _05374_ | _03635_;
  assign _05379_ = _05378_ | _03638_;
  assign _05395_ = _05394_ | _03650_;
  assign _05399_ = _05398_ | _03653_;
  assign _05403_ = _05402_ | _03656_;
  assign _05407_ = _05406_ | _03659_;
  assign _05411_ = _05410_ | _03662_;
  assign _05415_ = _05414_ | _03665_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_bgeu_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_bgeu_t0 <= 1'h0;
    else instr_bgeu_t0 <= _03696_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_bltu_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_bltu_t0 <= 1'h0;
    else instr_bltu_t0 <= _03700_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_bge_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_bge_t0 <= 1'h0;
    else instr_bge_t0 <= _03704_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_blt_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_blt_t0 <= 1'h0;
    else instr_blt_t0 <= _03708_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_bne_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_bne_t0 <= 1'h0;
    else instr_bne_t0 <= _03712_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_beq_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_beq_t0 <= 1'h0;
    else instr_beq_t0 <= _03716_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_timeout_counter_t0 */
  always_ff @(posedge clk)
    if (!_06607_) pcpi_timeout_counter_t0 <= 4'h0;
    else pcpi_timeout_counter_t0 <= _03740_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_is_lb_t0 */
  always_ff @(posedge clk)
    if (!resetn) latched_is_lb_t0 <= 1'h0;
    else latched_is_lb_t0 <= _03748_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_is_lh_t0 */
  always_ff @(posedge clk)
    if (!resetn) latched_is_lh_t0 <= 1'h0;
    else latched_is_lh_t0 <= _03752_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_branch_t0 */
  always_ff @(posedge clk)
    if (!resetn) latched_branch_t0 <= 1'h0;
    else latched_branch_t0 <= _03760_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_stalu_t0 */
  always_ff @(posedge clk)
    if (!resetn) latched_stalu_t0 <= 1'h0;
    else latched_stalu_t0 <= _03764_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_store_t0 */
  always_ff @(posedge clk)
    if (!resetn) latched_store_t0 <= 1'h0;
    else latched_store_t0 <= _03768_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME reg_pc_t0 */
  always_ff @(posedge clk)
    if (!resetn) reg_pc_t0 <= 32'd0;
    else reg_pc_t0 <= _03772_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME reg_next_pc_t0 */
  always_ff @(posedge clk)
    if (!resetn) reg_next_pc_t0 <= 32'd0;
    else reg_next_pc_t0 <= _03776_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_do_wdata_t0 */
  always_ff @(posedge clk)
    if (_00034_) mem_do_wdata_t0 <= 1'h0;
    else mem_do_wdata_t0 <= _03786_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_do_rdata_t0 */
  always_ff @(posedge clk)
    if (_00032_) mem_do_rdata_t0 <= 1'h0;
    else mem_do_rdata_t0 <= _03788_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_do_rinst_t0 */
  always_ff @(posedge clk)
    if (_00033_) mem_do_rinst_t0 <= 1'h0;
    else mem_do_rinst_t0 <= _03792_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sll_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_sll_t0 <= 1'h0;
    else instr_sll_t0 <= _03816_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rd_wdata_t0 */
  always_ff @(posedge clk)
    if (_01073_) rvfi_rd_wdata_t0 <= 32'd0;
    else rvfi_rd_wdata_t0 <= _03824_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rd_addr_t0 */
  always_ff @(posedge clk)
    if (_01073_) rvfi_rd_addr_t0 <= 5'h00;
    else rvfi_rd_addr_t0 <= _03828_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_do_prefetch_t0 */
  always_ff @(posedge clk)
    if (_06872_) mem_do_prefetch_t0 <= 1'h0;
    else mem_do_prefetch_t0 <= _03836_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME count_instr_t0 */
  always_ff @(posedge clk)
    if (!resetn) count_instr_t0 <= 64'h0000000000000000;
    else count_instr_t0 <= _03840_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_valid_t0 */
  always_ff @(posedge clk)
    if (!resetn) pcpi_valid_t0 <= 1'h0;
    else pcpi_valid_t0 <= _03844_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME prefetched_high_word_t0 */
  always_ff @(posedge clk)
    if (_01071_) prefetched_high_word_t0 <= 1'h0;
    else prefetched_high_word_t0 <= _05177_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_la_secondword_t0 */
  always_ff @(posedge clk)
    if (_06888_) mem_la_secondword_t0 <= 1'h0;
    else mem_la_secondword_t0 <= _05181_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_valid_insn_t0 */
  always_ff @(posedge clk)
    if (_06888_) dbg_valid_insn_t0 <= 1'h0;
    else dbg_valid_insn_t0 <= _05215_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_fence_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_fence_t0 <= 1'h0;
    else instr_fence_t0 <= _05227_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_beq_bne_blt_bge_bltu_bgeu_t0 */
  always_ff @(posedge clk)
    if (!resetn) is_beq_bne_blt_bge_bltu_bgeu_t0 <= 1'h0;
    else is_beq_bne_blt_bge_bltu_bgeu_t0 <= _05235_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_and_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_and_t0 <= 1'h0;
    else instr_and_t0 <= _05347_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_or_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_or_t0 <= 1'h0;
    else instr_or_t0 <= _05351_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sra_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_sra_t0 <= 1'h0;
    else instr_sra_t0 <= _05355_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_srl_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_srl_t0 <= 1'h0;
    else instr_srl_t0 <= _05359_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_xor_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_xor_t0 <= 1'h0;
    else instr_xor_t0 <= _05363_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sltu_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_sltu_t0 <= 1'h0;
    else instr_sltu_t0 <= _05367_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_slt_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_slt_t0 <= 1'h0;
    else instr_slt_t0 <= _05371_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sub_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_sub_t0 <= 1'h0;
    else instr_sub_t0 <= _05375_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_add_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_add_t0 <= 1'h0;
    else instr_add_t0 <= _05379_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_andi_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_andi_t0 <= 1'h0;
    else instr_andi_t0 <= _05395_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_ori_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_ori_t0 <= 1'h0;
    else instr_ori_t0 <= _05399_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_xori_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_xori_t0 <= 1'h0;
    else instr_xori_t0 <= _05403_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sltiu_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_sltiu_t0 <= 1'h0;
    else instr_sltiu_t0 <= _05407_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_slti_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_slti_t0 <= 1'h0;
    else instr_slti_t0 <= _05411_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_addi_t0 */
  always_ff @(posedge clk)
    if (!resetn) instr_addi_t0 <= 1'h0;
    else instr_addi_t0 <= _05415_;
  assign _06482_ = 4'h0 << pcpi_rs1[1:0];
  assign _07582_ = { _00224_, _00224_, _00224_, _00224_ } | _06482_;
  assign _00935_ = ~ { 28'h0000000, pcpi_timeout_counter_t0 };
  assign _00936_ = ~ { 27'h0000000, reg_sh_t0 };
  assign _03323_ = { 28'h0000000, pcpi_timeout_counter } & _00935_;
  assign _03324_ = { 27'h0000000, reg_sh } & _00936_;
  assign _05067_ = { 28'h0000000, pcpi_timeout_counter } | { 28'h0000000, pcpi_timeout_counter_t0 };
  assign _05068_ = { 27'h0000000, reg_sh } | { 27'h0000000, reg_sh_t0 };
  assign _06094_ = _05064_ - _03322_;
  assign _06096_ = _05067_ - 32'd1;
  assign _06098_ = _05068_ - 32'd4;
  assign _06100_ = _05068_ - 32'd1;
  assign _06095_ = _03321_ - _05065_;
  assign _06097_ = _03323_ - 32'd1;
  assign _06099_ = _03324_ - 32'd4;
  assign _06101_ = _03324_ - 32'd1;
  assign _05880_ = _06094_ ^ _06095_;
  assign _05881_ = _06096_ ^ _06097_;
  assign _05882_ = _06098_ ^ _06099_;
  assign _05883_ = _06100_ ^ _06101_;
  assign _05066_ = _05880_ | pcpi_rs1_t0;
  assign _07586_ = _05881_ | { 28'h0000000, pcpi_timeout_counter_t0 };
  assign _07588_ = _05882_ | { 27'h0000000, reg_sh_t0 };
  assign _07590_ = _05883_ | { 27'h0000000, reg_sh_t0 };
  assign _07584_ = _05066_ | pcpi_rs2_t0;
  assign alu_eq = pcpi_rs1 == /* src = "generated/out/vanilla.sv:1111.14-1111.32" */ pcpi_rs2;
  assign _06499_ = ! /* src = "generated/out/vanilla.sv:1579.10-1579.21" */ reg_sh;
  assign _06505_ = rvfi_insn[6:0] == /* src = "generated/out/vanilla.sv:1792.23-1792.51" */ 7'h73;
  assign _06507_ = rvfi_insn[13:12] == /* src = "generated/out/vanilla.sv:1792.58-1792.84" */ 2'h2;
  assign _06509_ = rvfi_insn[31:20] == /* src = "generated/out/vanilla.sv:1793.8-1793.35" */ 12'hc00;
  assign _06510_ = rvfi_insn[31:20] == /* src = "generated/out/vanilla.sv:1797.8-1797.35" */ 12'hc80;
  assign _06512_ = rvfi_insn[31:20] == /* src = "generated/out/vanilla.sv:1801.8-1801.35" */ 12'hc02;
  assign _06513_ = rvfi_insn[31:20] == /* src = "generated/out/vanilla.sv:1805.8-1805.35" */ 12'hc82;
  assign _06517_ = ! /* src = "generated/out/vanilla.sv:379.12-379.45" */ mem_rdata_latched[11:10];
  assign _06519_ = mem_rdata_latched[11:10] == /* src = "generated/out/vanilla.sv:383.12-383.45" */ 2'h1;
  assign _06527_ = mem_rdata_latched[6:5] == /* src = "generated/out/vanilla.sv:394.13-394.44" */ 2'h1;
  assign _06529_ = mem_rdata_latched[6:5] == /* src = "generated/out/vanilla.sv:396.13-396.44" */ 2'h2;
  assign _06531_ = mem_rdata_latched[6:5] == /* src = "generated/out/vanilla.sv:398.13-398.44" */ 2'h3;
  assign _06525_ = ! /* src = "generated/out/vanilla.sv:400.32-400.63" */ mem_rdata_latched[6:5];
  assign _06539_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:797.17-797.53" */ 7'h37;
  assign _06541_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:798.19-798.55" */ 7'h17;
  assign _06543_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:799.17-799.53" */ 7'h6f;
  assign _06545_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:800.19-800.55" */ 7'h67;
  assign _06547_ = ! /* src = "generated/out/vanilla.sv:800.61-800.95" */ mem_rdata_latched[14:12];
  assign _06549_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:803.36-803.72" */ 7'h63;
  assign _06551_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:804.27-804.63" */ 7'h03;
  assign _06553_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:805.19-805.55" */ 7'h23;
  assign _06555_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:806.22-806.58" */ 7'h13;
  assign _06557_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:807.22-807.58" */ 7'h33;
  assign _06515_ = mem_rdata_latched[11:7] == /* src = "generated/out/vanilla.sv:860.14-860.42" */ 5'h02;
  assign _06521_ = mem_rdata_latched[11:10] == /* src = "generated/out/vanilla.sv:877.13-877.46" */ 2'h2;
  assign _06523_ = mem_rdata_latched[12:10] == /* src = "generated/out/vanilla.sv:882.13-882.47" */ 3'h3;
  assign _06533_ = ! /* src = "generated/out/vanilla.sv:928.82-928.109" */ mem_rdata_latched[6:2];
  assign _06581_ = mem_rdata_q[31:20] == /* src = "generated/out/vanilla.sv:984.61-984.97" */ 12'hb00;
  assign _06583_ = mem_rdata_q[31:20] == /* src = "generated/out/vanilla.sv:984.174-984.210" */ 12'hb01;
  assign _06585_ = mem_rdata_q[31:20] == /* src = "generated/out/vanilla.sv:985.63-985.99" */ 12'hb80;
  assign _06587_ = mem_rdata_q[31:20] == /* src = "generated/out/vanilla.sv:985.176-985.212" */ 12'hb81;
  assign _06589_ = mem_rdata_q[31:20] == /* src = "generated/out/vanilla.sv:986.60-986.96" */ 12'hb02;
  assign _06591_ = mem_rdata_q[31:20] == /* src = "generated/out/vanilla.sv:987.62-987.98" */ 12'hb82;
  assign _06579_ = mem_rdata_q[6:0] == /* src = "generated/out/vanilla.sv:988.29-988.59" */ 7'h73;
  assign _06593_ = mem_rdata_q[15:0] == /* src = "generated/out/vanilla.sv:988.131-988.160" */ 16'h9002;
  assign _06595_ = mem_rdata_q[6:0] == /* src = "generated/out/vanilla.sv:989.20-989.50" */ 7'h0f;
  assign _06569_ = mem_rdata_q[14:12] == /* src = "generated/out/vanilla.sv:995.230-995.258" */ 3'h7;
  assign _06567_ = mem_rdata_q[14:12] == /* src = "generated/out/vanilla.sv:995.200-995.228" */ 3'h6;
  assign _06563_ = mem_rdata_q[14:12] == /* src = "generated/out/vanilla.sv:995.170-995.198" */ 3'h4;
  assign _06573_ = mem_rdata_q[14:12] == /* src = "generated/out/vanilla.sv:995.140-995.168" */ 3'h3;
  assign _06571_ = mem_rdata_q[14:12] == /* src = "generated/out/vanilla.sv:995.110-995.138" */ 3'h2;
  assign _06559_ = ! /* src = "generated/out/vanilla.sv:995.80-995.108" */ mem_rdata_q[14:12];
  assign _06577_ = mem_rdata_q[31:25] == /* src = "generated/out/vanilla.sv:996.217-996.249" */ 7'h20;
  assign _06565_ = mem_rdata_q[14:12] == /* src = "generated/out/vanilla.sv:996.113-996.141" */ 3'h5;
  assign _06561_ = mem_rdata_q[14:12] == /* src = "generated/out/vanilla.sv:996.43-996.71" */ 3'h1;
  assign _06575_ = ! /* src = "generated/out/vanilla.sv:996.77-996.109" */ mem_rdata_q[31:25];
  assign _06597_ = reg_sh >= /* src = "generated/out/vanilla.sv:1584.35-1584.46" */ 32'd4;
  assign _06599_ = latched_store && /* src = "generated/out/vanilla.sv:1080.20-1080.51" */ latched_branch;
  assign _06603_ = resetn && /* src = "generated/out/vanilla.sv:1181.8-1181.31" */ cpuregs_write;
  assign _06605_ = _06603_ && /* src = "generated/out/vanilla.sv:1181.7-1181.46" */ latched_rd;
  assign launch_next_insn = _06485_ && /* src = "generated/out/vanilla.sv:1195.29-1195.78" */ decoder_trigger;
  assign _06606_ = resetn && /* src = "generated/out/vanilla.sv:1214.9-1214.29" */ pcpi_valid;
  assign _06607_ = _06606_ && /* src = "generated/out/vanilla.sv:1214.8-1214.48" */ _06828_;
  assign _05738_ = mem_do_rinst && /* src = "generated/out/vanilla.sv:1234.22-1234.46" */ mem_done;
  assign _06601_ = latched_store && /* src = "generated/out/vanilla.sv:1281.7-1281.39" */ _06827_;
  assign _06613_ = is_lb_lh_lw_lbu_lhu && /* src = "generated/out/vanilla.sv:1454.7-1454.41" */ _06831_;
  assign _06615_ = _06832_ && /* src = "generated/out/vanilla.sv:1648.11-1648.39" */ mem_done;
  assign _06617_ = resetn && /* src = "generated/out/vanilla.sv:1668.7-1668.67" */ _06870_;
  assign _06619_ = _06501_ && /* src = "generated/out/vanilla.sv:1669.8-1669.50" */ _07087_;
  assign _06621_ = _06503_ && /* src = "generated/out/vanilla.sv:1674.8-1674.48" */ pcpi_rs1[0];
  assign _06623_ = resetn && /* src = "generated/out/vanilla.sv:1680.8-1680.50" */ mem_do_rinst;
  assign _06624_ = _06623_ && /* src = "generated/out/vanilla.sv:1680.7-1680.98" */ reg_pc[0];
  assign _06625_ = resetn && /* src = "generated/out/vanilla.sv:1715.18-1715.54" */ _06874_;
  assign _00030_ = _06625_ && /* src = "generated/out/vanilla.sv:1715.17-1715.73" */ dbg_valid_insn;
  assign _06627_ = mem_valid && /* src = "generated/out/vanilla.sv:1774.13-1774.43" */ mem_ready;
  assign _06629_ = rvfi_valid && /* src = "generated/out/vanilla.sv:1792.8-1792.52" */ _06505_;
  assign _06631_ = _06629_ && /* src = "generated/out/vanilla.sv:1792.7-1792.85" */ _06507_;
  assign _06635_ = _06633_ && /* src = "generated/out/vanilla.sv:286.27-286.94" */ next_pc[1];
  assign mem_la_firstword = _06635_ && /* src = "generated/out/vanilla.sv:286.26-286.117" */ _06833_;
  assign _06637_ = mem_la_firstword && /* src = "generated/out/vanilla.sv:293.42-293.102" */ prefetched_high_word;
  assign mem_la_use_prefetched_high_word = _06637_ && /* src = "generated/out/vanilla.sv:293.41-293.134" */ _06834_;
  assign _06639_ = mem_la_use_prefetched_high_word && /* src = "generated/out/vanilla.sv:294.49-294.96" */ mem_do_rinst;
  assign _06641_ = mem_xfer && /* src = "generated/out/vanilla.sv:296.32-296.54" */ _07572_;
  assign _06643_ = _06641_ && /* src = "generated/out/vanilla.sv:296.31-296.107" */ _06878_;
  assign _06645_ = _07561_ && /* src = "generated/out/vanilla.sv:296.113-296.139" */ mem_do_rinst;
  assign _06647_ = resetn && /* src = "generated/out/vanilla.sv:296.19-296.141" */ _06880_;
  assign _06649_ = _06821_ && /* src = "generated/out/vanilla.sv:296.169-296.205" */ mem_xfer;
  assign mem_done = _06647_ && /* src = "generated/out/vanilla.sv:296.18-296.207" */ _06882_;
  assign _06651_ = resetn && /* src = "generated/out/vanilla.sv:297.25-297.45" */ _06836_;
  assign mem_la_write = _06651_ && /* src = "generated/out/vanilla.sv:297.24-297.62" */ mem_do_wdata;
  assign _06653_ = _06838_ && /* src = "generated/out/vanilla.sv:298.36-298.82" */ _06836_;
  assign _06655_ = _06653_ && /* src = "generated/out/vanilla.sv:298.35-298.138" */ _06884_;
  assign mem_la_firstword_xfer = mem_xfer && /* src = "generated/out/vanilla.sv:298.146-298.237" */ _07559_;
  assign _06657_ = mem_la_firstword_xfer && /* src = "generated/out/vanilla.sv:298.145-298.260" */ _06833_;
  assign _06659_ = _06657_ && /* src = "generated/out/vanilla.sv:298.144-298.288" */ _07563_;
  assign mem_la_read = resetn && /* src = "generated/out/vanilla.sv:298.23-298.290" */ _06886_;
  assign _06661_ = mem_valid && /* src = "generated/out/vanilla.sv:310.22-310.45" */ _06839_;
  assign _06663_ = mem_done && /* src = "generated/out/vanilla.sv:344.7-344.72" */ _06633_;
  assign _06665_ = _00704_ && /* src = "generated/out/vanilla.sv:423.12-423.73" */ _06533_;
  assign _06675_ = _06545_ && /* src = "generated/out/vanilla.sv:800.18-800.96" */ _06547_;
  assign _06679_ = _06840_ && /* src = "generated/out/vanilla.sv:871.13-871.61" */ _06841_;
  assign _06681_ = _00704_ && /* src = "generated/out/vanilla.sv:917.14-917.76" */ _07090_;
  assign _06683_ = _06681_ && /* src = "generated/out/vanilla.sv:917.13-917.110" */ _06533_;
  assign _06667_ = _00704_ && /* src = "generated/out/vanilla.sv:922.13-922.74" */ _07089_;
  assign _06669_ = mem_rdata_latched[12] && /* src = "generated/out/vanilla.sv:928.14-928.76" */ _07090_;
  assign _06671_ = _06669_ && /* src = "generated/out/vanilla.sv:928.13-928.110" */ _06533_;
  assign _06673_ = mem_rdata_latched[12] && /* src = "generated/out/vanilla.sv:933.13-933.74" */ _07089_;
  assign _06685_ = decoder_trigger && /* src = "generated/out/vanilla.sv:949.7-949.49" */ _06842_;
  assign _06687_ = is_beq_bne_blt_bge_bltu_bgeu && /* src = "generated/out/vanilla.sv:951.17-951.79" */ _06559_;
  assign _06689_ = is_beq_bne_blt_bge_bltu_bgeu && /* src = "generated/out/vanilla.sv:952.17-952.79" */ _06561_;
  assign _06691_ = is_beq_bne_blt_bge_bltu_bgeu && /* src = "generated/out/vanilla.sv:953.17-953.79" */ _06563_;
  assign _06693_ = is_beq_bne_blt_bge_bltu_bgeu && /* src = "generated/out/vanilla.sv:954.17-954.79" */ _06565_;
  assign _06695_ = is_beq_bne_blt_bge_bltu_bgeu && /* src = "generated/out/vanilla.sv:955.18-955.80" */ _06567_;
  assign _06697_ = is_beq_bne_blt_bge_bltu_bgeu && /* src = "generated/out/vanilla.sv:956.18-956.80" */ _06569_;
  assign _06699_ = is_lb_lh_lw_lbu_lhu && /* src = "generated/out/vanilla.sv:957.16-957.69" */ _06559_;
  assign _06701_ = is_lb_lh_lw_lbu_lhu && /* src = "generated/out/vanilla.sv:958.16-958.69" */ _06561_;
  assign _06703_ = is_lb_lh_lw_lbu_lhu && /* src = "generated/out/vanilla.sv:959.16-959.69" */ _06571_;
  assign _06705_ = is_lb_lh_lw_lbu_lhu && /* src = "generated/out/vanilla.sv:960.17-960.70" */ _06563_;
  assign _06707_ = is_lb_lh_lw_lbu_lhu && /* src = "generated/out/vanilla.sv:961.17-961.70" */ _06565_;
  assign _06709_ = is_sb_sh_sw && /* src = "generated/out/vanilla.sv:962.16-962.61" */ _06559_;
  assign _06711_ = is_sb_sh_sw && /* src = "generated/out/vanilla.sv:963.16-963.61" */ _06561_;
  assign _06713_ = is_sb_sh_sw && /* src = "generated/out/vanilla.sv:964.16-964.61" */ _06571_;
  assign _06715_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:965.18-965.66" */ _06559_;
  assign _06717_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:966.18-966.66" */ _06571_;
  assign _06719_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:967.19-967.67" */ _06573_;
  assign _06721_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:968.18-968.66" */ _06563_;
  assign _06723_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:969.17-969.65" */ _06567_;
  assign _06725_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:970.18-970.66" */ _06569_;
  assign _06727_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:971.19-971.67" */ _06561_;
  assign _06729_ = _06727_ && /* src = "generated/out/vanilla.sv:971.18-971.106" */ _06575_;
  assign _06733_ = _06731_ && /* src = "generated/out/vanilla.sv:972.18-972.106" */ _06575_;
  assign _06731_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:973.19-973.67" */ _06565_;
  assign _06735_ = _06731_ && /* src = "generated/out/vanilla.sv:973.18-973.106" */ _06577_;
  assign _06739_ = _06737_ && /* src = "generated/out/vanilla.sv:974.17-974.105" */ _06575_;
  assign _06737_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:975.18-975.66" */ _06559_;
  assign _06741_ = _06737_ && /* src = "generated/out/vanilla.sv:975.17-975.105" */ _06577_;
  assign _06743_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:976.18-976.66" */ _06561_;
  assign _06745_ = _06743_ && /* src = "generated/out/vanilla.sv:976.17-976.105" */ _06575_;
  assign _06747_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:977.18-977.66" */ _06571_;
  assign _06749_ = _06747_ && /* src = "generated/out/vanilla.sv:977.17-977.105" */ _06575_;
  assign _06751_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:978.19-978.67" */ _06573_;
  assign _06753_ = _06751_ && /* src = "generated/out/vanilla.sv:978.18-978.106" */ _06575_;
  assign _06755_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:979.18-979.66" */ _06563_;
  assign _06757_ = _06755_ && /* src = "generated/out/vanilla.sv:979.17-979.105" */ _06575_;
  assign _06761_ = _06759_ && /* src = "generated/out/vanilla.sv:980.17-980.105" */ _06575_;
  assign _06759_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:981.18-981.66" */ _06565_;
  assign _06763_ = _06759_ && /* src = "generated/out/vanilla.sv:981.17-981.105" */ _06577_;
  assign _06765_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:982.17-982.65" */ _06567_;
  assign _06767_ = _06765_ && /* src = "generated/out/vanilla.sv:982.16-982.104" */ _06575_;
  assign _06769_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:983.18-983.66" */ _06569_;
  assign _06771_ = _06769_ && /* src = "generated/out/vanilla.sv:983.17-983.105" */ _06575_;
  assign _06773_ = _06579_ && /* src = "generated/out/vanilla.sv:984.24-984.98" */ _06581_;
  assign _06775_ = _06773_ && /* src = "generated/out/vanilla.sv:984.23-984.130" */ _07092_;
  assign _06777_ = _06579_ && /* src = "generated/out/vanilla.sv:984.137-984.211" */ _06583_;
  assign _06779_ = _06777_ && /* src = "generated/out/vanilla.sv:984.136-984.243" */ _07092_;
  assign _06783_ = _06579_ && /* src = "generated/out/vanilla.sv:985.26-985.100" */ _06585_;
  assign _06785_ = _06783_ && /* src = "generated/out/vanilla.sv:985.25-985.132" */ _07092_;
  assign _06787_ = _06579_ && /* src = "generated/out/vanilla.sv:985.139-985.213" */ _06587_;
  assign _06789_ = _06787_ && /* src = "generated/out/vanilla.sv:985.138-985.245" */ _07092_;
  assign _06793_ = _06579_ && /* src = "generated/out/vanilla.sv:986.23-986.97" */ _06589_;
  assign _06795_ = _06793_ && /* src = "generated/out/vanilla.sv:986.22-986.129" */ _07092_;
  assign _06797_ = _06579_ && /* src = "generated/out/vanilla.sv:987.25-987.99" */ _06591_;
  assign _06799_ = _06797_ && /* src = "generated/out/vanilla.sv:987.24-987.131" */ _07092_;
  assign _06801_ = _06579_ && /* src = "generated/out/vanilla.sv:988.28-988.83" */ _06843_;
  assign _06803_ = _06801_ && /* src = "generated/out/vanilla.sv:988.27-988.106" */ _06845_;
  assign _06805_ = _06595_ && /* src = "generated/out/vanilla.sv:989.19-989.74" */ _06847_;
  assign _06813_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:994.25-994.254" */ _07577_;
  assign _06815_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:995.60-995.259" */ _07579_;
  assign _06807_ = _06565_ && /* src = "generated/out/vanilla.sv:996.182-996.250" */ _06577_;
  assign _06809_ = _06565_ && /* src = "generated/out/vanilla.sv:996.112-996.180" */ _06575_;
  assign _06811_ = _06561_ && /* src = "generated/out/vanilla.sv:996.42-996.110" */ _06575_;
  assign _06817_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:996.22-996.251" */ _07577_;
  assign _06819_ = ! /* src = "generated/out/vanilla.sv:0.0-0.0" */ _00475_;
  assign _06821_ = ! /* src = "generated/out/vanilla.sv:0.0-0.0" */ _07563_;
  assign _06824_ = ! /* src = "generated/out/vanilla.sv:1124.27-1124.34" */ alu_eq;
  assign _06825_ = ! /* src = "generated/out/vanilla.sv:1125.27-1125.35" */ alu_lts;
  assign _06826_ = ! /* src = "generated/out/vanilla.sv:1126.28-1126.36" */ alu_ltu;
  assign _06828_ = ! /* src = "generated/out/vanilla.sv:1214.34-1214.48" */ pcpi_int_wait;
  assign _06829_ = ! /* src = "generated/out/vanilla.sv:1220.20-1220.41" */ pcpi_timeout_counter;
  assign _06609_ = ! /* src = "generated/out/vanilla.sv:1275.22-1275.38" */ decoder_trigger;
  assign _06827_ = ! /* src = "generated/out/vanilla.sv:1281.24-1281.39" */ latched_branch;
  assign _06610_ = ! /* src = "generated/out/vanilla.sv:1346.27-1346.38" */ instr_jalr;
  assign _06831_ = ! /* src = "generated/out/vanilla.sv:1454.30-1454.41" */ instr_trap;
  assign _06832_ = ! /* src = "generated/out/vanilla.sv:1648.11-1648.27" */ mem_do_prefetch;
  assign _06823_ = ! /* src = "generated/out/vanilla.sv:1740.7-1740.14" */ resetn;
  assign _06834_ = ! /* src = "generated/out/vanilla.sv:293.107-293.134" */ clear_prefetched_high_word;
  assign _06835_ = ! /* src = "generated/out/vanilla.sv:296.147-296.164" */ mem_la_firstword;
  assign _06833_ = ! /* src = "generated/out/vanilla.sv:298.242-298.260" */ mem_la_secondword;
  assign _06839_ = ! /* src = "generated/out/vanilla.sv:310.35-310.45" */ mem_ready;
  assign _06838_ = ! /* src = "generated/out/vanilla.sv:499.12-499.44" */ mem_la_use_prefetched_high_word;
  assign instr_trap = ! /* src = "generated/out/vanilla.sv:608.54-608.626" */ { instr_lui, instr_auipc, instr_jal, instr_jalr, instr_beq, instr_bne, instr_blt, instr_bge, instr_bltu, instr_bgeu, instr_lb, instr_lh, instr_lw, instr_lbu, instr_lhu, instr_sb, instr_sh, instr_sw, instr_addi, instr_slti, instr_sltiu, instr_xori, instr_ori, instr_andi, instr_slli, instr_srli, instr_srai, instr_add, instr_sub, instr_sll, instr_slt, instr_sltu, instr_xor, instr_srl, instr_sra, instr_or, instr_and, instr_rdcycle, instr_rdcycleh, instr_rdinstr, instr_rdinstrh, instr_fence, 6'h00 };
  assign _06840_ = ! /* src = "generated/out/vanilla.sv:871.13-871.35" */ mem_rdata_latched[11];
  assign _06841_ = ! /* src = "generated/out/vanilla.sv:904.13-904.35" */ mem_rdata_latched[12];
  assign _06842_ = ! /* src = "generated/out/vanilla.sv:949.26-949.49" */ decoder_pseudo_trigger;
  assign _06843_ = ! /* src = "generated/out/vanilla.sv:988.64-988.83" */ mem_rdata_q[31:21];
  assign _06845_ = ! /* src = "generated/out/vanilla.sv:988.88-988.106" */ mem_rdata_q[19:7];
  assign _06847_ = ! /* src = "generated/out/vanilla.sv:989.55-989.74" */ mem_rdata_q[15:12];
  assign _06849_ = instr_sra || /* src = "generated/out/vanilla.sv:1115.25-1115.48" */ instr_srai;
  assign _06851_ = instr_xori || /* src = "generated/out/vanilla.sv:1135.4-1135.27" */ instr_xor;
  assign _06853_ = instr_ori || /* src = "generated/out/vanilla.sv:1136.4-1136.25" */ instr_or;
  assign _06855_ = instr_andi || /* src = "generated/out/vanilla.sv:1137.4-1137.27" */ instr_and;
  assign _06861_ = latched_branch || /* src = "generated/out/vanilla.sv:1148.8-1148.35" */ 2'h0;
  assign _06863_ = _06861_ || /* src = "generated/out/vanilla.sv:1148.7-1148.47" */ _06823_;
  assign _06611_ = pcpi_timeout || /* src = "generated/out/vanilla.sv:1527.35-1527.69" */ instr_ecall_ebreak;
  assign _06857_ = instr_slli || /* src = "generated/out/vanilla.sv:1596.8-1596.31" */ instr_sll;
  assign _06859_ = instr_srli || /* src = "generated/out/vanilla.sv:1597.8-1597.31" */ instr_srl;
  assign _06865_ = _06832_ || /* src = "generated/out/vanilla.sv:1630.10-1630.38" */ mem_done;
  assign _06867_ = instr_lb || /* src = "generated/out/vanilla.sv:1634.9-1634.30" */ instr_lbu;
  assign _06869_ = instr_lh || /* src = "generated/out/vanilla.sv:1635.9-1635.30" */ instr_lhu;
  assign _06870_ = mem_do_rdata || /* src = "generated/out/vanilla.sv:1668.38-1668.66" */ mem_do_wdata;
  assign _06872_ = _06823_ || /* src = "generated/out/vanilla.sv:1687.7-1687.26" */ mem_done;
  assign _06874_ = launch_next_insn || /* src = "generated/out/vanilla.sv:1715.29-1715.53" */ trap;
  assign mem_xfer = _06627_ || /* src = "generated/out/vanilla.sv:294.20-294.97" */ _06639_;
  assign _06878_ = _06876_ || /* src = "generated/out/vanilla.sv:296.60-296.106" */ mem_do_wdata;
  assign _06880_ = _06643_ || /* src = "generated/out/vanilla.sv:296.30-296.140" */ _06645_;
  assign _06882_ = _06835_ || /* src = "generated/out/vanilla.sv:296.147-296.206" */ _06649_;
  assign _06886_ = _06655_ || /* src = "generated/out/vanilla.sv:298.34-298.289" */ _06659_;
  assign _06889_ = _06823_ || /* src = "generated/out/vanilla.sv:464.8-464.28" */ mem_ready;
  assign _06891_ = mem_la_read || /* src = "generated/out/vanilla.sv:470.8-470.35" */ mem_la_write;
  assign _06884_ = _06633_ || /* src = "generated/out/vanilla.sv:478.10-478.59" */ mem_do_rdata;
  assign _06633_ = mem_do_prefetch || /* src = "generated/out/vanilla.sv:480.20-480.51" */ mem_do_rinst;
  assign _06893_ = _06819_ || /* src = "generated/out/vanilla.sv:506.13-506.50" */ mem_la_secondword;
  assign _06876_ = mem_do_rinst || /* src = "generated/out/vanilla.sv:512.22-512.50" */ mem_do_rdata;
  assign _06888_ = _06823_ || /* src = "generated/out/vanilla.sv:743.7-743.22" */ trap;
  assign _06895_ = mem_rdata_latched[12] || /* src = "generated/out/vanilla.sv:859.13-859.60" */ mem_rdata_latched[6:2];
  assign _06781_ = _06775_ || /* src = "generated/out/vanilla.sv:984.22-984.244" */ _06779_;
  assign _06791_ = _06785_ || /* src = "generated/out/vanilla.sv:985.24-985.246" */ _06789_;
  assign _06897_ = _06803_ || /* src = "generated/out/vanilla.sv:988.26-988.162" */ _06593_;
  assign _06899_ = instr_jalr || /* src = "generated/out/vanilla.sv:995.45-995.260" */ _06815_;
  assign alu_lts = $signed(pcpi_rs1) < /* src = "generated/out/vanilla.sv:1112.15-1112.50" */ $signed(pcpi_rs2);
  assign alu_ltu = pcpi_rs1 < /* src = "generated/out/vanilla.sv:1113.15-1113.32" */ pcpi_rs2;
  assign _05887_ = _00080_[4] ? _06903_ : _06901_;
  assign _06901_ = _00080_[3] ? _06907_ : _06905_;
  assign _06903_ = _00080_[3] ? _06911_ : _06909_;
  assign _06905_ = _00080_[2] ? _06915_ : _06913_;
  assign _06907_ = _00080_[2] ? _06919_ : _06917_;
  assign _06909_ = _00080_[2] ? _06923_ : _06921_;
  assign _06911_ = _00080_[2] ? _06927_ : _06925_;
  assign _06913_ = _00080_[1] ? _06931_ : _06929_;
  assign _06915_ = _00080_[1] ? _06935_ : _06933_;
  assign _06917_ = _00080_[1] ? _06939_ : _06937_;
  assign _06919_ = _00080_[1] ? _06943_ : _06941_;
  assign _06921_ = _00080_[1] ? _06947_ : _06945_;
  assign _06923_ = _00080_[1] ? _06951_ : _06949_;
  assign _06925_ = _00080_[1] ? _06955_ : _06953_;
  assign _06927_ = _00080_[1] ? _06959_ : _06957_;
  assign _06929_ = _00080_[0] ? \cpuregs[1]  : \cpuregs[0] ;
  assign _06949_ = _00080_[0] ? \cpuregs[21]  : \cpuregs[20] ;
  assign _06951_ = _00080_[0] ? \cpuregs[23]  : \cpuregs[22] ;
  assign _06953_ = _00080_[0] ? \cpuregs[25]  : \cpuregs[24] ;
  assign _06955_ = _00080_[0] ? \cpuregs[27]  : \cpuregs[26] ;
  assign _06957_ = _00080_[0] ? \cpuregs[29]  : \cpuregs[28] ;
  assign _06959_ = _00080_[0] ? \cpuregs[31]  : \cpuregs[30] ;
  assign _06931_ = _00080_[0] ? \cpuregs[3]  : \cpuregs[2] ;
  assign _06933_ = _00080_[0] ? \cpuregs[5]  : \cpuregs[4] ;
  assign _06935_ = _00080_[0] ? \cpuregs[7]  : \cpuregs[6] ;
  assign _06937_ = _00080_[0] ? \cpuregs[9]  : \cpuregs[8] ;
  assign _06939_ = _00080_[0] ? \cpuregs[11]  : \cpuregs[10] ;
  assign _06941_ = _00080_[0] ? \cpuregs[13]  : \cpuregs[12] ;
  assign _06943_ = _00080_[0] ? \cpuregs[15]  : \cpuregs[14] ;
  assign _06945_ = _00080_[0] ? \cpuregs[17]  : \cpuregs[16] ;
  assign _06947_ = _00080_[0] ? \cpuregs[19]  : \cpuregs[18] ;
  assign _05886_ = _00082_[4] ? _06963_ : _06961_;
  assign _06961_ = _00082_[3] ? _06967_ : _06965_;
  assign _06963_ = _00082_[3] ? _06971_ : _06969_;
  assign _06965_ = _00082_[2] ? _06975_ : _06973_;
  assign _06967_ = _00082_[2] ? _06979_ : _06977_;
  assign _06969_ = _00082_[2] ? _06983_ : _06981_;
  assign _06971_ = _00082_[2] ? _06987_ : _06985_;
  assign _06973_ = _00082_[1] ? _06991_ : _06989_;
  assign _06975_ = _00082_[1] ? _06995_ : _06993_;
  assign _06977_ = _00082_[1] ? _06999_ : _06997_;
  assign _06979_ = _00082_[1] ? _07003_ : _07001_;
  assign _06981_ = _00082_[1] ? _07007_ : _07005_;
  assign _06983_ = _00082_[1] ? _07011_ : _07009_;
  assign _06985_ = _00082_[1] ? _07015_ : _07013_;
  assign _06987_ = _00082_[1] ? _07019_ : _07017_;
  assign _06989_ = _00082_[0] ? \cpuregs[1]  : \cpuregs[0] ;
  assign _07009_ = _00082_[0] ? \cpuregs[21]  : \cpuregs[20] ;
  assign _07011_ = _00082_[0] ? \cpuregs[23]  : \cpuregs[22] ;
  assign _07013_ = _00082_[0] ? \cpuregs[25]  : \cpuregs[24] ;
  assign _07015_ = _00082_[0] ? \cpuregs[27]  : \cpuregs[26] ;
  assign _07017_ = _00082_[0] ? \cpuregs[29]  : \cpuregs[28] ;
  assign _07019_ = _00082_[0] ? \cpuregs[31]  : \cpuregs[30] ;
  assign _06991_ = _00082_[0] ? \cpuregs[3]  : \cpuregs[2] ;
  assign _06993_ = _00082_[0] ? \cpuregs[5]  : \cpuregs[4] ;
  assign _06995_ = _00082_[0] ? \cpuregs[7]  : \cpuregs[6] ;
  assign _06997_ = _00082_[0] ? \cpuregs[9]  : \cpuregs[8] ;
  assign _06999_ = _00082_[0] ? \cpuregs[11]  : \cpuregs[10] ;
  assign _07001_ = _00082_[0] ? \cpuregs[13]  : \cpuregs[12] ;
  assign _07003_ = _00082_[0] ? \cpuregs[15]  : \cpuregs[14] ;
  assign _07005_ = _00082_[0] ? \cpuregs[17]  : \cpuregs[16] ;
  assign _07007_ = _00082_[0] ? \cpuregs[19]  : \cpuregs[18] ;
  assign _07021_ = _03366_ & _00004_[31];
  assign _07023_ = _03398_ & _00004_[31];
  assign _07025_ = _03400_ & _00004_[31];
  assign _07027_ = _03404_ & _00004_[31];
  assign _07029_ = _03406_ & _00004_[31];
  assign _07031_ = _03408_ & _00004_[31];
  assign _07033_ = _03410_ & _00004_[31];
  assign _07035_ = _03416_ & _00004_[31];
  assign _07037_ = _03418_ & _00004_[31];
  assign _07039_ = _03420_ & _00004_[31];
  assign _07041_ = _03422_ & _00004_[31];
  assign _07043_ = _03370_ & _00004_[31];
  assign _07045_ = _03426_ & _00004_[31];
  assign _07047_ = _03428_ & _00004_[31];
  assign _07049_ = _03430_ & _00004_[31];
  assign _07051_ = _03432_ & _00004_[31];
  assign _07053_ = _03438_ & _00004_[31];
  assign _07055_ = _03440_ & _00004_[31];
  assign _07057_ = _03442_ & _00004_[31];
  assign _07059_ = _03444_ & _00004_[31];
  assign _07061_ = _03448_ & _00004_[31];
  assign _07063_ = _03450_ & _00004_[31];
  assign _07065_ = _03374_ & _00004_[31];
  assign _07067_ = _03452_ & _00004_[31];
  assign _07069_ = _03454_ & _00004_[31];
  assign _07071_ = _03378_ & _00004_[31];
  assign _07073_ = _03382_ & _00004_[31];
  assign _07075_ = _03384_ & _00004_[31];
  assign _07077_ = _03386_ & _00004_[31];
  assign _07079_ = _03388_ & _00004_[31];
  assign _07081_ = _03394_ & _00004_[31];
  assign _07083_ = _03396_ & _00004_[31];
  assign _07087_ = | /* src = "generated/out/vanilla.sv:1669.32-1669.49" */ pcpi_rs1[1:0];
  assign _06677_ = mem_rdata_latched[1:0] != /* src = "generated/out/vanilla.sv:817.27-817.58" */ 2'h3;
  assign _07090_ = | /* src = "generated/out/vanilla.sv:928.47-928.75" */ mem_rdata_latched[11:7];
  assign _07089_ = | /* src = "generated/out/vanilla.sv:933.46-933.73" */ mem_rdata_latched[6:2];
  assign _07092_ = | /* src = "generated/out/vanilla.sv:987.105-987.130" */ mem_rdata_q[13:12];
  assign _07094_ = pcpi_rs1 | /* src = "generated/out/vanilla.sv:1136.37-1136.54" */ pcpi_rs2;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_valid */
  always_ff @(posedge clk)
    rvfi_valid <= _00030_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_halt */
  always_ff @(posedge clk)
    rvfi_halt <= trap;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_pc_rdata */
  always_ff @(posedge clk)
    rvfi_pc_rdata <= rvfi_pc_wdata;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME reg_out */
  always_ff @(posedge clk)
    reg_out <= _00026_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME reg_sh */
  always_ff @(posedge clk)
    reg_sh <= _00028_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoder_trigger */
  always_ff @(posedge clk)
    decoder_trigger <= _00012_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoder_trigger_q */
  always_ff @(posedge clk)
    decoder_trigger_q <= decoder_trigger;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME decoder_pseudo_trigger_q */
  always_ff @(posedge clk)
    decoder_pseudo_trigger_q <= decoder_pseudo_trigger;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_rs1val */
  always_ff @(posedge clk)
    dbg_rs1val <= _00006_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_rs2val */
  always_ff @(posedge clk)
    dbg_rs2val <= _00009_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_rs1val_valid */
  always_ff @(posedge clk)
    dbg_rs1val_valid <= _00008_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_rs2val_valid */
  always_ff @(posedge clk)
    dbg_rs2val_valid <= _00011_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME alu_out_q */
  always_ff @(posedge clk)
    alu_out_q <= alu_out;
  /* src = "generated/out/vanilla.sv:1143.2-1143.83" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME clear_prefetched_high_word_q */
  always_ff @(posedge clk)
    clear_prefetched_high_word_q <= clear_prefetched_high_word;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_lui_auipc_jal */
  always_ff @(posedge clk)
    is_lui_auipc_jal <= _00014_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_slti_blt_slt */
  always_ff @(posedge clk)
    is_slti_blt_slt <= _00016_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME is_sltiu_bltu_sltu */
  always_ff @(posedge clk)
    is_sltiu_bltu_sltu <= _00018_;
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME q_insn_rs1 */
  always_ff @(posedge clk)
    q_insn_rs1 <= dbg_insn_rs1;
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME q_insn_rs2 */
  always_ff @(posedge clk)
    q_insn_rs2 <= dbg_insn_rs2;
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_next */
  always_ff @(posedge clk)
    dbg_next <= launch_next_insn;
  assign _00051_ = _06509_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1793.8-1793.35|generated/out/vanilla.sv:1793.4-1796.7" */ 64'h00000000ffffffff : 64'h0000000000000000;
  assign rvfi_csr_minstret_rdata = _06631_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1792.7-1792.85|generated/out/vanilla.sv:1792.3-1809.6" */ _00070_ : 64'h0000000000000000;
  assign rvfi_csr_minstret_rmask = _06631_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1792.7-1792.85|generated/out/vanilla.sv:1792.3-1809.6" */ _00072_ : 64'h0000000000000000;
  assign rvfi_csr_mcycle_rdata = _06631_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1792.7-1792.85|generated/out/vanilla.sv:1792.3-1809.6" */ _00066_ : 64'h0000000000000000;
  assign rvfi_csr_mcycle_rmask = _06631_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1792.7-1792.85|generated/out/vanilla.sv:1792.3-1809.6" */ _00068_ : 64'h0000000000000000;
  assign _07096_ = { dbg_insn_opcode[31:25], dbg_insn_opcode[19:15], dbg_insn_opcode[11:0] } == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1752.3-1765.10" */ 24'h04000b;
  assign _07097_ = { dbg_insn_opcode[31:25], dbg_insn_opcode[19:17], dbg_insn_opcode[6:0] } == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1752.3-1765.10" */ 17'h0000b;
  assign _07098_ = _06627_ ? /* src = "generated/out/vanilla.sv:1774.13-1774.43|generated/out/vanilla.sv:1774.9-1780.7" */ mem_wdata : 32'hxxxxxxxx;
  assign _07100_ = _06627_ ? /* src = "generated/out/vanilla.sv:1774.13-1774.43|generated/out/vanilla.sv:1774.9-1780.7" */ mem_rdata : 32'hxxxxxxxx;
  assign _07102_ = _06627_ ? /* src = "generated/out/vanilla.sv:1774.13-1774.43|generated/out/vanilla.sv:1774.9-1780.7" */ mem_wstrb : 4'hx;
  assign _07104_ = _06627_ ? /* src = "generated/out/vanilla.sv:1774.13-1774.43|generated/out/vanilla.sv:1774.9-1780.7" */ _07601_[3:0] : 4'hx;
  assign _07106_ = _06627_ ? /* src = "generated/out/vanilla.sv:1774.13-1774.43|generated/out/vanilla.sv:1774.9-1780.7" */ mem_addr : 32'hxxxxxxxx;
  assign _07108_ = rvfi_valid ? /* src = "generated/out/vanilla.sv:1748.12-1748.22|generated/out/vanilla.sv:1748.8-1751.6" */ 32'd0 : 32'hxxxxxxxx;
  assign _07109_ = cpuregs_write ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1744.12-1744.39|generated/out/vanilla.sv:1744.8-1751.6" */ _07599_ : _07108_;
  assign _07112_ = rvfi_valid ? /* src = "generated/out/vanilla.sv:1748.12-1748.22|generated/out/vanilla.sv:1748.8-1751.6" */ 5'h00 : 5'hxx;
  assign _07113_ = cpuregs_write ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1744.12-1744.39|generated/out/vanilla.sv:1744.8-1751.6" */ latched_rd : _07112_;
  assign _07111_ = { dbg_insn_opcode[31:25], dbg_insn_opcode[11:9], dbg_insn_opcode[6:0] } == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1752.3-1765.10" */ 17'h0040b;
  assign _00074_ = _06865_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1630.10-1630.38|generated/out/vanilla.sv:1630.6-1659.9" */ _00077_ : 1'h0;
  assign _00076_ = _06865_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1606.10-1606.38|generated/out/vanilla.sv:1606.6-1626.9" */ _00078_ : 1'h0;
  assign _00075_ = is_beq_bne_blt_bge_bltu_bgeu ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1559.15-1559.43|generated/out/vanilla.sv:1559.11-1575.9" */ _00079_ : 1'h0;
  assign _00078_ = mem_do_wdata ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1607.11-1607.24|generated/out/vanilla.sv:1607.7-1620.10" */ 1'h0 : 1'h1;
  assign _00077_ = mem_do_rdata ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1631.11-1631.24|generated/out/vanilla.sv:1631.7-1647.10" */ 1'h0 : 1'h1;
  assign _00079_ = alu_out_0 ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1565.11-1565.56|generated/out/vanilla.sv:1565.7-1568.10" */ 1'h1 : 1'h0;
  assign _07115_ = latched_branch ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1279.6-1292.13" */ _07594_ : reg_next_pc;
  assign _07117_ = _06485_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ _07115_ : 32'hxxxxxxxx;
  assign _00060_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _07117_ : 32'hxxxxxxxx;
  assign _00034_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _00059_ : 1'h0;
  assign _00032_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _00057_ : 1'h0;
  assign _00033_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _00058_ : 1'h0;
  assign _07119_ = _06615_ ? /* src = "generated/out/vanilla.sv:1621.11-1621.39|generated/out/vanilla.sv:1621.7-1625.10" */ 1'h1 : 1'h0;
  assign _07120_ = _06615_ ? /* src = "generated/out/vanilla.sv:1621.11-1621.39|generated/out/vanilla.sv:1621.7-1625.10" */ 1'h1 : _05738_;
  assign _07122_ = _06865_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1606.10-1606.38|generated/out/vanilla.sv:1606.6-1626.9" */ _07120_ : _05738_;
  assign _07124_ = alu_out_0 ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1565.11-1565.56|generated/out/vanilla.sv:1565.7-1568.10" */ 1'h0 : _05738_;
  assign _07126_ = is_beq_bne_blt_bge_bltu_bgeu ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1559.15-1559.43|generated/out/vanilla.sv:1559.11-1575.9" */ _07124_ : _05738_;
  assign _00012_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _06108_ : _05738_;
  assign _07128_ = _06615_ ? /* src = "generated/out/vanilla.sv:1648.11-1648.39|generated/out/vanilla.sv:1648.7-1658.10" */ _06112_ : 32'hxxxxxxxx;
  assign _07130_ = _06865_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1630.10-1630.38|generated/out/vanilla.sv:1630.6-1659.9" */ _07128_ : 32'hxxxxxxxx;
  assign _07132_ = _06499_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1579.10-1579.21|generated/out/vanilla.sv:1579.6-1601.9" */ pcpi_rs1 : 32'hxxxxxxxx;
  assign _07136_ = instr_trap ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1517.6-1551.13" */ _07134_ : 32'hxxxxxxxx;
  assign _07134_ = pcpi_int_ready ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1367.14-1367.28|generated/out/vanilla.sv:1367.10-1382.13" */ pcpi_int_rd : 32'hxxxxxxxx;
  assign _00026_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _06120_ : 32'hxxxxxxxx;
  assign _07138_ = _06597_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1584.15-1584.47|generated/out/vanilla.sv:1584.11-1601.9" */ _07587_[4:0] : _07589_[4:0];
  assign _07140_ = _06499_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1579.10-1579.21|generated/out/vanilla.sv:1579.6-1601.9" */ 5'hxx : _07138_;
  assign _00028_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _06132_ : 5'hxx;
  assign _07142_ = _06483_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 1'h1 : 1'h0;
  assign _06483_ = cpu_state == /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 8'h80;
  assign _07144_ = is_beq_bne_blt_bge_bltu_bgeu ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1559.15-1559.43|generated/out/vanilla.sv:1559.11-1575.9" */ 5'h00 : 5'hxx;
  assign _07145_ = mem_do_rdata ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1631.11-1631.24|generated/out/vanilla.sv:1631.7-1647.10" */ 1'hx : instr_lb;
  assign _05526_ = _06865_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1630.10-1630.38|generated/out/vanilla.sv:1630.6-1659.9" */ _07145_ : 1'hx;
  assign _07148_ = mem_do_rdata ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1631.11-1631.24|generated/out/vanilla.sv:1631.7-1647.10" */ 1'hx : instr_lh;
  assign _05527_ = _06865_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1630.10-1630.38|generated/out/vanilla.sv:1630.6-1659.9" */ _07148_ : 1'hx;
  assign _07151_ = is_beq_bne_blt_bge_bltu_bgeu ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1559.15-1559.43|generated/out/vanilla.sv:1559.11-1575.9" */ alu_out_0 : instr_jalr;
  assign _05742_ = instr_jal ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1339.11-1339.20|generated/out/vanilla.sv:1339.7-1348.10" */ 1'h1 : 1'h0;
  assign _07153_ = decoder_trigger ? /* src = "generated/out/vanilla.sv:1329.15-1329.30|generated/out/vanilla.sv:1329.11-1349.9" */ _05742_ : 1'h0;
  assign _05529_ = is_beq_bne_blt_bge_bltu_bgeu ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1559.15-1559.43|generated/out/vanilla.sv:1559.11-1575.9" */ 1'hx : 1'h1;
  assign _07155_ = is_beq_bne_blt_bge_bltu_bgeu ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1559.15-1559.43|generated/out/vanilla.sv:1559.11-1575.9" */ alu_out_0 : 1'h1;
  assign _07159_ = instr_trap ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1517.6-1551.13" */ _07157_ : 1'hx;
  assign _07157_ = pcpi_int_ready ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1367.14-1367.28|generated/out/vanilla.sv:1367.10-1382.13" */ pcpi_int_wr : latched_store;
  assign _07161_ = _06615_ ? /* src = "generated/out/vanilla.sv:1621.11-1621.39|generated/out/vanilla.sv:1621.7-1625.10" */ 8'h40 : cpu_state;
  assign _07163_ = _06865_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1606.10-1606.38|generated/out/vanilla.sv:1606.6-1626.9" */ _07161_ : cpu_state;
  assign _07165_ = _06499_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1579.10-1579.21|generated/out/vanilla.sv:1579.6-1601.9" */ 8'h40 : cpu_state;
  assign { _05745_[7], _07167_[6], _05745_[5:0] } = mem_done ? /* src = "generated/out/vanilla.sv:1563.11-1563.19|generated/out/vanilla.sv:1563.7-1564.37" */ 8'h40 : cpu_state;
  assign _07169_ = is_beq_bne_blt_bge_bltu_bgeu ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1559.15-1559.43|generated/out/vanilla.sv:1559.11-1575.9" */ { _05745_[7], _07167_[6], _05745_[5:0] } : 8'h40;
  assign { _05746_[7], _07171_[6], _05746_[5:0] } = _06611_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1374.19-1374.72|generated/out/vanilla.sv:1374.15-1382.13" */ 8'h80 : cpu_state;
  assign { _05539_[7:4], _07173_[3], _05539_[2:0] } = pcpi_int_ready ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1367.14-1367.28|generated/out/vanilla.sv:1367.10-1382.13" */ 8'h40 : { _05746_[7], _07171_[6], _05746_[5:0] };
  assign _07175_ = instr_jal ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1339.11-1339.20|generated/out/vanilla.sv:1339.7-1348.10" */ cpu_state : 8'h20;
  assign _07177_ = decoder_trigger ? /* src = "generated/out/vanilla.sv:1329.15-1329.30|generated/out/vanilla.sv:1329.11-1349.9" */ _07175_ : cpu_state;
  assign { _07179_[7], _05749_[6:0] } = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ { _05748_[7], _06167_[6], _05748_[5:0] } : 8'h40;
  assign { _07181_[7], _05750_[6:0] } = _06619_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1669.8-1669.50|generated/out/vanilla.sv:1669.4-1673.34" */ 8'h80 : { _07179_[7], _05749_[6:0] };
  assign _07183_ = _06621_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1674.8-1674.48|generated/out/vanilla.sv:1674.4-1678.34" */ 8'h80 : { _07181_[7], _05750_[6:0] };
  assign _07185_ = _06617_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1668.7-1668.67|generated/out/vanilla.sv:1668.3-1679.6" */ _07183_ : { _07179_[7], _05749_[6:0] };
  assign _07187_ = launch_next_insn ? /* src = "generated/out/vanilla.sv:1207.7-1207.23|generated/out/vanilla.sv:1207.3-1212.6" */ 1'h0 : dbg_rs2val_valid;
  assign _07188_ = _00855_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1355.6-1509.13" */ _07187_ : 1'h1;
  assign _00011_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _06187_ : _07187_;
  assign _07189_ = launch_next_insn ? /* src = "generated/out/vanilla.sv:1207.7-1207.23|generated/out/vanilla.sv:1207.3-1212.6" */ 1'h0 : dbg_rs1val_valid;
  assign _07190_ = _00859_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1355.6-1509.13" */ _07189_ : 1'h1;
  assign _07191_ = _06487_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ _07190_ : _07189_;
  assign _00008_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _07191_ : _07189_;
  assign _07192_ = launch_next_insn ? /* src = "generated/out/vanilla.sv:1207.7-1207.23|generated/out/vanilla.sv:1207.3-1212.6" */ 32'hxxxxxxxx : dbg_rs2val;
  assign _07194_ = _00855_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1355.6-1509.13" */ _07192_ : cpuregs_rs2;
  assign _00009_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _06190_ : _07192_;
  assign _07196_ = launch_next_insn ? /* src = "generated/out/vanilla.sv:1207.7-1207.23|generated/out/vanilla.sv:1207.3-1212.6" */ 32'hxxxxxxxx : dbg_rs1val;
  assign _07198_ = _00859_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1355.6-1509.13" */ _07196_ : cpuregs_rs1;
  assign _07200_ = _06487_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ _07198_ : _07196_;
  assign _00006_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _07200_ : _07196_;
  assign _07202_ = _06499_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1579.10-1579.21|generated/out/vanilla.sv:1579.6-1601.9" */ mem_do_prefetch : 1'hx;
  assign _06491_ = cpu_state == /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 8'h08;
  assign _07204_ = pcpi_int_ready ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1367.14-1367.28|generated/out/vanilla.sv:1367.10-1382.13" */ 1'h1 : mem_do_rinst;
  assign _07206_ = decoder_trigger ? /* src = "generated/out/vanilla.sv:1329.15-1329.30|generated/out/vanilla.sv:1329.11-1349.9" */ _05742_ : _06609_;
  assign _05756_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _06196_ : 1'hx;
  assign _07209_ = _06872_ ? /* src = "generated/out/vanilla.sv:1687.7-1687.26|generated/out/vanilla.sv:1687.3-1692.6" */ 1'h0 : _05756_;
  assign _07211_ = mem_do_rdata ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1631.11-1631.24|generated/out/vanilla.sv:1631.7-1647.10" */ 2'hx : _06216_;
  assign _07213_ = _06865_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1630.10-1630.38|generated/out/vanilla.sv:1630.6-1659.9" */ _07211_ : 2'hx;
  assign _07215_ = mem_do_wdata ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1607.11-1607.24|generated/out/vanilla.sv:1607.7-1620.10" */ 2'hx : _06222_;
  assign _05556_ = _06865_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1606.10-1606.38|generated/out/vanilla.sv:1606.6-1626.9" */ _07215_ : 2'hx;
  assign _07218_ = mem_do_rdata ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1631.11-1631.24|generated/out/vanilla.sv:1631.7-1647.10" */ 32'hxxxxxxxx : _00098_;
  assign _07220_ = _06865_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1630.10-1630.38|generated/out/vanilla.sv:1630.6-1659.9" */ _07218_ : 32'hxxxxxxxx;
  assign _06497_ = cpu_state == /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 8'h01;
  assign _07222_ = mem_do_wdata ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1607.11-1607.24|generated/out/vanilla.sv:1607.7-1620.10" */ 32'hxxxxxxxx : _00098_;
  assign _07224_ = _06865_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1606.10-1606.38|generated/out/vanilla.sv:1606.6-1626.9" */ _07222_ : 32'hxxxxxxxx;
  assign _06495_ = cpu_state == /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 8'h02;
  assign _07226_ = _06597_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1584.15-1584.47|generated/out/vanilla.sv:1584.11-1601.9" */ _06242_ : _06238_;
  assign _07228_ = _06499_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1579.10-1579.21|generated/out/vanilla.sv:1579.6-1601.9" */ 32'hxxxxxxxx : _07226_;
  assign _06493_ = cpu_state == /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 8'h04;
  assign _07230_ = instr_jal ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1339.11-1339.20|generated/out/vanilla.sv:1339.7-1348.10" */ _00094_ : _00090_;
  assign _07232_ = decoder_trigger ? /* src = "generated/out/vanilla.sv:1329.15-1329.30|generated/out/vanilla.sv:1329.11-1349.9" */ _07230_ : _00060_;
  assign _06485_ = cpu_state == /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 8'h40;
  assign _07238_ = _00857_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ _07236_ : 1'hx;
  assign _06489_ = cpu_state == /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 8'h10;
  assign _05760_ = _06611_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1374.19-1374.72|generated/out/vanilla.sv:1374.15-1382.13" */ 1'h0 : 1'h1;
  assign _07234_ = pcpi_int_ready ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1367.14-1367.28|generated/out/vanilla.sv:1367.10-1382.13" */ 1'h0 : _05760_;
  assign _07236_ = instr_trap ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1355.6-1509.13" */ _07234_ : 1'hx;
  assign _06487_ = cpu_state == /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 8'h20;
  assign _00004_[31] = _06605_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1181.7-1181.46|generated/out/vanilla.sv:1181.3-1182.42" */ 1'h1 : 1'h0;
  assign _00002_ = _06605_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1181.7-1181.46|generated/out/vanilla.sv:1181.3-1182.42" */ cpuregs_wrdata : 32'hxxxxxxxx;
  assign _00000_ = _06605_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1181.7-1181.46|generated/out/vanilla.sv:1181.3-1182.42" */ latched_rd : 5'hxx;
  assign _00039_ = _01094_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1161.4-1178.11" */ 1'h1 : 1'h0;
  assign cpuregs_wrdata = _06485_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1159.7-1159.35|generated/out/vanilla.sv:1159.3-1178.11" */ _00037_ : 32'hxxxxxxxx;
  assign cpuregs_write = _06485_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1159.7-1159.35|generated/out/vanilla.sv:1159.3-1178.11" */ _00039_ : 1'h0;
  assign clear_prefetched_high_word = _06863_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1148.7-1148.47|generated/out/vanilla.sv:1148.3-1149.48" */ 1'h1 : _00035_;
  assign _00035_ = prefetched_high_word ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1146.7-1146.28|generated/out/vanilla.sv:1146.3-1147.35" */ clear_prefetched_high_word_q : 1'h0;
  assign _05761_ = _06683_ ? /* src = "generated/out/vanilla.sv:917.13-917.110|generated/out/vanilla.sv:917.9-921.12" */ mem_rdata_latched[11] : 1'h0;
  assign _07241_ = _06667_ ? /* src = "generated/out/vanilla.sv:922.13-922.74|generated/out/vanilla.sv:922.9-927.12" */ 1'h0 : _05761_;
  assign _07243_ = _06671_ ? /* src = "generated/out/vanilla.sv:928.13-928.110|generated/out/vanilla.sv:928.9-932.12" */ mem_rdata_latched[11] : _07241_;
  assign _07245_ = _06673_ ? /* src = "generated/out/vanilla.sv:933.13-933.74|generated/out/vanilla.sv:933.9-938.12" */ mem_rdata_latched[11] : _07243_;
  assign _05579_ = mem_rdata_latched[12] ? /* src = "generated/out/vanilla.sv:904.13-904.35|generated/out/vanilla.sv:904.9-909.12" */ 1'h0 : mem_rdata_latched[11];
  assign _07256_ = _06679_ ? /* src = "generated/out/vanilla.sv:871.13-871.61|generated/out/vanilla.sv:871.9-876.12" */ _00106_[4] : 1'h0;
  assign _07258_ = _06521_ ? /* src = "generated/out/vanilla.sv:877.13-877.46|generated/out/vanilla.sv:877.9-881.12" */ _00106_[4] : _07256_;
  assign _07260_ = _06523_ ? /* src = "generated/out/vanilla.sv:882.13-882.47|generated/out/vanilla.sv:882.9-887.12" */ _00106_[4] : _07258_;
  assign _05766_ = _06515_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:860.14-860.42|generated/out/vanilla.sv:860.10-869.13" */ mem_rdata_latched[11] : 1'h0;
  assign _07263_ = _06895_ ? /* src = "generated/out/vanilla.sv:859.13-859.60|generated/out/vanilla.sv:859.9-869.13" */ _05766_ : 1'h0;
  assign _05582_ = _01076_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ _00106_[4] : 1'h0;
  assign _07274_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _06270_ : mem_rdata_latched[19];
  assign _07276_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ mem_rdata_latched[8] : mem_rdata_latched[30];
  assign _07278_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ mem_rdata_latched[6] : mem_rdata_latched[27];
  assign _07280_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ mem_rdata_latched[7] : mem_rdata_latched[26];
  assign _07282_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ mem_rdata_latched[5:3] : mem_rdata_latched[23:21];
  assign _07284_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ mem_rdata_latched[2] : mem_rdata_latched[25];
  assign _07286_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ mem_rdata_latched[10:9] : mem_rdata_latched[29:28];
  assign _07288_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] } : { mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31] };
  assign _07290_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ mem_rdata_latched[11] : mem_rdata_latched[24];
  assign _07292_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ mem_rdata_latched[12] : mem_rdata_latched[20];
  assign _05777_ = _06683_ ? /* src = "generated/out/vanilla.sv:917.13-917.110|generated/out/vanilla.sv:917.9-921.12" */ mem_rdata_latched[10:7] : 4'h0;
  assign _07295_ = _06667_ ? /* src = "generated/out/vanilla.sv:922.13-922.74|generated/out/vanilla.sv:922.9-927.12" */ 4'h0 : _05777_;
  assign _07297_ = _06671_ ? /* src = "generated/out/vanilla.sv:928.13-928.110|generated/out/vanilla.sv:928.9-932.12" */ mem_rdata_latched[10:7] : _07295_;
  assign { _05587_[3:2], _07299_[1], _05587_[0] } = _06673_ ? /* src = "generated/out/vanilla.sv:933.13-933.74|generated/out/vanilla.sv:933.9-938.12" */ mem_rdata_latched[10:7] : _07297_;
  assign _07301_ = _07090_ ? /* src = "generated/out/vanilla.sv:911.13-911.36|generated/out/vanilla.sv:911.9-915.12" */ 4'h2 : 4'h0;
  assign _05588_ = mem_rdata_latched[12] ? /* src = "generated/out/vanilla.sv:904.13-904.35|generated/out/vanilla.sv:904.9-909.12" */ 4'h0 : mem_rdata_latched[10:7];
  assign _07303_ = _06679_ ? /* src = "generated/out/vanilla.sv:871.13-871.61|generated/out/vanilla.sv:871.9-876.12" */ _00106_[3:0] : 4'h0;
  assign _07305_ = _06521_ ? /* src = "generated/out/vanilla.sv:877.13-877.46|generated/out/vanilla.sv:877.9-881.12" */ _00106_[3:0] : _07303_;
  assign _07307_ = _06523_ ? /* src = "generated/out/vanilla.sv:882.13-882.47|generated/out/vanilla.sv:882.9-887.12" */ _00106_[3:0] : _07305_;
  assign _05782_ = _06515_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:860.14-860.42|generated/out/vanilla.sv:860.10-869.13" */ mem_rdata_latched[10:7] : 4'h0;
  assign _07310_ = _06895_ ? /* src = "generated/out/vanilla.sv:859.13-859.60|generated/out/vanilla.sv:859.9-869.13" */ _05782_ : 4'h0;
  assign _07312_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _06292_ : mem_rdata_latched[18:15];
  assign _07314_ = _06667_ ? /* src = "generated/out/vanilla.sv:922.13-922.74|generated/out/vanilla.sv:922.9-927.12" */ 1'h1 : _06557_;
  assign _07316_ = _06673_ ? /* src = "generated/out/vanilla.sv:933.13-933.74|generated/out/vanilla.sv:933.9-938.12" */ 1'h1 : _07314_;
  assign _07318_ = _07247_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:902.7-945.14" */ _07316_ : _06557_;
  assign _07320_ = _06523_ ? /* src = "generated/out/vanilla.sv:882.13-882.47|generated/out/vanilla.sv:882.9-887.12" */ 1'h1 : _06557_;
  assign _07322_ = _07247_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:843.7-900.14" */ _07320_ : _06557_;
  assign _07324_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _06307_ : _06557_;
  assign _07326_ = mem_rdata_latched[12] ? /* src = "generated/out/vanilla.sv:904.13-904.35|generated/out/vanilla.sv:904.9-909.12" */ _06555_ : 1'h1;
  assign _07328_ = _07250_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:902.7-945.14" */ _07326_ : _06555_;
  assign _07330_ = _06679_ ? /* src = "generated/out/vanilla.sv:871.13-871.61|generated/out/vanilla.sv:871.9-876.12" */ 1'h1 : _06555_;
  assign _07332_ = _06521_ ? /* src = "generated/out/vanilla.sv:877.13-877.46|generated/out/vanilla.sv:877.9-881.12" */ 1'h1 : _07330_;
  assign _07334_ = _06515_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:860.14-860.42|generated/out/vanilla.sv:860.10-869.13" */ 1'h1 : _06555_;
  assign _07336_ = _06895_ ? /* src = "generated/out/vanilla.sv:859.13-859.60|generated/out/vanilla.sv:859.9-869.13" */ _07334_ : _06555_;
  assign _07338_ = _07250_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ _07575_ : _06555_;
  assign _07340_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _06313_ : _06555_;
  assign _07342_ = _01078_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:843.7-900.14" */ 1'h1 : _06549_;
  assign _07344_ = _07267_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:823.5-946.12" */ _07342_ : _06549_;
  assign _07346_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _07344_ : _06549_;
  assign _07350_ = _00863_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:823.5-946.12" */ _07348_ : _06553_;
  assign _07348_ = _07254_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ 1'h1 : _06553_;
  assign _07352_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _07350_ : _06553_;
  assign _07354_ = _07090_ ? /* src = "generated/out/vanilla.sv:911.13-911.36|generated/out/vanilla.sv:911.9-915.12" */ 1'h1 : _06551_;
  assign _07356_ = _07270_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:902.7-945.14" */ _07354_ : _06551_;
  assign _07358_ = _07270_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ 1'h1 : _06551_;
  assign _07360_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _06323_ : _06551_;
  assign _07362_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ 1'h1 : 1'h0;
  assign _07365_ = _06667_ ? /* src = "generated/out/vanilla.sv:922.13-922.74|generated/out/vanilla.sv:922.9-927.12" */ mem_rdata_latched[6:2] : 5'h00;
  assign _07367_ = _06673_ ? /* src = "generated/out/vanilla.sv:933.13-933.74|generated/out/vanilla.sv:933.9-938.12" */ mem_rdata_latched[6:2] : _07365_;
  assign _05612_ = mem_rdata_latched[12] ? /* src = "generated/out/vanilla.sv:904.13-904.35|generated/out/vanilla.sv:904.9-909.12" */ 5'h00 : mem_rdata_latched[6:2];
  assign _07370_ = _06679_ ? /* src = "generated/out/vanilla.sv:871.13-871.61|generated/out/vanilla.sv:871.9-876.12" */ mem_rdata_latched[6:2] : 5'h00;
  assign _05799_ = _06523_ ? /* src = "generated/out/vanilla.sv:882.13-882.47|generated/out/vanilla.sv:882.9-887.12" */ _00104_[4:0] : _07370_;
  assign _07373_ = _07247_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:843.7-900.14" */ _05799_ : 5'h00;
  assign _05615_ = _07254_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ _00104_[4:0] : 5'h00;
  assign _07254_ = mem_rdata_latched[15:13] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ 3'h6;
  assign _07376_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _06345_ : mem_rdata_latched[24:20];
  assign _07378_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] } : mem_rdata_latched[19:12];
  assign { _05802_[4:1], _07380_[0] } = _06667_ ? /* src = "generated/out/vanilla.sv:922.13-922.74|generated/out/vanilla.sv:922.9-927.12" */ mem_rdata_latched[11:7] : 5'h00;
  assign _07382_ = _06671_ ? /* src = "generated/out/vanilla.sv:928.13-928.110|generated/out/vanilla.sv:928.9-932.12" */ 5'h01 : { _05802_[4:1], _07380_[0] };
  assign _07384_ = _06673_ ? /* src = "generated/out/vanilla.sv:933.13-933.74|generated/out/vanilla.sv:933.9-938.12" */ mem_rdata_latched[11:7] : _07382_;
  assign _07386_ = _07090_ ? /* src = "generated/out/vanilla.sv:911.13-911.36|generated/out/vanilla.sv:911.9-915.12" */ mem_rdata_latched[11:7] : 5'h00;
  assign _05618_ = mem_rdata_latched[12] ? /* src = "generated/out/vanilla.sv:904.13-904.35|generated/out/vanilla.sv:904.9-909.12" */ 5'h00 : mem_rdata_latched[11:7];
  assign _07389_ = _06679_ ? /* src = "generated/out/vanilla.sv:871.13-871.61|generated/out/vanilla.sv:871.9-876.12" */ _00106_[4:0] : 5'h00;
  assign _07391_ = _06521_ ? /* src = "generated/out/vanilla.sv:877.13-877.46|generated/out/vanilla.sv:877.9-881.12" */ _00106_[4:0] : _07389_;
  assign _07393_ = _06523_ ? /* src = "generated/out/vanilla.sv:882.13-882.47|generated/out/vanilla.sv:882.9-887.12" */ _00106_[4:0] : _07391_;
  assign _07395_ = _06895_ ? /* src = "generated/out/vanilla.sv:859.13-859.60|generated/out/vanilla.sv:859.9-869.13" */ mem_rdata_latched[11:7] : 5'h00;
  assign _05621_ = _00865_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ _00104_[4:0] : 5'h00;
  assign _07270_ = mem_rdata_latched[15:13] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ 3'h2;
  assign _07250_ = ! /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ mem_rdata_latched[15:13];
  assign _07272_ = ! /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:823.5-946.12" */ mem_rdata_latched[1:0];
  assign _07399_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _06357_ : mem_rdata_latched[11:7];
  assign _07401_ = _06683_ ? /* src = "generated/out/vanilla.sv:917.13-917.110|generated/out/vanilla.sv:917.9-921.12" */ 1'h1 : _06675_;
  assign _07403_ = _06671_ ? /* src = "generated/out/vanilla.sv:928.13-928.110|generated/out/vanilla.sv:928.9-932.12" */ 1'h1 : _07401_;
  assign _07405_ = _07247_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:902.7-945.14" */ _07403_ : _06675_;
  assign _07247_ = mem_rdata_latched[15:13] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:902.7-945.14" */ 3'h4;
  assign _07407_ = _07251_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:823.5-946.12" */ _07405_ : _06675_;
  assign _07251_ = mem_rdata_latched[1:0] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:823.5-946.12" */ 2'h2;
  assign _07409_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _07407_ : _06675_;
  assign _07411_ = _01088_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:843.7-900.14" */ 1'h1 : _06543_;
  assign _07413_ = mem_rdata_latched[15:13] == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:843.7-900.14" */ 3'h5;
  assign _07397_ = mem_rdata_latched[15:13] == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:843.7-900.14" */ 3'h1;
  assign _07415_ = _07267_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:823.5-946.12" */ _07411_ : _06543_;
  assign _07417_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _07415_ : _06543_;
  assign _07419_ = _06515_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:860.14-860.42|generated/out/vanilla.sv:860.10-869.13" */ _06539_ : 1'h1;
  assign _07421_ = _06895_ ? /* src = "generated/out/vanilla.sv:859.13-859.60|generated/out/vanilla.sv:859.9-869.13" */ _07419_ : _06539_;
  assign _07423_ = _07265_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:843.7-900.14" */ _07421_ : _06539_;
  assign _07265_ = mem_rdata_latched[15:13] == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:843.7-900.14" */ 3'h3;
  assign _07425_ = _07267_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:823.5-946.12" */ _07423_ : _06539_;
  assign _07267_ = mem_rdata_latched[1:0] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:823.5-946.12" */ 2'h1;
  assign _07427_ = _06677_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _07425_ : _06539_;
  assign _00045_ = decoder_pseudo_trigger_q ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:769.8-769.32|generated/out/vanilla.sv:769.4-787.7" */ cached_insn_rs2 : decoded_rs2;
  assign _00043_ = decoder_pseudo_trigger_q ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:769.8-769.32|generated/out/vanilla.sv:769.4-787.7" */ cached_insn_rs1 : decoded_rs1;
  assign _00041_ = decoder_pseudo_trigger_q ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:769.8-769.32|generated/out/vanilla.sv:769.4-787.7" */ cached_insn_opcode : _00062_;
  assign dbg_insn_rs2 = dbg_next ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:768.7-768.15|generated/out/vanilla.sv:768.3-787.7" */ _00045_ : q_insn_rs2;
  assign dbg_insn_rs1 = dbg_next ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:768.7-768.15|generated/out/vanilla.sv:768.3-787.7" */ _00043_ : q_insn_rs1;
  assign dbg_insn_opcode = dbg_next ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:768.7-768.15|generated/out/vanilla.sv:768.3-787.7" */ _00041_ : { rvfi_insn[31:25], 5'hxx, rvfi_insn[19:15], 3'hx, rvfi_insn[11:0] };
  assign _00062_ = _07429_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:750.8-750.30|generated/out/vanilla.sv:750.4-753.74" */ next_insn_opcode : { 16'h0000, next_insn_opcode[15:0] };
  assign _07431_ = _06893_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:506.13-506.50|generated/out/vanilla.sv:506.9-511.36" */ mem_rdata[31:16] : 16'hxxxx;
  assign _07433_ = mem_do_rdata ? /* src = "generated/out/vanilla.sv:505.12-505.43|generated/out/vanilla.sv:505.8-511.36" */ 16'hxxxx : _07431_;
  assign _07435_ = mem_la_use_prefetched_high_word ? /* src = "generated/out/vanilla.sv:499.12-499.44|generated/out/vanilla.sv:499.8-500.46" */ 16'hxxxx : mem_rdata[31:16];
  assign _07437_ = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:496.11-496.40|generated/out/vanilla.sv:496.7-513.10" */ _07435_ : _07433_;
  assign _07439_ = mem_state == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:476.4-529.11" */ 2'h1;
  assign _07441_ = _06893_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:506.13-506.50|generated/out/vanilla.sv:506.9-511.36" */ 1'h1 : 1'h0;
  assign _07442_ = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:496.11-496.40|generated/out/vanilla.sv:496.7-513.10" */ 1'h1 : 1'h0;
  assign _07443_ = mem_do_rinst ? /* src = "generated/out/vanilla.sv:526.10-526.22|generated/out/vanilla.sv:526.6-527.22" */ 2'h0 : 2'hx;
  assign _06537_ = mem_state == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:476.4-529.11" */ 2'h3;
  assign _07444_ = mem_xfer ? /* src = "generated/out/vanilla.sv:518.10-518.18|generated/out/vanilla.sv:518.6-521.9" */ 2'h0 : 2'hx;
  assign _06535_ = mem_state == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:476.4-529.11" */ 2'h2;
  assign _07445_ = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:496.11-496.40|generated/out/vanilla.sv:496.7-513.10" */ 2'hx : _07608_[1:0];
  assign _07447_ = mem_xfer ? /* src = "generated/out/vanilla.sv:495.10-495.18|generated/out/vanilla.sv:495.6-513.10" */ _07445_ : 2'hx;
  assign { _07449_[1], _05824_[0] } = _06884_ ? /* src = "generated/out/vanilla.sv:478.10-478.59|generated/out/vanilla.sv:478.6-483.9" */ 2'h1 : 2'hx;
  assign _07450_ = mem_do_wdata ? /* src = "generated/out/vanilla.sv:484.10-484.22|generated/out/vanilla.sv:484.6-488.9" */ 2'h2 : { _07449_[1], _05824_[0] };
  assign _07452_ = resetn ? /* src = "generated/out/vanilla.sv:462.8-462.15|generated/out/vanilla.sv:462.4-463.20" */ 2'hx : 2'h0;
  assign _00022_ = _06888_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:461.7-461.22|generated/out/vanilla.sv:461.3-530.6" */ _07452_ : _06371_;
  assign _05827_ = _06891_ ? /* src = "generated/out/vanilla.sv:470.8-470.35|generated/out/vanilla.sv:470.4-473.7" */ _00112_ : mem_wstrb;
  assign _07454_ = _06884_ ? /* src = "generated/out/vanilla.sv:478.10-478.59|generated/out/vanilla.sv:478.6-483.9" */ 4'h0 : _05827_;
  assign _07456_ = _06836_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:476.4-529.11" */ _07454_ : _05827_;
  assign _06836_ = ! /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:476.4-529.11" */ mem_state;
  assign _07458_ = _06884_ ? /* src = "generated/out/vanilla.sv:478.10-478.59|generated/out/vanilla.sv:478.6-483.9" */ _06633_ : 1'hx;
  assign _07460_ = mem_xfer ? /* src = "generated/out/vanilla.sv:518.10-518.18|generated/out/vanilla.sv:518.6-521.9" */ 1'h0 : 1'hx;
  assign _07461_ = mem_xfer ? /* src = "generated/out/vanilla.sv:495.10-495.18|generated/out/vanilla.sv:495.6-513.10" */ _07442_ : 1'hx;
  assign _07463_ = _06884_ ? /* src = "generated/out/vanilla.sv:478.10-478.59|generated/out/vanilla.sv:478.6-483.9" */ _06838_ : 1'hx;
  assign _07465_ = mem_do_wdata ? /* src = "generated/out/vanilla.sv:484.10-484.22|generated/out/vanilla.sv:484.6-488.9" */ 1'h1 : _07463_;
  assign _07467_ = _06889_ ? /* src = "generated/out/vanilla.sv:464.8-464.28|generated/out/vanilla.sv:464.4-465.20" */ 1'h0 : 1'hx;
  assign _00024_ = _06888_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:461.7-461.22|generated/out/vanilla.sv:461.3-530.6" */ _07467_ : _06375_;
  assign _05831_ = mem_xfer ? /* src = "generated/out/vanilla.sv:340.7-340.15|generated/out/vanilla.sv:340.3-343.6" */ mem_rdata_latched[31] : mem_rdata_q[31];
  assign _05832_ = _06665_ ? /* src = "generated/out/vanilla.sv:423.12-423.73|generated/out/vanilla.sv:423.8-426.11" */ 1'h0 : _05831_;
  assign _05833_ = _06667_ ? /* src = "generated/out/vanilla.sv:427.12-427.73|generated/out/vanilla.sv:427.8-430.11" */ 1'h0 : _05832_;
  assign _05834_ = _06671_ ? /* src = "generated/out/vanilla.sv:431.12-431.109|generated/out/vanilla.sv:431.8-434.11" */ 1'h0 : _05833_;
  assign _07472_ = _06673_ ? /* src = "generated/out/vanilla.sv:435.12-435.73|generated/out/vanilla.sv:435.8-438.11" */ 1'h0 : _05834_;
  assign _05835_ = _06517_ ? /* src = "generated/out/vanilla.sv:379.12-379.45|generated/out/vanilla.sv:379.8-382.11" */ 1'h0 : _05831_;
  assign _07475_ = _06519_ ? /* src = "generated/out/vanilla.sv:383.12-383.45|generated/out/vanilla.sv:383.8-386.11" */ 1'h0 : _05835_;
  assign _07477_ = _06521_ ? /* src = "generated/out/vanilla.sv:387.12-387.45|generated/out/vanilla.sv:387.8-390.11" */ mem_rdata_latched[12] : _07475_;
  assign _07479_ = _06523_ ? /* src = "generated/out/vanilla.sv:391.12-391.46|generated/out/vanilla.sv:391.8-401.11" */ _07607_[6] : _07477_;
  assign _07481_ = _00861_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:347.6-360.13" */ 1'h0 : _05831_;
  assign _00020_[31] = _06663_ ? /* src = "generated/out/vanilla.sv:344.7-344.72|generated/out/vanilla.sv:344.3-445.11" */ _06384_ : _05831_;
  assign _05840_ = mem_xfer ? /* src = "generated/out/vanilla.sv:340.7-340.15|generated/out/vanilla.sv:340.3-343.6" */ mem_rdata_latched[7] : mem_rdata_q[7];
  assign _07484_ = _07254_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:413.6-444.13" */ 1'h0 : _05840_;
  assign _07486_ = _01078_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:362.6-411.13" */ mem_rdata_latched[12] : _05840_;
  assign _07253_ = mem_rdata_latched[15:13] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:362.6-411.13" */ 3'h7;
  assign _00020_[7] = _06663_ ? /* src = "generated/out/vanilla.sv:344.7-344.72|generated/out/vanilla.sv:344.3-445.11" */ _06392_ : _05840_;
  assign _05844_ = mem_xfer ? /* src = "generated/out/vanilla.sv:340.7-340.15|generated/out/vanilla.sv:340.3-343.6" */ mem_rdata_latched[24:20] : mem_rdata_q[24:20];
  assign _05845_ = _06665_ ? /* src = "generated/out/vanilla.sv:423.12-423.73|generated/out/vanilla.sv:423.8-426.11" */ 5'h00 : _05844_;
  assign _07490_ = _06671_ ? /* src = "generated/out/vanilla.sv:431.12-431.109|generated/out/vanilla.sv:431.8-434.11" */ 5'h00 : _05845_;
  assign _07492_ = _06521_ ? /* src = "generated/out/vanilla.sv:387.12-387.45|generated/out/vanilla.sv:387.8-390.11" */ mem_rdata_latched[6:2] : _05844_;
  assign _07494_ = _06515_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:372.12-372.40|generated/out/vanilla.sv:372.8-377.88" */ { mem_rdata_latched[6], 4'h0 } : { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] };
  assign _00020_[24:20] = _06663_ ? /* src = "generated/out/vanilla.sv:344.7-344.72|generated/out/vanilla.sv:344.3-445.11" */ _06402_ : _05844_;
  assign _07496_ = mem_xfer ? /* src = "generated/out/vanilla.sv:340.7-340.15|generated/out/vanilla.sv:340.3-343.6" */ mem_rdata_latched[19:15] : mem_rdata_q[19:15];
  assign _07498_ = _06515_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:372.12-372.40|generated/out/vanilla.sv:372.8-377.88" */ _07496_ : { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[6:5] };
  assign _07500_ = _07265_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:362.6-411.13" */ _07498_ : _07496_;
  assign _07502_ = _07267_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:345.4-445.11" */ _07500_ : _07496_;
  assign _00020_[19:15] = _06663_ ? /* src = "generated/out/vanilla.sv:344.7-344.72|generated/out/vanilla.sv:344.3-445.11" */ _07502_ : _07496_;
  assign { _05651_[2:1], _05659_[0] } = mem_xfer ? /* src = "generated/out/vanilla.sv:340.7-340.15|generated/out/vanilla.sv:340.3-343.6" */ mem_rdata_latched[14:12] : mem_rdata_q[14:12];
  assign _05854_ = _06665_ ? /* src = "generated/out/vanilla.sv:423.12-423.73|generated/out/vanilla.sv:423.8-426.11" */ 3'h0 : { _05651_[2:1], _05659_[0] };
  assign _05855_ = _06667_ ? /* src = "generated/out/vanilla.sv:427.12-427.73|generated/out/vanilla.sv:427.8-430.11" */ 3'h0 : _05854_;
  assign _05856_ = _06671_ ? /* src = "generated/out/vanilla.sv:431.12-431.109|generated/out/vanilla.sv:431.8-434.11" */ 3'h0 : _05855_;
  assign { _05650_[2], _07508_[1], _05650_[0] } = _06673_ ? /* src = "generated/out/vanilla.sv:435.12-435.73|generated/out/vanilla.sv:435.8-438.11" */ 3'h0 : _05856_;
  assign { _07510_[2], _05857_[1], _07510_[0] } = _06517_ ? /* src = "generated/out/vanilla.sv:379.12-379.45|generated/out/vanilla.sv:379.8-382.11" */ 3'h5 : { _05651_[2:1], _05659_[0] };
  assign _07512_ = _06519_ ? /* src = "generated/out/vanilla.sv:383.12-383.45|generated/out/vanilla.sv:383.8-386.11" */ 3'h5 : { _07510_[2], _05857_[1], _07510_[0] };
  assign _05858_ = _06521_ ? /* src = "generated/out/vanilla.sv:387.12-387.45|generated/out/vanilla.sv:387.8-390.11" */ 3'h7 : _07512_;
  assign { _07515_[2], _05859_[1:0] } = _06525_ ? /* src = "generated/out/vanilla.sv:392.13-392.44|generated/out/vanilla.sv:392.9-393.39" */ 3'h0 : _05858_;
  assign { _07517_[2:1], _05860_[0] } = _06527_ ? /* src = "generated/out/vanilla.sv:394.13-394.44|generated/out/vanilla.sv:394.9-395.39" */ 3'h4 : { _07515_[2], _05859_[1:0] };
  assign _07519_ = _06529_ ? /* src = "generated/out/vanilla.sv:396.13-396.44|generated/out/vanilla.sv:396.9-397.39" */ 3'h6 : { _07517_[2:1], _05860_[0] };
  assign _07521_ = _06531_ ? /* src = "generated/out/vanilla.sv:398.13-398.44|generated/out/vanilla.sv:398.9-399.39" */ 3'h7 : _07519_;
  assign _07523_ = _06523_ ? /* src = "generated/out/vanilla.sv:391.12-391.46|generated/out/vanilla.sv:391.8-401.11" */ _07521_ : _05858_;
  assign _07525_ = _06515_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:372.12-372.40|generated/out/vanilla.sv:372.8-377.88" */ 3'h0 : mem_rdata_latched[4:2];
  assign _00020_[14:12] = _06663_ ? /* src = "generated/out/vanilla.sv:344.7-344.72|generated/out/vanilla.sv:344.3-445.11" */ _06424_ : { _05651_[2:1], _05659_[0] };
  assign _07527_ = mem_xfer ? /* src = "generated/out/vanilla.sv:340.7-340.15|generated/out/vanilla.sv:340.3-343.6" */ mem_rdata_latched[11:8] : mem_rdata_q[11:8];
  assign _07529_ = _07254_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:413.6-444.13" */ { mem_rdata_latched[11:9], 1'h0 } : _07527_;
  assign _07531_ = _01078_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:362.6-411.13" */ { mem_rdata_latched[11:10], mem_rdata_latched[4:3] } : _07527_;
  assign _07533_ = _07254_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:347.6-360.13" */ { mem_rdata_latched[11:10], mem_rdata_latched[6], 1'h0 } : _07527_;
  assign _00020_[11:8] = _06663_ ? /* src = "generated/out/vanilla.sv:344.7-344.72|generated/out/vanilla.sv:344.3-445.11" */ _06442_ : _07527_;
  assign _05665_ = mem_xfer ? /* src = "generated/out/vanilla.sv:340.7-340.15|generated/out/vanilla.sv:340.3-343.6" */ mem_rdata_latched[30:25] : mem_rdata_q[30:25];
  assign _05869_ = _06665_ ? /* src = "generated/out/vanilla.sv:423.12-423.73|generated/out/vanilla.sv:423.8-426.11" */ 6'h00 : _05665_;
  assign _05870_ = _06667_ ? /* src = "generated/out/vanilla.sv:427.12-427.73|generated/out/vanilla.sv:427.8-430.11" */ 6'h00 : _05869_;
  assign _05871_ = _06671_ ? /* src = "generated/out/vanilla.sv:431.12-431.109|generated/out/vanilla.sv:431.8-434.11" */ 6'h00 : _05870_;
  assign _07539_ = _06673_ ? /* src = "generated/out/vanilla.sv:435.12-435.73|generated/out/vanilla.sv:435.8-438.11" */ 6'h00 : _05871_;
  assign { _07541_[5], _05872_[4:0] } = _06517_ ? /* src = "generated/out/vanilla.sv:379.12-379.45|generated/out/vanilla.sv:379.8-382.11" */ 6'h00 : _05665_;
  assign _07543_ = _06519_ ? /* src = "generated/out/vanilla.sv:383.12-383.45|generated/out/vanilla.sv:383.8-386.11" */ 6'h20 : { _07541_[5], _05872_[4:0] };
  assign _07545_ = _06521_ ? /* src = "generated/out/vanilla.sv:387.12-387.45|generated/out/vanilla.sv:387.8-390.11" */ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] } : _07543_;
  assign _07547_ = _06523_ ? /* src = "generated/out/vanilla.sv:391.12-391.46|generated/out/vanilla.sv:391.8-401.11" */ _07607_[5:0] : _07545_;
  assign _07549_ = _06515_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:372.12-372.40|generated/out/vanilla.sv:372.8-377.88" */ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[4:3], mem_rdata_latched[5], mem_rdata_latched[2] } : { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] };
  assign _00020_[30:25] = _06663_ ? /* src = "generated/out/vanilla.sv:344.7-344.72|generated/out/vanilla.sv:344.3-445.11" */ _06456_ : _05665_;
  assign _07551_ = pcpi_rs1[1:0] == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:331.5-336.12" */ 2'h3;
  assign _07553_ = pcpi_rs1[1:0] == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:331.5-336.12" */ 2'h2;
  assign _07555_ = pcpi_rs1[1:0] == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:331.5-336.12" */ 2'h1;
  assign _07557_ = mem_wordsize == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:314.3-338.10" */ 2'h2;
  assign _06503_ = mem_wordsize == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:314.3-338.10" */ 2'h1;
  assign _06501_ = ! /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:314.3-338.10" */ mem_wordsize;
  assign _07559_ = last_mem_valid ? /* src = "generated/out/vanilla.sv:308.8-308.23|generated/out/vanilla.sv:308.4-309.46" */ mem_la_firstword_reg : mem_la_firstword;
  assign _00070_ = _06513_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1805.8-1805.35|generated/out/vanilla.sv:1805.4-1808.7" */ { rvfi_rd_wdata, 32'h00000000 } : _00053_;
  assign _00072_ = _06513_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1805.8-1805.35|generated/out/vanilla.sv:1805.4-1808.7" */ 64'hffffffff00000000 : _00055_;
  assign _00053_ = _06512_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1801.8-1801.35|generated/out/vanilla.sv:1801.4-1804.7" */ { 32'h00000000, rvfi_rd_wdata } : 64'h0000000000000000;
  assign _00055_ = _06512_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1801.8-1801.35|generated/out/vanilla.sv:1801.4-1804.7" */ 64'h00000000ffffffff : 64'h0000000000000000;
  assign _00066_ = _06510_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1797.8-1797.35|generated/out/vanilla.sv:1797.4-1800.7" */ { rvfi_rd_wdata, 32'h00000000 } : _00049_;
  assign _00068_ = _06510_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1797.8-1797.35|generated/out/vanilla.sv:1797.4-1800.7" */ 64'hffffffff00000000 : _00051_;
  assign _00049_ = _06509_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1793.8-1793.35|generated/out/vanilla.sv:1793.4-1796.7" */ { 32'h00000000, rvfi_rd_wdata } : 64'h0000000000000000;
  assign _07561_ = & /* src = "generated/out/vanilla.sv:296.113-296.123" */ mem_state;
  assign _07563_ = & /* src = "generated/out/vanilla.sv:298.265-298.288" */ mem_rdata_latched[1:0];
  assign _00475_ = & /* src = "generated/out/vanilla.sv:506.13-506.29" */ mem_rdata[1:0];
  assign _07429_ = & /* src = "generated/out/vanilla.sv:779.9-779.31" */ next_insn_opcode[1:0];
  assign _07143_ = | /* src = "generated/out/vanilla.sv:0.0-0.0" */ pcpi_timeout_counter;
  assign _07564_ = | /* src = "generated/out/vanilla.sv:1186.19-1186.57" */ decoded_rs1;
  assign _07566_ = | /* src = "generated/out/vanilla.sv:1187.19-1187.57" */ decoded_rs2;
  assign _07568_ = | /* src = "generated/out/vanilla.sv:1746.22-1746.53" */ latched_rd;
  assign _07570_ = | /* src = "generated/out/vanilla.sv:1776.24-1776.46" */ mem_wstrb;
  assign _07363_ = | /* src = "generated/out/vanilla.sv:1002.5-1002.30" */ { instr_auipc, instr_lui };
  assign pcpi_int_wait = | /* src = "generated/out/vanilla.sv:256.19-256.125" */ { pcpi_div_wait, pcpi_mul_wait };
  assign _07572_ = | /* src = "generated/out/vanilla.sv:296.44-296.54" */ mem_state;
  assign is_rdcycle_rdcycleh_rdinstr_rdinstrh = | /* src = "generated/out/vanilla.sv:610.48-610.111" */ { instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle };
  assign _00014_ = | /* src = "generated/out/vanilla.sv:790.23-790.59" */ { instr_jal, instr_auipc, instr_lui };
  assign _00016_ = | /* src = "generated/out/vanilla.sv:792.22-792.57" */ { instr_slt, instr_slti, instr_blt };
  assign _00018_ = | /* src = "generated/out/vanilla.sv:793.25-793.63" */ { instr_sltu, instr_sltiu, instr_bltu };
  assign _07573_ = | /* src = "generated/out/vanilla.sv:795.17-795.96" */ { is_beq_bne_blt_bge_bltu_bgeu, instr_sltu, instr_slt, instr_sltiu, instr_slti };
  assign _07575_ = | /* src = "generated/out/vanilla.sv:827.27-827.51" */ mem_rdata_latched[12:5];
  assign _07579_ = | /* src = "generated/out/vanilla.sv:995.78-995.259" */ { _06573_, _06571_, _06569_, _06567_, _06563_, _06559_ };
  assign _07577_ = | /* src = "generated/out/vanilla.sv:996.40-996.251" */ { _06811_, _06809_, _06807_ };
  assign _07581_ = 4'h1 << /* src = "generated/out/vanilla.sv:330.20-330.43" */ pcpi_rs1[1:0];
  assign _07583_ = pcpi_rs1 - /* src = "generated/out/vanilla.sv:1110.32-1110.49" */ pcpi_rs2;
  assign _07585_ = pcpi_timeout_counter - /* src = "generated/out/vanilla.sv:1216.30-1216.54" */ 32'd1;
  assign _07587_ = reg_sh - /* src = "generated/out/vanilla.sv:1591.17-1591.27" */ 32'd4;
  assign _07589_ = reg_sh - /* src = "generated/out/vanilla.sv:1600.17-1600.27" */ 32'd1;
  assign next_pc = _06599_ ? /* src = "generated/out/vanilla.sv:1080.20-1080.80" */ { reg_out[31:1], 1'h0 } : reg_next_pc;
  assign alu_add_sub = instr_sub ? /* src = "generated/out/vanilla.sv:1110.20-1110.69" */ _07583_ : _00084_;
  assign _07591_ = latched_compr ? /* src = "generated/out/vanilla.sv:1163.33-1163.54" */ 32'd2 : 32'd4;
  assign cpuregs_rs1 = _07564_ ? /* src = "generated/out/vanilla.sv:1186.19-1186.57" */ _05886_ : 32'd0;
  assign cpuregs_rs2 = _07566_ ? /* src = "generated/out/vanilla.sv:1187.19-1187.57" */ _05887_ : 32'd0;
  assign _07594_ = latched_store ? /* src = "generated/out/vanilla.sv:1280.37-1280.109" */ { _00110_[31:1], 1'h0 } : reg_next_pc;
  assign { _00110_[31:1], _07592_[0] } = latched_stalu ? /* src = "generated/out/vanilla.sv:1299.54-1299.89" */ alu_out_q : reg_out;
  assign _07596_ = compressed_instr ? /* src = "generated/out/vanilla.sv:1331.36-1331.60" */ 32'd2 : 32'd4;
  assign _07597_ = instr_lui ? /* src = "generated/out/vanilla.sv:1405.20-1405.42" */ 32'd0 : reg_pc;
  assign _07599_ = _07568_ ? /* src = "generated/out/vanilla.sv:1746.22-1746.53" */ cpuregs_wrdata : 32'd0;
  assign _07601_ = _07570_ ? /* src = "generated/out/vanilla.sv:1776.24-1776.46" */ 32'd0 : 32'd4294967295;
  assign mem_la_addr = _06633_ ? /* src = "generated/out/vanilla.sv:299.24-299.129" */ { _00102_, 2'h0 } : { pcpi_rs1[31:2], 2'h0 };
  assign mem_rdata_latched_noshuffle = mem_xfer ? /* src = "generated/out/vanilla.sv:300.40-300.95" */ mem_rdata : mem_rdata_q;
  assign mem_rdata_latched = mem_la_use_prefetched_high_word ? /* src = "generated/out/vanilla.sv:301.30-301.348" */ { 16'hxxxx, mem_16bit_buffer } : _07604_;
  assign _07602_ = mem_la_firstword ? /* src = "generated/out/vanilla.sv:301.221-301.346" */ { 16'hxxxx, mem_rdata_latched_noshuffle[31:16] } : mem_rdata_latched_noshuffle;
  assign _07604_ = mem_la_secondword ? /* src = "generated/out/vanilla.sv:301.126-301.347" */ { mem_rdata_latched_noshuffle[15:0], mem_16bit_buffer } : _07602_;
  assign _07606_ = pcpi_rs1[1] ? /* src = "generated/out/vanilla.sv:322.21-322.51" */ 4'hc : 4'h3;
  assign _07607_ = _06525_ ? /* src = "generated/out/vanilla.sv:400.32-400.89" */ 7'h20 : 7'h00;
  assign _07608_ = _06876_ ? /* src = "generated/out/vanilla.sv:512.22-512.58" */ 32'd0 : 32'd3;
  assign _07609_ = pcpi_rs1 ^ /* src = "generated/out/vanilla.sv:1135.39-1135.56" */ pcpi_rs2;
  /* module_not_derived = 32'd1 */
  /* src = "generated/out/vanilla.sv:213.22-224.5" */
  picorv32_pcpi_mul \genblk1.genblk1.pcpi_mul  (
    .clk(clk),
    .pcpi_insn(pcpi_insn),
    .pcpi_insn_t0(pcpi_insn_t0),
    .pcpi_rd(pcpi_mul_rd),
    .pcpi_rd_t0(pcpi_mul_rd_t0),
    .pcpi_ready(pcpi_mul_ready),
    .pcpi_ready_t0(pcpi_mul_ready_t0),
    .pcpi_rs1(pcpi_rs1),
    .pcpi_rs1_t0(pcpi_rs1_t0),
    .pcpi_rs2(pcpi_rs2),
    .pcpi_rs2_t0(pcpi_rs2_t0),
    .pcpi_valid(pcpi_valid),
    .pcpi_valid_t0(pcpi_valid_t0),
    .pcpi_wait(pcpi_mul_wait),
    .pcpi_wait_t0(pcpi_mul_wait_t0),
    .pcpi_wr(pcpi_mul_wr),
    .pcpi_wr_t0(pcpi_mul_wr_t0),
    .resetn(resetn)
  );
  /* module_not_derived = 32'd1 */
  /* src = "generated/out/vanilla.sv:233.22-244.5" */
  picorv32_pcpi_div \genblk2.pcpi_div  (
    .clk(clk),
    .pcpi_insn(pcpi_insn),
    .pcpi_insn_t0(pcpi_insn_t0),
    .pcpi_rd(pcpi_div_rd),
    .pcpi_rd_t0(pcpi_div_rd_t0),
    .pcpi_ready(pcpi_div_ready),
    .pcpi_ready_t0(pcpi_div_ready_t0),
    .pcpi_rs1(pcpi_rs1),
    .pcpi_rs1_t0(pcpi_rs1_t0),
    .pcpi_rs2(pcpi_rs2),
    .pcpi_rs2_t0(pcpi_rs2_t0),
    .pcpi_valid(pcpi_valid),
    .pcpi_valid_t0(pcpi_valid_t0),
    .pcpi_wait(pcpi_div_wait),
    .pcpi_wait_t0(pcpi_div_wait_t0),
    .pcpi_wr(pcpi_div_wr),
    .pcpi_wr_t0(pcpi_div_wr_t0),
    .resetn(resetn)
  );
  assign _00004_[30:0] = { _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31], _00004_[31] };
  assign _00005_[30:0] = { _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31], _00005_[31] };
  assign { _00052_[63:32], _00052_[30:0] } = { 32'h00000000, _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31], _00052_[31] };
  assign { _00056_[63:32], _00056_[30:0] } = { 32'h00000000, _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31], _00056_[31] };
  assign _00110_[0] = 1'h0;
  assign _00111_[0] = 1'h0;
  assign _05539_[3] = _00827_;
  assign _05541_[2] = _00822_;
  assign _05542_[3] = _00826_;
  assign _05544_[6] = _00825_;
  assign _05587_[1] = _00818_;
  assign _05650_[1] = _00829_;
  assign _05651_[0] = _00830_;
  assign _05659_[2:1] = _05651_[2:1];
  assign _05660_[1] = _00837_;
  assign _05745_[6] = _00821_;
  assign _05746_[6] = _00824_;
  assign _05749_[7] = _00841_;
  assign _05750_[7] = _00842_;
  assign _05802_[0] = _00819_;
  assign _05824_[1] = _00817_;
  assign { _05857_[2], _05857_[0] } = _00832_;
  assign _05859_[2] = _00834_;
  assign _05860_[2:1] = _00835_;
  assign _05872_[5] = _00838_;
  assign { _06167_[7], _06167_[5:0] } = { _05748_[7], _05748_[5:0] };
  assign { _06174_[7:3], _06174_[1:0] } = { _05541_[7:3], _05541_[1:0] };
  assign { _06177_[7:4], _06177_[2:0] } = { _05542_[7:4], _05542_[2:0] };
  assign { _06180_[7], _06180_[5:0] } = { _05544_[7], _05544_[5:0] };
  assign _06215_[0] = _06215_[1];
  assign { _06303_[3:2], _06303_[0] } = 3'h0;
  assign _06362_[4:1] = 4'h0;
  assign _06427_[2:1] = 2'h0;
  assign { _06434_[2], _06434_[0] } = { _05660_[2], _05660_[0] };
  assign { _07167_[7], _07167_[5:0] } = { _05745_[7], _05745_[5:0] };
  assign { _07171_[7], _07171_[5:0] } = { _05746_[7], _05746_[5:0] };
  assign { _07173_[7:4], _07173_[2:0] } = { _05539_[7:4], _05539_[2:0] };
  assign _07179_[6:0] = _05749_[6:0];
  assign _07181_[6:0] = _05750_[6:0];
  assign { _07299_[3:2], _07299_[0] } = { _05587_[3:2], _05587_[0] };
  assign _07380_[4:1] = _05802_[4:1];
  assign _07449_[0] = _05824_[0];
  assign { _07508_[2], _07508_[0] } = { _05650_[2], _05650_[0] };
  assign _07510_[1] = _05857_[1];
  assign _07515_[1:0] = _05859_[1:0];
  assign _07517_[0] = _05860_[0];
  assign _07541_[4:0] = _05872_[4:0];
  assign _07592_[31:1] = _00110_[31:1];
  assign _07593_[31:1] = _00111_[31:1];
  assign decoded_imm_j[0] = 1'h0;
  assign decoded_imm_j_t0[0] = 1'h0;
  assign eoi = 32'd0;
  assign eoi_t0 = 32'd0;
  assign rvfi_csr_mcycle_wdata = 64'h0000000000000000;
  assign rvfi_csr_mcycle_wdata_t0 = 64'h0000000000000000;
  assign rvfi_csr_mcycle_wmask = 64'h0000000000000000;
  assign rvfi_csr_mcycle_wmask_t0 = 64'h0000000000000000;
  assign rvfi_csr_minstret_wdata = 64'h0000000000000000;
  assign rvfi_csr_minstret_wdata_t0 = 64'h0000000000000000;
  assign rvfi_csr_minstret_wmask = 64'h0000000000000000;
  assign rvfi_csr_minstret_wmask_t0 = 64'h0000000000000000;
  assign rvfi_intr = 1'h0;
  assign rvfi_intr_t0 = 1'h0;
  assign rvfi_ixl = 2'h1;
  assign rvfi_ixl_t0 = 2'h0;
  assign rvfi_mode = 2'h3;
  assign rvfi_mode_t0 = 2'h0;
  assign rvfi_trap = rvfi_halt;
  assign rvfi_trap_t0 = rvfi_halt_t0;
  assign trace_data = 36'hxxxxxxxxx;
  assign trace_data_t0 = 36'h000000000;
  assign trace_valid = 1'h0;
  assign trace_valid_t0 = 1'h0;
endmodule

/* cellift =  1  */
/* hdlname = "\\picorv32_mem_top" */
/* top =  1  */
/* src = "generated/out/vanilla.sv:2703.1-2890.10" */
module picorv32_mem_top(clk, resetn, trap, instr_mem_req, instr_mem_gnt, instr_mem_addr, instr_mem_wdata, instr_mem_strb, instr_mem_we, instr_mem_rdata, data_mem_req, data_mem_gnt, data_mem_addr, data_mem_wdata, data_mem_strb, data_mem_we, data_mem_rdata, mem_la_read, mem_la_write, mem_la_addr, mem_la_wdata
, mem_la_wstrb, pcpi_valid, pcpi_insn, pcpi_rs1, pcpi_rs2, pcpi_wr, pcpi_rd, pcpi_wait, pcpi_ready, irq, eoi, trace_valid, trace_data, trap_t0, trace_valid_t0, trace_data_t0, pcpi_insn_t0, pcpi_rd_t0, pcpi_ready_t0, pcpi_rs1_t0, pcpi_rs2_t0
, pcpi_valid_t0, pcpi_wait_t0, pcpi_wr_t0, mem_la_wstrb_t0, mem_la_write_t0, mem_la_wdata_t0, mem_la_read_t0, mem_la_addr_t0, irq_t0, eoi_t0, data_mem_addr_t0, data_mem_gnt_t0, data_mem_rdata_t0, data_mem_req_t0, data_mem_strb_t0, data_mem_wdata_t0, data_mem_we_t0, instr_mem_addr_t0, instr_mem_gnt_t0, instr_mem_rdata_t0, instr_mem_req_t0
, instr_mem_strb_t0, instr_mem_wdata_t0, instr_mem_we_t0);
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _000_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _001_;
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire _002_;
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [3:0] _003_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [3:0] _004_;
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _005_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _006_;
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _007_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _008_;
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _009_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _010_;
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _011_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _012_;
  wire [31:0] _013_;
  wire [31:0] _014_;
  wire _015_;
  wire [3:0] _016_;
  wire [31:0] _017_;
  wire _018_;
  wire [31:0] _019_;
  wire [31:0] _020_;
  wire [31:0] _021_;
  wire [31:0] _022_;
  wire [31:0] _023_;
  wire [3:0] _024_;
  wire [3:0] _025_;
  wire [31:0] _026_;
  wire [31:0] _027_;
  wire [31:0] _028_;
  wire [31:0] _029_;
  wire [31:0] _030_;
  wire [31:0] _031_;
  wire _032_;
  wire _033_;
  wire [3:0] _034_;
  wire [3:0] _035_;
  wire [3:0] _036_;
  wire [31:0] _037_;
  wire [31:0] _038_;
  wire [31:0] _039_;
  wire [31:0] _040_;
  wire [31:0] _041_;
  wire [31:0] _042_;
  wire _043_;
  wire [3:0] _044_;
  wire [31:0] _045_;
  wire [31:0] _046_;
  wire [31:0] _047_;
  wire [31:0] _048_;
  wire [31:0] _049_;
  wire [31:0] _050_;
  wire [31:0] _051_;
  wire [31:0] _052_;
  wire [3:0] _053_;
  wire [31:0] _054_;
  wire [31:0] _055_;
  wire _056_;
  wire [3:0] _057_;
  wire [3:0] _058_;
  wire [3:0] _059_;
  wire [31:0] _060_;
  wire [31:0] _061_;
  wire [31:0] _062_;
  wire [31:0] _063_;
  wire [31:0] _064_;
  wire [3:0] _065_;
  wire [31:0] _066_;
  wire [31:0] _067_;
  /* src = "generated/out/vanilla.sv:2739.8-2739.11" */
  input clk;
  wire clk;
  /* src = "generated/out/vanilla.sv:2751.20-2751.33" */
  output [31:0] data_mem_addr;
  wire [31:0] data_mem_addr;
  /* cellift = 32'd1 */
  output [31:0] data_mem_addr_t0;
  wire [31:0] data_mem_addr_t0;
  /* src = "generated/out/vanilla.sv:2750.13-2750.25" */
  input data_mem_gnt;
  wire data_mem_gnt;
  /* cellift = 32'd1 */
  input data_mem_gnt_t0;
  wire data_mem_gnt_t0;
  /* src = "generated/out/vanilla.sv:2755.20-2755.34" */
  input [31:0] data_mem_rdata;
  wire [31:0] data_mem_rdata;
  /* cellift = 32'd1 */
  input [31:0] data_mem_rdata_t0;
  wire [31:0] data_mem_rdata_t0;
  /* src = "generated/out/vanilla.sv:2749.13-2749.25" */
  output data_mem_req;
  wire data_mem_req;
  /* cellift = 32'd1 */
  output data_mem_req_t0;
  wire data_mem_req_t0;
  /* src = "generated/out/vanilla.sv:2753.19-2753.32" */
  output [3:0] data_mem_strb;
  wire [3:0] data_mem_strb;
  /* cellift = 32'd1 */
  output [3:0] data_mem_strb_t0;
  wire [3:0] data_mem_strb_t0;
  /* src = "generated/out/vanilla.sv:2752.20-2752.34" */
  output [31:0] data_mem_wdata;
  wire [31:0] data_mem_wdata;
  /* cellift = 32'd1 */
  output [31:0] data_mem_wdata_t0;
  wire [31:0] data_mem_wdata_t0;
  /* src = "generated/out/vanilla.sv:2754.13-2754.24" */
  output data_mem_we;
  wire data_mem_we;
  /* cellift = 32'd1 */
  output data_mem_we_t0;
  wire data_mem_we_t0;
  /* src = "generated/out/vanilla.sv:2770.20-2770.23" */
  output [31:0] eoi;
  wire [31:0] eoi;
  /* cellift = 32'd1 */
  output [31:0] eoi_t0;
  wire [31:0] eoi_t0;
  /* src = "generated/out/vanilla.sv:2744.20-2744.34" */
  output [31:0] instr_mem_addr;
  wire [31:0] instr_mem_addr;
  /* cellift = 32'd1 */
  output [31:0] instr_mem_addr_t0;
  wire [31:0] instr_mem_addr_t0;
  /* src = "generated/out/vanilla.sv:2743.13-2743.26" */
  input instr_mem_gnt;
  wire instr_mem_gnt;
  /* cellift = 32'd1 */
  input instr_mem_gnt_t0;
  wire instr_mem_gnt_t0;
  /* src = "generated/out/vanilla.sv:2748.20-2748.35" */
  input [31:0] instr_mem_rdata;
  wire [31:0] instr_mem_rdata;
  /* cellift = 32'd1 */
  input [31:0] instr_mem_rdata_t0;
  wire [31:0] instr_mem_rdata_t0;
  /* src = "generated/out/vanilla.sv:2742.13-2742.26" */
  output instr_mem_req;
  wire instr_mem_req;
  /* cellift = 32'd1 */
  output instr_mem_req_t0;
  wire instr_mem_req_t0;
  /* src = "generated/out/vanilla.sv:2746.19-2746.33" */
  output [3:0] instr_mem_strb;
  wire [3:0] instr_mem_strb;
  /* cellift = 32'd1 */
  output [3:0] instr_mem_strb_t0;
  wire [3:0] instr_mem_strb_t0;
  /* src = "generated/out/vanilla.sv:2745.20-2745.35" */
  output [31:0] instr_mem_wdata;
  wire [31:0] instr_mem_wdata;
  /* cellift = 32'd1 */
  output [31:0] instr_mem_wdata_t0;
  wire [31:0] instr_mem_wdata_t0;
  /* src = "generated/out/vanilla.sv:2747.13-2747.25" */
  output instr_mem_we;
  wire instr_mem_we;
  /* cellift = 32'd1 */
  output instr_mem_we_t0;
  wire instr_mem_we_t0;
  /* src = "generated/out/vanilla.sv:2769.15-2769.18" */
  input [31:0] irq;
  wire [31:0] irq;
  /* cellift = 32'd1 */
  input [31:0] irq_t0;
  wire [31:0] irq_t0;
  /* src = "generated/out/vanilla.sv:2776.14-2776.22" */
  /* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] mem_addr;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2776.14-2776.22" */
  /* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] mem_addr_t0;
  /* src = "generated/out/vanilla.sv:2774.7-2774.16" */
  wire mem_instr;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2774.7-2774.16" */
  wire mem_instr_t0;
  /* src = "generated/out/vanilla.sv:2758.21-2758.32" */
  output [31:0] mem_la_addr;
  wire [31:0] mem_la_addr;
  /* cellift = 32'd1 */
  output [31:0] mem_la_addr_t0;
  wire [31:0] mem_la_addr_t0;
  /* src = "generated/out/vanilla.sv:2756.14-2756.25" */
  output mem_la_read;
  wire mem_la_read;
  /* cellift = 32'd1 */
  output mem_la_read_t0;
  wire mem_la_read_t0;
  /* src = "generated/out/vanilla.sv:2759.20-2759.32" */
  output [31:0] mem_la_wdata;
  wire [31:0] mem_la_wdata;
  /* cellift = 32'd1 */
  output [31:0] mem_la_wdata_t0;
  wire [31:0] mem_la_wdata_t0;
  /* src = "generated/out/vanilla.sv:2757.14-2757.26" */
  output mem_la_write;
  wire mem_la_write;
  /* cellift = 32'd1 */
  output mem_la_write_t0;
  wire mem_la_write_t0;
  /* src = "generated/out/vanilla.sv:2760.19-2760.31" */
  output [3:0] mem_la_wstrb;
  wire [3:0] mem_la_wstrb;
  /* cellift = 32'd1 */
  output [3:0] mem_la_wstrb_t0;
  wire [3:0] mem_la_wstrb_t0;
  /* src = "generated/out/vanilla.sv:2779.13-2779.22" */
  wire [31:0] mem_rdata;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2779.13-2779.22" */
  wire [31:0] mem_rdata_t0;
  /* src = "generated/out/vanilla.sv:2775.7-2775.16" */
  wire mem_ready;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2775.7-2775.16" */
  wire mem_ready_t0;
  /* src = "generated/out/vanilla.sv:2777.14-2777.23" */
  /* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] mem_wdata;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2777.14-2777.23" */
  /* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] mem_wdata_t0;
  /* src = "generated/out/vanilla.sv:2778.13-2778.22" */
  /* unused_bits = "0 1 2 3" */
  wire [3:0] mem_wstrb;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2778.13-2778.22" */
  /* unused_bits = "0 1 2 3" */
  wire [3:0] mem_wstrb_t0;
  /* src = "generated/out/vanilla.sv:2762.20-2762.29" */
  output [31:0] pcpi_insn;
  wire [31:0] pcpi_insn;
  /* cellift = 32'd1 */
  output [31:0] pcpi_insn_t0;
  wire [31:0] pcpi_insn_t0;
  /* src = "generated/out/vanilla.sv:2766.15-2766.22" */
  input [31:0] pcpi_rd;
  wire [31:0] pcpi_rd;
  /* cellift = 32'd1 */
  input [31:0] pcpi_rd_t0;
  wire [31:0] pcpi_rd_t0;
  /* src = "generated/out/vanilla.sv:2768.8-2768.18" */
  input pcpi_ready;
  wire pcpi_ready;
  /* cellift = 32'd1 */
  input pcpi_ready_t0;
  wire pcpi_ready_t0;
  /* src = "generated/out/vanilla.sv:2763.21-2763.29" */
  output [31:0] pcpi_rs1;
  wire [31:0] pcpi_rs1;
  /* cellift = 32'd1 */
  output [31:0] pcpi_rs1_t0;
  wire [31:0] pcpi_rs1_t0;
  /* src = "generated/out/vanilla.sv:2764.21-2764.29" */
  output [31:0] pcpi_rs2;
  wire [31:0] pcpi_rs2;
  /* cellift = 32'd1 */
  output [31:0] pcpi_rs2_t0;
  wire [31:0] pcpi_rs2_t0;
  /* src = "generated/out/vanilla.sv:2761.13-2761.23" */
  output pcpi_valid;
  wire pcpi_valid;
  /* cellift = 32'd1 */
  output pcpi_valid_t0;
  wire pcpi_valid_t0;
  /* src = "generated/out/vanilla.sv:2767.8-2767.17" */
  input pcpi_wait;
  wire pcpi_wait;
  /* cellift = 32'd1 */
  input pcpi_wait_t0;
  wire pcpi_wait_t0;
  /* src = "generated/out/vanilla.sv:2765.8-2765.15" */
  input pcpi_wr;
  wire pcpi_wr;
  /* cellift = 32'd1 */
  input pcpi_wr_t0;
  wire pcpi_wr_t0;
  /* src = "generated/out/vanilla.sv:2740.8-2740.14" */
  input resetn;
  wire resetn;
  /* src = "generated/out/vanilla.sv:2772.20-2772.30" */
  output [35:0] trace_data;
  wire [35:0] trace_data;
  /* cellift = 32'd1 */
  output [35:0] trace_data_t0;
  wire [35:0] trace_data_t0;
  /* src = "generated/out/vanilla.sv:2771.13-2771.24" */
  output trace_valid;
  wire trace_valid;
  /* cellift = 32'd1 */
  output trace_valid_t0;
  wire trace_valid_t0;
  /* src = "generated/out/vanilla.sv:2741.13-2741.17" */
  output trap;
  wire trap;
  /* cellift = 32'd1 */
  output trap_t0;
  wire trap_t0;
  assign _013_ = ~ { mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr };
  assign _014_ = ~ { mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write };
  assign _015_ = ~ mem_la_read;
  assign _017_ = ~ { mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read };
  assign _016_ = ~ { mem_la_read, mem_la_read, mem_la_read, mem_la_read };
  assign _049_ = { mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0 } | _013_;
  assign _054_ = { mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0 } | _014_;
  assign _056_ = instr_mem_req_t0 | _015_;
  assign _057_ = { instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0 } | _016_;
  assign _060_ = { instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0 } | _017_;
  assign _050_ = { mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0 } | { mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr };
  assign _052_ = { mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0 } | { mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready };
  assign _053_ = { mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0 } | { mem_la_write, mem_la_write, mem_la_write, mem_la_write };
  assign _055_ = { mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0 } | { mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write };
  assign _061_ = { instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0 } | { mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read };
  assign _058_ = { instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0 } | { mem_la_read, mem_la_read, mem_la_read, mem_la_read };
  assign _019_ = data_mem_rdata_t0 & _049_;
  assign _030_ = _010_ & _054_;
  assign _032_ = mem_la_write_t0 & _056_;
  assign _034_ = _004_ & _057_;
  assign _037_ = _006_ & _060_;
  assign _040_ = _001_ & _060_;
  assign _047_ = _008_ & _060_;
  assign _020_ = instr_mem_rdata_t0 & _050_;
  assign _022_ = _012_ & _052_;
  assign _024_ = mem_la_wstrb_t0 & _053_;
  assign _026_ = mem_la_wdata_t0 & _055_;
  assign _028_ = mem_la_addr_t0 & _055_;
  assign _035_ = mem_la_wstrb_t0 & _058_;
  assign _038_ = mem_la_wdata_t0 & _061_;
  assign _041_ = mem_la_addr_t0 & _061_;
  assign _051_ = _019_ | _020_;
  assign _059_ = _034_ | _035_;
  assign _062_ = _037_ | _038_;
  assign _063_ = _040_ | _041_;
  assign _064_ = data_mem_rdata ^ instr_mem_rdata;
  assign _065_ = _003_ ^ mem_la_wstrb;
  assign _066_ = _005_ ^ mem_la_wdata;
  assign _067_ = _000_ ^ mem_la_addr;
  assign _021_ = { mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0, mem_instr_t0 } & _064_;
  assign _023_ = { mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0, mem_ready_t0 } & _011_;
  assign _025_ = { mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0 } & mem_la_wstrb;
  assign _027_ = { mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0 } & mem_la_wdata;
  assign _029_ = { mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0 } & mem_la_addr;
  assign _031_ = { mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0, mem_la_write_t0 } & _009_;
  assign _033_ = instr_mem_req_t0 & _002_;
  assign _036_ = { instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0 } & _065_;
  assign _039_ = { instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0 } & _066_;
  assign _042_ = { instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0 } & _067_;
  assign _043_ = instr_mem_req_t0 & _018_;
  assign _044_ = { instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0 } & mem_la_wstrb;
  assign _045_ = { instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0 } & mem_la_wdata;
  assign _046_ = { instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0 } & mem_la_addr;
  assign _048_ = { instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0, instr_mem_req_t0 } & _007_;
  assign _012_ = _021_ | _051_;
  assign _010_ = _023_ | _022_;
  assign _004_ = _025_ | _024_;
  assign _006_ = _027_ | _026_;
  assign _001_ = _029_ | _028_;
  assign _008_ = _031_ | _030_;
  assign data_mem_we_t0 = _033_ | _032_;
  assign data_mem_strb_t0 = _036_ | _059_;
  assign data_mem_wdata_t0 = _039_ | _062_;
  assign data_mem_addr_t0 = _042_ | _063_;
  assign data_mem_req_t0 = _043_ | _032_;
  assign instr_mem_strb_t0 = _044_ | _035_;
  assign instr_mem_wdata_t0 = _045_ | _038_;
  assign instr_mem_addr_t0 = _046_ | _041_;
  assign mem_rdata_t0 = _048_ | _047_;
  assign _018_ = ~ _002_;
  assign _011_ = mem_instr ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2813.8-2813.17|generated/out/vanilla.sv:2813.4-2816.32" */ instr_mem_rdata : data_mem_rdata;
  assign _009_ = mem_ready ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2812.12-2812.21|generated/out/vanilla.sv:2812.8-2816.32" */ _011_ : 32'd0;
  assign _003_ = mem_la_write ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2805.12-2805.24|generated/out/vanilla.sv:2805.8-2816.32" */ mem_la_wstrb : 4'h0;
  assign _005_ = mem_la_write ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2805.12-2805.24|generated/out/vanilla.sv:2805.8-2816.32" */ mem_la_wdata : 32'd0;
  assign _000_ = mem_la_write ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2805.12-2805.24|generated/out/vanilla.sv:2805.8-2816.32" */ mem_la_addr : 32'd0;
  assign _002_ = mem_la_write ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2805.12-2805.24|generated/out/vanilla.sv:2805.8-2816.32" */ 1'h1 : 1'h0;
  assign _007_ = mem_la_write ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2805.12-2805.24|generated/out/vanilla.sv:2805.8-2816.32" */ 32'd0 : _009_;
  assign data_mem_we = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ 1'h0 : _002_;
  assign data_mem_strb = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ mem_la_wstrb : _003_;
  assign data_mem_wdata = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ mem_la_wdata : _005_;
  assign data_mem_addr = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ mem_la_addr : _000_;
  assign data_mem_req = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ 1'h1 : _002_;
  assign instr_mem_strb = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ mem_la_wstrb : 4'h0;
  assign instr_mem_wdata = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ mem_la_wdata : 32'd0;
  assign instr_mem_addr = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ mem_la_addr : 32'd0;
  assign instr_mem_req = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ 1'h1 : 1'h0;
  assign mem_rdata = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ 32'd0 : _007_;
  /* module_not_derived = 32'd1 */
  /* src = "generated/out/vanilla.sv:2861.4-2889.3" */
  \$paramod$47f4aa12d94f6638b23e6ab3bef6a1a82f6ab57b\picorv32  i_picorv32 (
    .clk(clk),
    .eoi(eoi),
    .eoi_t0(eoi_t0),
    .irq(irq),
    .irq_t0(irq_t0),
    .mem_addr(mem_addr),
    .mem_addr_t0(mem_addr_t0),
    .mem_instr(mem_instr),
    .mem_instr_t0(mem_instr_t0),
    .mem_la_addr(mem_la_addr),
    .mem_la_addr_t0(mem_la_addr_t0),
    .mem_la_read(mem_la_read),
    .mem_la_read_t0(instr_mem_req_t0),
    .mem_la_wdata(mem_la_wdata),
    .mem_la_wdata_t0(mem_la_wdata_t0),
    .mem_la_write(mem_la_write),
    .mem_la_write_t0(mem_la_write_t0),
    .mem_la_wstrb(mem_la_wstrb),
    .mem_la_wstrb_t0(mem_la_wstrb_t0),
    .mem_rdata(mem_rdata),
    .mem_rdata_t0(mem_rdata_t0),
    .mem_ready(mem_ready),
    .mem_ready_t0(mem_ready_t0),
    .mem_valid(mem_ready),
    .mem_valid_t0(mem_ready_t0),
    .mem_wdata(mem_wdata),
    .mem_wdata_t0(mem_wdata_t0),
    .mem_wstrb(mem_wstrb),
    .mem_wstrb_t0(mem_wstrb_t0),
    .pcpi_insn(pcpi_insn),
    .pcpi_insn_t0(pcpi_insn_t0),
    .pcpi_rd(pcpi_rd),
    .pcpi_rd_t0(pcpi_rd_t0),
    .pcpi_ready(pcpi_ready),
    .pcpi_ready_t0(pcpi_ready_t0),
    .pcpi_rs1(pcpi_rs1),
    .pcpi_rs1_t0(pcpi_rs1_t0),
    .pcpi_rs2(pcpi_rs2),
    .pcpi_rs2_t0(pcpi_rs2_t0),
    .pcpi_valid(pcpi_valid),
    .pcpi_valid_t0(pcpi_valid_t0),
    .pcpi_wait(pcpi_wait),
    .pcpi_wait_t0(pcpi_wait_t0),
    .pcpi_wr(pcpi_wr),
    .pcpi_wr_t0(pcpi_wr_t0),
    .resetn(resetn),
    .trace_data(trace_data),
    .trace_data_t0(trace_data_t0),
    .trace_valid(trace_valid),
    .trace_valid_t0(trace_valid_t0),
    .trap(trap),
    .trap_t0(trap_t0)
  );
  assign instr_mem_we = 1'h0;
  assign instr_mem_we_t0 = 1'h0;
  assign mem_la_read_t0 = instr_mem_req_t0;
endmodule

/* cellift =  1  */
/* hdlname = "\\picorv32_pcpi_div" */
/* src = "generated/out/vanilla.sv:2055.1-2137.10" */
module picorv32_pcpi_div(clk, resetn, pcpi_valid, pcpi_insn, pcpi_rs1, pcpi_rs2, pcpi_wr, pcpi_rd, pcpi_wait, pcpi_ready, pcpi_insn_t0, pcpi_rd_t0, pcpi_ready_t0, pcpi_rs1_t0, pcpi_rs2_t0, pcpi_valid_t0, pcpi_wait_t0, pcpi_wr_t0);
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
  wire [31:0] _000_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
  wire [31:0] _001_;
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
  wire _002_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
  wire _003_;
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
  wire _004_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire [1:0] _012_;
  wire _013_;
  wire [2:0] _014_;
  wire [61:0] _015_;
  wire _016_;
  wire [61:0] _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire [2:0] _022_;
  wire [31:0] _023_;
  wire [3:0] _024_;
  wire [31:0] _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire [31:0] _036_;
  wire [31:0] _037_;
  wire [31:0] _038_;
  wire [62:0] _039_;
  wire [62:0] _040_;
  wire [31:0] _041_;
  wire [62:0] _042_;
  wire [31:0] _043_;
  wire [31:0] _044_;
  wire [62:0] _045_;
  wire [31:0] _046_;
  wire [31:0] _047_;
  wire [31:0] _048_;
  wire [62:0] _049_;
  wire [31:0] _050_;
  wire [31:0] _051_;
  wire [31:0] _052_;
  wire [62:0] _053_;
  wire [31:0] _054_;
  wire [31:0] _055_;
  wire _056_;
  wire _057_;
  wire [31:0] _058_;
  wire [31:0] _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire [62:0] _065_;
  wire [62:0] _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  /* cellift = 32'd1 */
  wire _070_;
  wire _071_;
  /* cellift = 32'd1 */
  wire _072_;
  wire _073_;
  /* cellift = 32'd1 */
  wire _074_;
  wire _075_;
  /* cellift = 32'd1 */
  wire _076_;
  wire _077_;
  /* cellift = 32'd1 */
  wire _078_;
  wire _079_;
  /* cellift = 32'd1 */
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire [31:0] _088_;
  wire [31:0] _089_;
  wire [31:0] _090_;
  wire [31:0] _091_;
  wire [31:0] _092_;
  wire [31:0] _093_;
  wire [31:0] _094_;
  wire [31:0] _095_;
  wire [31:0] _096_;
  wire [30:0] _097_;
  wire [30:0] _098_;
  wire [30:0] _099_;
  wire [31:0] _100_;
  wire [31:0] _101_;
  wire [31:0] _102_;
  wire [1:0] _103_;
  wire [2:0] _104_;
  wire _105_;
  wire [61:0] _106_;
  wire [61:0] _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire [31:0] _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire [31:0] _141_;
  wire [62:0] _142_;
  wire [31:0] _143_;
  wire [31:0] _144_;
  wire [31:0] _145_;
  wire [31:0] _146_;
  wire [31:0] _147_;
  wire [31:0] _148_;
  wire [31:0] _149_;
  wire [31:0] _150_;
  wire [62:0] _151_;
  wire [62:0] _152_;
  wire [62:0] _153_;
  wire [31:0] _154_;
  wire [31:0] _155_;
  wire [31:0] _156_;
  wire [2:0] _157_;
  wire [3:0] _158_;
  wire [31:0] _159_;
  wire [62:0] _160_;
  wire [62:0] _161_;
  wire [31:0] _162_;
  wire [31:0] _163_;
  wire [31:0] _164_;
  wire [62:0] _165_;
  wire [62:0] _166_;
  wire [62:0] _167_;
  wire [31:0] _168_;
  wire [31:0] _169_;
  wire [31:0] _170_;
  wire [31:0] _171_;
  wire [31:0] _172_;
  wire [31:0] _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire [31:0] _182_;
  wire [31:0] _183_;
  wire [31:0] _184_;
  wire [31:0] _185_;
  wire [31:0] _186_;
  wire [31:0] _187_;
  wire [31:0] _188_;
  wire [31:0] _189_;
  wire [31:0] _190_;
  wire [31:0] _191_;
  wire [31:0] _192_;
  wire [31:0] _193_;
  wire [30:0] _194_;
  wire [30:0] _195_;
  wire [30:0] _196_;
  wire [30:0] _197_;
  wire [31:0] _198_;
  wire [31:0] _199_;
  wire [31:0] _200_;
  wire [31:0] _201_;
  wire [1:0] _202_;
  wire [1:0] _203_;
  wire [2:0] _204_;
  wire _205_;
  wire [61:0] _206_;
  wire [61:0] _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire [31:0] _219_;
  wire [62:0] _220_;
  wire [31:0] _221_;
  wire [31:0] _222_;
  wire [31:0] _223_;
  wire [31:0] _224_;
  wire [31:0] _225_;
  wire [31:0] _226_;
  wire [31:0] _227_;
  wire [31:0] _228_;
  wire [31:0] _229_;
  wire [31:0] _230_;
  wire [31:0] _231_;
  wire [62:0] _232_;
  wire [62:0] _233_;
  wire [62:0] _234_;
  wire [62:0] _235_;
  wire [31:0] _236_;
  wire [62:0] _237_;
  wire [62:0] _238_;
  wire [62:0] _239_;
  wire [31:0] _240_;
  wire [31:0] _241_;
  wire [31:0] _242_;
  wire [62:0] _243_;
  wire [62:0] _244_;
  wire [62:0] _245_;
  wire [31:0] _246_;
  wire [31:0] _247_;
  wire [31:0] _248_;
  wire [31:0] _249_;
  wire _250_;
  wire _251_;
  wire [31:0] _252_;
  wire [31:0] _253_;
  wire [31:0] _254_;
  wire [30:0] _255_;
  wire [31:0] _256_;
  wire [31:0] _257_;
  wire [62:0] _258_;
  wire [31:0] _259_;
  wire [31:0] _260_;
  wire [31:0] _261_;
  wire [62:0] _262_;
  wire [31:0] _263_;
  wire [62:0] _264_;
  wire [31:0] _265_;
  wire [62:0] _266_;
  wire [31:0] _267_;
  wire [31:0] _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire [62:0] _275_;
  wire [62:0] _276_;
  /* src = "generated/out/vanilla.sv:2089.52-2089.80" */
  wire _277_;
  /* src = "generated/out/vanilla.sv:2089.87-2089.117" */
  wire _278_;
  /* src = "generated/out/vanilla.sv:2129.8-2129.27" */
  wire _279_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2129.8-2129.27" */
  wire _280_;
  /* src = "generated/out/vanilla.sv:2089.10-2089.30" */
  wire _281_;
  /* src = "generated/out/vanilla.sv:2089.9-2089.46" */
  wire _282_;
  /* src = "generated/out/vanilla.sv:2089.8-2089.81" */
  wire _283_;
  /* src = "generated/out/vanilla.sv:2089.7-2089.118" */
  wire _284_;
  /* src = "generated/out/vanilla.sv:2113.17-2113.57" */
  wire _285_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2113.17-2113.57" */
  wire _286_;
  /* src = "generated/out/vanilla.sv:2114.16-2114.56" */
  wire _287_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2114.16-2114.56" */
  wire _288_;
  /* src = "generated/out/vanilla.sv:2115.17-2115.60" */
  wire _289_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2115.17-2115.60" */
  wire _290_;
  /* src = "generated/out/vanilla.sv:2115.16-2115.74" */
  wire _291_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2115.16-2115.74" */
  wire _292_;
  /* src = "generated/out/vanilla.sv:2115.80-2115.105" */
  wire _293_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2115.80-2115.105" */
  wire _294_;
  /* src = "generated/out/vanilla.sv:2119.12-2119.36" */
  wire _295_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2119.12-2119.36" */
  wire _296_;
  /* src = "generated/out/vanilla.sv:2083.28-2083.40" */
  wire _297_;
  /* src = "generated/out/vanilla.sv:2089.35-2089.46" */
  wire _298_;
  /* src = "generated/out/vanilla.sv:2119.12-2119.25" */
  wire _299_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2119.12-2119.25" */
  wire _300_;
  /* src = "generated/out/vanilla.sv:2113.18-2113.40" */
  wire _301_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2113.18-2113.40" */
  wire _302_;
  /* src = "generated/out/vanilla.sv:2115.15-2115.106" */
  wire _303_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2115.15-2115.106" */
  wire _304_;
  /* src = "generated/out/vanilla.sv:2123.8-2123.31" */
  wire _305_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2123.8-2123.31" */
  wire _306_;
  /* src = "generated/out/vanilla.sv:2115.31-2115.59" */
  wire _307_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2115.31-2115.59" */
  wire _308_;
  /* src = "generated/out/vanilla.sv:2113.60-2113.69" */
  wire [31:0] _309_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2113.60-2113.69" */
  wire [31:0] _310_;
  /* src = "generated/out/vanilla.sv:2114.59-2114.68" */
  wire [62:0] _311_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2114.59-2114.68" */
  wire [62:0] _312_;
  /* src = "generated/out/vanilla.sv:2124.27-2124.36" */
  wire [31:0] _313_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2124.27-2124.36" */
  wire [31:0] _314_;
  /* src = "generated/out/vanilla.sv:2126.27-2126.36" */
  wire [31:0] _315_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2126.27-2126.36" */
  wire [31:0] _316_;
  /* src = "generated/out/vanilla.sv:2131.17-2131.40" */
  wire [31:0] _317_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2131.17-2131.40" */
  wire [31:0] _318_;
  wire [31:0] _319_;
  /* cellift = 32'd1 */
  wire [31:0] _320_;
  wire [31:0] _321_;
  /* cellift = 32'd1 */
  wire [31:0] _322_;
  wire [31:0] _323_;
  /* cellift = 32'd1 */
  wire [31:0] _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  /* cellift = 32'd1 */
  wire _328_;
  wire [31:0] _329_;
  /* cellift = 32'd1 */
  wire [31:0] _330_;
  wire [31:0] _331_;
  /* cellift = 32'd1 */
  wire [31:0] _332_;
  wire [31:0] _333_;
  /* cellift = 32'd1 */
  wire [31:0] _334_;
  wire [62:0] _335_;
  /* cellift = 32'd1 */
  wire [62:0] _336_;
  /* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30" */
  wire [62:0] _337_;
  /* cellift = 32'd1 */
  /* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30" */
  wire [62:0] _338_;
  wire [31:0] _339_;
  /* cellift = 32'd1 */
  wire [31:0] _340_;
  wire [31:0] _341_;
  /* cellift = 32'd1 */
  wire [31:0] _342_;
  wire [31:0] _343_;
  /* cellift = 32'd1 */
  wire [31:0] _344_;
  wire _345_;
  /* cellift = 32'd1 */
  wire _346_;
  wire _347_;
  wire _348_;
  /* cellift = 32'd1 */
  wire _349_;
  wire _350_;
  wire _351_;
  /* cellift = 32'd1 */
  wire _352_;
  wire _353_;
  wire _354_;
  /* cellift = 32'd1 */
  wire _355_;
  wire _356_;
  /* src = "generated/out/vanilla.sv:2115.65-2115.74" */
  wire _357_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2115.65-2115.74" */
  wire _358_;
  /* src = "generated/out/vanilla.sv:2114.15-2114.86" */
  wire [62:0] _359_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2114.15-2114.86" */
  wire [62:0] _360_;
  /* src = "generated/out/vanilla.sv:2130.17-2130.35" */
  /* unused_bits = "32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62" */
  wire [62:0] _361_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2130.17-2130.35" */
  /* unused_bits = "32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62" */
  wire [62:0] _362_;
  /* src = "generated/out/vanilla.sv:2113.17-2113.80" */
  wire [31:0] _363_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2113.17-2113.80" */
  wire [31:0] _364_;
  /* src = "generated/out/vanilla.sv:2114.16-2114.79" */
  /* unused_bits = "32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62" */
  wire [62:0] _365_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2114.16-2114.79" */
  /* unused_bits = "32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62" */
  wire [62:0] _366_;
  /* src = "generated/out/vanilla.sv:2124.17-2124.47" */
  wire [31:0] _367_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2124.17-2124.47" */
  wire [31:0] _368_;
  /* src = "generated/out/vanilla.sv:2126.17-2126.47" */
  wire [31:0] _369_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2126.17-2126.47" */
  wire [31:0] _370_;
  /* src = "generated/out/vanilla.sv:2067.8-2067.11" */
  input clk;
  wire clk;
  /* src = "generated/out/vanilla.sv:2099.13-2099.21" */
  reg [31:0] dividend;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2099.13-2099.21" */
  reg [31:0] dividend_t0;
  /* src = "generated/out/vanilla.sv:2100.13-2100.20" */
  reg [62:0] divisor;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2100.13-2100.20" */
  reg [62:0] divisor_t0;
  /* src = "generated/out/vanilla.sv:2081.7-2081.24" */
  wire instr_any_div_rem;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2081.7-2081.24" */
  wire instr_any_div_rem_t0;
  /* src = "generated/out/vanilla.sv:2077.6-2077.15" */
  reg instr_div;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2077.6-2077.15" */
  reg instr_div_t0;
  /* src = "generated/out/vanilla.sv:2078.6-2078.16" */
  reg instr_divu;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2078.6-2078.16" */
  reg instr_divu_t0;
  /* src = "generated/out/vanilla.sv:2079.6-2079.15" */
  reg instr_rem;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2079.6-2079.15" */
  reg instr_rem_t0;
  /* src = "generated/out/vanilla.sv:2080.6-2080.16" */
  reg instr_remu;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2080.6-2080.16" */
  reg instr_remu_t0;
  /* src = "generated/out/vanilla.sv:2104.6-2104.13" */
  reg outsign;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2104.6-2104.13" */
  reg outsign_t0;
  /* src = "generated/out/vanilla.sv:2070.15-2070.24" */
  input [31:0] pcpi_insn;
  wire [31:0] pcpi_insn;
  /* cellift = 32'd1 */
  input [31:0] pcpi_insn_t0;
  wire [31:0] pcpi_insn_t0;
  /* src = "generated/out/vanilla.sv:2074.20-2074.27" */
  output [31:0] pcpi_rd;
  reg [31:0] pcpi_rd;
  /* cellift = 32'd1 */
  output [31:0] pcpi_rd_t0;
  reg [31:0] pcpi_rd_t0;
  /* src = "generated/out/vanilla.sv:2076.13-2076.23" */
  output pcpi_ready;
  reg pcpi_ready;
  /* cellift = 32'd1 */
  output pcpi_ready_t0;
  reg pcpi_ready_t0;
  /* src = "generated/out/vanilla.sv:2071.15-2071.23" */
  input [31:0] pcpi_rs1;
  wire [31:0] pcpi_rs1;
  /* cellift = 32'd1 */
  input [31:0] pcpi_rs1_t0;
  wire [31:0] pcpi_rs1_t0;
  /* src = "generated/out/vanilla.sv:2072.15-2072.23" */
  input [31:0] pcpi_rs2;
  wire [31:0] pcpi_rs2;
  /* cellift = 32'd1 */
  input [31:0] pcpi_rs2_t0;
  wire [31:0] pcpi_rs2_t0;
  /* src = "generated/out/vanilla.sv:2069.8-2069.18" */
  input pcpi_valid;
  wire pcpi_valid;
  /* cellift = 32'd1 */
  input pcpi_valid_t0;
  wire pcpi_valid_t0;
  /* src = "generated/out/vanilla.sv:2075.13-2075.22" */
  output pcpi_wait;
  reg pcpi_wait;
  /* src = "generated/out/vanilla.sv:2082.6-2082.17" */
  reg pcpi_wait_q;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2082.6-2082.17" */
  reg pcpi_wait_q_t0;
  /* cellift = 32'd1 */
  output pcpi_wait_t0;
  reg pcpi_wait_t0;
  /* src = "generated/out/vanilla.sv:2073.13-2073.20" */
  output pcpi_wr;
  wire pcpi_wr;
  /* cellift = 32'd1 */
  output pcpi_wr_t0;
  wire pcpi_wr_t0;
  /* src = "generated/out/vanilla.sv:2101.13-2101.21" */
  reg [31:0] quotient;
  /* src = "generated/out/vanilla.sv:2102.13-2102.25" */
  reg [31:0] quotient_msk;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2102.13-2102.25" */
  reg [31:0] quotient_msk_t0;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2101.13-2101.21" */
  reg [31:0] quotient_t0;
  /* src = "generated/out/vanilla.sv:2068.8-2068.14" */
  input resetn;
  wire resetn;
  /* src = "generated/out/vanilla.sv:2103.6-2103.13" */
  reg running;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2103.6-2103.13" */
  reg running_t0;
  /* src = "generated/out/vanilla.sv:2083.7-2083.12" */
  wire start;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2083.7-2083.12" */
  wire start_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME pcpi_rd_t0 */
  always_ff @(posedge clk)
    pcpi_rd_t0 <= _001_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME pcpi_wait_t0 */
  always_ff @(posedge clk)
    pcpi_wait_t0 <= _003_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME pcpi_wait_q_t0 */
  always_ff @(posedge clk)
    pcpi_wait_q_t0 <= _005_;
  assign _250_ = _303_ ^ outsign;
  assign _253_ = _343_ ^ dividend;
  assign _256_ = _337_[62:31] ^ divisor[62:31];
  assign _006_ = ~ _075_;
  assign _007_ = ~ _079_;
  assign _008_ = ~ _077_;
  assign _174_ = _304_ | outsign_t0;
  assign _186_ = _344_ | dividend_t0;
  assign _198_ = _338_[62:31] | divisor_t0[62:31];
  assign _175_ = _250_ | _174_;
  assign _187_ = _253_ | _186_;
  assign _199_ = _256_ | _198_;
  assign _082_ = _075_ & _304_;
  assign _091_ = { _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_ } & _344_;
  assign _100_ = { _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_ } & _338_[62:31];
  assign _083_ = _006_ & outsign_t0;
  assign _092_ = { _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_ } & dividend_t0;
  assign _101_ = { _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_ } & divisor_t0[62:31];
  assign _084_ = _175_ & _076_;
  assign _093_ = _187_ & { _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_ };
  assign _102_ = _199_ & { _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_ };
  assign _176_ = _082_ | _083_;
  assign _188_ = _091_ | _092_;
  assign _200_ = _100_ | _101_;
  assign _177_ = _176_ | _084_;
  assign _189_ = _188_ | _093_;
  assign _201_ = _200_ | _102_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME outsign_t0 */
  always_ff @(posedge clk)
    outsign_t0 <= _177_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME dividend_t0 */
  always_ff @(posedge clk)
    dividend_t0 <= _189_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME divisor_t0[62:31] */
  always_ff @(posedge clk)
    divisor_t0[62:31] <= _201_;
  assign _010_ = | { pcpi_rs2_t0[31], pcpi_rs1_t0[31] };
  assign _011_ = | pcpi_insn_t0[14:12];
  assign _218_ = pcpi_rs1_t0[31] | pcpi_rs2_t0[31];
  assign _013_ = ~ _218_;
  assign _014_ = ~ pcpi_insn_t0[14:12];
  assign _139_ = pcpi_rs1[31] & _013_;
  assign _157_ = pcpi_insn[14:12] & _014_;
  assign _140_ = pcpi_rs2[31] & _013_;
  assign _269_ = _103_ == { _012_[1], 1'h0 };
  assign _270_ = _139_ == _140_;
  assign _271_ = _157_ == _014_;
  assign _272_ = _157_ == { _014_[2:1], 1'h0 };
  assign _273_ = _157_ == { _014_[2], 1'h0, _014_[0] };
  assign _274_ = _157_ == { _014_[2], 2'h0 };
  assign _072_ = _269_ & _009_;
  assign _308_ = _270_ & _010_;
  assign _346_ = _271_ & _011_;
  assign _349_ = _272_ & _011_;
  assign _352_ = _273_ & _011_;
  assign _355_ = _274_ & _011_;
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME instr_div */
  always_ff @(posedge clk)
    if (!_284_) instr_div <= 1'h0;
    else instr_div <= _354_;
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME instr_divu */
  always_ff @(posedge clk)
    if (!_284_) instr_divu <= 1'h0;
    else instr_divu <= _351_;
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME instr_remu */
  always_ff @(posedge clk)
    if (!_284_) instr_remu <= 1'h0;
    else instr_remu <= _345_;
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME instr_rem */
  always_ff @(posedge clk)
    if (!_284_) instr_rem <= 1'h0;
    else instr_rem <= _348_;
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME outsign */
  always_ff @(posedge clk)
    if (_075_) outsign <= _303_;
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME running */
  always_ff @(posedge clk)
    if (!resetn) running <= 1'h0;
    else if (_069_) running <= _327_;
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME quotient_msk */
  always_ff @(posedge clk)
    if (_077_)
      if (start) quotient_msk <= 32'd2147483648;
      else quotient_msk <= _329_;
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME pcpi_ready */
  always_ff @(posedge clk)
    if (_081_) pcpi_ready <= 1'h0;
    else pcpi_ready <= _325_;
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME dividend */
  always_ff @(posedge clk)
    if (_079_) dividend <= _343_;
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME quotient */
  always_ff @(posedge clk)
    if (_079_)
      if (start) quotient <= 32'd0;
      else quotient <= _333_;
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME divisor[30:0] */
  always_ff @(posedge clk)
    if (_077_)
      if (start) divisor[30:0] <= 31'h00000000;
      else divisor[30:0] <= _335_[30:0];
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME divisor[62:31] */
  always_ff @(posedge clk)
    if (_077_) divisor[62:31] <= _337_[62:31];
  assign _067_ = { _105_, _106_ } <= { 1'h0, _207_ };
  assign _068_ = { _205_, _206_ } <= { 1'h0, _107_ };
  assign _280_ = _067_ ^ _068_;
  assign _015_ = ~ divisor_t0[61:0];
  assign _016_ = ~ divisor_t0[62];
  assign _017_ = ~ { 30'h00000000, dividend_t0 };
  assign _105_ = divisor[62] & _016_;
  assign _205_ = divisor[62] | divisor_t0[62];
  assign _106_ = divisor[61:0] & _015_;
  assign _107_ = { 30'h00000000, dividend } & _017_;
  assign _206_ = divisor[61:0] | divisor_t0[61:0];
  assign _207_ = { 30'h00000000, dividend } | { 30'h00000000, dividend_t0 };
  assign _108_ = pcpi_wait_t0 & _297_;
  assign _003_ = instr_any_div_rem_t0 & resetn;
  assign _005_ = pcpi_wait_t0 & resetn;
  assign _111_ = _302_ & pcpi_rs1[31];
  assign _114_ = _302_ & pcpi_rs2[31];
  assign _117_ = instr_div_t0 & _307_;
  assign _120_ = _290_ & _357_;
  assign _123_ = instr_rem_t0 & pcpi_rs1[31];
  assign _126_ = _300_ & running;
  assign _109_ = pcpi_wait_q_t0 & pcpi_wait;
  assign _112_ = pcpi_rs1_t0[31] & _301_;
  assign _115_ = pcpi_rs2_t0[31] & _301_;
  assign _118_ = _308_ & instr_div;
  assign _121_ = _358_ & _289_;
  assign _124_ = pcpi_rs1_t0[31] & instr_rem;
  assign _127_ = running_t0 & _299_;
  assign _110_ = pcpi_wait_t0 & pcpi_wait_q_t0;
  assign _113_ = _302_ & pcpi_rs1_t0[31];
  assign _116_ = _302_ & pcpi_rs2_t0[31];
  assign _119_ = instr_div_t0 & _308_;
  assign _122_ = _290_ & _358_;
  assign _125_ = instr_rem_t0 & pcpi_rs1_t0[31];
  assign _128_ = _300_ & running_t0;
  assign _208_ = _108_ | _109_;
  assign _209_ = _111_ | _112_;
  assign _210_ = _114_ | _115_;
  assign _211_ = _117_ | _118_;
  assign _212_ = _120_ | _121_;
  assign _213_ = _123_ | _124_;
  assign _214_ = _126_ | _127_;
  assign start_t0 = _208_ | _110_;
  assign _286_ = _209_ | _113_;
  assign _288_ = _210_ | _116_;
  assign _290_ = _211_ | _119_;
  assign _292_ = _212_ | _122_;
  assign _294_ = _213_ | _125_;
  assign _296_ = _214_ | _128_;
  assign _009_ = | { start_t0, _296_ };
  assign _018_ = | { start_t0, _296_, _280_ };
  assign _019_ = | quotient_msk_t0;
  assign _020_ = | { instr_div_t0, instr_divu_t0, instr_remu_t0, instr_rem_t0 };
  assign _021_ = | pcpi_rs2_t0;
  assign _012_ = ~ { _296_, start_t0 };
  assign _022_ = ~ { _280_, _296_, start_t0 };
  assign _023_ = ~ quotient_msk_t0;
  assign _024_ = ~ { instr_remu_t0, instr_rem_t0, instr_divu_t0, instr_div_t0 };
  assign _025_ = ~ pcpi_rs2_t0;
  assign _103_ = { _295_, start } & _012_;
  assign _104_ = { _279_, _295_, start } & _022_;
  assign _129_ = quotient_msk & _023_;
  assign _158_ = { instr_remu, instr_rem, instr_divu, instr_div } & _024_;
  assign _159_ = pcpi_rs2 & _025_;
  assign _026_ = ! _103_;
  assign _027_ = ! _104_;
  assign _028_ = ! _129_;
  assign _029_ = ! _158_;
  assign _030_ = ! _159_;
  assign _070_ = _026_ & _009_;
  assign _074_ = _027_ & _018_;
  assign _300_ = _028_ & _019_;
  assign instr_any_div_rem_t0 = _029_ & _020_;
  assign _358_ = _030_ & _021_;
  assign _031_ = ~ instr_div;
  assign _032_ = ~ _291_;
  assign _033_ = ~ instr_rem;
  assign _034_ = ~ _293_;
  assign _035_ = ~ instr_divu;
  assign _130_ = instr_div_t0 & _033_;
  assign _133_ = _292_ & _034_;
  assign _136_ = instr_div_t0 & _035_;
  assign _131_ = instr_rem_t0 & _031_;
  assign _134_ = _294_ & _032_;
  assign _137_ = instr_divu_t0 & _031_;
  assign _132_ = instr_div_t0 & instr_rem_t0;
  assign _135_ = _292_ & _294_;
  assign _138_ = instr_div_t0 & instr_divu_t0;
  assign _215_ = _130_ | _131_;
  assign _216_ = _133_ | _134_;
  assign _217_ = _136_ | _137_;
  assign _302_ = _215_ | _132_;
  assign _304_ = _216_ | _135_;
  assign _306_ = _217_ | _138_;
  assign _036_ = ~ { _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_ };
  assign _037_ = ~ { _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_ };
  assign _038_ = ~ { start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start };
  assign _039_ = ~ { _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_ };
  assign _040_ = ~ { start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start };
  assign _041_ = ~ { _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_ };
  assign _042_ = ~ { _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_ };
  assign _043_ = ~ { outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign };
  assign _224_ = { _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_ } | _036_;
  assign _227_ = { _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_ } | _037_;
  assign _229_ = { start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0 } | _038_;
  assign _232_ = { _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_ } | _039_;
  assign _233_ = { start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0 } | _040_;
  assign _240_ = { _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_ } | _041_;
  assign _243_ = { _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_ } | _042_;
  assign _246_ = { outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0 } | _043_;
  assign _225_ = { _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_ } | { _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_ };
  assign _228_ = { _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_, _296_ } | { _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_, _295_ };
  assign _230_ = { start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0 } | { start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start };
  assign _231_ = { _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_ } | { _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_ };
  assign _234_ = { start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0 } | { start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start };
  assign _241_ = { _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_ } | { _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_ };
  assign _244_ = { _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_ } | { _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_, _287_ };
  assign _247_ = { outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0 } | { outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign };
  assign _148_ = _370_ & _224_;
  assign _324_ = _322_ & _229_;
  assign _330_ = { 1'h0, quotient_msk_t0[31:1] } & _227_;
  assign _334_ = _332_ & _227_;
  assign _336_ = { 1'h0, divisor_t0[62:1] } & _232_;
  assign _151_ = _336_ & _233_;
  assign _342_ = _340_ & _227_;
  assign _154_ = _342_ & _229_;
  assign _162_ = pcpi_rs1_t0 & _240_;
  assign _165_ = { 31'h00000000, pcpi_rs2_t0 } & _243_;
  assign _168_ = quotient_t0 & _246_;
  assign _171_ = dividend_t0 & _246_;
  assign _149_ = _368_ & _225_;
  assign _322_ = _320_ & _228_;
  assign _001_ = _324_ & { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn };
  assign _332_ = _318_ & _231_;
  assign _152_ = { _360_[62:31], 31'h00000000 } & _234_;
  assign _340_ = _362_[31:0] & _231_;
  assign _155_ = _364_ & _230_;
  assign _163_ = _310_ & _241_;
  assign _166_ = _312_ & _244_;
  assign _169_ = _314_ & _247_;
  assign _172_ = _316_ & _247_;
  assign _226_ = _148_ | _149_;
  assign _235_ = _151_ | _152_;
  assign _236_ = _154_ | _155_;
  assign _242_ = _162_ | _163_;
  assign _245_ = _165_ | _166_;
  assign _248_ = _168_ | _169_;
  assign _249_ = _171_ | _172_;
  assign _261_ = _369_ ^ _367_;
  assign _262_ = _335_ ^ { _359_[62:31], 31'h00000000 };
  assign _263_ = _341_ ^ _363_;
  assign _265_ = pcpi_rs1 ^ _309_;
  assign _266_ = { 31'h00000000, pcpi_rs2 } ^ _311_;
  assign _267_ = quotient ^ _313_;
  assign _268_ = dividend ^ _315_;
  assign _150_ = { _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_ } & _261_;
  assign _328_ = start_t0 & _057_;
  assign _153_ = { start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0 } & _262_;
  assign _156_ = { start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0, start_t0 } & _263_;
  assign _164_ = { _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_ } & _265_;
  assign _167_ = { _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_ } & _266_;
  assign _170_ = { outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0 } & _267_;
  assign _173_ = { outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0, outsign_t0 } & _268_;
  assign _320_ = _150_ | _226_;
  assign _338_ = _153_ | _235_;
  assign _344_ = _156_ | _236_;
  assign _364_ = _164_ | _242_;
  assign { _366_[62:32], _360_[62:31] } = _167_ | _245_;
  assign _368_ = _170_ | _248_;
  assign _370_ = _173_ | _249_;
  assign _044_ = ~ pcpi_rs1_t0;
  assign _045_ = ~ { 31'h00000000, pcpi_rs2_t0 };
  assign _046_ = ~ quotient_t0;
  assign _047_ = ~ dividend_t0;
  assign _141_ = pcpi_rs1 & _044_;
  assign _142_ = { 31'h00000000, pcpi_rs2 } & _045_;
  assign _143_ = quotient & _046_;
  assign _144_ = dividend & _047_;
  assign _219_ = pcpi_rs1 | pcpi_rs1_t0;
  assign _220_ = { 31'h00000000, pcpi_rs2 } | { 31'h00000000, pcpi_rs2_t0 };
  assign _221_ = quotient | quotient_t0;
  assign _222_ = dividend | dividend_t0;
  assign _048_ = - _141_;
  assign _049_ = - _142_;
  assign _050_ = - _143_;
  assign _051_ = - _144_;
  assign _052_ = - _219_;
  assign _053_ = - _220_;
  assign _054_ = - _221_;
  assign _055_ = - _222_;
  assign _257_ = _048_ ^ _052_;
  assign _258_ = _049_ ^ _053_;
  assign _259_ = _050_ ^ _054_;
  assign _260_ = _051_ ^ _055_;
  assign _310_ = _257_ | pcpi_rs1_t0;
  assign _312_ = _258_ | { 31'h00000000, pcpi_rs2_t0 };
  assign _314_ = _259_ | quotient_t0;
  assign _316_ = _260_ | dividend_t0;
  assign _069_ = | { _295_, start };
  assign _071_ = { _295_, start } != 2'h2;
  assign _073_ = | { _279_, _295_, start };
  assign _075_ = & { start, resetn };
  assign _077_ = & { _071_, resetn };
  assign _079_ = & { _071_, _073_, resetn };
  assign _056_ = ~ resetn;
  assign _081_ = | { _056_, start };
  assign _057_ = ~ _326_;
  assign _058_ = ~ quotient;
  assign _059_ = ~ quotient_msk;
  assign _145_ = quotient_t0 & _059_;
  assign _146_ = quotient_msk_t0 & _058_;
  assign _147_ = quotient_t0 & quotient_msk_t0;
  assign _223_ = _145_ | _146_;
  assign _318_ = _223_ | _147_;
  assign _060_ = | { _072_, _074_ };
  assign _202_ = { start, resetn } | { start_t0, 1'h0 };
  assign _203_ = { _071_, resetn } | { _072_, 1'h0 };
  assign _204_ = { _071_, _073_, resetn } | { _072_, _074_, 1'h0 };
  assign _061_ = & _202_;
  assign _062_ = & _203_;
  assign _063_ = & _204_;
  assign _076_ = start_t0 & _061_;
  assign _078_ = _072_ & _062_;
  assign _080_ = _060_ & _063_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME instr_div_t0 */
  always_ff @(posedge clk)
    if (!_284_) instr_div_t0 <= 1'h0;
    else instr_div_t0 <= _355_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME instr_divu_t0 */
  always_ff @(posedge clk)
    if (!_284_) instr_divu_t0 <= 1'h0;
    else instr_divu_t0 <= _352_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME instr_remu_t0 */
  always_ff @(posedge clk)
    if (!_284_) instr_remu_t0 <= 1'h0;
    else instr_remu_t0 <= _346_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME instr_rem_t0 */
  always_ff @(posedge clk)
    if (!_284_) instr_rem_t0 <= 1'h0;
    else instr_rem_t0 <= _349_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME pcpi_ready_t0 */
  always_ff @(posedge clk)
    if (_081_) pcpi_ready_t0 <= 1'h0;
    else pcpi_ready_t0 <= _296_;
  assign _252_ = _329_ ^ quotient_msk;
  assign _254_ = _333_ ^ quotient;
  assign _255_ = _335_[30:0] ^ divisor[30:0];
  assign _182_ = _330_ | quotient_msk_t0;
  assign _190_ = _334_ | quotient_t0;
  assign _194_ = _336_[30:0] | divisor_t0[30:0];
  assign _183_ = _252_ | _182_;
  assign _191_ = _254_ | _190_;
  assign _195_ = _255_ | _194_;
  assign _088_ = { _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_ } & _330_;
  assign _094_ = { _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_ } & _334_;
  assign _097_ = { _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_ } & _336_[30:0];
  assign _089_ = { _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_ } & quotient_msk_t0;
  assign _095_ = { _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_, _007_ } & quotient_t0;
  assign _098_ = { _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_, _008_ } & divisor_t0[30:0];
  assign _090_ = _183_ & { _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_ };
  assign _096_ = _191_ & { _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_, _080_ };
  assign _099_ = _195_ & { _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_ };
  assign _184_ = _088_ | _089_;
  assign _192_ = _094_ | _095_;
  assign _196_ = _097_ | _098_;
  assign _185_ = _184_ | _090_;
  assign _193_ = _192_ | _096_;
  assign _197_ = _196_ | _099_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME quotient_msk_t0 */
  always_ff @(posedge clk)
    if (start) quotient_msk_t0 <= 32'd0;
    else quotient_msk_t0 <= _185_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME quotient_t0 */
  always_ff @(posedge clk)
    if (start) quotient_t0 <= 32'd0;
    else quotient_t0 <= _193_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME divisor_t0[30:0] */
  always_ff @(posedge clk)
    if (start) divisor_t0[30:0] <= 31'h00000000;
    else divisor_t0[30:0] <= _197_;
  assign _064_ = ~ _069_;
  assign _251_ = _327_ ^ running;
  assign _178_ = _328_ | running_t0;
  assign _179_ = _251_ | _178_;
  assign _085_ = _069_ & _328_;
  assign _086_ = _064_ & running_t0;
  assign _087_ = _179_ & _070_;
  assign _180_ = _085_ | _086_;
  assign _181_ = _180_ | _087_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME running_t0 */
  always_ff @(posedge clk)
    if (!resetn) running_t0 <= 1'h0;
    else running_t0 <= _181_;
  assign _065_ = ~ { 31'h00000000, dividend_t0 };
  assign _066_ = ~ divisor_t0;
  assign _160_ = { 31'h00000000, dividend } & _065_;
  assign _161_ = divisor & _066_;
  assign _237_ = { 31'h00000000, dividend } | { 31'h00000000, dividend_t0 };
  assign _238_ = divisor | divisor_t0;
  assign _275_ = _237_ - _161_;
  assign _276_ = _160_ - _238_;
  assign _264_ = _275_ ^ _276_;
  assign _239_ = _264_ | { 31'h00000000, dividend_t0 };
  assign _362_ = _239_ | divisor_t0;
  assign _277_ = pcpi_insn[6:0] == /* src = "generated/out/vanilla.sv:2089.52-2089.80" */ 7'h33;
  assign _278_ = pcpi_insn[31:25] == /* src = "generated/out/vanilla.sv:2089.87-2089.117" */ 7'h01;
  assign _279_ = divisor <= /* src = "generated/out/vanilla.sv:2129.8-2129.27" */ dividend;
  assign start = pcpi_wait && /* src = "generated/out/vanilla.sv:2083.15-2083.40" */ _297_;
  assign _281_ = resetn && /* src = "generated/out/vanilla.sv:2089.10-2089.30" */ pcpi_valid;
  assign _282_ = _281_ && /* src = "generated/out/vanilla.sv:2089.9-2089.46" */ _298_;
  assign _283_ = _282_ && /* src = "generated/out/vanilla.sv:2089.8-2089.81" */ _277_;
  assign _284_ = _283_ && /* src = "generated/out/vanilla.sv:2089.7-2089.118" */ _278_;
  assign _002_ = instr_any_div_rem && /* src = "generated/out/vanilla.sv:2096.16-2096.43" */ resetn;
  assign _004_ = pcpi_wait && /* src = "generated/out/vanilla.sv:2097.18-2097.37" */ resetn;
  assign _285_ = _301_ && /* src = "generated/out/vanilla.sv:2113.17-2113.57" */ pcpi_rs1[31];
  assign _287_ = _301_ && /* src = "generated/out/vanilla.sv:2114.16-2114.56" */ pcpi_rs2[31];
  assign _289_ = instr_div && /* src = "generated/out/vanilla.sv:2115.17-2115.60" */ _307_;
  assign _291_ = _289_ && /* src = "generated/out/vanilla.sv:2115.16-2115.74" */ _357_;
  assign _293_ = instr_rem && /* src = "generated/out/vanilla.sv:2115.80-2115.105" */ pcpi_rs1[31];
  assign _295_ = _299_ && /* src = "generated/out/vanilla.sv:2119.12-2119.36" */ running;
  assign _297_ = ! /* src = "generated/out/vanilla.sv:2083.28-2083.40" */ pcpi_wait_q;
  assign _298_ = ! /* src = "generated/out/vanilla.sv:2089.35-2089.46" */ pcpi_ready;
  assign _299_ = ! /* src = "generated/out/vanilla.sv:2119.12-2119.25" */ quotient_msk;
  assign _301_ = instr_div || /* src = "generated/out/vanilla.sv:2114.17-2114.39" */ instr_rem;
  assign _303_ = _291_ || /* src = "generated/out/vanilla.sv:2115.15-2115.106" */ _293_;
  assign _305_ = instr_div || /* src = "generated/out/vanilla.sv:2123.8-2123.31" */ instr_divu;
  assign _307_ = pcpi_rs1[31] != /* src = "generated/out/vanilla.sv:2115.31-2115.59" */ pcpi_rs2[31];
  assign _309_ = - /* src = "generated/out/vanilla.sv:2113.60-2113.69" */ pcpi_rs1;
  assign _311_ = - /* src = "generated/out/vanilla.sv:2114.59-2114.68" */ { 31'h00000000, pcpi_rs2 };
  assign _313_ = - /* src = "generated/out/vanilla.sv:2124.27-2124.36" */ quotient;
  assign _315_ = - /* src = "generated/out/vanilla.sv:2126.27-2126.36" */ dividend;
  assign _317_ = quotient | /* src = "generated/out/vanilla.sv:2131.17-2131.40" */ quotient_msk;
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME pcpi_rd */
  always_ff @(posedge clk)
    pcpi_rd <= _000_;
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME pcpi_wait */
  always_ff @(posedge clk)
    pcpi_wait <= _002_;
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME pcpi_wait_q */
  always_ff @(posedge clk)
    pcpi_wait_q <= _004_;
  assign _319_ = _305_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2123.8-2123.31|generated/out/vanilla.sv:2123.4-2126.49" */ _367_ : _369_;
  assign _321_ = _295_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2119.12-2119.36|generated/out/vanilla.sv:2119.8-2135.6" */ _319_ : 32'hxxxxxxxx;
  assign _323_ = start ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2111.12-2111.17|generated/out/vanilla.sv:2111.8-2135.6" */ 32'hxxxxxxxx : _321_;
  assign _000_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2109.7-2109.14|generated/out/vanilla.sv:2109.3-2135.6" */ _323_ : 32'hxxxxxxxx;
  assign _325_ = _295_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2119.12-2119.36|generated/out/vanilla.sv:2119.8-2135.6" */ 1'h1 : 1'h0;
  assign _326_ = _295_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2119.12-2119.36|generated/out/vanilla.sv:2119.8-2135.6" */ 1'h0 : 1'hx;
  assign _327_ = start ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2111.12-2111.17|generated/out/vanilla.sv:2111.8-2135.6" */ 1'h1 : _326_;
  assign _329_ = _295_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2119.12-2119.36|generated/out/vanilla.sv:2119.8-2135.6" */ 32'hxxxxxxxx : { 1'h0, quotient_msk[31:1] };
  assign _331_ = _279_ ? /* src = "generated/out/vanilla.sv:2129.8-2129.27|generated/out/vanilla.sv:2129.4-2132.7" */ _317_ : 32'hxxxxxxxx;
  assign _333_ = _295_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2119.12-2119.36|generated/out/vanilla.sv:2119.8-2135.6" */ 32'hxxxxxxxx : _331_;
  assign _335_ = _295_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2119.12-2119.36|generated/out/vanilla.sv:2119.8-2135.6" */ 63'hxxxxxxxxxxxxxxxx : { 1'h0, divisor[62:1] };
  assign _337_ = start ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2111.12-2111.17|generated/out/vanilla.sv:2111.8-2135.6" */ { _359_[62:31], 31'h00000000 } : _335_;
  assign _339_ = _279_ ? /* src = "generated/out/vanilla.sv:2129.8-2129.27|generated/out/vanilla.sv:2129.4-2132.7" */ _361_[31:0] : 32'hxxxxxxxx;
  assign _341_ = _295_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2119.12-2119.36|generated/out/vanilla.sv:2119.8-2135.6" */ 32'hxxxxxxxx : _339_;
  assign _343_ = start ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2111.12-2111.17|generated/out/vanilla.sv:2111.8-2135.6" */ _363_ : _341_;
  assign _345_ = _347_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:2090.4-2095.11" */ 1'h1 : 1'h0;
  assign _347_ = pcpi_insn[14:12] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:2090.4-2095.11" */ 3'h7;
  assign _348_ = _350_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:2090.4-2095.11" */ 1'h1 : 1'h0;
  assign _350_ = pcpi_insn[14:12] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:2090.4-2095.11" */ 3'h6;
  assign _351_ = _353_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:2090.4-2095.11" */ 1'h1 : 1'h0;
  assign _353_ = pcpi_insn[14:12] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:2090.4-2095.11" */ 3'h5;
  assign _354_ = _356_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:2090.4-2095.11" */ 1'h1 : 1'h0;
  assign _356_ = pcpi_insn[14:12] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:2090.4-2095.11" */ 3'h4;
  assign instr_any_div_rem = | /* src = "generated/out/vanilla.sv:2081.27-2081.74" */ { instr_remu, instr_rem, instr_divu, instr_div };
  assign _357_ = | /* src = "generated/out/vanilla.sv:2115.65-2115.74" */ pcpi_rs2;
  assign _361_ = dividend - /* src = "generated/out/vanilla.sv:2130.17-2130.35" */ divisor;
  assign _363_ = _285_ ? /* src = "generated/out/vanilla.sv:2113.17-2113.80" */ _309_ : pcpi_rs1;
  assign { _365_[62:32], _359_[62:31] } = _287_ ? /* src = "generated/out/vanilla.sv:2114.16-2114.79" */ _311_ : { 31'h00000000, pcpi_rs2 };
  assign _367_ = outsign ? /* src = "generated/out/vanilla.sv:2124.17-2124.47" */ _313_ : quotient;
  assign _369_ = outsign ? /* src = "generated/out/vanilla.sv:2126.17-2126.47" */ _315_ : dividend;
  assign _359_[30:0] = 31'h00000000;
  assign _360_[30:0] = 31'h00000000;
  assign _365_[31:0] = _359_[62:31];
  assign _366_[31:0] = _360_[62:31];
  assign pcpi_wr = pcpi_ready;
  assign pcpi_wr_t0 = pcpi_ready_t0;
endmodule

/* cellift =  1  */
/* hdlname = "\\picorv32_pcpi_mul" */
/* src = "generated/out/vanilla.sv:1837.1-1963.10" */
module picorv32_pcpi_mul(clk, resetn, pcpi_valid, pcpi_insn, pcpi_rs1, pcpi_rs2, pcpi_wr, pcpi_rd, pcpi_wait, pcpi_ready, pcpi_insn_t0, pcpi_rd_t0, pcpi_ready_t0, pcpi_rs1_t0, pcpi_rs2_t0, pcpi_valid_t0, pcpi_wait_t0, pcpi_wr_t0);
  /* src = "generated/out/vanilla.sv:1954.2-1962.5" */
  wire _0000_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1954.2-1962.5" */
  wire _0001_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0002_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0003_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0004_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0005_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0006_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0007_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0008_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0009_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0010_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0011_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0012_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0013_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0014_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0015_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0016_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0017_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0018_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0019_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0020_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0021_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0022_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0023_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0024_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0025_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0026_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0027_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0028_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0029_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0030_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _0031_;
  wire [4:0] _0032_;
  wire [4:0] _0033_;
  wire [4:0] _0034_;
  wire [4:0] _0035_;
  wire [4:0] _0036_;
  wire [4:0] _0037_;
  wire [4:0] _0038_;
  wire [4:0] _0039_;
  wire [4:0] _0040_;
  wire [4:0] _0041_;
  wire [4:0] _0042_;
  wire [4:0] _0043_;
  wire [4:0] _0044_;
  wire [4:0] _0045_;
  wire [4:0] _0046_;
  wire [4:0] _0047_;
  wire [4:0] _0048_;
  wire [4:0] _0049_;
  wire [4:0] _0050_;
  wire [4:0] _0051_;
  wire [4:0] _0052_;
  wire [4:0] _0053_;
  wire [4:0] _0054_;
  wire [4:0] _0055_;
  wire [4:0] _0056_;
  wire [4:0] _0057_;
  wire [4:0] _0058_;
  wire [4:0] _0059_;
  wire [4:0] _0060_;
  wire [4:0] _0061_;
  wire [4:0] _0062_;
  wire [4:0] _0063_;
  wire [4:0] _0064_;
  wire [4:0] _0065_;
  wire [4:0] _0066_;
  wire [4:0] _0067_;
  wire [4:0] _0068_;
  wire [4:0] _0069_;
  wire [4:0] _0070_;
  wire [4:0] _0071_;
  wire [4:0] _0072_;
  wire [4:0] _0073_;
  wire [4:0] _0074_;
  wire [4:0] _0075_;
  wire [4:0] _0076_;
  wire [4:0] _0077_;
  wire [4:0] _0078_;
  wire [4:0] _0079_;
  wire [4:0] _0080_;
  wire [4:0] _0081_;
  wire [4:0] _0082_;
  wire [4:0] _0083_;
  wire [4:0] _0084_;
  wire [4:0] _0085_;
  wire [4:0] _0086_;
  wire [4:0] _0087_;
  wire [4:0] _0088_;
  wire [4:0] _0089_;
  wire [4:0] _0090_;
  wire [4:0] _0091_;
  wire [4:0] _0092_;
  wire [4:0] _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire [2:0] _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire [3:0] _0101_;
  wire [2:0] _0102_;
  wire [1:0] _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire [6:0] _0109_;
  wire [63:0] _0110_;
  wire [63:0] _0111_;
  wire [63:0] _0112_;
  wire [63:0] _0113_;
  wire [31:0] _0114_;
  wire _0115_;
  wire _0116_;
  wire [4:0] _0117_;
  wire [4:0] _0118_;
  wire [4:0] _0119_;
  wire [4:0] _0120_;
  wire [4:0] _0121_;
  wire [4:0] _0122_;
  wire [4:0] _0123_;
  wire [4:0] _0124_;
  wire [4:0] _0125_;
  wire [4:0] _0126_;
  wire [4:0] _0127_;
  wire [4:0] _0128_;
  wire [4:0] _0129_;
  wire [4:0] _0130_;
  wire [4:0] _0131_;
  wire [4:0] _0132_;
  wire [4:0] _0133_;
  wire [4:0] _0134_;
  wire [4:0] _0135_;
  wire [4:0] _0136_;
  wire [4:0] _0137_;
  wire [4:0] _0138_;
  wire [4:0] _0139_;
  wire [4:0] _0140_;
  wire [4:0] _0141_;
  wire [4:0] _0142_;
  wire [4:0] _0143_;
  wire [4:0] _0144_;
  wire [4:0] _0145_;
  wire [4:0] _0146_;
  wire [4:0] _0147_;
  wire [4:0] _0148_;
  wire [4:0] _0149_;
  wire [4:0] _0150_;
  wire [4:0] _0151_;
  wire [4:0] _0152_;
  wire [4:0] _0153_;
  wire [4:0] _0154_;
  wire [4:0] _0155_;
  wire [4:0] _0156_;
  wire [4:0] _0157_;
  wire [4:0] _0158_;
  wire [4:0] _0159_;
  wire [4:0] _0160_;
  wire [4:0] _0161_;
  wire [4:0] _0162_;
  wire [4:0] _0163_;
  wire [4:0] _0164_;
  wire [4:0] _0165_;
  wire [4:0] _0166_;
  wire [4:0] _0167_;
  wire [4:0] _0168_;
  wire [4:0] _0169_;
  wire [4:0] _0170_;
  wire [4:0] _0171_;
  wire [4:0] _0172_;
  wire [4:0] _0173_;
  wire [4:0] _0174_;
  wire [4:0] _0175_;
  wire [4:0] _0176_;
  wire [4:0] _0177_;
  wire [4:0] _0178_;
  wire [6:0] _0179_;
  wire [6:0] _0180_;
  wire [31:0] _0181_;
  wire [31:0] _0182_;
  wire [31:0] _0183_;
  wire [63:0] _0184_;
  wire [63:0] _0185_;
  wire _0186_;
  wire _0187_;
  wire [62:0] _0188_;
  wire [62:0] _0189_;
  wire _0190_;
  wire _0191_;
  wire [62:0] _0192_;
  wire [62:0] _0193_;
  wire [14:0] _0194_;
  wire [14:0] _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire [6:0] _0202_;
  wire [6:0] _0203_;
  wire [6:0] _0204_;
  wire [63:0] _0205_;
  wire [63:0] _0206_;
  wire [63:0] _0207_;
  wire [63:0] _0208_;
  wire [63:0] _0209_;
  wire [63:0] _0210_;
  wire [63:0] _0211_;
  wire [63:0] _0212_;
  wire [63:0] _0213_;
  wire [63:0] _0214_;
  wire [63:0] _0215_;
  wire [63:0] _0216_;
  wire [2:0] _0217_;
  wire [3:0] _0218_;
  wire [2:0] _0219_;
  wire [1:0] _0220_;
  wire [31:0] _0221_;
  wire [63:0] _0222_;
  wire [63:0] _0223_;
  wire [63:0] _0224_;
  wire [63:0] _0225_;
  wire [63:0] _0226_;
  wire [4:0] _0227_;
  wire [4:0] _0228_;
  wire [4:0] _0229_;
  wire [4:0] _0230_;
  wire [4:0] _0231_;
  wire [4:0] _0232_;
  wire [4:0] _0233_;
  wire [4:0] _0234_;
  wire [4:0] _0235_;
  wire [4:0] _0236_;
  wire [4:0] _0237_;
  wire [4:0] _0238_;
  wire [4:0] _0239_;
  wire [4:0] _0240_;
  wire [4:0] _0241_;
  wire [4:0] _0242_;
  wire [4:0] _0243_;
  wire [4:0] _0244_;
  wire [4:0] _0245_;
  wire [4:0] _0246_;
  wire [4:0] _0247_;
  wire [4:0] _0248_;
  wire [4:0] _0249_;
  wire [4:0] _0250_;
  wire [4:0] _0251_;
  wire [4:0] _0252_;
  wire [4:0] _0253_;
  wire [4:0] _0254_;
  wire [4:0] _0255_;
  wire [4:0] _0256_;
  wire [4:0] _0257_;
  wire [4:0] _0258_;
  wire [4:0] _0259_;
  wire [4:0] _0260_;
  wire [4:0] _0261_;
  wire [4:0] _0262_;
  wire [4:0] _0263_;
  wire [4:0] _0264_;
  wire [4:0] _0265_;
  wire [4:0] _0266_;
  wire [4:0] _0267_;
  wire [4:0] _0268_;
  wire [4:0] _0269_;
  wire [4:0] _0270_;
  wire [4:0] _0271_;
  wire [4:0] _0272_;
  wire [4:0] _0273_;
  wire [4:0] _0274_;
  wire [4:0] _0275_;
  wire [4:0] _0276_;
  wire [4:0] _0277_;
  wire [4:0] _0278_;
  wire [4:0] _0279_;
  wire [4:0] _0280_;
  wire [4:0] _0281_;
  wire [4:0] _0282_;
  wire [4:0] _0283_;
  wire [4:0] _0284_;
  wire [4:0] _0285_;
  wire [4:0] _0286_;
  wire [4:0] _0287_;
  wire [4:0] _0288_;
  wire [4:0] _0289_;
  wire [4:0] _0290_;
  wire [4:0] _0291_;
  wire [4:0] _0292_;
  wire [4:0] _0293_;
  wire [4:0] _0294_;
  wire [4:0] _0295_;
  wire [4:0] _0296_;
  wire [4:0] _0297_;
  wire [4:0] _0298_;
  wire [4:0] _0299_;
  wire [4:0] _0300_;
  wire [4:0] _0301_;
  wire [4:0] _0302_;
  wire [4:0] _0303_;
  wire [4:0] _0304_;
  wire [4:0] _0305_;
  wire [4:0] _0306_;
  wire [4:0] _0307_;
  wire [4:0] _0308_;
  wire [4:0] _0309_;
  wire [4:0] _0310_;
  wire [4:0] _0311_;
  wire [4:0] _0312_;
  wire [4:0] _0313_;
  wire [4:0] _0314_;
  wire [4:0] _0315_;
  wire [4:0] _0316_;
  wire [4:0] _0317_;
  wire [4:0] _0318_;
  wire [4:0] _0319_;
  wire [6:0] _0320_;
  wire [31:0] _0321_;
  wire [31:0] _0322_;
  wire [31:0] _0323_;
  wire [31:0] _0324_;
  wire [63:0] _0325_;
  wire _0326_;
  wire [62:0] _0327_;
  wire _0328_;
  wire [62:0] _0329_;
  wire [14:0] _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire [6:0] _0335_;
  wire [6:0] _0336_;
  wire [6:0] _0337_;
  wire [63:0] _0338_;
  wire [63:0] _0339_;
  wire [63:0] _0340_;
  wire [63:0] _0341_;
  wire [63:0] _0342_;
  wire [63:0] _0343_;
  wire [63:0] _0344_;
  wire [63:0] _0345_;
  wire [63:0] _0346_;
  wire [63:0] _0347_;
  wire [31:0] _0348_;
  wire [63:0] _0349_;
  wire [63:0] _0350_;
  wire [63:0] _0351_;
  wire [63:0] _0352_;
  wire [4:0] _0353_;
  wire [4:0] _0354_;
  wire [4:0] _0355_;
  wire [4:0] _0356_;
  wire [4:0] _0357_;
  wire [4:0] _0358_;
  wire [4:0] _0359_;
  wire [4:0] _0360_;
  wire [4:0] _0361_;
  wire [4:0] _0362_;
  wire [4:0] _0363_;
  wire [4:0] _0364_;
  wire [4:0] _0365_;
  wire [4:0] _0366_;
  wire [4:0] _0367_;
  wire [4:0] _0368_;
  wire [4:0] _0369_;
  wire [4:0] _0370_;
  wire [4:0] _0371_;
  wire [4:0] _0372_;
  wire [4:0] _0373_;
  wire [4:0] _0374_;
  wire [4:0] _0375_;
  wire [4:0] _0376_;
  wire [4:0] _0377_;
  wire [4:0] _0378_;
  wire [4:0] _0379_;
  wire [4:0] _0380_;
  wire [4:0] _0381_;
  wire [4:0] _0382_;
  wire [4:0] _0383_;
  wire [31:0] _0384_;
  wire _0385_;
  wire [6:0] _0386_;
  wire [63:0] _0387_;
  wire [63:0] _0388_;
  wire [63:0] _0389_;
  wire [63:0] _0390_;
  wire [31:0] _0391_;
  wire [63:0] _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire [4:0] _0396_;
  wire [4:0] _0397_;
  wire [4:0] _0398_;
  wire [4:0] _0399_;
  wire [4:0] _0400_;
  wire [4:0] _0401_;
  wire [4:0] _0402_;
  wire [4:0] _0403_;
  wire [4:0] _0404_;
  wire [4:0] _0405_;
  wire [4:0] _0406_;
  wire [4:0] _0407_;
  wire [4:0] _0408_;
  wire [4:0] _0409_;
  wire [4:0] _0410_;
  wire [4:0] _0411_;
  wire [4:0] _0412_;
  wire [4:0] _0413_;
  wire [4:0] _0414_;
  wire [4:0] _0415_;
  wire [4:0] _0416_;
  wire [4:0] _0417_;
  wire [4:0] _0418_;
  wire [4:0] _0419_;
  wire [4:0] _0420_;
  wire [4:0] _0421_;
  wire [4:0] _0422_;
  wire [4:0] _0423_;
  wire [4:0] _0424_;
  wire [4:0] _0425_;
  wire [4:0] _0426_;
  wire [4:0] _0427_;
  wire [4:0] _0428_;
  wire [4:0] _0429_;
  wire [4:0] _0430_;
  wire [4:0] _0431_;
  wire [4:0] _0432_;
  wire [4:0] _0433_;
  wire [4:0] _0434_;
  wire [4:0] _0435_;
  wire [4:0] _0436_;
  wire [4:0] _0437_;
  wire [4:0] _0438_;
  wire [4:0] _0439_;
  wire [4:0] _0440_;
  wire [4:0] _0441_;
  wire [4:0] _0442_;
  wire [4:0] _0443_;
  wire [4:0] _0444_;
  wire [4:0] _0445_;
  wire [4:0] _0446_;
  wire [4:0] _0447_;
  wire [4:0] _0448_;
  wire [4:0] _0449_;
  wire [4:0] _0450_;
  wire [4:0] _0451_;
  wire [4:0] _0452_;
  wire [4:0] _0453_;
  wire [4:0] _0454_;
  wire [4:0] _0455_;
  wire [4:0] _0456_;
  wire [4:0] _0457_;
  wire [31:0] _0458_;
  wire [31:0] _0459_;
  /* src = "generated/out/vanilla.sv:1876.35-1876.63" */
  wire _0460_;
  /* src = "generated/out/vanilla.sv:1876.70-1876.100" */
  wire _0461_;
  /* src = "generated/out/vanilla.sv:1876.9-1876.29" */
  wire _0462_;
  /* src = "generated/out/vanilla.sv:1876.8-1876.64" */
  wire _0463_;
  /* src = "generated/out/vanilla.sv:1876.7-1876.101" */
  wire _0464_;
  /* src = "generated/out/vanilla.sv:1957.7-1957.27" */
  wire _0465_;
  /* src = "generated/out/vanilla.sv:1870.32-1870.44" */
  wire _0466_;
  /* src = "generated/out/vanilla.sv:1940.19-1940.29" */
  wire _0467_;
  wire _0468_;
  wire _0469_;
  /* cellift = 32'd1 */
  wire _0470_;
  wire [6:0] _0471_;
  /* cellift = 32'd1 */
  wire [6:0] _0472_;
  wire [63:0] _0473_;
  /* cellift = 32'd1 */
  wire [63:0] _0474_;
  /* unused_bits = "0" */
  wire [63:0] _0475_;
  /* cellift = 32'd1 */
  /* unused_bits = "0" */
  wire [63:0] _0476_;
  wire [63:0] _0477_;
  /* cellift = 32'd1 */
  wire [63:0] _0478_;
  /* unused_bits = "63" */
  wire [63:0] _0479_;
  /* cellift = 32'd1 */
  /* unused_bits = "63" */
  wire [63:0] _0480_;
  wire _0481_;
  /* cellift = 32'd1 */
  wire _0482_;
  wire _0483_;
  wire _0484_;
  /* cellift = 32'd1 */
  wire _0485_;
  wire _0486_;
  wire _0487_;
  /* cellift = 32'd1 */
  wire _0488_;
  wire _0489_;
  wire _0490_;
  /* cellift = 32'd1 */
  wire _0491_;
  wire _0492_;
  /* src = "generated/out/vanilla.sv:1947.19-1947.46" */
  /* unused_bits = "7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _0493_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1947.19-1947.46" */
  /* unused_bits = "7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _0494_;
  /* src = "generated/out/vanilla.sv:1939.20-1939.76" */
  /* unused_bits = "7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _0495_;
  /* src = "generated/out/vanilla.sv:1960.16-1960.46" */
  /* unused_bits = "32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63" */
  wire [63:0] _0496_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1960.16-1960.46" */
  /* unused_bits = "32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63" */
  wire [63:0] _0497_;
  /* src = "generated/out/vanilla.sv:1851.8-1851.11" */
  input clk;
  wire clk;
  /* src = "generated/out/vanilla.sv:1865.7-1865.20" */
  wire instr_any_mul;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1865.7-1865.20" */
  wire instr_any_mul_t0;
  /* src = "generated/out/vanilla.sv:1866.7-1866.21" */
  wire instr_any_mulh;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1866.7-1866.21" */
  wire instr_any_mulh_t0;
  /* src = "generated/out/vanilla.sv:1861.6-1861.15" */
  reg instr_mul;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1861.6-1861.15" */
  reg instr_mul_t0;
  /* src = "generated/out/vanilla.sv:1862.6-1862.16" */
  reg instr_mulh;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1862.6-1862.16" */
  reg instr_mulh_t0;
  /* src = "generated/out/vanilla.sv:1863.6-1863.18" */
  reg instr_mulhsu;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1863.6-1863.18" */
  reg instr_mulhsu_t0;
  /* src = "generated/out/vanilla.sv:1864.6-1864.17" */
  reg instr_mulhu;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1864.6-1864.17" */
  reg instr_mulhu_t0;
  /* src = "generated/out/vanilla.sv:1867.7-1867.23" */
  wire instr_rs1_signed;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1867.7-1867.23" */
  wire instr_rs1_signed_t0;
  /* src = "generated/out/vanilla.sv:1896.12-1896.23" */
  reg [6:0] mul_counter;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1896.12-1896.23" */
  reg [6:0] mul_counter_t0;
  /* src = "generated/out/vanilla.sv:1898.6-1898.16" */
  reg mul_finish;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1898.6-1898.16" */
  reg mul_finish_t0;
  /* src = "generated/out/vanilla.sv:1870.7-1870.16" */
  wire mul_start;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1870.7-1870.16" */
  wire mul_start_t0;
  /* src = "generated/out/vanilla.sv:1897.6-1897.17" */
  reg mul_waiting;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1897.6-1897.17" */
  reg mul_waiting_t0;
  /* src = "generated/out/vanilla.sv:1893.13-1893.20" */
  wire [63:0] next_rd;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1893.13-1893.20" */
  wire [63:0] next_rd_t0;
  /* src = "generated/out/vanilla.sv:1895.13-1895.21" */
  /* unused_bits = "63" */
  wire [63:0] next_rdt;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1895.13-1895.21" */
  /* unused_bits = "63" */
  wire [63:0] next_rdt_t0;
  /* src = "generated/out/vanilla.sv:1854.15-1854.24" */
  input [31:0] pcpi_insn;
  wire [31:0] pcpi_insn;
  /* cellift = 32'd1 */
  input [31:0] pcpi_insn_t0;
  wire [31:0] pcpi_insn_t0;
  /* src = "generated/out/vanilla.sv:1858.20-1858.27" */
  output [31:0] pcpi_rd;
  reg [31:0] pcpi_rd;
  /* cellift = 32'd1 */
  output [31:0] pcpi_rd_t0;
  reg [31:0] pcpi_rd_t0;
  /* src = "generated/out/vanilla.sv:1860.13-1860.23" */
  output pcpi_ready;
  reg pcpi_ready;
  /* cellift = 32'd1 */
  output pcpi_ready_t0;
  reg pcpi_ready_t0;
  /* src = "generated/out/vanilla.sv:1855.15-1855.23" */
  input [31:0] pcpi_rs1;
  wire [31:0] pcpi_rs1;
  /* cellift = 32'd1 */
  input [31:0] pcpi_rs1_t0;
  wire [31:0] pcpi_rs1_t0;
  /* src = "generated/out/vanilla.sv:1856.15-1856.23" */
  input [31:0] pcpi_rs2;
  wire [31:0] pcpi_rs2;
  /* cellift = 32'd1 */
  input [31:0] pcpi_rs2_t0;
  wire [31:0] pcpi_rs2_t0;
  /* src = "generated/out/vanilla.sv:1853.8-1853.18" */
  input pcpi_valid;
  wire pcpi_valid;
  /* cellift = 32'd1 */
  input pcpi_valid_t0;
  wire pcpi_valid_t0;
  /* src = "generated/out/vanilla.sv:1859.13-1859.22" */
  output pcpi_wait;
  reg pcpi_wait;
  /* src = "generated/out/vanilla.sv:1869.6-1869.17" */
  reg pcpi_wait_q;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1869.6-1869.17" */
  reg pcpi_wait_q_t0;
  /* cellift = 32'd1 */
  output pcpi_wait_t0;
  reg pcpi_wait_t0;
  /* src = "generated/out/vanilla.sv:1857.13-1857.20" */
  output pcpi_wr;
  wire pcpi_wr;
  /* cellift = 32'd1 */
  output pcpi_wr_t0;
  wire pcpi_wr_t0;
  /* src = "generated/out/vanilla.sv:1888.13-1888.15" */
  reg [63:0] rd;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1888.13-1888.15" */
  reg [63:0] rd_t0;
  /* src = "generated/out/vanilla.sv:1889.13-1889.16" */
  wire [63:0] rdx;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1889.13-1889.16" */
  wire [63:0] rdx_t0;
  /* src = "generated/out/vanilla.sv:1852.8-1852.14" */
  input resetn;
  wire resetn;
  /* src = "generated/out/vanilla.sv:1886.13-1886.16" */
  reg [63:0] rs1;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1886.13-1886.16" */
  reg [63:0] rs1_t0;
  /* src = "generated/out/vanilla.sv:1887.13-1887.16" */
  reg [63:0] rs2;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1887.13-1887.16" */
  reg [63:0] rs2_t0;
  /* src = "generated/out/vanilla.sv:1892.13-1892.21" */
  wire [63:0] this_rs2;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1892.13-1892.21" */
  wire [63:0] this_rs2_t0;
  assign { next_rdt[3], next_rd[3:0] } = { 1'h0, rd[3:0] } + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[3:0];
  assign _0002_ = rd[7:4] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[4] };
  assign { next_rdt[7], next_rd[7:4] } = _0002_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[7:4];
  assign _0004_ = rd[11:8] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[8] };
  assign { next_rdt[11], next_rd[11:8] } = _0004_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[11:8];
  assign _0006_ = rd[15:12] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[12] };
  assign { next_rdt[15], next_rd[15:12] } = _0006_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[15:12];
  assign _0008_ = rd[19:16] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[16] };
  assign { next_rdt[19], next_rd[19:16] } = _0008_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[19:16];
  assign _0010_ = rd[23:20] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[20] };
  assign { next_rdt[23], next_rd[23:20] } = _0010_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[23:20];
  assign _0012_ = rd[27:24] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[24] };
  assign { next_rdt[27], next_rd[27:24] } = _0012_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[27:24];
  assign _0014_ = rd[31:28] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[28] };
  assign { next_rdt[31], next_rd[31:28] } = _0014_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[31:28];
  assign _0016_ = rd[35:32] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[32] };
  assign { next_rdt[35], next_rd[35:32] } = _0016_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[35:32];
  assign _0018_ = rd[39:36] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[36] };
  assign { next_rdt[39], next_rd[39:36] } = _0018_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[39:36];
  assign _0020_ = rd[43:40] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[40] };
  assign { next_rdt[43], next_rd[43:40] } = _0020_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[43:40];
  assign _0022_ = rd[47:44] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[44] };
  assign { next_rdt[47], next_rd[47:44] } = _0022_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[47:44];
  assign _0024_ = rd[51:48] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[48] };
  assign { next_rdt[51], next_rd[51:48] } = _0024_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[51:48];
  assign _0026_ = rd[55:52] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[52] };
  assign { next_rdt[55], next_rd[55:52] } = _0026_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[55:52];
  assign _0028_ = rd[59:56] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[56] };
  assign { next_rdt[59], next_rd[59:56] } = _0028_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[59:56];
  assign _0030_ = rd[63:60] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[60] };
  assign { next_rdt[63], next_rd[63:60] } = _0030_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[63:60];
  assign _0032_ = ~ { 1'h0, rd_t0[3:0] };
  assign _0033_ = ~ { 1'h0, rd_t0[7:4] };
  assign _0034_ = ~ _0003_;
  assign _0035_ = ~ { 1'h0, rd_t0[11:8] };
  assign _0036_ = ~ _0005_;
  assign _0037_ = ~ { 1'h0, rd_t0[15:12] };
  assign _0038_ = ~ _0007_;
  assign _0039_ = ~ { 1'h0, rd_t0[19:16] };
  assign _0040_ = ~ _0009_;
  assign _0041_ = ~ { 1'h0, rd_t0[23:20] };
  assign _0042_ = ~ _0011_;
  assign _0043_ = ~ { 1'h0, rd_t0[27:24] };
  assign _0044_ = ~ _0013_;
  assign _0045_ = ~ { 1'h0, rd_t0[31:28] };
  assign _0046_ = ~ _0015_;
  assign _0047_ = ~ { 1'h0, rd_t0[35:32] };
  assign _0048_ = ~ _0017_;
  assign _0049_ = ~ { 1'h0, rd_t0[39:36] };
  assign _0050_ = ~ _0019_;
  assign _0051_ = ~ { 1'h0, rd_t0[43:40] };
  assign _0052_ = ~ _0021_;
  assign _0053_ = ~ { 1'h0, rd_t0[47:44] };
  assign _0054_ = ~ _0023_;
  assign _0055_ = ~ { 1'h0, rd_t0[51:48] };
  assign _0056_ = ~ _0025_;
  assign _0057_ = ~ { 1'h0, rd_t0[55:52] };
  assign _0058_ = ~ _0027_;
  assign _0059_ = ~ { 1'h0, rd_t0[59:56] };
  assign _0060_ = ~ _0029_;
  assign _0061_ = ~ { 1'h0, rd_t0[63:60] };
  assign _0062_ = ~ _0031_;
  assign _0063_ = ~ { 1'h0, this_rs2_t0[3:0] };
  assign _0064_ = ~ { 4'h0, rdx_t0[4] };
  assign _0065_ = ~ { 1'h0, this_rs2_t0[7:4] };
  assign _0066_ = ~ { 4'h0, rdx_t0[8] };
  assign _0067_ = ~ { 1'h0, this_rs2_t0[11:8] };
  assign _0068_ = ~ { 4'h0, rdx_t0[12] };
  assign _0069_ = ~ { 1'h0, this_rs2_t0[15:12] };
  assign _0070_ = ~ { 4'h0, rdx_t0[16] };
  assign _0071_ = ~ { 1'h0, this_rs2_t0[19:16] };
  assign _0072_ = ~ { 4'h0, rdx_t0[20] };
  assign _0073_ = ~ { 1'h0, this_rs2_t0[23:20] };
  assign _0074_ = ~ { 4'h0, rdx_t0[24] };
  assign _0075_ = ~ { 1'h0, this_rs2_t0[27:24] };
  assign _0076_ = ~ { 4'h0, rdx_t0[28] };
  assign _0077_ = ~ { 1'h0, this_rs2_t0[31:28] };
  assign _0078_ = ~ { 4'h0, rdx_t0[32] };
  assign _0079_ = ~ { 1'h0, this_rs2_t0[35:32] };
  assign _0080_ = ~ { 4'h0, rdx_t0[36] };
  assign _0081_ = ~ { 1'h0, this_rs2_t0[39:36] };
  assign _0082_ = ~ { 4'h0, rdx_t0[40] };
  assign _0083_ = ~ { 1'h0, this_rs2_t0[43:40] };
  assign _0084_ = ~ { 4'h0, rdx_t0[44] };
  assign _0085_ = ~ { 1'h0, this_rs2_t0[47:44] };
  assign _0086_ = ~ { 4'h0, rdx_t0[48] };
  assign _0087_ = ~ { 1'h0, this_rs2_t0[51:48] };
  assign _0088_ = ~ { 4'h0, rdx_t0[52] };
  assign _0089_ = ~ { 1'h0, this_rs2_t0[55:52] };
  assign _0090_ = ~ { 4'h0, rdx_t0[56] };
  assign _0091_ = ~ { 1'h0, this_rs2_t0[59:56] };
  assign _0092_ = ~ { 4'h0, rdx_t0[60] };
  assign _0093_ = ~ { 1'h0, this_rs2_t0[63:60] };
  assign _0117_ = { 1'h0, rd[3:0] } & _0032_;
  assign _0119_ = { 1'h0, rd[7:4] } & _0033_;
  assign _0121_ = _0002_ & _0034_;
  assign _0123_ = { 1'h0, rd[11:8] } & _0035_;
  assign _0125_ = _0004_ & _0036_;
  assign _0127_ = { 1'h0, rd[15:12] } & _0037_;
  assign _0129_ = _0006_ & _0038_;
  assign _0131_ = { 1'h0, rd[19:16] } & _0039_;
  assign _0133_ = _0008_ & _0040_;
  assign _0135_ = { 1'h0, rd[23:20] } & _0041_;
  assign _0137_ = _0010_ & _0042_;
  assign _0139_ = { 1'h0, rd[27:24] } & _0043_;
  assign _0141_ = _0012_ & _0044_;
  assign _0143_ = { 1'h0, rd[31:28] } & _0045_;
  assign _0145_ = _0014_ & _0046_;
  assign _0147_ = { 1'h0, rd[35:32] } & _0047_;
  assign _0149_ = _0016_ & _0048_;
  assign _0151_ = { 1'h0, rd[39:36] } & _0049_;
  assign _0153_ = _0018_ & _0050_;
  assign _0155_ = { 1'h0, rd[43:40] } & _0051_;
  assign _0157_ = _0020_ & _0052_;
  assign _0159_ = { 1'h0, rd[47:44] } & _0053_;
  assign _0161_ = _0022_ & _0054_;
  assign _0163_ = { 1'h0, rd[51:48] } & _0055_;
  assign _0165_ = _0024_ & _0056_;
  assign _0167_ = { 1'h0, rd[55:52] } & _0057_;
  assign _0169_ = _0026_ & _0058_;
  assign _0171_ = { 1'h0, rd[59:56] } & _0059_;
  assign _0173_ = _0028_ & _0060_;
  assign _0175_ = { 1'h0, rd[63:60] } & _0061_;
  assign _0177_ = _0030_ & _0062_;
  assign _0118_ = { 1'h0, this_rs2[3:0] } & _0063_;
  assign _0120_ = { 4'h0, rdx[4] } & _0064_;
  assign _0122_ = { 1'h0, this_rs2[7:4] } & _0065_;
  assign _0124_ = { 4'h0, rdx[8] } & _0066_;
  assign _0126_ = { 1'h0, this_rs2[11:8] } & _0067_;
  assign _0128_ = { 4'h0, rdx[12] } & _0068_;
  assign _0130_ = { 1'h0, this_rs2[15:12] } & _0069_;
  assign _0132_ = { 4'h0, rdx[16] } & _0070_;
  assign _0134_ = { 1'h0, this_rs2[19:16] } & _0071_;
  assign _0136_ = { 4'h0, rdx[20] } & _0072_;
  assign _0138_ = { 1'h0, this_rs2[23:20] } & _0073_;
  assign _0140_ = { 4'h0, rdx[24] } & _0074_;
  assign _0142_ = { 1'h0, this_rs2[27:24] } & _0075_;
  assign _0144_ = { 4'h0, rdx[28] } & _0076_;
  assign _0146_ = { 1'h0, this_rs2[31:28] } & _0077_;
  assign _0148_ = { 4'h0, rdx[32] } & _0078_;
  assign _0150_ = { 1'h0, this_rs2[35:32] } & _0079_;
  assign _0152_ = { 4'h0, rdx[36] } & _0080_;
  assign _0154_ = { 1'h0, this_rs2[39:36] } & _0081_;
  assign _0156_ = { 4'h0, rdx[40] } & _0082_;
  assign _0158_ = { 1'h0, this_rs2[43:40] } & _0083_;
  assign _0160_ = { 4'h0, rdx[44] } & _0084_;
  assign _0162_ = { 1'h0, this_rs2[47:44] } & _0085_;
  assign _0164_ = { 4'h0, rdx[48] } & _0086_;
  assign _0166_ = { 1'h0, this_rs2[51:48] } & _0087_;
  assign _0168_ = { 4'h0, rdx[52] } & _0088_;
  assign _0170_ = { 1'h0, this_rs2[55:52] } & _0089_;
  assign _0172_ = { 4'h0, rdx[56] } & _0090_;
  assign _0174_ = { 1'h0, this_rs2[59:56] } & _0091_;
  assign _0176_ = { 4'h0, rdx[60] } & _0092_;
  assign _0178_ = { 1'h0, this_rs2[63:60] } & _0093_;
  assign _0396_ = _0117_ + _0118_;
  assign _0398_ = _0119_ + _0120_;
  assign _0400_ = _0121_ + _0122_;
  assign _0402_ = _0123_ + _0124_;
  assign _0404_ = _0125_ + _0126_;
  assign _0406_ = _0127_ + _0128_;
  assign _0408_ = _0129_ + _0130_;
  assign _0410_ = _0131_ + _0132_;
  assign _0412_ = _0133_ + _0134_;
  assign _0414_ = _0135_ + _0136_;
  assign _0416_ = _0137_ + _0138_;
  assign _0418_ = _0139_ + _0140_;
  assign _0420_ = _0141_ + _0142_;
  assign _0422_ = _0143_ + _0144_;
  assign _0424_ = _0145_ + _0146_;
  assign _0426_ = _0147_ + _0148_;
  assign _0428_ = _0149_ + _0150_;
  assign _0430_ = _0151_ + _0152_;
  assign _0432_ = _0153_ + _0154_;
  assign _0434_ = _0155_ + _0156_;
  assign _0436_ = _0157_ + _0158_;
  assign _0438_ = _0159_ + _0160_;
  assign _0440_ = _0161_ + _0162_;
  assign _0442_ = _0163_ + _0164_;
  assign _0444_ = _0165_ + _0166_;
  assign _0446_ = _0167_ + _0168_;
  assign _0448_ = _0169_ + _0170_;
  assign _0450_ = _0171_ + _0172_;
  assign _0452_ = _0173_ + _0174_;
  assign _0454_ = _0175_ + _0176_;
  assign _0456_ = _0177_ + _0178_;
  assign _0227_ = { 1'h0, rd[3:0] } | { 1'h0, rd_t0[3:0] };
  assign _0230_ = { 1'h0, rd[7:4] } | { 1'h0, rd_t0[7:4] };
  assign _0233_ = _0002_ | _0003_;
  assign _0236_ = { 1'h0, rd[11:8] } | { 1'h0, rd_t0[11:8] };
  assign _0239_ = _0004_ | _0005_;
  assign _0242_ = { 1'h0, rd[15:12] } | { 1'h0, rd_t0[15:12] };
  assign _0245_ = _0006_ | _0007_;
  assign _0248_ = { 1'h0, rd[19:16] } | { 1'h0, rd_t0[19:16] };
  assign _0251_ = _0008_ | _0009_;
  assign _0254_ = { 1'h0, rd[23:20] } | { 1'h0, rd_t0[23:20] };
  assign _0257_ = _0010_ | _0011_;
  assign _0260_ = { 1'h0, rd[27:24] } | { 1'h0, rd_t0[27:24] };
  assign _0263_ = _0012_ | _0013_;
  assign _0266_ = { 1'h0, rd[31:28] } | { 1'h0, rd_t0[31:28] };
  assign _0269_ = _0014_ | _0015_;
  assign _0272_ = { 1'h0, rd[35:32] } | { 1'h0, rd_t0[35:32] };
  assign _0275_ = _0016_ | _0017_;
  assign _0278_ = { 1'h0, rd[39:36] } | { 1'h0, rd_t0[39:36] };
  assign _0281_ = _0018_ | _0019_;
  assign _0284_ = { 1'h0, rd[43:40] } | { 1'h0, rd_t0[43:40] };
  assign _0287_ = _0020_ | _0021_;
  assign _0290_ = { 1'h0, rd[47:44] } | { 1'h0, rd_t0[47:44] };
  assign _0293_ = _0022_ | _0023_;
  assign _0296_ = { 1'h0, rd[51:48] } | { 1'h0, rd_t0[51:48] };
  assign _0299_ = _0024_ | _0025_;
  assign _0302_ = { 1'h0, rd[55:52] } | { 1'h0, rd_t0[55:52] };
  assign _0305_ = _0026_ | _0027_;
  assign _0308_ = { 1'h0, rd[59:56] } | { 1'h0, rd_t0[59:56] };
  assign _0311_ = _0028_ | _0029_;
  assign _0314_ = { 1'h0, rd[63:60] } | { 1'h0, rd_t0[63:60] };
  assign _0317_ = _0030_ | _0031_;
  assign _0228_ = { 1'h0, this_rs2[3:0] } | { 1'h0, this_rs2_t0[3:0] };
  assign _0231_ = { 4'h0, rdx[4] } | { 4'h0, rdx_t0[4] };
  assign _0234_ = { 1'h0, this_rs2[7:4] } | { 1'h0, this_rs2_t0[7:4] };
  assign _0237_ = { 4'h0, rdx[8] } | { 4'h0, rdx_t0[8] };
  assign _0240_ = { 1'h0, this_rs2[11:8] } | { 1'h0, this_rs2_t0[11:8] };
  assign _0243_ = { 4'h0, rdx[12] } | { 4'h0, rdx_t0[12] };
  assign _0246_ = { 1'h0, this_rs2[15:12] } | { 1'h0, this_rs2_t0[15:12] };
  assign _0249_ = { 4'h0, rdx[16] } | { 4'h0, rdx_t0[16] };
  assign _0252_ = { 1'h0, this_rs2[19:16] } | { 1'h0, this_rs2_t0[19:16] };
  assign _0255_ = { 4'h0, rdx[20] } | { 4'h0, rdx_t0[20] };
  assign _0258_ = { 1'h0, this_rs2[23:20] } | { 1'h0, this_rs2_t0[23:20] };
  assign _0261_ = { 4'h0, rdx[24] } | { 4'h0, rdx_t0[24] };
  assign _0264_ = { 1'h0, this_rs2[27:24] } | { 1'h0, this_rs2_t0[27:24] };
  assign _0267_ = { 4'h0, rdx[28] } | { 4'h0, rdx_t0[28] };
  assign _0270_ = { 1'h0, this_rs2[31:28] } | { 1'h0, this_rs2_t0[31:28] };
  assign _0273_ = { 4'h0, rdx[32] } | { 4'h0, rdx_t0[32] };
  assign _0276_ = { 1'h0, this_rs2[35:32] } | { 1'h0, this_rs2_t0[35:32] };
  assign _0279_ = { 4'h0, rdx[36] } | { 4'h0, rdx_t0[36] };
  assign _0282_ = { 1'h0, this_rs2[39:36] } | { 1'h0, this_rs2_t0[39:36] };
  assign _0285_ = { 4'h0, rdx[40] } | { 4'h0, rdx_t0[40] };
  assign _0288_ = { 1'h0, this_rs2[43:40] } | { 1'h0, this_rs2_t0[43:40] };
  assign _0291_ = { 4'h0, rdx[44] } | { 4'h0, rdx_t0[44] };
  assign _0294_ = { 1'h0, this_rs2[47:44] } | { 1'h0, this_rs2_t0[47:44] };
  assign _0297_ = { 4'h0, rdx[48] } | { 4'h0, rdx_t0[48] };
  assign _0300_ = { 1'h0, this_rs2[51:48] } | { 1'h0, this_rs2_t0[51:48] };
  assign _0303_ = { 4'h0, rdx[52] } | { 4'h0, rdx_t0[52] };
  assign _0306_ = { 1'h0, this_rs2[55:52] } | { 1'h0, this_rs2_t0[55:52] };
  assign _0309_ = { 4'h0, rdx[56] } | { 4'h0, rdx_t0[56] };
  assign _0312_ = { 1'h0, this_rs2[59:56] } | { 1'h0, this_rs2_t0[59:56] };
  assign _0315_ = { 4'h0, rdx[60] } | { 4'h0, rdx_t0[60] };
  assign _0318_ = { 1'h0, this_rs2[63:60] } | { 1'h0, this_rs2_t0[63:60] };
  assign _0397_ = _0227_ + _0228_;
  assign _0399_ = _0230_ + _0231_;
  assign _0401_ = _0233_ + _0234_;
  assign _0403_ = _0236_ + _0237_;
  assign _0405_ = _0239_ + _0240_;
  assign _0407_ = _0242_ + _0243_;
  assign _0409_ = _0245_ + _0246_;
  assign _0411_ = _0248_ + _0249_;
  assign _0413_ = _0251_ + _0252_;
  assign _0415_ = _0254_ + _0255_;
  assign _0417_ = _0257_ + _0258_;
  assign _0419_ = _0260_ + _0261_;
  assign _0421_ = _0263_ + _0264_;
  assign _0423_ = _0266_ + _0267_;
  assign _0425_ = _0269_ + _0270_;
  assign _0427_ = _0272_ + _0273_;
  assign _0429_ = _0275_ + _0276_;
  assign _0431_ = _0278_ + _0279_;
  assign _0433_ = _0281_ + _0282_;
  assign _0435_ = _0284_ + _0285_;
  assign _0437_ = _0287_ + _0288_;
  assign _0439_ = _0290_ + _0291_;
  assign _0441_ = _0293_ + _0294_;
  assign _0443_ = _0296_ + _0297_;
  assign _0445_ = _0299_ + _0300_;
  assign _0447_ = _0302_ + _0303_;
  assign _0449_ = _0305_ + _0306_;
  assign _0451_ = _0308_ + _0309_;
  assign _0453_ = _0311_ + _0312_;
  assign _0455_ = _0314_ + _0315_;
  assign _0457_ = _0317_ + _0318_;
  assign _0353_ = _0396_ ^ _0397_;
  assign _0354_ = _0398_ ^ _0399_;
  assign _0355_ = _0400_ ^ _0401_;
  assign _0356_ = _0402_ ^ _0403_;
  assign _0357_ = _0404_ ^ _0405_;
  assign _0358_ = _0406_ ^ _0407_;
  assign _0359_ = _0408_ ^ _0409_;
  assign _0360_ = _0410_ ^ _0411_;
  assign _0361_ = _0412_ ^ _0413_;
  assign _0362_ = _0414_ ^ _0415_;
  assign _0363_ = _0416_ ^ _0417_;
  assign _0364_ = _0418_ ^ _0419_;
  assign _0365_ = _0420_ ^ _0421_;
  assign _0366_ = _0422_ ^ _0423_;
  assign _0367_ = _0424_ ^ _0425_;
  assign _0368_ = _0426_ ^ _0427_;
  assign _0369_ = _0428_ ^ _0429_;
  assign _0370_ = _0430_ ^ _0431_;
  assign _0371_ = _0432_ ^ _0433_;
  assign _0372_ = _0434_ ^ _0435_;
  assign _0373_ = _0436_ ^ _0437_;
  assign _0374_ = _0438_ ^ _0439_;
  assign _0375_ = _0440_ ^ _0441_;
  assign _0376_ = _0442_ ^ _0443_;
  assign _0377_ = _0444_ ^ _0445_;
  assign _0378_ = _0446_ ^ _0447_;
  assign _0379_ = _0448_ ^ _0449_;
  assign _0380_ = _0450_ ^ _0451_;
  assign _0381_ = _0452_ ^ _0453_;
  assign _0382_ = _0454_ ^ _0455_;
  assign _0383_ = _0456_ ^ _0457_;
  assign _0229_ = _0353_ | { 1'h0, rd_t0[3:0] };
  assign _0232_ = _0354_ | { 1'h0, rd_t0[7:4] };
  assign _0235_ = _0355_ | _0003_;
  assign _0238_ = _0356_ | { 1'h0, rd_t0[11:8] };
  assign _0241_ = _0357_ | _0005_;
  assign _0244_ = _0358_ | { 1'h0, rd_t0[15:12] };
  assign _0247_ = _0359_ | _0007_;
  assign _0250_ = _0360_ | { 1'h0, rd_t0[19:16] };
  assign _0253_ = _0361_ | _0009_;
  assign _0256_ = _0362_ | { 1'h0, rd_t0[23:20] };
  assign _0259_ = _0363_ | _0011_;
  assign _0262_ = _0364_ | { 1'h0, rd_t0[27:24] };
  assign _0265_ = _0365_ | _0013_;
  assign _0268_ = _0366_ | { 1'h0, rd_t0[31:28] };
  assign _0271_ = _0367_ | _0015_;
  assign _0274_ = _0368_ | { 1'h0, rd_t0[35:32] };
  assign _0277_ = _0369_ | _0017_;
  assign _0280_ = _0370_ | { 1'h0, rd_t0[39:36] };
  assign _0283_ = _0371_ | _0019_;
  assign _0286_ = _0372_ | { 1'h0, rd_t0[43:40] };
  assign _0289_ = _0373_ | _0021_;
  assign _0292_ = _0374_ | { 1'h0, rd_t0[47:44] };
  assign _0295_ = _0375_ | _0023_;
  assign _0298_ = _0376_ | { 1'h0, rd_t0[51:48] };
  assign _0301_ = _0377_ | _0025_;
  assign _0304_ = _0378_ | { 1'h0, rd_t0[55:52] };
  assign _0307_ = _0379_ | _0027_;
  assign _0310_ = _0380_ | { 1'h0, rd_t0[59:56] };
  assign _0313_ = _0381_ | _0029_;
  assign _0316_ = _0382_ | { 1'h0, rd_t0[63:60] };
  assign _0319_ = _0383_ | _0031_;
  assign { next_rdt_t0[3], next_rd_t0[3:0] } = _0229_ | { 1'h0, this_rs2_t0[3:0] };
  assign _0003_ = _0232_ | { 4'h0, rdx_t0[4] };
  assign { next_rdt_t0[7], next_rd_t0[7:4] } = _0235_ | { 1'h0, this_rs2_t0[7:4] };
  assign _0005_ = _0238_ | { 4'h0, rdx_t0[8] };
  assign { next_rdt_t0[11], next_rd_t0[11:8] } = _0241_ | { 1'h0, this_rs2_t0[11:8] };
  assign _0007_ = _0244_ | { 4'h0, rdx_t0[12] };
  assign { next_rdt_t0[15], next_rd_t0[15:12] } = _0247_ | { 1'h0, this_rs2_t0[15:12] };
  assign _0009_ = _0250_ | { 4'h0, rdx_t0[16] };
  assign { next_rdt_t0[19], next_rd_t0[19:16] } = _0253_ | { 1'h0, this_rs2_t0[19:16] };
  assign _0011_ = _0256_ | { 4'h0, rdx_t0[20] };
  assign { next_rdt_t0[23], next_rd_t0[23:20] } = _0259_ | { 1'h0, this_rs2_t0[23:20] };
  assign _0013_ = _0262_ | { 4'h0, rdx_t0[24] };
  assign { next_rdt_t0[27], next_rd_t0[27:24] } = _0265_ | { 1'h0, this_rs2_t0[27:24] };
  assign _0015_ = _0268_ | { 4'h0, rdx_t0[28] };
  assign { next_rdt_t0[31], next_rd_t0[31:28] } = _0271_ | { 1'h0, this_rs2_t0[31:28] };
  assign _0017_ = _0274_ | { 4'h0, rdx_t0[32] };
  assign { next_rdt_t0[35], next_rd_t0[35:32] } = _0277_ | { 1'h0, this_rs2_t0[35:32] };
  assign _0019_ = _0280_ | { 4'h0, rdx_t0[36] };
  assign { next_rdt_t0[39], next_rd_t0[39:36] } = _0283_ | { 1'h0, this_rs2_t0[39:36] };
  assign _0021_ = _0286_ | { 4'h0, rdx_t0[40] };
  assign { next_rdt_t0[43], next_rd_t0[43:40] } = _0289_ | { 1'h0, this_rs2_t0[43:40] };
  assign _0023_ = _0292_ | { 4'h0, rdx_t0[44] };
  assign { next_rdt_t0[47], next_rd_t0[47:44] } = _0295_ | { 1'h0, this_rs2_t0[47:44] };
  assign _0025_ = _0298_ | { 4'h0, rdx_t0[48] };
  assign { next_rdt_t0[51], next_rd_t0[51:48] } = _0301_ | { 1'h0, this_rs2_t0[51:48] };
  assign _0027_ = _0304_ | { 4'h0, rdx_t0[52] };
  assign { next_rdt_t0[55], next_rd_t0[55:52] } = _0307_ | { 1'h0, this_rs2_t0[55:52] };
  assign _0029_ = _0310_ | { 4'h0, rdx_t0[56] };
  assign { next_rdt_t0[59], next_rd_t0[59:56] } = _0313_ | { 1'h0, this_rs2_t0[59:56] };
  assign _0031_ = _0316_ | { 4'h0, rdx_t0[60] };
  assign { next_rdt_t0[63], next_rd_t0[63:60] } = _0319_ | { 1'h0, this_rs2_t0[63:60] };
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME pcpi_ready_t0 */
  always_ff @(posedge clk)
    pcpi_ready_t0 <= _0001_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME pcpi_wait_t0 */
  always_ff @(posedge clk)
    pcpi_wait_t0 <= instr_any_mul_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME pcpi_wait_q_t0 */
  always_ff @(posedge clk)
    pcpi_wait_q_t0 <= pcpi_wait_t0;
  assign _0384_ = _0496_[31:0] ^ pcpi_rd;
  assign _0094_ = ~ resetn;
  assign _0095_ = ~ _0465_;
  assign _0321_ = _0497_[31:0] | pcpi_rd_t0;
  assign _0322_ = _0384_ | _0321_;
  assign _0179_ = { resetn, resetn, resetn, resetn, resetn, resetn, resetn } & _0472_;
  assign _0181_ = { _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_, _0465_ } & _0497_[31:0];
  assign _0188_ = { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn } & _0476_[63:1];
  assign _0192_ = { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn } & _0480_[62:0];
  assign _0180_ = { _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_ } & mul_counter_t0;
  assign _0182_ = { _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_ } & pcpi_rd_t0;
  assign _0189_ = { _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_ } & rs2_t0[63:1];
  assign _0193_ = { _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_ } & rs1_t0[62:0];
  assign _0183_ = _0322_ & { _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_ };
  assign _0320_ = _0179_ | _0180_;
  assign _0323_ = _0181_ | _0182_;
  assign _0327_ = _0188_ | _0189_;
  assign _0329_ = _0192_ | _0193_;
  assign _0324_ = _0323_ | _0183_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME mul_counter_t0 */
  always_ff @(posedge clk)
    mul_counter_t0 <= _0320_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME pcpi_rd_t0 */
  always_ff @(posedge clk)
    pcpi_rd_t0 <= _0324_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rs2_t0[63:1] */
  always_ff @(posedge clk)
    rs2_t0[63:1] <= _0327_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rs1_t0[62:0] */
  always_ff @(posedge clk)
    rs1_t0[62:0] <= _0329_;
  assign _0096_ = | pcpi_insn_t0[14:12];
  assign _0097_ = ~ pcpi_insn_t0[14:12];
  assign _0217_ = pcpi_insn[14:12] & _0097_;
  assign _0393_ = _0217_ == { 1'h0, _0097_[1:0] };
  assign _0394_ = _0217_ == { 1'h0, _0097_[1], 1'h0 };
  assign _0395_ = _0217_ == { 2'h0, _0097_[0] };
  assign _0482_ = _0393_ & _0096_;
  assign _0485_ = _0394_ & _0096_;
  assign _0488_ = _0395_ & _0096_;
  /* src = "generated/out/vanilla.sv:1871.2-1885.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME instr_mulhu */
  always_ff @(posedge clk)
    if (!_0464_) instr_mulhu <= 1'h0;
    else instr_mulhu <= _0481_;
  /* src = "generated/out/vanilla.sv:1871.2-1885.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME instr_mulhsu */
  always_ff @(posedge clk)
    if (!_0464_) instr_mulhsu <= 1'h0;
    else instr_mulhsu <= _0484_;
  /* src = "generated/out/vanilla.sv:1871.2-1885.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME instr_mulh */
  always_ff @(posedge clk)
    if (!_0464_) instr_mulh <= 1'h0;
    else instr_mulh <= _0487_;
  /* src = "generated/out/vanilla.sv:1871.2-1885.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME instr_mul */
  always_ff @(posedge clk)
    if (!_0464_) instr_mul <= 1'h0;
    else instr_mul <= _0490_;
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME mul_waiting */
  always_ff @(posedge clk)
    if (!resetn) mul_waiting <= 1'h1;
    else mul_waiting <= _0469_;
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME mul_finish */
  always_ff @(posedge clk)
    if (_0115_) mul_finish <= 1'h0;
    else mul_finish <= _0468_;
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME mul_counter */
  always_ff @(posedge clk)
    if (resetn) mul_counter <= _0471_;
  /* src = "generated/out/vanilla.sv:1954.2-1962.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME pcpi_rd */
  always_ff @(posedge clk)
    if (_0465_) pcpi_rd <= _0496_[31:0];
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rd */
  always_ff @(posedge clk)
    if (resetn)
      if (mul_waiting) rd <= 64'h0000000000000000;
      else rd <= next_rd;
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rs2[0] */
  always_ff @(posedge clk)
    if (resetn)
      if (!mul_waiting) rs2[0] <= 1'h0;
      else rs2[0] <= _0473_[0];
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rs2[63:1] */
  always_ff @(posedge clk)
    if (resetn) rs2[63:1] <= _0475_[63:1];
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rs1[63] */
  always_ff @(posedge clk)
    if (resetn)
      if (!_0116_) rs1[63] <= 1'h0;
      else rs1[63] <= pcpi_rs1[31];
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rs1[62:0] */
  always_ff @(posedge clk)
    if (resetn) rs1[62:0] <= _0479_[62:0];
  reg [14:0] _0918_;
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME _0918_ */
  always_ff @(posedge clk)
    if (resetn)
      if (mul_waiting) _0918_ <= 15'h0000;
      else _0918_ <= { next_rdt[59], next_rdt[55], next_rdt[51], next_rdt[47], next_rdt[43], next_rdt[39], next_rdt[35], next_rdt[31], next_rdt[27], next_rdt[23], next_rdt[19], next_rdt[15], next_rdt[11], next_rdt[7], next_rdt[3] };
  assign { rdx[60], rdx[56], rdx[52], rdx[48], rdx[44], rdx[40], rdx[36], rdx[32], rdx[28], rdx[24], rdx[20], rdx[16], rdx[12], rdx[8], rdx[4] } = _0918_;
  assign _0196_ = pcpi_wait_t0 & _0466_;
  assign _0001_ = mul_finish_t0 & resetn;
  assign _0197_ = pcpi_wait_q_t0 & pcpi_wait;
  assign _0198_ = pcpi_wait_t0 & pcpi_wait_q_t0;
  assign _0331_ = _0196_ | _0197_;
  assign mul_start_t0 = _0331_ | _0198_;
  assign _0098_ = | { instr_mulhu_t0, instr_mulhsu_t0, instr_mulh_t0, instr_mul_t0 };
  assign _0099_ = | { instr_mulhu_t0, instr_mulhsu_t0, instr_mulh_t0 };
  assign _0100_ = | { instr_mulhsu_t0, instr_mulh_t0 };
  assign _0101_ = ~ { instr_mulhu_t0, instr_mulhsu_t0, instr_mulh_t0, instr_mul_t0 };
  assign _0102_ = ~ { instr_mulhu_t0, instr_mulhsu_t0, instr_mulh_t0 };
  assign _0103_ = ~ { instr_mulhsu_t0, instr_mulh_t0 };
  assign _0218_ = { instr_mulhu, instr_mulhsu, instr_mulh, instr_mul } & _0101_;
  assign _0219_ = { instr_mulhu, instr_mulhsu, instr_mulh } & _0102_;
  assign _0220_ = { instr_mulhsu, instr_mulh } & _0103_;
  assign _0104_ = ! _0217_;
  assign _0105_ = ! _0218_;
  assign _0106_ = ! _0219_;
  assign _0107_ = ! _0220_;
  assign _0491_ = _0104_ & _0096_;
  assign instr_any_mul_t0 = _0105_ & _0098_;
  assign instr_any_mulh_t0 = _0106_ & _0099_;
  assign instr_rs1_signed_t0 = _0107_ & _0100_;
  assign _0108_ = ~ mul_waiting;
  assign _0109_ = ~ { mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting };
  assign _0110_ = ~ { instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh };
  assign _0111_ = ~ { mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting };
  assign _0112_ = ~ { instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed };
  assign _0113_ = ~ { instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh };
  assign _0332_ = mul_waiting_t0 | _0108_;
  assign _0335_ = { mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0 } | _0109_;
  assign _0338_ = { instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0 } | _0110_;
  assign _0341_ = { mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0 } | _0111_;
  assign _0344_ = { instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0 } | _0112_;
  assign _0350_ = { instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0 } | _0113_;
  assign _0333_ = mul_waiting_t0 | mul_waiting;
  assign _0336_ = { mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0 } | { mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting };
  assign _0339_ = { instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0 } | { instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh };
  assign _0342_ = { mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0 } | { mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting };
  assign _0345_ = { instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0 } | { instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed, instr_rs1_signed };
  assign _0349_ = { rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0] } | { rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0] };
  assign _0351_ = { instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0 } | { instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh };
  assign _0199_ = mul_counter_t0[6] & _0332_;
  assign _0202_ = _0494_[6:0] & _0335_;
  assign _0205_ = { 32'h00000000, pcpi_rs2_t0 } & _0338_;
  assign _0208_ = { rs2_t0[62:0], 1'h0 } & _0341_;
  assign _0211_ = { 32'h00000000, pcpi_rs1_t0 } & _0344_;
  assign _0214_ = { 1'h0, rs1_t0[63:1] } & _0341_;
  assign _0224_ = rd_t0 & _0350_;
  assign _0200_ = mul_start_t0 & _0333_;
  assign _0203_ = { 1'h0, instr_any_mulh_t0, 5'h00 } & _0336_;
  assign _0206_ = { pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0 } & _0339_;
  assign _0209_ = _0474_ & _0342_;
  assign _0212_ = { pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0 } & _0345_;
  assign _0215_ = _0478_ & _0342_;
  assign _0222_ = rs2_t0 & _0349_;
  assign _0225_ = { 32'h00000000, rd_t0[63:32] } & _0351_;
  assign _0334_ = _0199_ | _0200_;
  assign _0337_ = _0202_ | _0203_;
  assign _0340_ = _0205_ | _0206_;
  assign _0343_ = _0208_ | _0209_;
  assign _0346_ = _0211_ | _0212_;
  assign _0347_ = _0214_ | _0215_;
  assign _0352_ = _0224_ | _0225_;
  assign _0385_ = _0468_ ^ _0467_;
  assign _0386_ = _0493_[6:0] ^ _0495_[6:0];
  assign _0387_ = { 32'h00000000, pcpi_rs2 } ^ { pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2 };
  assign _0388_ = { rs2[62:0], 1'h0 } ^ _0473_;
  assign _0389_ = { 32'h00000000, pcpi_rs1 } ^ { pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1 };
  assign _0390_ = { 1'h0, rs1[63:1] } ^ _0477_;
  assign _0392_ = rd ^ { 32'h00000000, rd[63:32] };
  assign _0201_ = mul_waiting_t0 & _0385_;
  assign _0204_ = { mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0 } & _0386_;
  assign _0207_ = { instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0, instr_mulh_t0 } & _0387_;
  assign _0210_ = { mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0 } & _0388_;
  assign _0213_ = { instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0, instr_rs1_signed_t0 } & _0389_;
  assign _0216_ = { mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0, mul_waiting_t0 } & _0390_;
  assign _0223_ = { rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0], rs1_t0[0] } & rs2;
  assign _0226_ = { instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0, instr_any_mulh_t0 } & _0392_;
  assign _0470_ = _0201_ | _0334_;
  assign _0472_ = _0204_ | _0337_;
  assign _0474_ = _0207_ | _0340_;
  assign _0476_ = _0210_ | _0343_;
  assign _0478_ = _0213_ | _0346_;
  assign _0480_ = _0216_ | _0347_;
  assign this_rs2_t0 = _0223_ | _0222_;
  assign _0497_ = _0226_ | _0352_;
  assign _0115_ = | { _0094_, mul_waiting };
  assign _0116_ = & { mul_waiting, instr_rs1_signed };
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME instr_mulhu_t0 */
  always_ff @(posedge clk)
    if (!_0464_) instr_mulhu_t0 <= 1'h0;
    else instr_mulhu_t0 <= _0482_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME instr_mulhsu_t0 */
  always_ff @(posedge clk)
    if (!_0464_) instr_mulhsu_t0 <= 1'h0;
    else instr_mulhsu_t0 <= _0485_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME instr_mulh_t0 */
  always_ff @(posedge clk)
    if (!_0464_) instr_mulh_t0 <= 1'h0;
    else instr_mulh_t0 <= _0488_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME instr_mul_t0 */
  always_ff @(posedge clk)
    if (!_0464_) instr_mul_t0 <= 1'h0;
    else instr_mul_t0 <= _0491_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME mul_waiting_t0 */
  always_ff @(posedge clk)
    if (!resetn) mul_waiting_t0 <= 1'h0;
    else mul_waiting_t0 <= _0470_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME mul_finish_t0 */
  always_ff @(posedge clk)
    if (_0115_) mul_finish_t0 <= 1'h0;
    else mul_finish_t0 <= mul_counter_t0[6];
  assign _0184_ = { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn } & next_rd_t0;
  assign _0186_ = resetn & _0474_[0];
  assign _0190_ = resetn & pcpi_rs1_t0[31];
  assign _0194_ = { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn } & { next_rdt_t0[59], next_rdt_t0[55], next_rdt_t0[51], next_rdt_t0[47], next_rdt_t0[43], next_rdt_t0[39], next_rdt_t0[35], next_rdt_t0[31], next_rdt_t0[27], next_rdt_t0[23], next_rdt_t0[19], next_rdt_t0[15], next_rdt_t0[11], next_rdt_t0[7], next_rdt_t0[3] };
  assign _0185_ = { _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_ } & rd_t0;
  assign _0187_ = _0094_ & rs2_t0[0];
  assign _0191_ = _0094_ & rs1_t0[63];
  assign _0195_ = { _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_ } & { rdx_t0[60], rdx_t0[56], rdx_t0[52], rdx_t0[48], rdx_t0[44], rdx_t0[40], rdx_t0[36], rdx_t0[32], rdx_t0[28], rdx_t0[24], rdx_t0[20], rdx_t0[16], rdx_t0[12], rdx_t0[8], rdx_t0[4] };
  assign _0325_ = _0184_ | _0185_;
  assign _0326_ = _0186_ | _0187_;
  assign _0328_ = _0190_ | _0191_;
  assign _0330_ = _0194_ | _0195_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rd_t0 */
  always_ff @(posedge clk)
    if (mul_waiting) rd_t0 <= 64'h0000000000000000;
    else rd_t0 <= _0325_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rs2_t0[0] */
  always_ff @(posedge clk)
    if (!mul_waiting) rs2_t0[0] <= 1'h0;
    else rs2_t0[0] <= _0326_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rs1_t0[63] */
  always_ff @(posedge clk)
    if (!_0116_) rs1_t0[63] <= 1'h0;
    else rs1_t0[63] <= _0328_;
  reg [14:0] _1029_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME _1029_ */
  always_ff @(posedge clk)
    if (mul_waiting) _1029_ <= 15'h0000;
    else _1029_ <= _0330_;
  assign { rdx_t0[60], rdx_t0[56], rdx_t0[52], rdx_t0[48], rdx_t0[44], rdx_t0[40], rdx_t0[36], rdx_t0[32], rdx_t0[28], rdx_t0[24], rdx_t0[20], rdx_t0[16], rdx_t0[12], rdx_t0[8], rdx_t0[4] } = _1029_;
  assign _0114_ = ~ { 25'h0000000, mul_counter_t0 };
  assign _0221_ = { 25'h0000000, mul_counter } & _0114_;
  assign _0348_ = { 25'h0000000, mul_counter } | { 25'h0000000, mul_counter_t0 };
  assign _0458_ = _0348_ - 32'd1;
  assign _0459_ = _0221_ - 32'd1;
  assign _0391_ = _0458_ ^ _0459_;
  assign _0494_ = _0391_ | { 25'h0000000, mul_counter_t0 };
  assign _0460_ = pcpi_insn[6:0] == /* src = "generated/out/vanilla.sv:1876.35-1876.63" */ 7'h33;
  assign _0461_ = pcpi_insn[31:25] == /* src = "generated/out/vanilla.sv:1876.70-1876.100" */ 7'h01;
  assign mul_start = pcpi_wait && /* src = "generated/out/vanilla.sv:1870.19-1870.44" */ _0466_;
  assign _0462_ = resetn && /* src = "generated/out/vanilla.sv:1876.9-1876.29" */ pcpi_valid;
  assign _0463_ = _0462_ && /* src = "generated/out/vanilla.sv:1876.8-1876.64" */ _0460_;
  assign _0464_ = _0463_ && /* src = "generated/out/vanilla.sv:1876.7-1876.101" */ _0461_;
  assign _0465_ = mul_finish && /* src = "generated/out/vanilla.sv:1957.7-1957.27" */ resetn;
  assign _0466_ = ! /* src = "generated/out/vanilla.sv:1870.32-1870.44" */ pcpi_wait_q;
  assign _0467_ = ! /* src = "generated/out/vanilla.sv:1940.19-1940.29" */ mul_start;
  /* src = "generated/out/vanilla.sv:1954.2-1962.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME pcpi_ready */
  always_ff @(posedge clk)
    pcpi_ready <= _0000_;
  /* src = "generated/out/vanilla.sv:1871.2-1885.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME pcpi_wait */
  always_ff @(posedge clk)
    pcpi_wait <= instr_any_mul;
  /* src = "generated/out/vanilla.sv:1871.2-1885.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME pcpi_wait_q */
  always_ff @(posedge clk)
    pcpi_wait_q <= pcpi_wait;
  assign _0000_ = _0465_ ? /* src = "generated/out/vanilla.sv:1957.7-1957.27|generated/out/vanilla.sv:1957.3-1961.6" */ 1'h1 : 1'h0;
  assign _0468_ = mul_counter[6] ? /* src = "generated/out/vanilla.sv:1948.8-1948.22|generated/out/vanilla.sv:1948.4-1951.7" */ 1'h1 : 1'h0;
  assign _0469_ = mul_waiting ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1928.12-1928.23|generated/out/vanilla.sv:1928.8-1952.6" */ _0467_ : _0468_;
  assign _0471_ = mul_waiting ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1928.12-1928.23|generated/out/vanilla.sv:1928.8-1952.6" */ _0495_[6:0] : _0493_[6:0];
  assign _0473_ = instr_mulh ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1933.8-1933.24|generated/out/vanilla.sv:1933.4-1936.32" */ { pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2 } : { 32'h00000000, pcpi_rs2 };
  assign _0475_ = mul_waiting ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1928.12-1928.23|generated/out/vanilla.sv:1928.8-1952.6" */ _0473_ : { rs2[62:0], 1'h0 };
  assign _0477_ = instr_rs1_signed ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1929.8-1929.24|generated/out/vanilla.sv:1929.4-1932.32" */ { pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1 } : { 32'h00000000, pcpi_rs1 };
  assign _0479_ = mul_waiting ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1928.12-1928.23|generated/out/vanilla.sv:1928.8-1952.6" */ _0477_ : { 1'h0, rs1[63:1] };
  assign _0481_ = _0483_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1877.4-1882.11" */ 1'h1 : 1'h0;
  assign _0483_ = pcpi_insn[14:12] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1877.4-1882.11" */ 3'h3;
  assign _0484_ = _0486_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1877.4-1882.11" */ 1'h1 : 1'h0;
  assign _0486_ = pcpi_insn[14:12] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1877.4-1882.11" */ 3'h2;
  assign _0487_ = _0489_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1877.4-1882.11" */ 1'h1 : 1'h0;
  assign _0489_ = pcpi_insn[14:12] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1877.4-1882.11" */ 3'h1;
  assign _0490_ = _0492_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1877.4-1882.11" */ 1'h1 : 1'h0;
  assign _0492_ = ! /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1877.4-1882.11" */ pcpi_insn[14:12];
  assign instr_any_mul = | /* src = "generated/out/vanilla.sv:1865.23-1865.74" */ { instr_mulhu, instr_mulhsu, instr_mulh, instr_mul };
  assign instr_any_mulh = | /* src = "generated/out/vanilla.sv:1866.24-1866.64" */ { instr_mulhu, instr_mulhsu, instr_mulh };
  assign instr_rs1_signed = | /* src = "generated/out/vanilla.sv:1867.26-1867.53" */ { instr_mulhsu, instr_mulh };
  assign _0493_ = mul_counter - /* src = "generated/out/vanilla.sv:1947.19-1947.46" */ 32'd1;
  assign this_rs2 = rs1[0] ? /* src = "generated/out/vanilla.sv:1908.17-1908.43" */ rs2 : 64'h0000000000000000;
  assign _0495_ = instr_any_mulh ? /* src = "generated/out/vanilla.sv:1939.20-1939.76" */ 32'd62 : 32'd30;
  assign _0496_ = instr_any_mulh ? /* src = "generated/out/vanilla.sv:1960.16-1960.46" */ { 32'h00000000, rd[63:32] } : rd;
  assign { next_rdt[62:60], next_rdt[58:56], next_rdt[54:52], next_rdt[50:48], next_rdt[46:44], next_rdt[42:40], next_rdt[38:36], next_rdt[34:32], next_rdt[30:28], next_rdt[26:24], next_rdt[22:20], next_rdt[18:16], next_rdt[14:12], next_rdt[10:8], next_rdt[6:4], next_rdt[2:0] } = 48'h000000000000;
  assign { next_rdt_t0[62:60], next_rdt_t0[58:56], next_rdt_t0[54:52], next_rdt_t0[50:48], next_rdt_t0[46:44], next_rdt_t0[42:40], next_rdt_t0[38:36], next_rdt_t0[34:32], next_rdt_t0[30:28], next_rdt_t0[26:24], next_rdt_t0[22:20], next_rdt_t0[18:16], next_rdt_t0[14:12], next_rdt_t0[10:8], next_rdt_t0[6:4], next_rdt_t0[2:0] } = 48'h000000000000;
  assign pcpi_wr = pcpi_ready;
  assign pcpi_wr_t0 = pcpi_ready_t0;
  assign { rdx[63:61], rdx[59:57], rdx[55:53], rdx[51:49], rdx[47:45], rdx[43:41], rdx[39:37], rdx[35:33], rdx[31:29], rdx[27:25], rdx[23:21], rdx[19:17], rdx[15:13], rdx[11:9], rdx[7:5], rdx[3:0] } = 49'h0000000000000;
  assign { rdx_t0[63:61], rdx_t0[59:57], rdx_t0[55:53], rdx_t0[51:49], rdx_t0[47:45], rdx_t0[43:41], rdx_t0[39:37], rdx_t0[35:33], rdx_t0[31:29], rdx_t0[27:25], rdx_t0[23:21], rdx_t0[19:17], rdx_t0[15:13], rdx_t0[11:9], rdx_t0[7:5], rdx_t0[3:0] } = 49'h0000000000000;
endmodule
