bit gen_regrd_rs2;
assign gen_regrd_rs2 = 
 (((| { (i_pipeline__i_gprs__rs2_addr  ==  5'h1c), (i_pipeline__i_gprs__rs2_addr  ==  5'h18), (i_pipeline__i_gprs__rs2_addr  ==  5'h14), (i_pipeline__i_gprs__rs2_addr  ==  5'h10), (i_pipeline__i_gprs__rs2_addr  ==  5'h11), ((i_pipeline__i_gprs__rs2_addr  ==  5'h12) | (i_pipeline__i_gprs__rs2_addr  ==  5'h13)), (i_pipeline__i_gprs__rs2_addr  ==  5'h1d), ((i_pipeline__i_gprs__rs2_addr  ==  5'h1e) | (i_pipeline__i_gprs__rs2_addr  ==  5'h1f)), (i_pipeline__i_gprs__rs2_addr  ==  5'h19), (i_pipeline__i_gprs__rs2_addr  ==  5'h15), ((i_pipeline__i_gprs__rs2_addr  ==  5'h1a) | (i_pipeline__i_gprs__rs2_addr  ==  5'h1b)), ((i_pipeline__i_gprs__rs2_addr  ==  5'h16) | (i_pipeline__i_gprs__rs2_addr  ==  5'h17)) }) | ((~ (| { (i_pipeline__i_gprs__rs2_addr  ==  5'h1c), (i_pipeline__i_gprs__rs2_addr  ==  5'h18), (i_pipeline__i_gprs__rs2_addr  ==  5'h14), (i_pipeline__i_gprs__rs2_addr  ==  5'h10), (i_pipeline__i_gprs__rs2_addr  ==  5'h11), ((i_pipeline__i_gprs__rs2_addr  ==  5'h12) | (i_pipeline__i_gprs__rs2_addr  ==  5'h13)), (i_pipeline__i_gprs__rs2_addr  ==  5'h1d), ((i_pipeline__i_gprs__rs2_addr  ==  5'h1e) | (i_pipeline__i_gprs__rs2_addr  ==  5'h1f)), (i_pipeline__i_gprs__rs2_addr  ==  5'h19), (i_pipeline__i_gprs__rs2_addr  ==  5'h15), ((i_pipeline__i_gprs__rs2_addr  ==  5'h1a) | (i_pipeline__i_gprs__rs2_addr  ==  5'h1b)), ((i_pipeline__i_gprs__rs2_addr  ==  5'h16) | (i_pipeline__i_gprs__rs2_addr  ==  5'h17)) })) &
((| { (i_pipeline__i_gprs__rs2_addr  ==  5'h0c), (i_pipeline__i_gprs__rs2_addr  ==  5'h08), (i_pipeline__i_gprs__rs2_addr  ==  5'h09), ((i_pipeline__i_gprs__rs2_addr  ==  5'h0a) | (i_pipeline__i_gprs__rs2_addr  ==  5'h0b)), (i_pipeline__i_gprs__rs2_addr  ==  5'h0d), ((i_pipeline__i_gprs__rs2_addr  ==  5'h0e) | (i_pipeline__i_gprs__rs2_addr  ==  5'h0f)) }) | ((~ (| { (i_pipeline__i_gprs__rs2_addr  ==  5'h0c), (i_pipeline__i_gprs__rs2_addr  ==  5'h08), (i_pipeline__i_gprs__rs2_addr  ==  5'h09), ((i_pipeline__i_gprs__rs2_addr  ==  5'h0a) | (i_pipeline__i_gprs__rs2_addr  ==  5'h0b)), (i_pipeline__i_gprs__rs2_addr  ==  5'h0d), ((i_pipeline__i_gprs__rs2_addr  ==  5'h0e) | (i_pipeline__i_gprs__rs2_addr  ==  5'h0f)) })) &
((| { (i_pipeline__i_gprs__rs2_addr  ==  5'h04), (i_pipeline__i_gprs__rs2_addr  ==  5'h05), ((i_pipeline__i_gprs__rs2_addr  ==  5'h06) | (i_pipeline__i_gprs__rs2_addr  ==  5'h07)) }) | ((~ (| { (i_pipeline__i_gprs__rs2_addr  ==  5'h04), (i_pipeline__i_gprs__rs2_addr  ==  5'h05), ((i_pipeline__i_gprs__rs2_addr  ==  5'h06) | (i_pipeline__i_gprs__rs2_addr  ==  5'h07)) })) &
(((i_pipeline__i_gprs__rs2_addr  ==  5'h02) | (i_pipeline__i_gprs__rs2_addr  ==  5'h03)) | ((~ ((i_pipeline__i_gprs__rs2_addr  ==  5'h02) | (i_pipeline__i_gprs__rs2_addr  ==  5'h03))) &
(i_pipeline__i_gprs__rs2_addr  ==  5'h01))))))))));
;