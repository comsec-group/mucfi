`include "formal/assumptions/cellift_scarv_di_asm.sv"
`include "formal/assumptions/cellift_scarv_ti_asm.sv"
