module names
//   0bc5471c4599dca6379e3da212968f59ed7c2433kronos_EX: simplif_9e9afc4272f55a9beacc
//   0bc5471c4599dca6379e3da212968f59ed7c2433kronos_csr: simplif_23175af27fd2ffc5d196
//   7f28a733942cfa68708efb963cc03bff51aab720kronos_counter64: simplif_b656ed3944a4d79ba92b
//   18af26cedc4b6bb625254872dcfca9175553c879kronos_agu: simplif_8a2982a34f91f245ed13
//   3d7c8832d64513bf58d5683a07b8f397329345dckronos_IF: simplif_db7b5d87aea4226b70fe
//   56f4e880e76900c55ae6bcfa76aead2ec9aaa66ekronos_core: simplif_1b215dccbb32fdcc253c
//   7ba81c6d179a62ecfdf087977491187ed598ce2ekronos_ID: simplif_62dbb6e3107130a7cf75

/* Generated by Yosys 0.29+11 (git sha1 e3db31c02, gcc 9.4.0-1ubuntu1~20.04.1 -fPIC -Os) */

/* cellift =  1  */
/* hdlname = "\\kronos_EX" */
/* src = "generated/sv2v_out.v:589.1-839.10" */
module paramodsimplif_9e9afc4272f55a9beacc (clk, rstz, decode, decode_vld, decode_rdy, regwr_data, regwr_sel, regwr_en, regwr_pending, branch_target, branch, data_addr, data_rd_data, data_wr_data, data_mask, data_wr_en, data_req, data_ack, software_interrupt, timer_interrupt, external_interrupt
, clk_t0, timer_interrupt_t0, software_interrupt_t0, external_interrupt_t0, decode_t0, data_ack_t0, data_addr_t0, data_mask_t0, data_rd_data_t0, data_req_t0, data_wr_data_t0, data_wr_en_t0, branch_t0, branch_target_t0, decode_rdy_t0, decode_vld_t0, regwr_data_t0, regwr_en_t0, regwr_pending_t0, regwr_sel_t0);
/* src = "generated/sv2v_out.v:770.2-805.7" */
wire [31:0] _0000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:770.2-805.7" */
wire [31:0] _0001_;
/* src = "generated/sv2v_out.v:770.2-805.7" */
wire [31:0] _0002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:770.2-805.7" */
wire [31:0] _0003_;
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0004_;
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0005_;
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0006_;
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0007_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0008_;
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0009_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0010_;
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0011_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0012_;
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0013_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0014_;
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0015_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0016_;
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0017_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0018_;
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0019_;
/* src = "generated/sv2v_out.v:673.2-707.5" */
wire [2:0] _0020_;
wire _0021_;
/* cellift = 32'd1 */
wire _0022_;
wire _0023_;
/* cellift = 32'd1 */
wire _0024_;
wire _0025_;
/* cellift = 32'd1 */
wire _0026_;
wire _0027_;
/* cellift = 32'd1 */
wire _0028_;
wire _0029_;
/* cellift = 32'd1 */
wire _0030_;
wire _0031_;
/* cellift = 32'd1 */
wire _0032_;
wire _0033_;
/* cellift = 32'd1 */
wire _0034_;
wire _0035_;
/* cellift = 32'd1 */
wire _0036_;
wire _0037_;
/* cellift = 32'd1 */
wire _0038_;
wire _0039_;
/* cellift = 32'd1 */
wire _0040_;
wire _0041_;
/* cellift = 32'd1 */
wire _0042_;
wire _0043_;
/* cellift = 32'd1 */
wire _0044_;
wire _0045_;
/* cellift = 32'd1 */
wire _0046_;
wire _0047_;
/* cellift = 32'd1 */
wire _0048_;
wire _0049_;
/* cellift = 32'd1 */
wire _0050_;
wire [2:0] _0051_;
wire [1:0] _0052_;
wire _0053_;
wire _0054_;
wire _0055_;
wire [1:0] _0056_;
wire [1:0] _0057_;
wire [1:0] _0058_;
wire [1:0] _0059_;
wire _0060_;
wire _0061_;
wire _0062_;
wire _0063_;
wire _0064_;
wire _0065_;
wire [7:0] _0066_;
wire [2:0] _0067_;
wire [1:0] _0068_;
wire [2:0] _0069_;
wire [6:0] _0070_;
wire [1:0] _0071_;
wire [1:0] _0072_;
wire [1:0] _0073_;
wire [1:0] _0074_;
wire [1:0] _0075_;
wire [5:0] _0076_;
wire [1:0] _0077_;
wire [3:0] _0078_;
wire [2:0] _0079_;
wire [2:0] _0080_;
wire [2:0] _0081_;
wire [2:0] _0082_;
wire [2:0] _0083_;
wire _0084_;
wire _0085_;
wire _0086_;
wire _0087_;
wire _0088_;
wire _0089_;
wire _0090_;
wire _0091_;
wire _0092_;
wire _0093_;
wire _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire [31:0] _0107_;
wire [31:0] _0108_;
wire [31:0] _0109_;
wire [31:0] _0110_;
wire [31:0] _0111_;
wire [31:0] _0112_;
wire [31:0] _0113_;
wire _0114_;
wire _0115_;
wire _0116_;
wire [31:0] _0117_;
wire [31:0] _0118_;
wire [2:0] _0119_;
wire [1:0] _0120_;
wire [2:0] _0121_;
wire [2:0] _0122_;
wire [2:0] _0123_;
wire [2:0] _0124_;
wire [31:0] _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
/* cellift = 32'd1 */
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire _0139_;
wire _0140_;
wire _0141_;
wire _0142_;
wire _0143_;
wire _0144_;
wire _0145_;
wire _0146_;
wire _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
wire _0152_;
wire _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire [31:0] _0160_;
wire [31:0] _0161_;
wire [31:0] _0162_;
wire [31:0] _0163_;
wire [31:0] _0164_;
wire [31:0] _0165_;
wire [4:0] _0166_;
wire [4:0] _0167_;
wire [31:0] _0168_;
wire [31:0] _0169_;
wire [31:0] _0170_;
wire [2:0] _0171_;
wire [2:0] _0172_;
wire [2:0] _0173_;
wire [7:0] _0174_;
wire [2:0] _0175_;
wire [1:0] _0176_;
wire [2:0] _0177_;
wire [6:0] _0178_;
wire [1:0] _0179_;
wire [1:0] _0180_;
wire [1:0] _0181_;
wire [1:0] _0182_;
wire [1:0] _0183_;
wire [5:0] _0184_;
wire [1:0] _0185_;
wire [3:0] _0186_;
wire [2:0] _0187_;
wire [2:0] _0188_;
wire [2:0] _0189_;
wire [2:0] _0190_;
wire [2:0] _0191_;
wire [2:0] _0192_;
wire [2:0] _0193_;
wire [2:0] _0194_;
wire [2:0] _0195_;
wire [2:0] _0196_;
wire [2:0] _0197_;
wire _0198_;
wire _0199_;
wire _0200_;
wire _0201_;
wire _0202_;
wire _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
wire _0221_;
wire _0222_;
wire _0223_;
wire _0224_;
wire _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire _0241_;
wire _0242_;
wire _0243_;
wire _0244_;
wire _0245_;
wire _0246_;
wire _0247_;
wire _0248_;
wire _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire _0271_;
wire _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire _0276_;
wire _0277_;
wire [31:0] _0278_;
wire [31:0] _0279_;
wire [31:0] _0280_;
wire [31:0] _0281_;
wire [31:0] _0282_;
wire [31:0] _0283_;
wire [31:0] _0284_;
wire [31:0] _0285_;
wire [31:0] _0286_;
wire [31:0] _0287_;
wire [31:0] _0288_;
wire [31:0] _0289_;
wire [31:0] _0290_;
wire [31:0] _0291_;
wire [31:0] _0292_;
wire [31:0] _0293_;
wire [31:0] _0294_;
wire [31:0] _0295_;
wire [31:0] _0296_;
wire [31:0] _0297_;
wire [31:0] _0298_;
wire [31:0] _0299_;
wire [31:0] _0300_;
wire [31:0] _0301_;
wire [31:0] _0302_;
wire [31:0] _0303_;
wire [31:0] _0304_;
wire [31:0] _0305_;
wire [31:0] _0306_;
wire [31:0] _0307_;
wire [31:0] _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire [31:0] _0323_;
wire [31:0] _0324_;
wire [31:0] _0325_;
wire [31:0] _0326_;
wire [31:0] _0327_;
wire [31:0] _0328_;
wire [1:0] _0329_;
wire [2:0] _0330_;
wire [2:0] _0331_;
wire [2:0] _0332_;
wire [2:0] _0333_;
wire [2:0] _0334_;
wire [2:0] _0335_;
wire [2:0] _0336_;
wire [2:0] _0337_;
wire [2:0] _0338_;
wire [31:0] _0339_;
wire [31:0] _0340_;
wire [31:0] _0341_;
wire _0342_;
wire [31:0] _0343_;
wire [31:0] _0344_;
wire [31:0] _0345_;
wire [31:0] _0346_;
wire [31:0] _0347_;
wire [31:0] _0348_;
wire [31:0] _0349_;
wire [31:0] _0350_;
wire [4:0] _0351_;
wire [31:0] _0352_;
wire [31:0] _0353_;
wire [31:0] _0354_;
wire [31:0] _0355_;
wire [2:0] _0356_;
wire [2:0] _0357_;
wire [2:0] _0358_;
wire [2:0] _0359_;
wire [2:0] _0360_;
wire [1:0] _0361_;
wire [6:0] _0362_;
wire [2:0] _0363_;
wire [2:0] _0364_;
wire [2:0] _0365_;
wire [2:0] _0366_;
wire [2:0] _0367_;
wire [2:0] _0368_;
wire [2:0] _0369_;
wire _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire _0376_;
wire _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire _0382_;
wire _0383_;
wire _0384_;
wire _0385_;
wire _0386_;
wire _0387_;
wire _0388_;
wire _0389_;
wire _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire [31:0] _0398_;
wire [31:0] _0399_;
wire [31:0] _0400_;
wire [31:0] _0401_;
wire [31:0] _0402_;
wire [31:0] _0403_;
wire [31:0] _0404_;
wire [31:0] _0405_;
wire [31:0] _0406_;
wire [31:0] _0407_;
wire [31:0] _0408_;
wire [31:0] _0409_;
wire [31:0] _0410_;
wire [31:0] _0411_;
wire [31:0] _0412_;
wire [31:0] _0413_;
wire [31:0] _0414_;
wire [31:0] _0415_;
wire [31:0] _0416_;
wire [31:0] _0417_;
wire [31:0] _0418_;
wire _0419_;
wire _0420_;
wire _0421_;
wire _0422_;
wire _0423_;
wire _0424_;
wire _0425_;
wire _0426_;
wire [31:0] _0427_;
wire [31:0] _0428_;
wire [31:0] _0429_;
wire [31:0] _0430_;
wire [31:0] _0431_;
wire [31:0] _0432_;
wire [31:0] _0433_;
wire [2:0] _0434_;
wire [2:0] _0435_;
wire [2:0] _0436_;
wire [2:0] _0437_;
wire [2:0] _0438_;
wire [2:0] _0439_;
wire [31:0] _0440_;
wire [31:0] _0441_;
wire [31:0] _0442_;
wire [31:0] _0443_;
wire [31:0] _0444_;
wire [31:0] _0445_;
wire [2:0] _0446_;
wire [2:0] _0447_;
wire [2:0] _0448_;
wire [2:0] _0449_;
wire [2:0] _0450_;
wire [2:0] _0451_;
wire [31:0] _0452_;
wire [31:0] _0453_;
wire [31:0] _0454_;
wire [31:0] _0455_;
wire [31:0] _0456_;
wire [31:0] _0457_;
wire [31:0] _0458_;
wire [31:0] _0459_;
wire [31:0] _0460_;
wire [31:0] _0461_;
wire [31:0] _0462_;
wire [31:0] _0463_;
wire [31:0] _0464_;
wire [31:0] _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire _0469_;
wire [31:0] _0470_;
wire [31:0] _0471_;
wire [2:0] _0472_;
wire [31:0] _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire _0477_;
wire _0478_;
wire _0479_;
wire _0480_;
wire _0481_;
wire _0482_;
wire _0483_;
wire _0484_;
wire _0485_;
wire _0486_;
wire _0487_;
wire _0488_;
wire _0489_;
wire _0490_;
wire [2:0] _0491_;
/* cellift = 32'd1 */
wire [2:0] _0492_;
wire [2:0] _0493_;
/* cellift = 32'd1 */
wire [2:0] _0494_;
wire [2:0] _0495_;
/* cellift = 32'd1 */
wire [2:0] _0496_;
wire [2:0] _0497_;
/* cellift = 32'd1 */
wire [2:0] _0498_;
wire [2:0] _0499_;
/* cellift = 32'd1 */
wire [2:0] _0500_;
/* src = "generated/sv2v_out.v:708.38-708.51" */
wire _0501_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:708.38-708.51" */
wire _0502_;
/* src = "generated/sv2v_out.v:717.33-717.46" */
wire _0503_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:717.33-717.46" */
wire _0504_;
/* src = "generated/sv2v_out.v:792.13-792.47" */
wire _0505_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:792.13-792.47" */
wire _0506_;
/* src = "generated/sv2v_out.v:796.13-796.48" */
wire _0507_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:796.13-796.48" */
wire _0508_;
/* src = "generated/sv2v_out.v:801.12-801.25" */
wire _0509_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:801.12-801.25" */
wire _0510_;
/* src = "generated/sv2v_out.v:806.33-806.46" */
wire _0511_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:806.33-806.46" */
wire _0512_;
/* src = "generated/sv2v_out.v:708.22-708.67" */
wire _0513_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:708.22-708.67" */
wire _0514_;
/* src = "generated/sv2v_out.v:708.23-708.52" */
wire _0515_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:708.23-708.52" */
wire _0516_;
/* src = "generated/sv2v_out.v:732.37-732.61" */
wire _0517_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:732.37-732.61" */
wire _0518_;
/* src = "generated/sv2v_out.v:733.53-733.103" */
wire _0519_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:733.53-733.103" */
wire _0520_;
/* src = "generated/sv2v_out.v:742.29-742.50" */
wire _0521_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:742.29-742.50" */
wire _0522_;
/* src = "generated/sv2v_out.v:742.55-742.76" */
wire _0523_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:742.55-742.76" */
wire _0524_;
/* src = "generated/sv2v_out.v:743.8-743.31" */
wire _0525_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:743.8-743.31" */
wire _0526_;
/* src = "generated/sv2v_out.v:747.13-747.33" */
wire _0527_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:747.13-747.33" */
wire _0528_;
/* src = "generated/sv2v_out.v:752.13-752.33" */
wire _0529_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:752.13-752.33" */
wire _0530_;
/* src = "generated/sv2v_out.v:762.19-762.42" */
wire _0531_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:762.19-762.42" */
wire _0532_;
/* src = "generated/sv2v_out.v:763.50-763.73" */
wire _0533_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:763.50-763.73" */
wire _0534_;
/* src = "generated/sv2v_out.v:784.13-784.36" */
wire _0535_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:784.13-784.36" */
wire _0536_;
/* src = "generated/sv2v_out.v:788.13-788.36" */
wire _0537_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:788.13-788.36" */
wire _0538_;
/* src = "generated/sv2v_out.v:838.46-838.68" */
wire _0539_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:838.46-838.68" */
wire _0540_;
/* src = "generated/sv2v_out.v:688.15-688.39" */
wire _0541_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:688.15-688.39" */
wire _0542_;
/* src = "generated/sv2v_out.v:763.22-763.44" */
wire _0543_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:763.22-763.44" */
wire _0544_;
/* src = "generated/sv2v_out.v:838.15-838.69" */
wire _0545_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:838.15-838.69" */
wire _0546_;
/* src = "generated/sv2v_out.v:708.57-708.67" */
wire _0547_;
/* src = "generated/sv2v_out.v:708.72-708.87" */
wire _0548_;
/* src = "generated/sv2v_out.v:742.42-742.50" */
wire _0549_;
/* src = "generated/sv2v_out.v:742.68-742.76" */
wire _0550_;
/* src = "generated/sv2v_out.v:732.67-732.89" */
wire _0551_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:732.67-732.89" */
wire _0552_;
/* src = "generated/sv2v_out.v:732.66-732.102" */
wire _0553_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:732.66-732.102" */
wire _0554_;
/* src = "generated/sv2v_out.v:742.28-742.77" */
wire _0555_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:742.28-742.77" */
wire _0556_;
wire [31:0] _0557_;
wire [31:0] _0558_;
/* cellift = 32'd1 */
wire [31:0] _0559_;
wire [31:0] _0560_;
/* cellift = 32'd1 */
wire [31:0] _0561_;
wire [31:0] _0562_;
/* cellift = 32'd1 */
wire [31:0] _0563_;
wire [31:0] _0564_;
/* cellift = 32'd1 */
wire [31:0] _0565_;
wire [31:0] _0566_;
/* cellift = 32'd1 */
wire [31:0] _0567_;
/* cellift = 32'd1 */
wire [31:0] _0568_;
wire [31:0] _0569_;
/* cellift = 32'd1 */
wire [31:0] _0570_;
wire [31:0] _0571_;
/* cellift = 32'd1 */
wire [31:0] _0572_;
wire [31:0] _0573_;
/* cellift = 32'd1 */
wire [31:0] _0574_;
wire [31:0] _0575_;
wire [31:0] _0576_;
/* cellift = 32'd1 */
wire [31:0] _0577_;
wire [31:0] _0578_;
/* cellift = 32'd1 */
wire [31:0] _0579_;
/* cellift = 32'd1 */
wire [31:0] _0580_;
wire [31:0] _0581_;
/* cellift = 32'd1 */
wire [31:0] _0582_;
wire [31:0] _0583_;
/* cellift = 32'd1 */
wire [31:0] _0584_;
wire [31:0] _0585_;
/* cellift = 32'd1 */
wire [31:0] _0586_;
wire _0587_;
wire _0588_;
/* cellift = 32'd1 */
wire _0589_;
wire _0590_;
/* cellift = 32'd1 */
wire _0591_;
/* cellift = 32'd1 */
wire _0592_;
/* cellift = 32'd1 */
wire _0593_;
wire _0594_;
/* cellift = 32'd1 */
wire _0595_;
wire _0596_;
/* cellift = 32'd1 */
wire _0597_;
wire [31:0] _0598_;
/* cellift = 32'd1 */
wire [31:0] _0599_;
wire [31:0] _0600_;
/* cellift = 32'd1 */
wire [31:0] _0601_;
wire [31:0] _0602_;
/* cellift = 32'd1 */
wire [31:0] _0603_;
wire _0604_;
/* cellift = 32'd1 */
wire _0605_;
wire _0606_;
/* cellift = 32'd1 */
wire _0607_;
wire _0608_;
/* src = "generated/sv2v_out.v:653.7-653.20" */
wire activate_trap;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:653.7-653.20" */
wire activate_trap_t0;
/* src = "generated/sv2v_out.v:640.7-640.16" */
wire basic_rdy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:640.7-640.16" */
wire basic_rdy_t0;
/* src = "generated/sv2v_out.v:625.14-625.20" */
output branch;
wire branch;
/* cellift = 32'd1 */
output branch_t0;
wire branch_t0;
/* src = "generated/sv2v_out.v:624.21-624.34" */
output [31:0] branch_target;
wire [31:0] branch_target;
/* cellift = 32'd1 */
output [31:0] branch_target_t0;
wire [31:0] branch_target_t0;
/* src = "generated/sv2v_out.v:615.13-615.16" */
input clk;
wire clk;
/* cellift = 32'd1 */
input clk_t0;
wire clk_t0;
/* src = "generated/sv2v_out.v:650.7-650.21" */
wire core_interrupt;
/* src = "generated/sv2v_out.v:651.13-651.33" */
wire [3:0] core_interrupt_cause;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:651.13-651.33" */
wire [3:0] core_interrupt_cause_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:650.7-650.21" */
wire core_interrupt_t0;
/* src = "generated/sv2v_out.v:647.14-647.22" */
wire [31:0] csr_data;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:647.14-647.22" */
wire [31:0] csr_data_t0;
/* src = "generated/sv2v_out.v:646.7-646.14" */
wire csr_rdy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:646.7-646.14" */
wire csr_rdy_t0;
/* src = "generated/sv2v_out.v:645.7-645.14" */
wire csr_vld;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:645.7-645.14" */
wire csr_vld_t0;
/* src = "generated/sv2v_out.v:632.13-632.21" */
input data_ack;
wire data_ack;
/* cellift = 32'd1 */
input data_ack_t0;
wire data_ack_t0;
/* src = "generated/sv2v_out.v:626.21-626.30" */
output [31:0] data_addr;
wire [31:0] data_addr;
/* cellift = 32'd1 */
output [31:0] data_addr_t0;
wire [31:0] data_addr_t0;
/* src = "generated/sv2v_out.v:629.20-629.29" */
output [3:0] data_mask;
wire [3:0] data_mask;
/* cellift = 32'd1 */
output [3:0] data_mask_t0;
wire [3:0] data_mask_t0;
/* src = "generated/sv2v_out.v:627.20-627.32" */
input [31:0] data_rd_data;
wire [31:0] data_rd_data;
/* cellift = 32'd1 */
input [31:0] data_rd_data_t0;
wire [31:0] data_rd_data_t0;
/* src = "generated/sv2v_out.v:631.14-631.22" */
output data_req;
wire data_req;
/* cellift = 32'd1 */
output data_req_t0;
wire data_req_t0;
/* src = "generated/sv2v_out.v:628.21-628.33" */
output [31:0] data_wr_data;
wire [31:0] data_wr_data;
/* cellift = 32'd1 */
output [31:0] data_wr_data_t0;
wire [31:0] data_wr_data_t0;
/* src = "generated/sv2v_out.v:630.14-630.24" */
output data_wr_en;
wire data_wr_en;
/* cellift = 32'd1 */
output data_wr_en_t0;
wire data_wr_en_t0;
/* src = "generated/sv2v_out.v:617.21-617.27" */
input [180:0] decode;
wire [180:0] decode;
/* src = "generated/sv2v_out.v:619.14-619.24" */
output decode_rdy;
wire decode_rdy;
/* cellift = 32'd1 */
output decode_rdy_t0;
wire decode_rdy_t0;
/* cellift = 32'd1 */
input [180:0] decode_t0;
wire [180:0] decode_t0;
/* src = "generated/sv2v_out.v:618.13-618.23" */
input decode_vld;
wire decode_vld;
/* cellift = 32'd1 */
input decode_vld_t0;
wire decode_vld_t0;
/* src = "generated/sv2v_out.v:652.7-652.16" */
wire exception;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:652.7-652.16" */
wire exception_t0;
/* src = "generated/sv2v_out.v:635.13-635.31" */
input external_interrupt;
wire external_interrupt;
/* cellift = 32'd1 */
input external_interrupt_t0;
wire external_interrupt_t0;
/* src = "generated/sv2v_out.v:639.7-639.17" */
wire instr_jump;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:639.7-639.17" */
wire instr_jump_t0;
/* src = "generated/sv2v_out.v:638.7-638.16" */
wire instr_vld;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:638.7-638.16" */
wire instr_vld_t0;
/* src = "generated/sv2v_out.v:649.6-649.13" */
reg instret;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:649.6-649.13" */
reg instret_t0;
/* src = "generated/sv2v_out.v:643.14-643.23" */
wire [31:0] load_data;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:643.14-643.23" */
wire [31:0] load_data_t0;
/* src = "generated/sv2v_out.v:642.7-642.14" */
wire lsu_rdy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:642.7-642.14" */
wire lsu_rdy_t0;
/* src = "generated/sv2v_out.v:641.7-641.14" */
wire lsu_vld;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:641.7-641.14" */
wire lsu_vld_t0;
/* src = "generated/sv2v_out.v:662.12-662.22" */
wire [2:0] next_state;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:662.12-662.22" */
wire [2:0] next_state_t0;
/* src = "generated/sv2v_out.v:648.7-648.16" */
wire regwr_csr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:648.7-648.16" */
wire regwr_csr_t0;
/* src = "generated/sv2v_out.v:620.20-620.30" */
output [31:0] regwr_data;
reg [31:0] regwr_data;
/* cellift = 32'd1 */
output [31:0] regwr_data_t0;
reg [31:0] regwr_data_t0;
/* src = "generated/sv2v_out.v:622.13-622.21" */
output regwr_en;
reg regwr_en;
/* cellift = 32'd1 */
output regwr_en_t0;
reg regwr_en_t0;
/* src = "generated/sv2v_out.v:644.7-644.16" */
wire regwr_lsu;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:644.7-644.16" */
wire regwr_lsu_t0;
/* src = "generated/sv2v_out.v:623.14-623.27" */
output regwr_pending;
wire regwr_pending;
/* src = "generated/sv2v_out.v:659.7-659.31" */
wire regwr_pending_firstcycle;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:659.7-659.31" */
wire regwr_pending_firstcycle_t0;
/* src = "generated/sv2v_out.v:660.6-660.25" */
reg regwr_pending_later;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:660.6-660.25" */
reg regwr_pending_later_t0;
/* cellift = 32'd1 */
output regwr_pending_t0;
wire regwr_pending_t0;
/* src = "generated/sv2v_out.v:621.19-621.28" */
output [4:0] regwr_sel;
reg [4:0] regwr_sel;
/* cellift = 32'd1 */
output [4:0] regwr_sel_t0;
reg [4:0] regwr_sel_t0;
/* src = "generated/sv2v_out.v:636.14-636.20" */
wire [31:0] result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:636.14-636.20" */
wire [31:0] result_t0;
/* src = "generated/sv2v_out.v:654.7-654.18" */
wire return_trap;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:654.7-654.18" */
wire return_trap_t0;
/* src = "generated/sv2v_out.v:616.13-616.17" */
input rstz;
wire rstz;
/* src = "generated/sv2v_out.v:633.13-633.31" */
input software_interrupt;
wire software_interrupt;
/* cellift = 32'd1 */
input software_interrupt_t0;
wire software_interrupt_t0;
/* src = "generated/sv2v_out.v:661.12-661.17" */
reg [2:0] state;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:661.12-661.17" */
reg [2:0] state_t0;
/* src = "generated/sv2v_out.v:634.13-634.28" */
input timer_interrupt;
wire timer_interrupt;
/* cellift = 32'd1 */
input timer_interrupt_t0;
wire timer_interrupt_t0;
/* src = "generated/sv2v_out.v:655.13-655.23" */
reg [31:0] trap_cause;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:655.13-655.23" */
reg [31:0] trap_cause_t0;
/* src = "generated/sv2v_out.v:656.14-656.25" */
wire [31:0] trap_handle;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:656.14-656.25" */
wire [31:0] trap_handle_t0;
/* src = "generated/sv2v_out.v:658.7-658.16" */
wire trap_jump;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:658.7-658.16" */
wire trap_jump_t0;
/* src = "generated/sv2v_out.v:657.13-657.23" */
reg [31:0] trap_value;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:657.13-657.23" */
reg [31:0] trap_value_t0;
assign regwr_pending_firstcycle = _0517_ & /* src = "generated/sv2v_out.v:732.36-732.103" */ _0553_;
assign _0157_ = _0518_ & _0553_;
assign _0158_ = _0554_ & _0517_;
assign _0159_ = _0518_ & _0554_;
assign _0342_ = _0157_ | _0158_;
assign regwr_pending_firstcycle_t0 = _0342_ | _0159_;
assign _0443_ = _0000_ ^ trap_cause;
assign _0444_ = _0602_ ^ regwr_data;
assign _0445_ = _0002_ ^ trap_value;
assign _0063_ = ~ _0045_;
assign _0064_ = ~ rstz;
assign _0062_ = ~ _0043_;
assign _0343_ = _0001_ | trap_cause_t0;
assign _0347_ = _0603_ | regwr_data_t0;
assign _0352_ = _0003_ | trap_value_t0;
assign _0344_ = _0443_ | _0343_;
assign _0348_ = _0444_ | _0347_;
assign _0353_ = _0445_ | _0352_;
assign _0160_ = { _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_ } & _0001_;
assign _0163_ = { _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_, _0045_ } & _0603_;
assign _0166_ = { rstz, rstz, rstz, rstz, rstz } & decode_t0[128:124];
assign _0168_ = { _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_, _0043_ } & _0003_;
assign _0161_ = { _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_ } & trap_cause_t0;
assign _0164_ = { _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_ } & regwr_data_t0;
assign _0167_ = { _0064_, _0064_, _0064_, _0064_, _0064_ } & regwr_sel_t0;
assign _0169_ = { _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_ } & trap_value_t0;
assign _0162_ = _0344_ & { _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_ };
assign _0165_ = _0348_ & { _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_ };
assign _0170_ = _0353_ & { _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_, _0044_ };
assign _0345_ = _0160_ | _0161_;
assign _0349_ = _0163_ | _0164_;
assign _0351_ = _0166_ | _0167_;
assign _0354_ = _0168_ | _0169_;
assign _0346_ = _0345_ | _0162_;
assign _0350_ = _0349_ | _0165_;
assign _0355_ = _0354_ | _0170_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_9e9afc4272f55a9beacc  */
/* PC_TAINT_INFO STATE_NAME trap_cause_t0 */
always_ff @(posedge clk)
trap_cause_t0 <= _0346_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_9e9afc4272f55a9beacc  */
/* PC_TAINT_INFO STATE_NAME regwr_data_t0 */
always_ff @(posedge clk)
regwr_data_t0 <= _0350_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_9e9afc4272f55a9beacc  */
/* PC_TAINT_INFO STATE_NAME regwr_sel_t0 */
always_ff @(posedge clk)
regwr_sel_t0 <= _0351_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_9e9afc4272f55a9beacc  */
/* PC_TAINT_INFO STATE_NAME trap_value_t0 */
always_ff @(posedge clk)
trap_value_t0 <= _0355_;
assign _0131_ = | { _0508_, _0506_, _0538_, _0536_, _0534_, _0516_, core_interrupt_t0, decode_t0[2] };
assign _0132_ = | { _0510_, _0516_, core_interrupt_t0 };
assign _0135_ = | { _0502_, _0542_, exception_t0, decode_vld_t0, core_interrupt_t0, decode_t0[6:5] };
assign _0136_ = | { _0502_, decode_vld_t0 };
assign _0137_ = | { _0504_, lsu_rdy_t0 };
assign _0138_ = | { _0512_, csr_rdy_t0 };
assign _0139_ = | { _0510_, core_interrupt_t0 };
assign _0140_ = | { _0605_, trap_jump_t0 };
assign _0146_ = | decode_t0[4:3];
assign _0066_ = ~ { _0508_, _0506_, _0538_, _0536_, _0534_, _0516_, core_interrupt_t0, decode_t0[2] };
assign _0067_ = ~ { _0510_, _0516_, core_interrupt_t0 };
assign _0070_ = ~ { _0502_, _0542_, exception_t0, core_interrupt_t0, decode_vld_t0, decode_t0[6:5] };
assign _0071_ = ~ { _0502_, decode_vld_t0 };
assign _0072_ = ~ { _0504_, lsu_rdy_t0 };
assign _0073_ = ~ { _0512_, csr_rdy_t0 };
assign _0074_ = ~ { _0510_, core_interrupt_t0 };
assign _0075_ = ~ { _0605_, trap_jump_t0 };
assign _0123_ = ~ state_t0;
assign _0174_ = { _0507_, _0505_, _0537_, _0535_, _0533_, _0515_, core_interrupt, decode[2] } & _0066_;
assign _0175_ = { _0509_, _0515_, core_interrupt } & _0067_;
assign _0178_ = { _0501_, _0541_, exception, core_interrupt, decode_vld, decode[6:5] } & _0070_;
assign _0179_ = { _0501_, decode_vld } & _0071_;
assign _0180_ = { _0503_, lsu_rdy } & _0072_;
assign _0181_ = { _0511_, csr_rdy } & _0073_;
assign _0182_ = { _0509_, core_interrupt } & _0074_;
assign _0183_ = { _0604_, trap_jump } & _0075_;
assign _0329_ = decode[4:3] & _0120_;
assign _0337_ = state & _0123_;
assign _0474_ = _0174_ == { 5'h00, _0066_[2], 2'h0 };
assign _0475_ = _0175_ == { _0067_[2], 2'h0 };
assign _0476_ = _0178_ == { _0070_[6], 3'h0, _0070_[2], 2'h0 };
assign _0477_ = _0179_ == { _0071_[1], 1'h0 };
assign _0478_ = _0180_ == { _0072_[1], 1'h0 };
assign _0479_ = _0181_ == { _0073_[1], 1'h0 };
assign _0480_ = _0182_ == { _0074_[1], 1'h0 };
assign _0481_ = _0183_ == { _0075_[1], 1'h0 };
assign _0482_ = _0329_ == _0120_;
assign _0483_ = _0329_ == { _0120_[1], 1'h0 };
assign _0484_ = _0329_ == { 1'h0, _0120_[0] };
assign _0485_ = _0337_ == { _0123_[2:1], 1'h0 };
assign _0486_ = _0337_ == { _0123_[2], 2'h0 };
assign _0487_ = _0337_ == { 1'h0, _0123_[1:0] };
assign _0488_ = _0337_ == { _0123_[2], 1'h0, _0123_[0] };
assign _0489_ = _0337_ == { 1'h0, _0123_[1], 1'h0 };
assign _0490_ = _0337_ == { 2'h0, _0123_[0] };
assign _0022_ = _0474_ & _0131_;
assign _0024_ = _0475_ & _0132_;
assign _0030_ = _0476_ & _0135_;
assign _0032_ = _0477_ & _0136_;
assign _0034_ = _0478_ & _0137_;
assign _0036_ = _0479_ & _0138_;
assign _0038_ = _0480_ & _0139_;
assign _0040_ = _0481_ & _0140_;
assign _0607_ = _0482_ & _0146_;
assign _0492_[2] = _0483_ & _0146_;
assign _0508_ = _0484_ & _0146_;
assign _0605_ = _0485_ & _0147_;
assign return_trap_t0 = _0486_ & _0147_;
assign activate_trap_t0 = _0487_ & _0147_;
assign _0510_ = _0488_ & _0147_;
assign _0512_ = _0489_ & _0147_;
assign _0504_ = _0490_ & _0147_;
/* src = "generated/sv2v_out.v:734.2-759.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_9e9afc4272f55a9beacc  */
/* PC_TAINT_INFO STATE_NAME regwr_en */
always_ff @(posedge clk)
if (!rstz) regwr_en <= 1'h0;
else regwr_en <= _0590_;
/* src = "generated/sv2v_out.v:770.2-805.7" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_9e9afc4272f55a9beacc  */
/* PC_TAINT_INFO STATE_NAME trap_cause */
always_ff @(posedge clk)
if (_0043_) trap_cause <= _0000_;
/* src = "generated/sv2v_out.v:734.2-759.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_9e9afc4272f55a9beacc  */
/* PC_TAINT_INFO STATE_NAME regwr_pending_later */
always_ff @(posedge clk)
if (!rstz) regwr_pending_later <= 1'h0;
else regwr_pending_later <= _0596_;
/* src = "generated/sv2v_out.v:734.2-759.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_9e9afc4272f55a9beacc  */
/* PC_TAINT_INFO STATE_NAME regwr_data */
always_ff @(posedge clk)
if (_0045_) regwr_data <= _0602_;
/* src = "generated/sv2v_out.v:734.2-759.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_9e9afc4272f55a9beacc  */
/* PC_TAINT_INFO STATE_NAME regwr_sel */
always_ff @(posedge clk)
if (rstz) regwr_sel <= decode[128:124];
/* src = "generated/sv2v_out.v:834.2-838.70" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_9e9afc4272f55a9beacc  */
/* PC_TAINT_INFO STATE_NAME instret */
always_ff @(posedge clk)
if (!rstz) instret <= 1'h0;
else instret <= _0545_;
/* src = "generated/sv2v_out.v:770.2-805.7" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_9e9afc4272f55a9beacc  */
/* PC_TAINT_INFO STATE_NAME trap_value */
always_ff @(posedge clk)
if (_0043_) trap_value <= _0002_;
/* src = "generated/sv2v_out.v:664.2-668.24" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_9e9afc4272f55a9beacc  */
/* PC_TAINT_INFO STATE_NAME state */
always_ff @(posedge clk)
if (!rstz) state <= 3'h0;
else if (_0047_) state <= next_state;
assign _0198_ = _0516_ & _0547_;
assign _0201_ = _0514_ & _0548_;
assign _0204_ = instr_vld_t0 & decode[20];
assign _0207_ = _0518_ & regwr_pending_later;
assign _0210_ = regwr_lsu_t0 & _0549_;
assign _0213_ = regwr_csr_t0 & _0550_;
assign _0216_ = instr_vld_t0 & decode[15];
assign _0211_ = lsu_rdy_t0 & regwr_lsu;
assign _0214_ = csr_rdy_t0 & regwr_csr;
assign _0221_ = instr_vld_t0 & instr_jump;
assign _0224_ = decode_vld_t0 & _0501_;
assign _0227_ = decode_t0[1] & instr_jump;
assign _0230_ = decode_t0[0] & decode[12];
assign _0233_ = decode_t0[0] & decode[11];
assign _0236_ = decode_vld_t0 & decode_rdy;
assign _0239_ = decode_t0[5] & trap_jump;
assign _0199_ = exception_t0 & _0515_;
assign _0202_ = core_interrupt_t0 & _0513_;
assign _0205_ = decode_t0[20] & instr_vld;
assign _0208_ = regwr_pending_later_t0 & _0097_;
assign _0217_ = decode_t0[15] & instr_vld;
assign _0219_ = regwr_lsu_t0 & lsu_rdy;
assign _0220_ = regwr_csr_t0 & csr_rdy;
assign _0222_ = instr_jump_t0 & instr_vld;
assign _0225_ = _0502_ & decode_vld;
assign _0228_ = instr_jump_t0 & decode[1];
assign _0231_ = decode_t0[12] & decode[0];
assign _0234_ = decode_t0[11] & decode[0];
assign _0237_ = decode_rdy_t0 & decode_vld;
assign _0240_ = trap_jump_t0 & decode[5];
assign _0200_ = _0516_ & exception_t0;
assign _0203_ = _0514_ & core_interrupt_t0;
assign _0206_ = instr_vld_t0 & decode_t0[20];
assign _0209_ = _0518_ & regwr_pending_later_t0;
assign _0218_ = instr_vld_t0 & decode_t0[15];
assign _0212_ = lsu_rdy_t0 & regwr_lsu_t0;
assign _0215_ = csr_rdy_t0 & regwr_csr_t0;
assign _0223_ = instr_vld_t0 & instr_jump_t0;
assign _0226_ = decode_vld_t0 & _0502_;
assign _0229_ = decode_t0[1] & instr_jump_t0;
assign _0232_ = decode_t0[0] & decode_t0[12];
assign _0235_ = decode_t0[0] & decode_t0[11];
assign _0238_ = decode_vld_t0 & decode_rdy_t0;
assign _0241_ = decode_t0[5] & trap_jump_t0;
assign _0370_ = _0198_ | _0199_;
assign _0371_ = _0201_ | _0202_;
assign _0372_ = _0204_ | _0205_;
assign _0373_ = _0207_ | _0208_;
assign _0374_ = _0210_ | _0211_;
assign _0375_ = _0213_ | _0214_;
assign _0376_ = _0216_ | _0217_;
assign _0377_ = _0211_ | _0219_;
assign _0378_ = _0214_ | _0220_;
assign _0379_ = _0221_ | _0222_;
assign _0380_ = _0224_ | _0225_;
assign _0381_ = _0227_ | _0228_;
assign _0382_ = _0230_ | _0231_;
assign _0383_ = _0233_ | _0234_;
assign _0384_ = _0236_ | _0237_;
assign _0385_ = _0239_ | _0240_;
assign _0514_ = _0370_ | _0200_;
assign instr_vld_t0 = _0371_ | _0203_;
assign basic_rdy_t0 = _0372_ | _0206_;
assign _0520_ = _0373_ | _0209_;
assign _0522_ = _0374_ | _0212_;
assign _0524_ = _0375_ | _0215_;
assign _0526_ = _0376_ | _0218_;
assign _0528_ = _0377_ | _0212_;
assign _0530_ = _0378_ | _0215_;
assign _0532_ = _0379_ | _0223_;
assign _0516_ = _0380_ | _0226_;
assign _0534_ = _0381_ | _0229_;
assign _0536_ = _0382_ | _0232_;
assign _0538_ = _0383_ | _0235_;
assign _0518_ = _0384_ | _0238_;
assign _0540_ = _0385_ | _0241_;
assign _0133_ = | { _0510_, _0516_ };
assign _0134_ = | { _0530_, _0528_, _0526_ };
assign _0141_ = | { _0050_, _0605_, _0512_, _0504_, _0502_, _0510_ };
assign _0144_ = | { activate_trap_t0, return_trap_t0 };
assign _0145_ = | { _0605_, _0510_, activate_trap_t0, return_trap_t0 };
assign _0147_ = | state_t0;
assign _0148_ = | { basic_rdy_t0, lsu_rdy_t0, csr_rdy_t0 };
assign _0068_ = ~ { _0510_, _0516_ };
assign _0069_ = ~ { _0530_, _0528_, _0526_ };
assign _0076_ = ~ { _0050_, _0605_, _0512_, _0510_, _0504_, _0502_ };
assign _0077_ = ~ { return_trap_t0, activate_trap_t0 };
assign _0078_ = ~ { _0605_, _0510_, return_trap_t0, activate_trap_t0 };
assign _0120_ = ~ decode_t0[4:3];
assign _0124_ = ~ { csr_rdy_t0, lsu_rdy_t0, basic_rdy_t0 };
assign _0176_ = { _0509_, _0515_ } & _0068_;
assign _0177_ = { _0529_, _0527_, _0525_ } & _0069_;
assign _0184_ = { _0049_, _0604_, _0511_, _0509_, _0503_, _0501_ } & _0076_;
assign _0185_ = { return_trap, activate_trap } & _0077_;
assign _0186_ = { _0604_, _0509_, return_trap, activate_trap } & _0078_;
assign _0338_ = { csr_rdy, lsu_rdy, basic_rdy } & _0124_;
assign _0149_ = ! _0176_;
assign _0150_ = ! _0177_;
assign _0151_ = ! _0184_;
assign _0152_ = ! _0185_;
assign _0153_ = ! _0186_;
assign _0154_ = ! _0329_;
assign _0155_ = ! _0337_;
assign _0156_ = ! _0338_;
assign _0026_ = _0149_ & _0133_;
assign _0028_ = _0150_ & _0134_;
assign _0042_ = _0151_ & _0141_;
assign _0050_ = _0152_ & _0144_;
assign _0130_ = _0153_ & _0145_;
assign _0506_ = _0154_ & _0146_;
assign _0502_ = _0155_ & _0147_;
assign decode_rdy_t0 = _0156_ & _0148_;
assign _0084_ = ~ decode[12];
assign _0088_ = ~ decode[14];
assign _0090_ = ~ _0531_;
assign _0092_ = ~ decode[2];
assign _0094_ = ~ _0543_;
assign _0086_ = ~ instr_vld;
assign _0085_ = ~ decode[11];
assign _0087_ = ~ _0503_;
assign _0089_ = ~ decode[13];
assign _0091_ = ~ trap_jump;
assign _0093_ = ~ decode[0];
assign _0095_ = ~ _0533_;
assign _0096_ = ~ _0511_;
assign _0098_ = ~ _0539_;
assign _0242_ = decode_t0[12] & _0085_;
assign _0245_ = instr_vld_t0 & _0087_;
assign _0248_ = decode_t0[14] & _0089_;
assign _0251_ = _0532_ & _0091_;
assign _0254_ = decode_t0[2] & _0093_;
assign _0257_ = _0544_ & _0095_;
assign _0260_ = instr_vld_t0 & _0096_;
assign _0263_ = _0518_ & _0098_;
assign _0243_ = decode_t0[11] & _0084_;
assign _0246_ = _0504_ & _0086_;
assign _0249_ = decode_t0[13] & _0088_;
assign _0252_ = trap_jump_t0 & _0090_;
assign _0255_ = decode_t0[0] & _0092_;
assign _0258_ = _0534_ & _0094_;
assign _0261_ = _0512_ & _0086_;
assign _0264_ = _0540_ & _0097_;
assign _0244_ = decode_t0[12] & decode_t0[11];
assign _0247_ = instr_vld_t0 & _0504_;
assign _0250_ = decode_t0[14] & decode_t0[13];
assign _0253_ = _0532_ & trap_jump_t0;
assign _0256_ = decode_t0[2] & decode_t0[0];
assign _0259_ = _0544_ & _0534_;
assign _0262_ = instr_vld_t0 & _0512_;
assign _0265_ = _0518_ & _0540_;
assign _0386_ = _0242_ | _0243_;
assign _0387_ = _0245_ | _0246_;
assign _0388_ = _0248_ | _0249_;
assign _0389_ = _0251_ | _0252_;
assign _0390_ = _0254_ | _0255_;
assign _0391_ = _0257_ | _0258_;
assign _0392_ = _0260_ | _0261_;
assign _0393_ = _0263_ | _0264_;
assign _0542_ = _0386_ | _0244_;
assign lsu_vld_t0 = _0387_ | _0247_;
assign instr_jump_t0 = _0388_ | _0250_;
assign branch_t0 = _0389_ | _0253_;
assign _0544_ = _0390_ | _0256_;
assign exception_t0 = _0391_ | _0259_;
assign csr_vld_t0 = _0392_ | _0262_;
assign _0546_ = _0393_ | _0265_;
assign _0079_ = ~ { _0606_, _0606_, _0606_ };
assign _0080_ = ~ { _0604_, _0604_, _0604_ };
assign _0081_ = ~ { _0503_, _0503_, _0503_ };
assign _0082_ = ~ { _0511_, _0511_, _0511_ };
assign _0083_ = ~ { _0129_, _0129_, _0129_ };
assign _0108_ = ~ { _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_ };
assign _0109_ = ~ { _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_ };
assign _0110_ = ~ { _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_ };
assign _0111_ = ~ { _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_ };
assign _0112_ = ~ { decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2] };
assign _0107_ = ~ { core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt };
assign _0113_ = ~ { _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_ };
assign _0097_ = ~ _0517_;
assign _0114_ = ~ _0529_;
assign _0115_ = ~ _0527_;
assign _0116_ = ~ _0525_;
assign _0117_ = ~ { _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_ };
assign _0118_ = ~ { _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_ };
assign _0119_ = ~ { core_interrupt, core_interrupt, core_interrupt };
assign _0121_ = ~ { decode[5], decode[5], decode[5] };
assign _0122_ = ~ { exception, exception, exception };
assign _0125_ = ~ { trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump };
assign _0363_ = { _0607_, _0607_, _0607_ } | _0079_;
assign _0364_ = { _0605_, _0605_, _0605_ } | _0080_;
assign _0365_ = { _0504_, _0504_, _0504_ } | _0081_;
assign _0366_ = { _0512_, _0512_, _0512_ } | _0082_;
assign _0367_ = { _0130_, _0130_, _0130_ } | _0083_;
assign _0402_ = { _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_ } | _0108_;
assign _0403_ = { _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_ } | _0109_;
assign _0406_ = { _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_ } | _0110_;
assign _0409_ = { _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_ } | _0111_;
assign _0412_ = { decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2] } | _0112_;
assign _0398_ = { core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0 } | _0107_;
assign _0415_ = { _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_ } | _0113_;
assign _0419_ = _0530_ | _0114_;
assign _0420_ = _0528_ | _0115_;
assign _0421_ = _0526_ | _0116_;
assign _0423_ = _0518_ | _0097_;
assign _0428_ = { _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_ } | _0117_;
assign _0431_ = { _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_ } | _0118_;
assign _0434_ = { core_interrupt_t0, core_interrupt_t0, core_interrupt_t0 } | _0119_;
assign _0435_ = { decode_t0[5], decode_t0[5], decode_t0[5] } | _0121_;
assign _0438_ = { exception_t0, exception_t0, exception_t0 } | _0122_;
assign _0440_ = { trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0 } | _0125_;
assign _0368_ = { _0130_, _0130_, _0130_ } | { _0129_, _0129_, _0129_ };
assign _0400_ = { _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_ } | { _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_ };
assign _0401_ = { _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_ } | { _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_ };
assign _0404_ = { _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_ } | { _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_ };
assign _0407_ = { _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_ } | { _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_ };
assign _0410_ = { _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_ } | { _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_ };
assign _0413_ = { decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2] } | { decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2], decode[2] };
assign _0399_ = { core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0 } | { core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt, core_interrupt };
assign _0416_ = { _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_ } | { _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_ };
assign _0424_ = _0518_ | _0517_;
assign _0422_ = _0526_ | _0525_;
assign _0427_ = { _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_, _0530_ } | { _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_ };
assign _0429_ = { _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_ } | { _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_ };
assign _0432_ = { _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_ } | { _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_ };
assign _0436_ = { decode_t0[5], decode_t0[5], decode_t0[5] } | { decode[5], decode[5], decode[5] };
assign _0439_ = { decode_vld_t0, decode_vld_t0, decode_vld_t0 } | { decode_vld, decode_vld, decode_vld };
assign _0441_ = { trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0 } | { trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump, trap_jump };
assign _0187_ = { _0492_[2], _0492_[2], _0492_[2] } & _0363_;
assign _0189_ = _0494_ & _0364_;
assign _0191_ = _0008_ & _0365_;
assign _0193_ = _0498_ & _0366_;
assign _0195_ = _0500_ & _0367_;
assign _0278_ = _0559_ & _0402_;
assign _0280_ = _0561_ & _0403_;
assign _0283_ = _0563_ & _0406_;
assign _0286_ = _0565_ & _0409_;
assign _0289_ = _0567_ & _0412_;
assign _0292_ = _0568_ & _0398_;
assign _0296_ = _0577_ & _0403_;
assign _0298_ = _0579_ & _0406_;
assign _0300_ = _0580_ & _0409_;
assign _0302_ = _0582_ & _0412_;
assign _0304_ = _0584_ & _0398_;
assign _0306_ = _0574_ & _0415_;
assign _0309_ = _0530_ & _0420_;
assign _0311_ = _0589_ & _0421_;
assign _0313_ = regwr_pending_later_t0 & _0423_;
assign _0316_ = _0592_ & _0419_;
assign _0318_ = _0593_ & _0420_;
assign _0320_ = _0595_ & _0421_;
assign _0323_ = _0599_ & _0428_;
assign _0326_ = _0601_ & _0431_;
assign _0330_ = _0018_ & _0435_;
assign _0333_ = _0014_ & _0438_;
assign _0335_ = _0012_ & _0434_;
assign _0339_ = decode_t0[52:21] & _0440_;
assign _0196_ = _0496_ & _0368_;
assign _0559_ = decode_t0[180:149] & _0401_;
assign _0281_ = decode_t0[52:21] & _0404_;
assign _0284_ = decode_t0[52:21] & _0407_;
assign _0287_ = decode_t0[52:21] & _0410_;
assign _0290_ = decode_t0[148:117] & _0413_;
assign _0294_ = _0570_ & _0416_;
assign _0574_ = _0572_ & _0400_;
assign _0572_ = { 28'h0000000, core_interrupt_cause_t0 } & _0399_;
assign _0307_ = _0586_ & _0416_;
assign _0314_ = _0556_ & _0424_;
assign _0321_ = _0592_ & _0422_;
assign _0599_ = csr_data_t0 & _0427_;
assign _0324_ = load_data_t0 & _0429_;
assign _0327_ = result_t0 & _0432_;
assign _0331_ = _0016_ & _0436_;
assign _0008_ = _0010_ & _0439_;
assign _0340_ = trap_handle_t0 & _0441_;
assign _0369_ = _0195_ | _0196_;
assign _0405_ = _0280_ | _0281_;
assign _0408_ = _0283_ | _0284_;
assign _0411_ = _0286_ | _0287_;
assign _0414_ = _0289_ | _0290_;
assign _0417_ = _0304_ | _0572_;
assign _0418_ = _0306_ | _0307_;
assign _0425_ = _0313_ | _0314_;
assign _0426_ = _0320_ | _0321_;
assign _0430_ = _0323_ | _0324_;
assign _0433_ = _0326_ | _0327_;
assign _0437_ = _0330_ | _0331_;
assign _0442_ = _0339_ | _0340_;
assign _0448_ = _0493_ ^ _0006_;
assign _0449_ = _0007_ ^ _0020_;
assign _0450_ = _0497_ ^ _0004_;
assign _0451_ = _0499_ ^ _0495_;
assign _0453_ = _0560_ ^ decode[52:21];
assign _0454_ = _0562_ ^ decode[52:21];
assign _0455_ = _0564_ ^ decode[52:21];
assign _0456_ = _0566_ ^ decode[148:117];
assign _0458_ = _0558_ ^ _0569_;
assign _0464_ = _0583_ ^ { 28'h8000000, core_interrupt_cause };
assign _0465_ = _0573_ ^ _0585_;
assign _0466_ = regwr_pending_later ^ _0555_;
assign _0469_ = _0594_ ^ _0467_;
assign _0470_ = _0598_ ^ load_data;
assign _0471_ = _0600_ ^ result;
assign _0472_ = _0017_ ^ _0015_;
assign _0473_ = decode[52:21] ^ trap_handle;
assign _0188_ = { _0607_, _0607_, _0607_ } & { _0056_[1], _0447_[1], _0056_[0] };
assign _0494_ = { _0050_, _0050_, _0050_ } & { _0059_, _0005_[0] };
assign _0190_ = { _0605_, _0605_, _0605_ } & _0448_;
assign _0192_ = { _0504_, _0504_, _0504_ } & _0449_;
assign _0194_ = { _0512_, _0512_, _0512_ } & _0450_;
assign _0197_ = { _0130_, _0130_, _0130_ } & _0451_;
assign _0279_ = { _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_ } & _0452_;
assign _0282_ = { _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_ } & _0453_;
assign _0285_ = { _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_ } & _0454_;
assign _0288_ = { _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_ } & _0455_;
assign _0291_ = { decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2] } & _0456_;
assign _0293_ = { core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0 } & _0457_;
assign _0295_ = { _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_ } & _0458_;
assign _0577_ = { _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_ } & { _0459_[31:4], _0051_[2], _0459_[2], _0051_[1:0] };
assign _0297_ = { _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_, _0538_ } & { _0460_[31:3], _0052_, _0460_[0] };
assign _0299_ = { _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_, _0536_ } & { _0461_[31:3], _0053_, _0461_[1:0] };
assign _0301_ = { _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_, _0534_ } & _0462_;
assign _0303_ = { decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2], decode_t0[2] } & { _0463_[31:2], _0054_, _0463_[0] };
assign _0305_ = { core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0, core_interrupt_t0 } & _0464_;
assign _0308_ = { _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_ } & _0465_;
assign _0310_ = _0528_ & _0060_;
assign _0312_ = _0526_ & _0061_;
assign _0315_ = _0518_ & _0466_;
assign _0317_ = _0530_ & _0467_;
assign _0319_ = _0528_ & _0468_;
assign _0322_ = _0526_ & _0469_;
assign _0325_ = { _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_, _0528_ } & _0470_;
assign _0328_ = { _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_ } & _0471_;
assign _0018_ = { _0542_, _0542_, _0542_ } & { _0019_[2:1], _0055_ };
assign _0332_ = { decode_t0[5], decode_t0[5], decode_t0[5] } & _0472_;
assign _0334_ = { exception_t0, exception_t0, exception_t0 } & { _0013_[2], _0057_ };
assign _0336_ = { core_interrupt_t0, core_interrupt_t0, core_interrupt_t0 } & { _0011_[2], _0058_ };
assign _0341_ = { trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0, trap_jump_t0 } & _0473_;
assign _0016_ = _0188_ | _0187_;
assign _0496_ = _0190_ | _0189_;
assign _0498_ = _0192_ | _0191_;
assign _0500_ = _0194_ | _0193_;
assign next_state_t0 = _0197_ | _0369_;
assign _0561_ = _0279_ | _0278_;
assign _0563_ = _0282_ | _0405_;
assign _0565_ = _0285_ | _0408_;
assign _0567_ = _0288_ | _0411_;
assign _0568_ = _0291_ | _0414_;
assign _0570_ = _0293_ | _0292_;
assign _0003_ = _0295_ | _0294_;
assign _0579_ = _0297_ | _0296_;
assign _0580_ = _0299_ | _0298_;
assign _0582_ = _0301_ | _0300_;
assign _0584_ = _0303_ | _0302_;
assign _0586_ = _0305_ | _0417_;
assign _0001_ = _0308_ | _0418_;
assign _0589_ = _0310_ | _0309_;
assign _0591_ = _0312_ | _0311_;
assign _0592_ = _0315_ | _0425_;
assign _0593_ = _0317_ | _0316_;
assign _0595_ = _0319_ | _0318_;
assign _0597_ = _0322_ | _0426_;
assign _0601_ = _0325_ | _0430_;
assign _0603_ = _0328_ | _0433_;
assign _0014_ = _0332_ | _0437_;
assign _0012_ = _0334_ | _0333_;
assign _0010_ = _0336_ | _0335_;
assign branch_target_t0 = _0341_ | _0442_;
assign _0021_ = { _0507_, _0505_, _0537_, _0535_, _0533_, _0515_, core_interrupt, decode[2] } != 8'h04;
assign _0023_ = { _0509_, _0515_, core_interrupt } != 3'h4;
assign _0025_ = | { _0509_, _0515_ };
assign _0027_ = | { _0529_, _0527_, _0525_ };
assign _0029_ = { _0501_, _0541_, exception, core_interrupt, decode_vld, decode[6:5] } != 7'h44;
assign _0031_ = { _0501_, decode_vld } != 2'h2;
assign _0033_ = { _0503_, lsu_rdy } != 2'h2;
assign _0035_ = { _0511_, csr_rdy } != 2'h2;
assign _0037_ = { _0509_, core_interrupt } != 2'h2;
assign _0039_ = { _0604_, trap_jump } != 2'h2;
assign _0041_ = | { _0049_, _0604_, _0511_, _0509_, _0503_, _0501_ };
assign _0043_ = & { _0025_, _0023_, _0021_ };
assign _0045_ = & { _0027_, rstz };
assign _0047_ = & { _0029_, _0031_, _0033_, _0035_, _0037_, _0039_, _0041_ };
assign _0060_ = ~ _0587_;
assign _0061_ = ~ _0588_;
assign _0051_ = ~ { _0575_[3], _0575_[1:0] };
assign _0052_ = ~ _0576_[2:1];
assign _0053_ = ~ _0578_[2];
assign _0054_ = ~ _0581_[1];
assign _0055_ = ~ _0019_[0];
assign _0056_ = ~ { _0491_[2], _0491_[0] };
assign _0057_ = ~ _0013_[1:0];
assign _0058_ = ~ _0011_[1:0];
assign _0059_ = ~ _0005_[2:1];
assign _0049_ = | { return_trap, activate_trap };
assign _0099_ = ~ decode[15];
assign _0101_ = ~ _0551_;
assign _0103_ = ~ regwr_pending_firstcycle;
assign _0105_ = ~ _0521_;
assign _0100_ = ~ regwr_lsu;
assign _0102_ = ~ regwr_csr;
assign _0104_ = ~ _0519_;
assign _0106_ = ~ _0523_;
assign _0266_ = decode_t0[15] & _0100_;
assign _0269_ = _0552_ & _0102_;
assign _0272_ = regwr_pending_firstcycle_t0 & _0104_;
assign _0275_ = _0522_ & _0106_;
assign _0267_ = regwr_lsu_t0 & _0099_;
assign _0270_ = regwr_csr_t0 & _0101_;
assign _0273_ = _0520_ & _0103_;
assign _0276_ = _0524_ & _0105_;
assign _0268_ = decode_t0[15] & regwr_lsu_t0;
assign _0271_ = _0552_ & regwr_csr_t0;
assign _0274_ = regwr_pending_firstcycle_t0 & _0520_;
assign _0277_ = _0522_ & _0524_;
assign _0394_ = _0266_ | _0267_;
assign _0395_ = _0269_ | _0270_;
assign _0396_ = _0272_ | _0273_;
assign _0397_ = _0275_ | _0276_;
assign _0552_ = _0394_ | _0268_;
assign _0554_ = _0395_ | _0271_;
assign regwr_pending_t0 = _0396_ | _0274_;
assign _0556_ = _0397_ | _0277_;
assign _0129_ = | { _0604_, _0509_, return_trap, activate_trap };
assign { _0491_[2], _0447_[1], _0491_[0] } = _0608_ ? 3'h4 : 3'h3;
assign _0015_ = _0606_ ? 3'h5 : { _0491_[2], _0447_[1], _0491_[0] };
assign _0493_ = _0049_ ? 3'h6 : _0005_;
assign _0495_ = _0604_ ? _0006_ : _0493_;
assign _0497_ = _0503_ ? _0020_ : _0007_;
assign _0499_ = _0511_ ? _0004_ : _0497_;
assign next_state = _0129_ ? _0495_ : _0499_;
assign _0142_ = | { _0026_, _0024_, _0022_ };
assign _0143_ = | { _0042_, _0040_, _0038_, _0036_, _0034_, _0032_, _0030_ };
assign _0360_ = { _0025_, _0023_, _0021_ } | { _0026_, _0024_, _0022_ };
assign _0361_ = { _0027_, rstz } | { _0028_, 1'h0 };
assign _0362_ = { _0029_, _0031_, _0033_, _0035_, _0037_, _0039_, _0041_ } | { _0030_, _0032_, _0034_, _0036_, _0038_, _0040_, _0042_ };
assign _0126_ = & _0360_;
assign _0127_ = & _0361_;
assign _0128_ = & _0362_;
assign _0044_ = _0142_ & _0126_;
assign _0046_ = _0028_ & _0127_;
assign _0048_ = _0143_ & _0128_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_9e9afc4272f55a9beacc  */
/* PC_TAINT_INFO STATE_NAME regwr_en_t0 */
always_ff @(posedge clk)
if (!rstz) regwr_en_t0 <= 1'h0;
else regwr_en_t0 <= _0591_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_9e9afc4272f55a9beacc  */
/* PC_TAINT_INFO STATE_NAME regwr_pending_later_t0 */
always_ff @(posedge clk)
if (!rstz) regwr_pending_later_t0 <= 1'h0;
else regwr_pending_later_t0 <= _0597_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_9e9afc4272f55a9beacc  */
/* PC_TAINT_INFO STATE_NAME instret_t0 */
always_ff @(posedge clk)
if (!rstz) instret_t0 <= 1'h0;
else instret_t0 <= _0546_;
assign _0065_ = ~ _0047_;
assign _0446_ = next_state ^ state;
assign _0356_ = next_state_t0 | state_t0;
assign _0357_ = _0446_ | _0356_;
assign _0171_ = { _0047_, _0047_, _0047_ } & next_state_t0;
assign _0172_ = { _0065_, _0065_, _0065_ } & state_t0;
assign _0173_ = _0357_ & { _0048_, _0048_, _0048_ };
assign _0358_ = _0171_ | _0172_;
assign _0359_ = _0358_ | _0173_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_9e9afc4272f55a9beacc  */
/* PC_TAINT_INFO STATE_NAME state_t0 */
always_ff @(posedge clk)
if (!rstz) state_t0 <= 3'h0;
else state_t0 <= _0359_;
assign _0513_ = _0515_ && /* src = "generated/sv2v_out.v:708.22-708.67" */ _0547_;
assign instr_vld = _0513_ && /* src = "generated/sv2v_out.v:708.21-708.87" */ _0548_;
assign basic_rdy = instr_vld && /* src = "generated/sv2v_out.v:709.21-709.44" */ decode[20];
assign _0519_ = _0097_ && /* src = "generated/sv2v_out.v:733.53-733.103" */ regwr_pending_later;
assign _0521_ = regwr_lsu && /* src = "generated/sv2v_out.v:742.29-742.50" */ _0549_;
assign _0523_ = regwr_csr && /* src = "generated/sv2v_out.v:742.55-742.76" */ _0550_;
assign _0525_ = instr_vld && /* src = "generated/sv2v_out.v:743.8-743.31" */ decode[15];
assign _0527_ = lsu_rdy && /* src = "generated/sv2v_out.v:747.13-747.33" */ regwr_lsu;
assign _0529_ = csr_rdy && /* src = "generated/sv2v_out.v:752.13-752.33" */ regwr_csr;
assign _0531_ = instr_vld && /* src = "generated/sv2v_out.v:762.19-762.42" */ instr_jump;
assign _0515_ = decode_vld && /* src = "generated/sv2v_out.v:771.7-771.36" */ _0501_;
assign _0533_ = decode[1] && /* src = "generated/sv2v_out.v:780.13-780.36" */ instr_jump;
assign _0535_ = decode[0] && /* src = "generated/sv2v_out.v:784.13-784.36" */ decode[12];
assign _0537_ = decode[0] && /* src = "generated/sv2v_out.v:788.13-788.36" */ decode[11];
assign _0517_ = decode_vld && /* src = "generated/sv2v_out.v:838.16-838.40" */ decode_rdy;
assign _0539_ = decode[5] && /* src = "generated/sv2v_out.v:838.46-838.68" */ trap_jump;
assign _0541_ = decode[12] || /* src = "generated/sv2v_out.v:688.15-688.39" */ decode[11];
assign lsu_vld = instr_vld || /* src = "generated/sv2v_out.v:717.19-717.47" */ _0503_;
assign instr_jump = decode[14] || /* src = "generated/sv2v_out.v:761.22-761.46" */ decode[13];
assign branch = _0531_ || /* src = "generated/sv2v_out.v:762.18-762.56" */ trap_jump;
assign _0543_ = decode[2] || /* src = "generated/sv2v_out.v:763.22-763.44" */ decode[0];
assign exception = _0543_ || /* src = "generated/sv2v_out.v:763.21-763.74" */ _0533_;
assign csr_vld = instr_vld || /* src = "generated/sv2v_out.v:806.19-806.47" */ _0511_;
assign _0545_ = _0517_ || /* src = "generated/sv2v_out.v:838.15-838.69" */ _0539_;
assign _0547_ = ~ /* src = "generated/sv2v_out.v:708.57-708.67" */ exception;
assign _0548_ = ~ /* src = "generated/sv2v_out.v:708.72-708.87" */ core_interrupt;
assign _0549_ = ~ /* src = "generated/sv2v_out.v:742.42-742.50" */ lsu_rdy;
assign _0550_ = ~ /* src = "generated/sv2v_out.v:742.68-742.76" */ csr_rdy;
assign _0551_ = decode[15] | /* src = "generated/sv2v_out.v:732.67-732.89" */ regwr_lsu;
assign _0553_ = _0551_ | /* src = "generated/sv2v_out.v:732.66-732.102" */ regwr_csr;
assign regwr_pending = regwr_pending_firstcycle | /* src = "generated/sv2v_out.v:733.25-733.104" */ _0519_;
assign _0555_ = _0521_ | /* src = "generated/sv2v_out.v:742.28-742.77" */ _0523_;
assign _0557_ = core_interrupt ? /* src = "generated/sv2v_out.v:802.8-802.22|generated/sv2v_out.v:802.4-805.7" */ 32'd0 : 32'hxxxxxxxx;
assign _0558_ = _0509_ ? /* src = "generated/sv2v_out.v:801.12-801.25|generated/sv2v_out.v:801.8-805.7" */ _0557_ : 32'hxxxxxxxx;
assign _0452_ = _0507_ ? /* src = "generated/sv2v_out.v:796.13-796.48|generated/sv2v_out.v:796.9-799.7" */ decode[180:149] : 32'hxxxxxxxx;
assign _0560_ = _0505_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:792.13-792.47|generated/sv2v_out.v:792.9-799.7" */ 32'd0 : _0452_;
assign _0562_ = _0537_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:788.13-788.36|generated/sv2v_out.v:788.9-799.7" */ decode[52:21] : _0560_;
assign _0564_ = _0535_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:784.13-784.36|generated/sv2v_out.v:784.9-799.7" */ decode[52:21] : _0562_;
assign _0566_ = _0533_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:780.13-780.36|generated/sv2v_out.v:780.9-799.7" */ decode[52:21] : _0564_;
assign _0457_ = decode[2] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:776.13-776.22|generated/sv2v_out.v:776.9-799.7" */ decode[148:117] : _0566_;
assign _0569_ = core_interrupt ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:772.8-772.22|generated/sv2v_out.v:772.4-799.7" */ 32'd0 : _0457_;
assign _0002_ = _0515_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:771.7-771.36|generated/sv2v_out.v:771.3-805.7" */ _0569_ : _0558_;
assign _0571_ = core_interrupt ? /* src = "generated/sv2v_out.v:802.8-802.22|generated/sv2v_out.v:802.4-805.7" */ { 28'h8000000, core_interrupt_cause } : 32'hxxxxxxxx;
assign _0573_ = _0509_ ? /* src = "generated/sv2v_out.v:801.12-801.25|generated/sv2v_out.v:801.8-805.7" */ _0571_ : 32'hxxxxxxxx;
assign { _0459_[31:4], _0575_[3], _0459_[2], _0575_[1:0] } = _0507_ ? /* src = "generated/sv2v_out.v:796.13-796.48|generated/sv2v_out.v:796.9-799.7" */ 32'd3 : 32'hxxxxxxxx;
assign { _0460_[31:3], _0576_[2:1], _0460_[0] } = _0505_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:792.13-792.47|generated/sv2v_out.v:792.9-799.7" */ 32'd11 : { _0459_[31:4], _0575_[3], _0459_[2], _0575_[1:0] };
assign { _0461_[31:3], _0578_[2], _0461_[1:0] } = _0537_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:788.13-788.36|generated/sv2v_out.v:788.9-799.7" */ 32'd6 : { _0460_[31:3], _0576_[2:1], _0460_[0] };
assign _0462_ = _0535_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:784.13-784.36|generated/sv2v_out.v:784.9-799.7" */ 32'd4 : { _0461_[31:3], _0578_[2], _0461_[1:0] };
assign { _0463_[31:2], _0581_[1], _0463_[0] } = _0533_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:780.13-780.36|generated/sv2v_out.v:780.9-799.7" */ 32'd0 : _0462_;
assign _0583_ = decode[2] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:776.13-776.22|generated/sv2v_out.v:776.9-799.7" */ 32'd2 : { _0463_[31:2], _0581_[1], _0463_[0] };
assign _0585_ = core_interrupt ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:772.8-772.22|generated/sv2v_out.v:772.4-799.7" */ { 28'h8000000, core_interrupt_cause } : _0583_;
assign _0000_ = _0515_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:771.7-771.36|generated/sv2v_out.v:771.3-805.7" */ _0585_ : _0573_;
assign _0587_ = _0529_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:752.13-752.33|generated/sv2v_out.v:752.9-758.22" */ 1'h1 : 1'h0;
assign _0588_ = _0527_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:747.13-747.33|generated/sv2v_out.v:747.9-758.22" */ 1'h1 : _0587_;
assign _0590_ = _0525_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:743.8-743.31|generated/sv2v_out.v:743.4-758.22" */ 1'h1 : _0588_;
assign _0467_ = _0517_ ? /* src = "generated/sv2v_out.v:741.8-741.32|generated/sv2v_out.v:741.4-742.78" */ _0555_ : regwr_pending_later;
assign _0468_ = _0529_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:752.13-752.33|generated/sv2v_out.v:752.9-758.22" */ 1'h0 : _0467_;
assign _0594_ = _0527_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:747.13-747.33|generated/sv2v_out.v:747.9-758.22" */ 1'h0 : _0468_;
assign _0596_ = _0525_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:743.8-743.31|generated/sv2v_out.v:743.4-758.22" */ _0467_ : _0594_;
assign _0598_ = _0529_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:752.13-752.33|generated/sv2v_out.v:752.9-758.22" */ csr_data : 32'hxxxxxxxx;
assign _0600_ = _0527_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:747.13-747.33|generated/sv2v_out.v:747.9-758.22" */ load_data : _0598_;
assign _0602_ = _0525_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:743.8-743.31|generated/sv2v_out.v:743.4-758.22" */ result : _0600_;
assign _0006_ = trap_jump ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:704.9-704.18|generated/sv2v_out.v:704.5-705.24" */ 3'h0 : 3'hx;
assign _0005_ = core_interrupt ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:699.9-699.23|generated/sv2v_out.v:699.5-700.24" */ 3'h3 : 3'hx;
assign _0004_ = csr_rdy ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:696.9-696.16|generated/sv2v_out.v:696.5-697.24" */ 3'h0 : 3'hx;
assign _0020_ = lsu_rdy ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:693.9-693.16|generated/sv2v_out.v:693.5-694.24" */ 3'h0 : 3'hx;
assign _0019_ = decode[6] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:690.15-690.24|generated/sv2v_out.v:690.11-691.25" */ 3'h2 : 3'hx;
assign _0017_ = _0541_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:688.15-688.39|generated/sv2v_out.v:688.11-691.25" */ 3'h1 : _0019_;
assign _0606_ = decode[4:3] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:683.7-687.14" */ 2'h3;
assign _0608_ = decode[4:3] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:683.7-687.14" */ 2'h2;
assign _0505_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:683.7-687.14" */ decode[4:3];
assign _0507_ = decode[4:3] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:683.7-687.14" */ 2'h1;
assign _0013_ = decode[5] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:682.15-682.24|generated/sv2v_out.v:682.11-691.25" */ _0015_ : _0017_;
assign _0011_ = exception ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:680.15-680.24|generated/sv2v_out.v:680.11-691.25" */ 3'h3 : _0013_;
assign _0009_ = core_interrupt ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:678.10-678.24|generated/sv2v_out.v:678.6-691.25" */ 3'h3 : _0011_;
assign _0007_ = decode_vld ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:677.9-677.19|generated/sv2v_out.v:677.5-691.25" */ _0009_ : 3'hx;
assign _0604_ = state == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:675.3-706.10" */ 3'h6;
assign return_trap = state == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:675.3-706.10" */ 3'h4;
assign activate_trap = state == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:675.3-706.10" */ 3'h3;
assign _0509_ = state == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:675.3-706.10" */ 3'h5;
assign _0511_ = state == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:675.3-706.10" */ 3'h2;
assign _0503_ = state == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:675.3-706.10" */ 3'h1;
assign _0501_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:675.3-706.10" */ state;
assign decode_rdy = | /* src = "generated/sv2v_out.v:710.22-710.52" */ { csr_rdy, lsu_rdy, basic_rdy };
assign branch_target = trap_jump ? /* src = "generated/sv2v_out.v:760.26-760.66" */ trap_handle : decode[52:21];
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:711.13-716.3" */
kronos_alu u_alu (
.aluop(decode[19:16]),
.aluop_t0(decode_t0[19:16]),
.op1(decode[116:85]),
.op1_t0(decode_t0[116:85]),
.op2(decode[84:53]),
.op2_t0(decode_t0[84:53]),
.result(result),
.result_t0(result_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:811.4-831.3" */
paramodsimplif_23175af27fd2ffc5d196  u_csr (
.activate_trap(activate_trap),
.activate_trap_t0(activate_trap_t0),
.clk(clk),
.clk_t0(clk_t0),
.core_interrupt(core_interrupt),
.core_interrupt_cause(core_interrupt_cause),
.core_interrupt_cause_t0(core_interrupt_cause_t0),
.core_interrupt_t0(core_interrupt_t0),
.csr_data(csr_data),
.csr_data_t0(csr_data_t0),
.csr_rdy(csr_rdy),
.csr_rdy_t0(csr_rdy_t0),
.csr_vld(csr_vld),
.csr_vld_t0(csr_vld_t0),
.decode(decode),
.decode_t0(decode_t0),
.external_interrupt(external_interrupt),
.external_interrupt_t0(external_interrupt_t0),
.instret(instret),
.instret_t0(instret_t0),
.regwr_csr(regwr_csr),
.regwr_csr_t0(regwr_csr_t0),
.return_trap(return_trap),
.return_trap_t0(return_trap_t0),
.rstz(rstz),
.software_interrupt(software_interrupt),
.software_interrupt_t0(software_interrupt_t0),
.timer_interrupt(timer_interrupt),
.timer_interrupt_t0(timer_interrupt_t0),
.trap_cause(trap_cause),
.trap_cause_t0(trap_cause_t0),
.trap_handle(trap_handle),
.trap_handle_t0(trap_handle_t0),
.trap_jump(trap_jump),
.trap_jump_t0(trap_jump_t0),
.trap_value(trap_value),
.trap_value_t0(trap_value_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:718.13-731.3" */
kronos_lsu u_lsu (
.data_ack(data_ack),
.data_ack_t0(data_ack_t0),
.data_addr(data_addr),
.data_addr_t0(data_addr_t0),
.data_mask(data_mask),
.data_mask_t0(data_mask_t0),
.data_rd_data(data_rd_data),
.data_rd_data_t0(data_rd_data_t0),
.data_req(data_req),
.data_req_t0(data_req_t0),
.data_wr_data(data_wr_data),
.data_wr_data_t0(data_wr_data_t0),
.data_wr_en(data_wr_en),
.data_wr_en_t0(data_wr_en_t0),
.decode(decode),
.decode_t0(decode_t0),
.load_data(load_data),
.load_data_t0(load_data_t0),
.lsu_rdy(lsu_rdy),
.lsu_rdy_t0(lsu_rdy_t0),
.lsu_vld(lsu_vld),
.lsu_vld_t0(lsu_vld_t0),
.regwr_lsu(regwr_lsu),
.regwr_lsu_t0(regwr_lsu_t0)
);
assign { _0447_[2], _0447_[0] } = _0056_;
assign { _0459_[3], _0459_[1:0] } = _0051_;
assign _0460_[2:1] = _0052_;
assign _0461_[2] = _0053_;
assign _0463_[1] = _0054_;
assign _0491_[1] = _0447_[1];
assign _0492_[1:0] = { _0492_[2], _0492_[2] };
assign { _0575_[31:4], _0575_[2] } = { _0459_[31:4], _0459_[2] };
assign { _0576_[31:3], _0576_[0] } = { _0460_[31:3], _0460_[0] };
assign { _0578_[31:3], _0578_[1:0] } = { _0461_[31:3], _0461_[1:0] };
assign { _0581_[31:2], _0581_[0] } = { _0463_[31:2], _0463_[0] };
// Added block to randomize initial values.
`ifdef RANDOMIZE_INIT
  initial begin
    trap_cause_t0 = '0;
    regwr_data_t0 = '0;
    regwr_sel_t0 = '0;
    trap_value_t0 = '0;
    regwr_en = '0;
    trap_cause = '0;
    regwr_pending_later = '0;
    regwr_data = '0;
    regwr_sel = '0;
    instret = '0;
    trap_value = '0;
    state = '0;
    regwr_en_t0 = '0;
    regwr_pending_later_t0 = '0;
    instret_t0 = '0;
    state_t0 = '0;
  end
`endif // RANDOMIZE_INIT
endmodule

module paramodsimplif_23175af27fd2ffc5d196 (clk, rstz, decode, csr_vld, csr_rdy, csr_data, regwr_csr, instret, activate_trap, return_trap, trap_cause, trap_value, trap_handle, trap_jump, software_interrupt, timer_interrupt, external_interrupt, core_interrupt, core_interrupt_cause, clk_t0, trap_value_t0
, trap_jump_t0, trap_handle_t0, trap_cause_t0, timer_interrupt_t0, software_interrupt_t0, return_trap_t0, regwr_csr_t0, instret_t0, external_interrupt_t0, decode_t0, csr_vld_t0, csr_rdy_t0, csr_data_t0, core_interrupt_cause_t0, core_interrupt_t0, activate_trap_t0);
/* src = "generated/sv2v_out.v:407.2-418.5" */
wire [1:0] _0000_;
/* src = "generated/sv2v_out.v:407.2-418.5" */
wire [1:0] _0001_;
/* src = "generated/sv2v_out.v:495.39-495.58" */
wire [31:0] _0002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:495.39-495.58" */
wire [31:0] _0003_;
/* src = "generated/sv2v_out.v:539.15-539.46" */
wire _0004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:539.15-539.46" */
wire _0005_;
/* src = "generated/sv2v_out.v:539.14-539.56" */
wire _0006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:539.14-539.56" */
wire _0007_;
/* src = "generated/sv2v_out.v:540.15-540.43" */
wire _0008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:540.15-540.43" */
wire _0009_;
/* src = "generated/sv2v_out.v:540.14-540.53" */
wire _0010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:540.14-540.53" */
wire _0011_;
/* src = "generated/sv2v_out.v:541.15-541.46" */
wire _0012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:541.15-541.46" */
wire _0013_;
/* src = "generated/sv2v_out.v:541.14-541.56" */
wire _0014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:541.14-541.56" */
wire _0015_;
wire _0016_;
/* cellift = 32'd1 */
wire _0017_;
wire _0018_;
/* cellift = 32'd1 */
wire _0019_;
wire _0020_;
/* cellift = 32'd1 */
wire _0021_;
wire _0022_;
/* cellift = 32'd1 */
wire _0023_;
wire _0024_;
/* cellift = 32'd1 */
wire _0025_;
wire _0026_;
/* cellift = 32'd1 */
wire _0027_;
wire _0028_;
/* cellift = 32'd1 */
wire _0029_;
wire _0030_;
/* cellift = 32'd1 */
wire _0031_;
wire _0032_;
/* cellift = 32'd1 */
wire _0033_;
wire _0034_;
/* cellift = 32'd1 */
wire _0035_;
wire _0036_;
/* cellift = 32'd1 */
wire _0037_;
wire _0038_;
/* cellift = 32'd1 */
wire _0039_;
wire _0040_;
/* cellift = 32'd1 */
wire _0041_;
wire _0042_;
/* cellift = 32'd1 */
wire _0043_;
wire _0044_;
/* cellift = 32'd1 */
wire _0045_;
wire _0046_;
/* cellift = 32'd1 */
wire _0047_;
wire _0048_;
/* cellift = 32'd1 */
wire _0049_;
wire _0050_;
/* cellift = 32'd1 */
wire _0051_;
wire _0052_;
/* cellift = 32'd1 */
wire _0053_;
wire _0054_;
/* cellift = 32'd1 */
wire _0055_;
wire _0056_;
/* cellift = 32'd1 */
wire _0057_;
wire _0058_;
/* cellift = 32'd1 */
wire _0059_;
wire _0060_;
wire [1:0] _0061_;
wire _0062_;
wire _0063_;
wire _0064_;
wire _0065_;
wire _0066_;
wire _0067_;
wire _0068_;
wire _0069_;
wire _0070_;
wire _0071_;
wire _0072_;
wire _0073_;
wire _0074_;
wire _0075_;
wire [2:0] _0076_;
wire [2:0] _0077_;
wire [1:0] _0078_;
wire [1:0] _0079_;
wire [1:0] _0080_;
wire [1:0] _0081_;
wire [1:0] _0082_;
wire [1:0] _0083_;
wire [1:0] _0084_;
wire [2:0] _0085_;
wire [1:0] _0086_;
wire [1:0] _0087_;
wire _0088_;
wire _0089_;
wire _0090_;
wire _0091_;
wire _0092_;
wire _0093_;
wire [3:0] _0094_;
wire [2:0] _0095_;
wire [2:0] _0096_;
wire [5:0] _0097_;
wire [31:0] _0098_;
wire [31:0] _0099_;
wire [18:0] _0100_;
wire [18:0] _0101_;
wire [18:0] _0102_;
wire [18:0] _0103_;
wire [18:0] _0104_;
wire [18:0] _0105_;
wire [18:0] _0106_;
wire [18:0] _0107_;
wire [2:0] _0108_;
wire [2:0] _0109_;
wire [2:0] _0110_;
wire [2:0] _0111_;
wire [2:0] _0112_;
wire [2:0] _0113_;
wire [2:0] _0114_;
wire [2:0] _0115_;
wire _0116_;
wire _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire [1:0] _0125_;
wire [2:0] _0126_;
wire [4:0] _0127_;
wire _0128_;
wire _0129_;
wire [4:0] _0130_;
wire [31:0] _0131_;
wire [31:0] _0132_;
wire _0133_;
wire _0134_;
wire [31:0] _0135_;
wire [31:0] _0136_;
wire [1:0] _0137_;
wire [11:0] _0138_;
wire [1:0] _0139_;
wire [31:0] _0140_;
wire _0141_;
wire _0142_;
wire _0143_;
wire _0144_;
wire _0145_;
wire _0146_;
wire _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
/* cellift = 32'd1 */
wire _0152_;
wire _0153_;
/* cellift = 32'd1 */
wire _0154_;
wire _0155_;
/* cellift = 32'd1 */
wire _0156_;
wire _0157_;
/* cellift = 32'd1 */
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire _0186_;
wire _0187_;
wire _0188_;
wire _0189_;
wire _0190_;
wire _0191_;
wire _0192_;
wire _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire _0199_;
wire _0200_;
wire _0201_;
wire [31:0] _0202_;
wire [31:0] _0203_;
wire [31:0] _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
wire _0221_;
wire _0222_;
wire _0223_;
wire _0224_;
wire _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire [1:0] _0231_;
wire [1:0] _0232_;
wire [1:0] _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire _0241_;
wire _0242_;
wire [29:0] _0243_;
wire [29:0] _0244_;
wire [29:0] _0245_;
wire [31:0] _0246_;
wire [31:0] _0247_;
wire [31:0] _0248_;
wire [31:0] _0249_;
wire [31:0] _0250_;
wire [31:0] _0251_;
wire [31:0] _0252_;
wire [31:0] _0253_;
wire [31:0] _0254_;
wire [31:0] _0255_;
wire [31:0] _0256_;
wire [31:0] _0257_;
wire [31:0] _0258_;
wire [31:0] _0259_;
wire [31:0] _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire [1:0] _0264_;
wire [1:0] _0265_;
wire [1:0] _0266_;
wire [29:0] _0267_;
wire [29:0] _0268_;
wire [29:0] _0269_;
wire [1:0] _0270_;
wire [1:0] _0271_;
wire [1:0] _0272_;
wire [2:0] _0273_;
wire [2:0] _0274_;
wire [1:0] _0275_;
wire [1:0] _0276_;
wire [1:0] _0277_;
wire [1:0] _0278_;
wire [1:0] _0279_;
wire [1:0] _0280_;
wire [1:0] _0281_;
wire [2:0] _0282_;
wire [1:0] _0283_;
wire [1:0] _0284_;
wire _0285_;
wire _0286_;
wire _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire [3:0] _0294_;
wire [2:0] _0295_;
wire [2:0] _0296_;
wire [5:0] _0297_;
wire [31:0] _0298_;
wire [31:0] _0299_;
wire [31:0] _0300_;
wire [31:0] _0301_;
wire [31:0] _0302_;
wire [31:0] _0303_;
wire [18:0] _0304_;
wire [18:0] _0305_;
wire [18:0] _0306_;
wire [18:0] _0307_;
wire [18:0] _0308_;
wire [18:0] _0309_;
wire [18:0] _0310_;
wire [18:0] _0311_;
wire [18:0] _0312_;
wire [18:0] _0313_;
wire [18:0] _0314_;
wire [18:0] _0315_;
wire [18:0] _0316_;
wire [18:0] _0317_;
wire [18:0] _0318_;
wire [18:0] _0319_;
wire [18:0] _0320_;
wire [18:0] _0321_;
wire [18:0] _0322_;
wire [18:0] _0323_;
wire [18:0] _0324_;
wire [18:0] _0325_;
wire [18:0] _0326_;
wire [18:0] _0327_;
wire [18:0] _0328_;
wire [18:0] _0329_;
wire [2:0] _0330_;
wire [2:0] _0331_;
wire [2:0] _0332_;
wire [2:0] _0333_;
wire [2:0] _0334_;
wire [2:0] _0335_;
wire [2:0] _0336_;
wire [2:0] _0337_;
wire [2:0] _0338_;
wire [2:0] _0339_;
wire [2:0] _0340_;
wire [2:0] _0341_;
wire [2:0] _0342_;
wire [2:0] _0343_;
wire [2:0] _0344_;
wire [2:0] _0345_;
wire [2:0] _0346_;
wire [2:0] _0347_;
wire [2:0] _0348_;
wire [2:0] _0349_;
wire [2:0] _0350_;
wire [2:0] _0351_;
wire [2:0] _0352_;
wire [2:0] _0353_;
wire [2:0] _0354_;
wire [2:0] _0355_;
wire _0356_;
wire _0357_;
wire _0358_;
wire _0359_;
wire _0360_;
wire _0361_;
wire _0362_;
wire _0363_;
wire _0364_;
wire _0365_;
wire _0366_;
wire _0367_;
wire _0368_;
wire _0369_;
wire _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire _0376_;
wire _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire _0382_;
wire _0383_;
wire _0384_;
wire _0385_;
wire _0386_;
wire _0387_;
wire _0388_;
wire _0389_;
wire _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire _0398_;
wire _0399_;
wire _0400_;
wire _0401_;
wire _0402_;
wire _0403_;
wire _0404_;
wire _0405_;
wire _0406_;
wire _0407_;
wire _0408_;
wire _0409_;
wire _0410_;
wire _0411_;
wire _0412_;
wire _0413_;
wire _0414_;
wire _0415_;
wire _0416_;
wire _0417_;
wire _0418_;
wire _0419_;
wire _0420_;
wire _0421_;
wire _0422_;
wire _0423_;
wire [2:0] _0424_;
wire [2:0] _0425_;
wire [2:0] _0426_;
wire [2:0] _0427_;
wire [2:0] _0428_;
wire [2:0] _0429_;
wire [2:0] _0430_;
wire [2:0] _0431_;
wire [2:0] _0432_;
wire [2:0] _0433_;
wire [2:0] _0434_;
wire [2:0] _0435_;
wire [2:0] _0436_;
wire [2:0] _0437_;
wire [2:0] _0438_;
wire [2:0] _0439_;
wire [2:0] _0440_;
wire [2:0] _0441_;
wire [2:0] _0442_;
wire [2:0] _0443_;
wire [2:0] _0444_;
wire [2:0] _0445_;
wire [2:0] _0446_;
wire [2:0] _0447_;
wire [2:0] _0448_;
wire [2:0] _0449_;
wire _0450_;
wire _0451_;
wire _0452_;
wire _0453_;
wire _0454_;
wire _0455_;
wire _0456_;
wire _0457_;
wire _0458_;
wire _0459_;
wire _0460_;
wire _0461_;
wire _0462_;
wire _0463_;
wire _0464_;
wire _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire _0469_;
wire _0470_;
wire _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire [2:0] _0477_;
wire [2:0] _0478_;
wire [2:0] _0479_;
wire [2:0] _0480_;
wire [2:0] _0481_;
wire [2:0] _0482_;
wire [2:0] _0483_;
wire [2:0] _0484_;
wire [2:0] _0485_;
wire [2:0] _0486_;
wire [2:0] _0487_;
wire [2:0] _0488_;
wire [2:0] _0489_;
wire [2:0] _0490_;
wire [2:0] _0491_;
wire [2:0] _0492_;
wire [2:0] _0493_;
wire [2:0] _0494_;
wire [2:0] _0495_;
wire [2:0] _0496_;
wire [2:0] _0497_;
wire [2:0] _0498_;
wire [2:0] _0499_;
wire [2:0] _0500_;
wire [2:0] _0501_;
wire [2:0] _0502_;
wire _0503_;
wire _0504_;
wire _0505_;
wire _0506_;
wire _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0517_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
wire _0525_;
wire _0526_;
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire _0534_;
wire _0535_;
wire _0536_;
wire _0537_;
wire [1:0] _0538_;
wire [1:0] _0539_;
wire [2:0] _0540_;
wire [4:0] _0541_;
wire _0542_;
wire _0543_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire _0560_;
wire _0561_;
wire _0562_;
wire _0563_;
wire _0564_;
wire _0565_;
wire _0566_;
wire _0567_;
wire _0568_;
wire _0569_;
wire _0570_;
wire _0571_;
wire _0572_;
wire _0573_;
wire _0574_;
wire _0575_;
wire _0576_;
wire _0577_;
wire [4:0] _0578_;
wire [31:0] _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire [31:0] _0590_;
wire [31:0] _0591_;
wire [31:0] _0592_;
wire [31:0] _0593_;
wire [31:0] _0594_;
wire [31:0] _0595_;
wire [31:0] _0596_;
wire [31:0] _0597_;
wire [31:0] _0598_;
wire [1:0] _0599_;
wire [11:0] _0600_;
wire _0601_;
wire _0602_;
wire [31:0] _0603_;
wire [31:0] _0604_;
wire [31:0] _0605_;
wire _0606_;
wire _0607_;
wire [1:0] _0608_;
wire [31:0] _0609_;
wire [31:0] _0610_;
wire [31:0] _0611_;
wire _0612_;
/* cellift = 32'd1 */
wire _0613_;
wire _0614_;
/* cellift = 32'd1 */
wire _0615_;
wire _0616_;
/* cellift = 32'd1 */
wire _0617_;
wire [31:0] _0618_;
wire _0619_;
wire _0620_;
wire _0621_;
wire _0622_;
wire _0623_;
wire _0624_;
wire _0625_;
wire _0626_;
wire _0627_;
wire _0628_;
wire _0629_;
wire _0630_;
wire _0631_;
wire _0632_;
wire _0633_;
wire _0634_;
wire [1:0] _0635_;
wire [1:0] _0636_;
wire [1:0] _0637_;
wire [1:0] _0638_;
wire _0639_;
wire _0640_;
wire _0641_;
wire _0642_;
wire _0643_;
wire _0644_;
wire _0645_;
wire _0646_;
wire _0647_;
wire _0648_;
wire _0649_;
wire _0650_;
wire [29:0] _0651_;
wire [29:0] _0652_;
wire [29:0] _0653_;
wire [29:0] _0654_;
wire [31:0] _0655_;
wire [31:0] _0656_;
wire [31:0] _0657_;
wire [31:0] _0658_;
wire [31:0] _0659_;
wire [31:0] _0660_;
wire [31:0] _0661_;
wire [31:0] _0662_;
wire [31:0] _0663_;
wire [31:0] _0664_;
wire [31:0] _0665_;
wire [31:0] _0666_;
wire [31:0] _0667_;
wire [31:0] _0668_;
wire [31:0] _0669_;
wire [31:0] _0670_;
wire [31:0] _0671_;
wire [31:0] _0672_;
wire [31:0] _0673_;
wire [31:0] _0674_;
wire _0675_;
wire _0676_;
wire _0677_;
wire _0678_;
wire [1:0] _0679_;
wire [1:0] _0680_;
wire [1:0] _0681_;
wire [1:0] _0682_;
wire [29:0] _0683_;
wire [29:0] _0684_;
wire [29:0] _0685_;
wire [29:0] _0686_;
wire [1:0] _0687_;
wire [1:0] _0688_;
wire [1:0] _0689_;
wire [1:0] _0690_;
wire [1:0] _0691_;
wire [1:0] _0692_;
wire [1:0] _0693_;
wire [1:0] _0694_;
wire [2:0] _0695_;
wire [2:0] _0696_;
wire [2:0] _0697_;
wire [2:0] _0698_;
wire [1:0] _0699_;
wire [2:0] _0700_;
wire _0701_;
wire _0702_;
wire _0703_;
wire [31:0] _0704_;
wire [31:0] _0705_;
wire [31:0] _0706_;
wire [31:0] _0707_;
wire [31:0] _0708_;
wire [31:0] _0709_;
wire [18:0] _0710_;
wire [18:0] _0711_;
wire [18:0] _0712_;
wire [18:0] _0713_;
wire [18:0] _0714_;
wire [18:0] _0715_;
wire [18:0] _0716_;
wire [18:0] _0717_;
wire [18:0] _0718_;
wire [18:0] _0719_;
wire [18:0] _0720_;
wire [18:0] _0721_;
wire [18:0] _0722_;
wire [18:0] _0723_;
wire [18:0] _0724_;
wire [18:0] _0725_;
wire [18:0] _0726_;
wire [18:0] _0727_;
wire [18:0] _0728_;
wire [18:0] _0729_;
wire [18:0] _0730_;
wire [18:0] _0731_;
wire [18:0] _0732_;
wire [18:0] _0733_;
wire [18:0] _0734_;
wire [2:0] _0735_;
wire [2:0] _0736_;
wire [2:0] _0737_;
wire [2:0] _0738_;
wire [2:0] _0739_;
wire [2:0] _0740_;
wire [2:0] _0741_;
wire [2:0] _0742_;
wire [2:0] _0743_;
wire [2:0] _0744_;
wire [2:0] _0745_;
wire [2:0] _0746_;
wire [2:0] _0747_;
wire [2:0] _0748_;
wire [2:0] _0749_;
wire [2:0] _0750_;
wire [2:0] _0751_;
wire [2:0] _0752_;
wire [2:0] _0753_;
wire [2:0] _0754_;
wire [2:0] _0755_;
wire [2:0] _0756_;
wire [2:0] _0757_;
wire [2:0] _0758_;
wire [2:0] _0759_;
wire _0760_;
wire _0761_;
wire _0762_;
wire _0763_;
wire _0764_;
wire _0765_;
wire _0766_;
wire _0767_;
wire _0768_;
wire _0769_;
wire _0770_;
wire _0771_;
wire _0772_;
wire _0773_;
wire _0774_;
wire _0775_;
wire _0776_;
wire _0777_;
wire _0778_;
wire _0779_;
wire _0780_;
wire _0781_;
wire _0782_;
wire _0783_;
wire _0784_;
wire _0785_;
wire _0786_;
wire _0787_;
wire _0788_;
wire _0789_;
wire _0790_;
wire _0791_;
wire _0792_;
wire _0793_;
wire _0794_;
wire _0795_;
wire _0796_;
wire _0797_;
wire _0798_;
wire _0799_;
wire _0800_;
wire _0801_;
wire _0802_;
wire _0803_;
wire _0804_;
wire [2:0] _0805_;
wire [2:0] _0806_;
wire [2:0] _0807_;
wire [2:0] _0808_;
wire [2:0] _0809_;
wire [2:0] _0810_;
wire [2:0] _0811_;
wire [2:0] _0812_;
wire _0813_;
wire _0814_;
wire _0815_;
wire _0816_;
wire _0817_;
wire _0818_;
wire _0819_;
wire _0820_;
wire _0821_;
wire _0822_;
wire _0823_;
wire _0824_;
wire _0825_;
wire _0826_;
wire _0827_;
wire [2:0] _0828_;
wire [2:0] _0829_;
wire [2:0] _0830_;
wire [2:0] _0831_;
wire [2:0] _0832_;
wire [2:0] _0833_;
wire [2:0] _0834_;
wire [2:0] _0835_;
wire _0836_;
wire _0837_;
wire _0838_;
wire _0839_;
wire _0840_;
wire _0841_;
wire _0842_;
wire _0843_;
wire _0844_;
wire _0845_;
wire _0846_;
wire [1:0] _0847_;
wire _0848_;
wire _0849_;
wire _0850_;
wire _0851_;
wire _0852_;
wire _0853_;
wire _0854_;
wire _0855_;
wire _0856_;
wire _0857_;
wire _0858_;
wire _0859_;
wire [31:0] _0860_;
wire _0861_;
wire _0862_;
wire _0863_;
wire _0864_;
wire _0865_;
wire _0866_;
wire _0867_;
wire [31:0] _0868_;
wire [31:0] _0869_;
wire [31:0] _0870_;
wire [31:0] _0871_;
wire [31:0] _0872_;
wire [31:0] _0873_;
wire [31:0] _0874_;
wire [31:0] _0875_;
wire [31:0] _0876_;
wire [31:0] _0877_;
wire [31:0] _0878_;
wire [31:0] _0879_;
wire _0880_;
wire [31:0] _0881_;
wire [31:0] _0882_;
wire [31:0] _0883_;
wire _0884_;
wire _0885_;
wire _0886_;
wire [1:0] _0887_;
wire _0888_;
wire _0889_;
wire _0890_;
wire [29:0] _0891_;
wire [31:0] _0892_;
wire [31:0] _0893_;
wire [31:0] _0894_;
wire [31:0] _0895_;
wire [31:0] _0896_;
wire _0897_;
wire [1:0] _0898_;
wire [29:0] _0899_;
wire [1:0] _0900_;
wire [31:0] _0901_;
wire [31:0] _0902_;
wire [18:0] _0903_;
wire [18:0] _0904_;
wire [18:0] _0905_;
wire [18:0] _0906_;
wire [18:0] _0907_;
wire [18:0] _0908_;
wire [18:0] _0909_;
wire [18:0] _0910_;
wire [2:0] _0911_;
wire [2:0] _0912_;
wire [2:0] _0913_;
wire [2:0] _0914_;
wire [2:0] _0915_;
wire [2:0] _0916_;
wire [2:0] _0917_;
wire [2:0] _0918_;
wire _0919_;
wire _0920_;
wire _0921_;
wire _0922_;
wire _0923_;
wire _0924_;
wire _0925_;
wire _0926_;
wire _0927_;
wire _0928_;
wire _0929_;
wire _0930_;
wire _0931_;
wire _0932_;
wire _0933_;
wire _0934_;
wire _0935_;
wire _0936_;
wire _0937_;
wire _0938_;
wire _0939_;
wire _0940_;
wire [2:0] _0941_;
wire [2:0] _0942_;
wire [2:0] _0943_;
wire [2:0] _0944_;
wire [2:0] _0945_;
wire [2:0] _0946_;
wire [2:0] _0947_;
wire [2:0] _0948_;
wire _0949_;
wire _0950_;
wire _0951_;
wire _0952_;
wire _0953_;
wire _0954_;
wire _0955_;
wire _0956_;
wire _0957_;
wire [2:0] _0958_;
wire [2:0] _0959_;
wire [2:0] _0960_;
wire [2:0] _0961_;
wire [2:0] _0962_;
wire [2:0] _0963_;
wire [2:0] _0964_;
wire [2:0] _0965_;
wire _0966_;
wire _0967_;
wire _0968_;
wire _0969_;
wire _0970_;
wire _0971_;
wire _0972_;
wire _0973_;
wire _0974_;
wire _0975_;
wire _0976_;
wire [1:0] _0977_;
wire [1:0] _0978_;
wire [3:0] _0979_;
wire _0980_;
wire _0981_;
wire _0982_;
wire _0983_;
wire [31:0] _0984_;
wire [31:0] _0985_;
wire [31:0] _0986_;
wire [31:0] _0987_;
wire _0988_;
wire [31:0] _0989_;
wire _0990_;
wire _0991_;
wire _0992_;
wire _0993_;
wire _0994_;
wire _0995_;
wire _0996_;
wire _0997_;
wire _0998_;
wire _0999_;
wire _1000_;
wire _1001_;
wire _1002_;
wire _1003_;
wire _1004_;
wire _1005_;
wire _1006_;
wire _1007_;
wire _1008_;
wire _1009_;
wire _1010_;
wire _1011_;
wire _1012_;
wire _1013_;
wire [31:0] _1014_;
/* cellift = 32'd1 */
wire [31:0] _1015_;
wire [18:0] _1016_;
/* cellift = 32'd1 */
wire [18:0] _1017_;
wire [18:0] _1018_;
/* cellift = 32'd1 */
wire [18:0] _1019_;
wire [18:0] _1020_;
/* cellift = 32'd1 */
wire [18:0] _1021_;
wire [18:0] _1022_;
/* cellift = 32'd1 */
wire [18:0] _1023_;
wire [18:0] _1024_;
/* cellift = 32'd1 */
wire [18:0] _1025_;
wire [18:0] _1026_;
/* cellift = 32'd1 */
wire [18:0] _1027_;
wire [18:0] _1028_;
/* cellift = 32'd1 */
wire [18:0] _1029_;
wire [18:0] _1030_;
/* cellift = 32'd1 */
wire [18:0] _1031_;
wire [2:0] _1032_;
/* cellift = 32'd1 */
wire [2:0] _1033_;
wire [2:0] _1034_;
/* cellift = 32'd1 */
wire [2:0] _1035_;
wire [2:0] _1036_;
/* cellift = 32'd1 */
wire [2:0] _1037_;
wire [2:0] _1038_;
/* cellift = 32'd1 */
wire [2:0] _1039_;
wire [2:0] _1040_;
/* cellift = 32'd1 */
wire [2:0] _1041_;
wire [2:0] _1042_;
/* cellift = 32'd1 */
wire [2:0] _1043_;
wire [2:0] _1044_;
/* cellift = 32'd1 */
wire [2:0] _1045_;
wire [2:0] _1046_;
/* cellift = 32'd1 */
wire [2:0] _1047_;
wire _1048_;
/* cellift = 32'd1 */
wire _1049_;
wire _1050_;
/* cellift = 32'd1 */
wire _1051_;
wire _1052_;
/* cellift = 32'd1 */
wire _1053_;
wire _1054_;
/* cellift = 32'd1 */
wire _1055_;
wire _1056_;
/* cellift = 32'd1 */
wire _1057_;
wire _1058_;
/* cellift = 32'd1 */
wire _1059_;
wire _1060_;
/* cellift = 32'd1 */
wire _1061_;
wire _1062_;
/* cellift = 32'd1 */
wire _1063_;
wire _1064_;
/* cellift = 32'd1 */
wire _1065_;
wire _1066_;
/* cellift = 32'd1 */
wire _1067_;
wire _1068_;
/* cellift = 32'd1 */
wire _1069_;
wire _1070_;
/* cellift = 32'd1 */
wire _1071_;
wire _1072_;
/* cellift = 32'd1 */
wire _1073_;
wire _1074_;
/* cellift = 32'd1 */
wire _1075_;
wire _1076_;
/* cellift = 32'd1 */
wire _1077_;
wire _1078_;
/* cellift = 32'd1 */
wire _1079_;
wire _1080_;
/* cellift = 32'd1 */
wire _1081_;
wire _1082_;
/* cellift = 32'd1 */
wire _1083_;
wire _1084_;
/* cellift = 32'd1 */
wire _1085_;
wire _1086_;
/* cellift = 32'd1 */
wire _1087_;
wire _1088_;
/* cellift = 32'd1 */
wire _1089_;
wire _1090_;
/* cellift = 32'd1 */
wire _1091_;
wire [2:0] _1092_;
/* cellift = 32'd1 */
wire [2:0] _1093_;
wire [2:0] _1094_;
/* cellift = 32'd1 */
wire [2:0] _1095_;
wire [2:0] _1096_;
/* cellift = 32'd1 */
wire [2:0] _1097_;
wire [2:0] _1098_;
/* cellift = 32'd1 */
wire [2:0] _1099_;
wire [2:0] _1100_;
/* cellift = 32'd1 */
wire [2:0] _1101_;
wire [2:0] _1102_;
/* cellift = 32'd1 */
wire [2:0] _1103_;
wire [2:0] _1104_;
/* cellift = 32'd1 */
wire [2:0] _1105_;
wire [2:0] _1106_;
/* cellift = 32'd1 */
wire [2:0] _1107_;
wire _1108_;
/* cellift = 32'd1 */
wire _1109_;
wire _1110_;
/* cellift = 32'd1 */
wire _1111_;
wire _1112_;
/* cellift = 32'd1 */
wire _1113_;
wire _1114_;
/* cellift = 32'd1 */
wire _1115_;
wire _1116_;
/* cellift = 32'd1 */
wire _1117_;
wire _1118_;
/* cellift = 32'd1 */
wire _1119_;
wire _1120_;
/* cellift = 32'd1 */
wire _1121_;
wire _1122_;
/* cellift = 32'd1 */
wire _1123_;
wire [2:0] _1124_;
/* cellift = 32'd1 */
wire [2:0] _1125_;
wire [2:0] _1126_;
/* cellift = 32'd1 */
wire [2:0] _1127_;
wire [2:0] _1128_;
/* cellift = 32'd1 */
wire [2:0] _1129_;
wire [2:0] _1130_;
/* cellift = 32'd1 */
wire [2:0] _1131_;
wire [2:0] _1132_;
/* cellift = 32'd1 */
wire [2:0] _1133_;
wire [2:0] _1134_;
/* cellift = 32'd1 */
wire [2:0] _1135_;
wire [2:0] _1136_;
/* cellift = 32'd1 */
wire [2:0] _1137_;
wire [2:0] _1138_;
/* cellift = 32'd1 */
wire [2:0] _1139_;
wire _1140_;
/* cellift = 32'd1 */
wire _1141_;
wire _1142_;
/* cellift = 32'd1 */
wire _1143_;
wire _1144_;
/* cellift = 32'd1 */
wire _1145_;
wire _1146_;
/* cellift = 32'd1 */
wire _1147_;
wire _1148_;
/* cellift = 32'd1 */
wire _1149_;
wire _1150_;
/* cellift = 32'd1 */
wire _1151_;
wire _1152_;
/* cellift = 32'd1 */
wire _1153_;
wire _1154_;
/* cellift = 32'd1 */
wire _1155_;
wire _1156_;
/* cellift = 32'd1 */
wire _1157_;
wire _1158_;
/* cellift = 32'd1 */
wire _1159_;
wire _1160_;
/* cellift = 32'd1 */
wire _1161_;
/* cellift = 32'd1 */
wire [1:0] _1162_;
/* src = "generated/sv2v_out.v:424.14-424.27" */
wire _1163_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:424.14-424.27" */
wire _1164_;
/* src = "generated/sv2v_out.v:425.22-425.38" */
wire _1165_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:425.22-425.38" */
wire _1166_;
/* src = "generated/sv2v_out.v:425.44-425.60" */
wire _1167_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:425.44-425.60" */
wire _1168_;
/* src = "generated/sv2v_out.v:425.67-425.86" */
wire _1169_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:425.67-425.86" */
wire _1170_;
/* src = "generated/sv2v_out.v:431.22-431.35" */
wire _1171_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:431.22-431.35" */
wire _1172_;
/* src = "generated/sv2v_out.v:558.38-558.65" */
wire _1173_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:558.38-558.65" */
wire _1174_;
/* src = "generated/sv2v_out.v:559.38-559.66" */
wire _1175_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:559.38-559.66" */
wire _1176_;
/* src = "generated/sv2v_out.v:573.40-573.69" */
wire _1177_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:573.40-573.69" */
wire _1178_;
/* src = "generated/sv2v_out.v:574.40-574.70" */
wire _1179_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:574.40-574.70" */
wire _1180_;
/* src = "generated/sv2v_out.v:411.9-411.29" */
wire _1181_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:411.9-411.29" */
wire _1182_;
/* src = "generated/sv2v_out.v:424.13-424.39" */
wire _1183_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:424.13-424.39" */
wire _1184_;
/* src = "generated/sv2v_out.v:424.12-424.53" */
wire _1185_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:424.12-424.53" */
wire _1186_;
/* src = "generated/sv2v_out.v:425.20-425.87" */
wire _1187_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:425.20-425.87" */
wire _1188_;
/* src = "generated/sv2v_out.v:425.21-425.61" */
wire _1189_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:425.21-425.61" */
wire _1190_;
/* src = "generated/sv2v_out.v:426.17-426.34" */
wire _1191_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:426.17-426.34" */
wire _1192_;
/* src = "generated/sv2v_out.v:425.18-425.88" */
wire _1193_;
/* src = "generated/sv2v_out.v:494.39-494.57" */
wire [31:0] _1194_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:494.39-494.57" */
wire [31:0] _1195_;
wire [3:0] _1196_;
/* unused_bits = "0 1 2" */
wire [3:0] _1197_;
/* cellift = 32'd1 */
/* unused_bits = "0 1 2" */
wire [3:0] _1198_;
wire _1199_;
/* cellift = 32'd1 */
wire _1200_;
wire _1201_;
wire _1202_;
/* cellift = 32'd1 */
wire _1203_;
wire _1204_;
/* cellift = 32'd1 */
wire _1205_;
wire _1206_;
wire _1207_;
/* cellift = 32'd1 */
wire _1208_;
/* cellift = 32'd1 */
wire _1209_;
wire _1210_;
/* cellift = 32'd1 */
wire _1211_;
wire _1212_;
/* cellift = 32'd1 */
wire _1213_;
wire _1214_;
/* cellift = 32'd1 */
wire _1215_;
wire [31:0] _1216_;
/* cellift = 32'd1 */
wire [31:0] _1217_;
wire [31:0] _1218_;
/* cellift = 32'd1 */
wire [31:0] _1219_;
wire _1220_;
/* cellift = 32'd1 */
wire _1221_;
wire [31:0] _1222_;
/* cellift = 32'd1 */
wire [31:0] _1223_;
wire [31:0] _1224_;
/* cellift = 32'd1 */
wire [31:0] _1225_;
wire [31:0] _1226_;
/* cellift = 32'd1 */
wire [31:0] _1227_;
wire _1228_;
/* cellift = 32'd1 */
wire _1229_;
wire [31:0] _1230_;
/* cellift = 32'd1 */
wire [31:0] _1231_;
wire _1232_;
/* cellift = 32'd1 */
wire _1233_;
wire _1234_;
/* cellift = 32'd1 */
wire _1235_;
wire [31:0] _1236_;
/* cellift = 32'd1 */
wire [31:0] _1237_;
wire [31:0] _1238_;
/* cellift = 32'd1 */
wire [31:0] _1239_;
wire _1240_;
/* cellift = 32'd1 */
wire _1241_;
wire [31:0] _1242_;
/* cellift = 32'd1 */
wire [31:0] _1243_;
wire _1244_;
/* cellift = 32'd1 */
wire _1245_;
wire _1246_;
/* cellift = 32'd1 */
wire _1247_;
wire _1248_;
/* cellift = 32'd1 */
wire _1249_;
wire _1250_;
wire _1251_;
/* cellift = 32'd1 */
wire _1252_;
wire [31:0] _1253_;
/* cellift = 32'd1 */
wire [31:0] _1254_;
/* unused_bits = "0 1" */
wire [31:0] _1255_;
/* cellift = 32'd1 */
/* unused_bits = "0 1" */
wire [31:0] _1256_;
wire _1257_;
wire _1258_;
/* cellift = 32'd1 */
wire _1259_;
/* src = "generated/sv2v_out.v:550.22-550.28" */
wire _1260_;
/* src = "generated/sv2v_out.v:356.13-356.26" */
input activate_trap;
wire activate_trap;
/* cellift = 32'd1 */
input activate_trap_t0;
wire activate_trap_t0;
/* src = "generated/sv2v_out.v:348.13-348.16" */
input clk;
wire clk;
/* cellift = 32'd1 */
input clk_t0;
wire clk_t0;
/* src = "generated/sv2v_out.v:365.13-365.27" */
output core_interrupt;
reg core_interrupt;
/* src = "generated/sv2v_out.v:366.19-366.39" */
output [3:0] core_interrupt_cause;
wire [3:0] core_interrupt_cause;
/* cellift = 32'd1 */
output [3:0] core_interrupt_cause_t0;
wire [3:0] core_interrupt_cause_t0;
/* cellift = 32'd1 */
output core_interrupt_t0;
reg core_interrupt_t0;
/* src = "generated/sv2v_out.v:353.20-353.28" */
output [31:0] csr_data;
reg [31:0] csr_data;
/* cellift = 32'd1 */
output [31:0] csr_data_t0;
reg [31:0] csr_data_t0;
/* src = "generated/sv2v_out.v:372.13-372.24" */
wire [31:0] csr_rd_data;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:372.13-372.24" */
wire [31:0] csr_rd_data_t0;
/* src = "generated/sv2v_out.v:376.7-376.16" */
wire csr_rd_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:376.7-376.16" */
wire csr_rd_en_t0;
/* src = "generated/sv2v_out.v:374.7-374.17" */
wire csr_rd_vld;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:374.7-374.17" */
wire csr_rd_vld_t0;
/* src = "generated/sv2v_out.v:352.14-352.21" */
output csr_rdy;
wire csr_rdy;
/* cellift = 32'd1 */
output csr_rdy_t0;
wire csr_rdy_t0;
/* src = "generated/sv2v_out.v:351.13-351.20" */
input csr_vld;
wire csr_vld;
/* cellift = 32'd1 */
input csr_vld_t0;
wire csr_vld_t0;
/* src = "generated/sv2v_out.v:373.13-373.24" */
wire [31:0] csr_wr_data;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:373.13-373.24" */
wire [31:0] csr_wr_data_t0;
/* src = "generated/sv2v_out.v:377.7-377.16" */
wire csr_wr_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:377.7-377.16" */
wire csr_wr_en_t0;
/* src = "generated/sv2v_out.v:375.6-375.16" */
reg csr_wr_vld;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:375.6-375.16" */
reg csr_wr_vld_t0;
/* src = "generated/sv2v_out.v:350.21-350.27" */
input [180:0] decode;
wire [180:0] decode;
/* cellift = 32'd1 */
input [180:0] decode_t0;
wire [180:0] decode_t0;
/* src = "generated/sv2v_out.v:364.13-364.31" */
input external_interrupt;
wire external_interrupt;
/* cellift = 32'd1 */
input external_interrupt_t0;
wire external_interrupt_t0;
/* src = "generated/sv2v_out.v:355.13-355.20" */
input instret;
wire instret;
/* cellift = 32'd1 */
input instret_t0;
wire instret_t0;
/* src = "generated/sv2v_out.v:384.13-384.19" */
reg [31:0] mcause;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:384.13-384.19" */
reg [31:0] mcause_t0;
/* src = "generated/sv2v_out.v:389.14-389.20" */
wire [63:0] mcycle;
/* src = "generated/sv2v_out.v:388.7-388.20" */
wire mcycle_rd_vld;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:388.7-388.20" */
wire mcycle_rd_vld_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:389.14-389.20" */
wire [63:0] mcycle_t0;
/* src = "generated/sv2v_out.v:387.7-387.19" */
wire mcycle_wrenh;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:387.7-387.19" */
wire mcycle_wrenh_t0;
/* src = "generated/sv2v_out.v:386.7-386.19" */
wire mcycle_wrenl;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:386.7-386.19" */
wire mcycle_wrenl_t0;
/* src = "generated/sv2v_out.v:383.13-383.17" */
reg [31:0] mepc;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:383.13-383.17" */
reg [31:0] mepc_t0;
/* src = "generated/sv2v_out.v:379.12-379.15" */
reg [2:0] mie;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:379.12-379.15" */
reg [2:0] mie_t0;
/* src = "generated/sv2v_out.v:393.14-393.22" */
wire [63:0] minstret;
/* src = "generated/sv2v_out.v:392.7-392.22" */
wire minstret_rd_vld;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:392.7-392.22" */
wire minstret_rd_vld_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:393.14-393.22" */
wire [63:0] minstret_t0;
/* src = "generated/sv2v_out.v:391.7-391.21" */
wire minstret_wrenh;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:391.7-391.21" */
wire minstret_wrenh_t0;
/* src = "generated/sv2v_out.v:390.7-390.21" */
wire minstret_wrenl;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:390.7-390.21" */
wire minstret_wrenl_t0;
/* src = "generated/sv2v_out.v:380.12-380.15" */
reg [2:0] mip;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:380.12-380.15" */
reg [2:0] mip_t0;
/* src = "generated/sv2v_out.v:382.13-382.21" */
reg [31:0] mscratch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:382.13-382.21" */
reg [31:0] mscratch_t0;
/* src = "generated/sv2v_out.v:378.12-378.19" */
wire [3:0] mstatus;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:378.12-378.19" */
wire [3:0] mstatus_t0;
/* src = "generated/sv2v_out.v:385.13-385.18" */
reg [31:0] mtval;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:385.13-385.18" */
reg [31:0] mtval_t0;
/* src = "generated/sv2v_out.v:381.13-381.18" */
wire [31:0] mtvec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:381.13-381.18" */
wire [31:0] mtvec_t0;
/* src = "generated/sv2v_out.v:395.12-395.22" */
wire [1:0] next_state;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:395.12-395.22" */
wire [1:0] next_state_t0;
/* src = "generated/sv2v_out.v:354.13-354.22" */
output regwr_csr;
reg regwr_csr;
/* cellift = 32'd1 */
output regwr_csr_t0;
reg regwr_csr_t0;
/* src = "generated/sv2v_out.v:357.13-357.24" */
input return_trap;
wire return_trap;
/* cellift = 32'd1 */
input return_trap_t0;
wire return_trap_t0;
/* src = "generated/sv2v_out.v:349.13-349.17" */
input rstz;
wire rstz;
/* src = "generated/sv2v_out.v:362.13-362.31" */
input software_interrupt;
wire software_interrupt;
/* cellift = 32'd1 */
input software_interrupt_t0;
wire software_interrupt_t0;
/* src = "generated/sv2v_out.v:394.12-394.17" */
reg [1:0] state;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:394.12-394.17" */
reg [1:0] state_t0;
/* src = "generated/sv2v_out.v:363.13-363.28" */
input timer_interrupt;
wire timer_interrupt;
/* cellift = 32'd1 */
input timer_interrupt_t0;
wire timer_interrupt_t0;
/* src = "generated/sv2v_out.v:358.20-358.30" */
input [31:0] trap_cause;
wire [31:0] trap_cause;
/* cellift = 32'd1 */
input [31:0] trap_cause_t0;
wire [31:0] trap_cause_t0;
/* src = "generated/sv2v_out.v:360.20-360.31" */
output [31:0] trap_handle;
reg [31:0] trap_handle;
/* cellift = 32'd1 */
output [31:0] trap_handle_t0;
reg [31:0] trap_handle_t0;
/* src = "generated/sv2v_out.v:361.13-361.22" */
output trap_jump;
reg trap_jump;
/* cellift = 32'd1 */
output trap_jump_t0;
reg trap_jump_t0;
/* src = "generated/sv2v_out.v:359.20-359.30" */
input [31:0] trap_value;
wire [31:0] trap_value;
/* cellift = 32'd1 */
input [31:0] trap_value_t0;
wire [31:0] trap_value_t0;
/* src = "generated/sv2v_out.v:371.14-371.21" */
wire [31:0] wr_data;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:371.14-371.21" */
wire [31:0] wr_data_t0;
assign _0002_ = csr_data & /* src = "generated/sv2v_out.v:495.39-495.58" */ _0132_;
assign _0004_ = software_interrupt & /* src = "generated/sv2v_out.v:539.15-539.46" */ mstatus[0];
assign _0006_ = _0004_ & /* src = "generated/sv2v_out.v:539.14-539.56" */ mie[0];
assign _0008_ = timer_interrupt & /* src = "generated/sv2v_out.v:540.15-540.43" */ mstatus[0];
assign _0010_ = _0008_ & /* src = "generated/sv2v_out.v:540.14-540.53" */ mie[1];
assign _0012_ = external_interrupt & /* src = "generated/sv2v_out.v:541.15-541.46" */ mstatus[0];
assign _0014_ = _0012_ & /* src = "generated/sv2v_out.v:541.14-541.56" */ mie[2];
assign _0205_ = software_interrupt_t0 & mstatus[0];
assign _0208_ = _0005_ & mie[0];
assign _0211_ = timer_interrupt_t0 & mstatus[0];
assign _0214_ = _0009_ & mie[1];
assign _0217_ = external_interrupt_t0 & mstatus[0];
assign _0220_ = _0013_ & mie[2];
assign _0203_ = wr_data_t0 & csr_data;
assign _0206_ = mstatus_t0[0] & software_interrupt;
assign _0209_ = mie_t0[0] & _0004_;
assign _0212_ = mstatus_t0[0] & timer_interrupt;
assign _0215_ = mie_t0[1] & _0008_;
assign _0218_ = mstatus_t0[0] & external_interrupt;
assign _0221_ = mie_t0[2] & _0012_;
assign _0207_ = software_interrupt_t0 & mstatus_t0[0];
assign _0210_ = _0005_ & mie_t0[0];
assign _0213_ = timer_interrupt_t0 & mstatus_t0[0];
assign _0216_ = _0009_ & mie_t0[1];
assign _0219_ = external_interrupt_t0 & mstatus_t0[0];
assign _0222_ = _0013_ & mie_t0[2];
assign _0618_ = _0202_ | _0203_;
assign _0619_ = _0205_ | _0206_;
assign _0620_ = _0208_ | _0209_;
assign _0621_ = _0211_ | _0212_;
assign _0622_ = _0214_ | _0215_;
assign _0623_ = _0217_ | _0218_;
assign _0624_ = _0220_ | _0221_;
assign _0003_ = _0618_ | _0204_;
assign _0005_ = _0619_ | _0207_;
assign _0007_ = _0620_ | _0210_;
assign _0009_ = _0621_ | _0213_;
assign _0011_ = _0622_ | _0216_;
assign _0013_ = _0623_ | _0219_;
assign _0015_ = _0624_ | _0222_;
assign _0892_ = csr_wr_data ^ mscratch;
assign _0893_ = _1230_ ^ mepc;
assign _0894_ = _1222_ ^ mcause;
assign _0895_ = _1242_ ^ mtval;
assign _0896_ = csr_rd_data ^ csr_data;
assign _0899_ = _1255_[31:2] ^ trap_handle[31:2];
assign _0068_ = ~ _0048_;
assign _0069_ = ~ _0050_;
assign _0070_ = ~ _0052_;
assign _0071_ = ~ _0054_;
assign _0072_ = ~ csr_rd_en;
assign _0074_ = ~ _0056_;
assign _0655_ = csr_wr_data_t0 | mscratch_t0;
assign _0659_ = _1231_ | mepc_t0;
assign _0663_ = _1223_ | mcause_t0;
assign _0667_ = _1243_ | mtval_t0;
assign _0671_ = csr_rd_data_t0 | csr_data_t0;
assign _0683_ = _1256_[31:2] | trap_handle_t0[31:2];
assign _0656_ = _0892_ | _0655_;
assign _0660_ = _0893_ | _0659_;
assign _0664_ = _0894_ | _0663_;
assign _0668_ = _0895_ | _0667_;
assign _0672_ = _0896_ | _0671_;
assign _0684_ = _0899_ | _0683_;
assign _0246_ = { _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_, _0048_ } & csr_wr_data_t0;
assign _0249_ = { _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_, _0050_ } & _1231_;
assign _0252_ = { _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_, _0052_ } & _1223_;
assign _0255_ = { _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_ } & _1243_;
assign _0258_ = { csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en, csr_rd_en } & csr_rd_data_t0;
assign _0267_ = { _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_, _0056_ } & _1256_[31:2];
assign _0247_ = { _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_ } & mscratch_t0;
assign _0250_ = { _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_, _0069_ } & mepc_t0;
assign _0253_ = { _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_, _0070_ } & mcause_t0;
assign _0256_ = { _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_ } & mtval_t0;
assign _0259_ = { _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_ } & csr_data_t0;
assign _0268_ = { _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_, _0074_ } & trap_handle_t0[31:2];
assign _0248_ = _0656_ & { _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_, _0049_ };
assign _0251_ = _0660_ & { _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_, _0051_ };
assign _0254_ = _0664_ & { _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_ };
assign _0257_ = _0668_ & { _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_ };
assign _0260_ = _0672_ & { csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0, csr_rd_en_t0 };
assign _0269_ = _0684_ & { _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_, _0057_ };
assign _0657_ = _0246_ | _0247_;
assign _0661_ = _0249_ | _0250_;
assign _0665_ = _0252_ | _0253_;
assign _0669_ = _0255_ | _0256_;
assign _0673_ = _0258_ | _0259_;
assign _0685_ = _0267_ | _0268_;
assign _0658_ = _0657_ | _0248_;
assign _0662_ = _0661_ | _0251_;
assign _0666_ = _0665_ | _0254_;
assign _0670_ = _0669_ | _0257_;
assign _0674_ = _0673_ | _0260_;
assign _0686_ = _0685_ | _0269_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME mscratch_t0 */
always_ff @(posedge clk)
mscratch_t0 <= _0658_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME mepc_t0 */
always_ff @(posedge clk)
mepc_t0 <= _0662_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME mcause_t0 */
always_ff @(posedge clk)
mcause_t0 <= _0666_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME mtval_t0 */
always_ff @(posedge clk)
mtval_t0 <= _0670_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME csr_data_t0 */
always_ff @(posedge clk)
csr_data_t0 <= _0674_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME trap_handle_t0[31:2] */
always_ff @(posedge clk)
trap_handle_t0[31:2] <= _0686_;
assign _0161_ = | { _1065_, csr_wr_en_t0 };
assign _0163_ = | { _1229_, csr_wr_en_t0 };
assign _0164_ = | { _1221_, csr_wr_en_t0 };
assign _0165_ = | { _1241_, csr_wr_en_t0 };
assign _0169_ = | { _1172_, csr_rd_vld_t0 };
assign _0170_ = | { _1164_, _1182_ };
assign _0183_ = | decode_t0[131:129];
assign _0186_ = | decode_t0[130:129];
assign _0187_ = | decode_t0[148:137];
assign _0078_ = ~ { _1065_, csr_wr_en_t0 };
assign _0080_ = ~ { _1229_, csr_wr_en_t0 };
assign _0081_ = ~ { _1221_, csr_wr_en_t0 };
assign _0082_ = ~ { _1241_, csr_wr_en_t0 };
assign _0086_ = ~ { _1172_, csr_rd_vld_t0 };
assign _0087_ = ~ { _1164_, _1182_ };
assign _0126_ = ~ decode_t0[131:129];
assign _0137_ = ~ decode_t0[130:129];
assign _0138_ = ~ decode_t0[148:137];
assign _0139_ = ~ state_t0;
assign _0275_ = { _1206_, csr_wr_en } & _0078_;
assign _0277_ = { _1228_, csr_wr_en } & _0080_;
assign _0278_ = { _1220_, csr_wr_en } & _0081_;
assign _0279_ = { _1240_, csr_wr_en } & _0082_;
assign _0283_ = { _1171_, csr_rd_vld } & _0086_;
assign _0284_ = { _1163_, _1181_ } & _0087_;
assign _0540_ = decode[131:129] & _0126_;
assign _0599_ = decode[130:129] & _0137_;
assign _0600_ = decode[148:137] & _0138_;
assign _0608_ = state & _0139_;
assign _0990_ = _0275_ == { 1'h0, _0078_[0] };
assign _0991_ = _0277_ == { 1'h0, _0080_[0] };
assign _0992_ = _0278_ == { 1'h0, _0081_[0] };
assign _0993_ = _0279_ == { 1'h0, _0082_[0] };
assign _0994_ = _0283_ == { _0086_[1], 1'h0 };
assign _0995_ = _0284_ == { _0087_[1], 1'h0 };
assign _0996_ = _0540_ == { 1'h0, _0126_[1], 1'h0 };
assign _0997_ = _0540_ == { 1'h0, _0126_[1:0] };
assign _0998_ = _0599_ == _0137_;
assign _0999_ = _0599_ == { _0137_[1], 1'h0 };
assign _1000_ = _0600_ == { _0138_[11], 1'h0, _0138_[9:7], 5'h00, _0138_[1], 1'h0 };
assign _1001_ = _0600_ == { _0138_[11], 1'h0, _0138_[9:7], 7'h00 };
assign _1002_ = _0600_ == { _0138_[11], 1'h0, _0138_[9:8], 6'h00, _0138_[1], 1'h0 };
assign _1003_ = _0600_ == { _0138_[11], 1'h0, _0138_[9:8], 8'h00 };
assign _1004_ = _0600_ == { 2'h0, _0138_[9:8], 1'h0, _0138_[6], 3'h0, _0138_[2], 2'h0 };
assign _1005_ = _0600_ == { 2'h0, _0138_[9:8], 1'h0, _0138_[6], 4'h0, _0138_[1:0] };
assign _1006_ = _0600_ == { 2'h0, _0138_[9:8], 1'h0, _0138_[6], 4'h0, _0138_[1], 1'h0 };
assign _1007_ = _0600_ == { 2'h0, _0138_[9:8], 1'h0, _0138_[6], 5'h00, _0138_[0] };
assign _1008_ = _0600_ == { 2'h0, _0138_[9:8], 1'h0, _0138_[6], 6'h00 };
assign _1009_ = _0600_ == { 2'h0, _0138_[9:8], 5'h00, _0138_[2], 1'h0, _0138_[0] };
assign _1010_ = _0600_ == { 2'h0, _0138_[9:8], 5'h00, _0138_[2], 2'h0 };
assign _1011_ = _0600_ == { 2'h0, _0138_[9:8], 8'h00 };
assign _1012_ = _0608_ == { _0139_[1], 1'h0 };
assign _1013_ = _0608_ == { 1'h0, _0139_[0] };
assign _0021_ = _0990_ & _0161_;
assign _0025_ = _0991_ & _0163_;
assign _0027_ = _0992_ & _0164_;
assign _0029_ = _0993_ & _0165_;
assign _0037_ = _0994_ & _0169_;
assign _0039_ = _0995_ & _0170_;
assign _1166_ = _0996_ & _0183_;
assign _1168_ = _0997_ & _0183_;
assign _1245_ = _0998_ & _0186_;
assign _1247_ = _0999_ & _0186_;
assign _1180_ = _1000_ & _0187_;
assign _1176_ = _1001_ & _0187_;
assign _1178_ = _1002_ & _0187_;
assign _1174_ = _1003_ & _0187_;
assign _1249_ = _1004_ & _0187_;
assign _1241_ = _1005_ & _0187_;
assign _1221_ = _1006_ & _0187_;
assign _1229_ = _1007_ & _0187_;
assign _1233_ = _1008_ & _0187_;
assign _1235_ = _1009_ & _0187_;
assign _1200_ = _1010_ & _0187_;
assign _1065_ = _1011_ & _0187_;
assign csr_rdy_t0 = _1012_ & _0188_;
assign _1172_ = _1013_ & _0188_;
/* src = "generated/sv2v_out.v:419.2-429.22" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME csr_wr_vld */
always_ff @(posedge clk)
if (!rstz) csr_wr_vld <= 1'h0;
else if (_1185_) csr_wr_vld <= _1193_;
/* src = "generated/sv2v_out.v:546.2-557.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME core_interrupt */
always_ff @(posedge clk)
if (!rstz) core_interrupt <= 1'h0;
else core_interrupt <= _1260_;
reg core_interrupt_cause_reg__2_ ;
/* src = "generated/sv2v_out.v:546.2-557.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME core_interrupt_cause_reg__2_  */
always_ff @(posedge clk)
if (_0040_)
if (_0060_) core_interrupt_cause_reg__2_  <= 1'h0;
else core_interrupt_cause_reg__2_  <= _0979_[2];
assign core_interrupt_cause[2] = core_interrupt_cause_reg__2_ ;
reg core_interrupt_cause_reg__3_ ;
/* src = "generated/sv2v_out.v:546.2-557.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME core_interrupt_cause_reg__3_  */
always_ff @(posedge clk)
if (_0040_)
if (mip[2]) core_interrupt_cause_reg__3_  <= 1'h1;
else core_interrupt_cause_reg__3_  <= _1197_[3];
assign core_interrupt_cause[3] = core_interrupt_cause_reg__3_ ;
reg [1:0] _1442_;
/* src = "generated/sv2v_out.v:500.2-542.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME _1442_ */
always_ff @(posedge clk)
if (!rstz) _1442_ <= 2'h0;
else if (_0042_) _1442_ <= { _1207_, _1214_ };
assign mstatus[1:0] = _1442_;
/* src = "generated/sv2v_out.v:500.2-542.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME mie[2] */
always_ff @(posedge clk)
if (!rstz) mie[2] <= 1'h0;
else if (_0044_) mie[2] <= csr_wr_data[11];
/* src = "generated/sv2v_out.v:500.2-542.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME mie[1] */
always_ff @(posedge clk)
if (!rstz) mie[1] <= 1'h0;
else if (_0044_) mie[1] <= csr_wr_data[7];
/* src = "generated/sv2v_out.v:500.2-542.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME mie[0] */
always_ff @(posedge clk)
if (!rstz) mie[0] <= 1'h0;
else if (_0044_) mie[0] <= csr_wr_data[3];
/* src = "generated/sv2v_out.v:500.2-542.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME mip */
always_ff @(posedge clk)
if (!rstz) mip <= 3'h0;
else mip <= { _0014_, _0010_, _0006_ };
reg [29:0] _1447_;
/* src = "generated/sv2v_out.v:500.2-542.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME _1447_ */
always_ff @(posedge clk)
if (!rstz) _1447_ <= 30'h20000000;
else if (_0046_) _1447_ <= csr_wr_data[31:2];
assign mtvec[31:2] = _1447_;
/* src = "generated/sv2v_out.v:500.2-542.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME mscratch */
always_ff @(posedge clk)
if (_0048_) mscratch <= csr_wr_data;
/* src = "generated/sv2v_out.v:500.2-542.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME mepc */
always_ff @(posedge clk)
if (_0050_) mepc <= _1230_;
/* src = "generated/sv2v_out.v:500.2-542.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME mcause */
always_ff @(posedge clk)
if (_0052_) mcause <= _1222_;
/* src = "generated/sv2v_out.v:500.2-542.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME mtval */
always_ff @(posedge clk)
if (_0054_) mtval <= _1242_;
/* src = "generated/sv2v_out.v:436.2-448.22" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME trap_jump */
always_ff @(posedge clk)
if (!rstz) trap_jump <= 1'h0;
else trap_jump <= _1251_;
/* src = "generated/sv2v_out.v:433.2-435.28" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME csr_data */
always_ff @(posedge clk)
if (csr_rd_en) csr_data <= csr_rd_data;
/* src = "generated/sv2v_out.v:419.2-429.22" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME regwr_csr */
always_ff @(posedge clk)
if (!rstz) regwr_csr <= 1'h0;
else if (_0032_) regwr_csr <= _1258_;
/* src = "generated/sv2v_out.v:436.2-448.22" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME trap_handle[1:0] */
always_ff @(posedge clk)
if (_0056_)
if (activate_trap) trap_handle[1:0] <= 2'h0;
else trap_handle[1:0] <= _1253_[1:0];
/* src = "generated/sv2v_out.v:436.2-448.22" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME trap_handle[31:2] */
always_ff @(posedge clk)
if (_0056_) trap_handle[31:2] <= _1255_[31:2];
/* src = "generated/sv2v_out.v:402.2-406.24" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME state */
always_ff @(posedge clk)
if (!rstz) state <= 2'h0;
else if (_0058_) state <= next_state;
assign _0542_ = csr_vld_t0 & decode[6];
assign _0545_ = _1164_ & csr_vld;
assign _0548_ = _1184_ & decode[6];
assign _0551_ = _1190_ & _1169_;
assign _0554_ = mcycle_rd_vld_t0 & minstret_rd_vld;
assign _0557_ = _1172_ & csr_rd_vld;
assign _0560_ = csr_rdy_t0 & csr_wr_vld;
assign _0563_ = csr_wr_en_t0 & _1173_;
assign _0566_ = csr_wr_en_t0 & _1175_;
assign _0569_ = csr_wr_en_t0 & _1177_;
assign _0572_ = csr_wr_en_t0 & _1179_;
assign _0543_ = decode_t0[6] & csr_vld;
assign _0546_ = csr_vld_t0 & _1163_;
assign _0549_ = decode_t0[6] & _1183_;
assign _0552_ = _1170_ & _1189_;
assign _0555_ = minstret_rd_vld_t0 & mcycle_rd_vld;
assign _0558_ = csr_rd_vld_t0 & _1171_;
assign _0561_ = csr_wr_vld_t0 & csr_rdy;
assign _0564_ = _1174_ & csr_wr_en;
assign _0567_ = _1176_ & csr_wr_en;
assign _0570_ = _1178_ & csr_wr_en;
assign _0573_ = _1180_ & csr_wr_en;
assign _0544_ = csr_vld_t0 & decode_t0[6];
assign _0547_ = _1164_ & csr_vld_t0;
assign _0550_ = _1184_ & decode_t0[6];
assign _0553_ = _1190_ & _1170_;
assign _0556_ = mcycle_rd_vld_t0 & minstret_rd_vld_t0;
assign _0559_ = _1172_ & csr_rd_vld_t0;
assign _0562_ = csr_rdy_t0 & csr_wr_vld_t0;
assign _0565_ = csr_wr_en_t0 & _1174_;
assign _0568_ = csr_wr_en_t0 & _1176_;
assign _0571_ = csr_wr_en_t0 & _1178_;
assign _0574_ = csr_wr_en_t0 & _1180_;
assign _0848_ = _0542_ | _0543_;
assign _0849_ = _0545_ | _0546_;
assign _0850_ = _0548_ | _0549_;
assign _0851_ = _0551_ | _0552_;
assign _0852_ = _0554_ | _0555_;
assign _0853_ = _0557_ | _0558_;
assign _0854_ = _0560_ | _0561_;
assign _0855_ = _0563_ | _0564_;
assign _0856_ = _0566_ | _0567_;
assign _0857_ = _0569_ | _0570_;
assign _0858_ = _0572_ | _0573_;
assign _1182_ = _0848_ | _0544_;
assign _1184_ = _0849_ | _0547_;
assign _1186_ = _0850_ | _0550_;
assign _1188_ = _0851_ | _0553_;
assign csr_rd_vld_t0 = _0852_ | _0556_;
assign csr_rd_en_t0 = _0853_ | _0559_;
assign csr_wr_en_t0 = _0854_ | _0562_;
assign mcycle_wrenl_t0 = _0855_ | _0565_;
assign mcycle_wrenh_t0 = _0856_ | _0568_;
assign minstret_wrenl_t0 = _0857_ | _0571_;
assign minstret_wrenh_t0 = _0858_ | _0574_;
assign _0160_ = | { activate_trap_t0, return_trap_t0, csr_wr_en_t0 };
assign _0162_ = | { activate_trap_t0, csr_wr_en_t0 };
assign _0166_ = | { activate_trap_t0, return_trap_t0 };
assign _0167_ = | { csr_rdy_t0, _1186_ };
assign _0168_ = | { csr_rdy_t0, _1164_, _1172_ };
assign _0179_ = | { _1241_, _0613_, _1174_, _1178_ };
assign _0180_ = | { _1176_, _1180_, _1178_ };
assign _0181_ = | { _1229_, _1221_, _1233_ };
assign _0182_ = | { _1249_, _1241_, _1176_, _1180_, _1174_, _1178_ };
assign _0184_ = | decode_t0[136:132];
assign _0185_ = | decode_t0[128:124];
assign _0188_ = | state_t0;
assign _0159_ = | mip_t0;
assign _0077_ = ~ { csr_wr_en_t0, return_trap_t0, activate_trap_t0 };
assign _0079_ = ~ { csr_wr_en_t0, activate_trap_t0 };
assign _0083_ = ~ { return_trap_t0, activate_trap_t0 };
assign _0084_ = ~ { csr_rdy_t0, _1186_ };
assign _0085_ = ~ { _1172_, _1164_, csr_rdy_t0 };
assign _0094_ = ~ { _0613_, _1241_, _1178_, _1174_ };
assign _0095_ = ~ { _1180_, _1178_, _1176_ };
assign _0096_ = ~ { _1233_, _1229_, _1221_ };
assign _0097_ = ~ { _1249_, _1241_, _1180_, _1178_, _1176_, _1174_ };
assign _0127_ = ~ decode_t0[136:132];
assign _0130_ = ~ decode_t0[128:124];
assign _0076_ = ~ mip_t0;
assign _0274_ = { csr_wr_en, return_trap, activate_trap } & _0077_;
assign _0276_ = { csr_wr_en, activate_trap } & _0079_;
assign _0280_ = { return_trap, activate_trap } & _0083_;
assign _0281_ = { csr_rdy, _1185_ } & _0084_;
assign _0282_ = { _1171_, _1163_, csr_rdy } & _0085_;
assign _0294_ = { _0612_, _1240_, _1177_, _1173_ } & _0094_;
assign _0295_ = { _1179_, _1177_, _1175_ } & _0095_;
assign _0296_ = { _1232_, _1228_, _1220_ } & _0096_;
assign _0297_ = { _1248_, _1240_, _1179_, _1177_, _1175_, _1173_ } & _0097_;
assign _0541_ = decode[136:132] & _0127_;
assign _0578_ = decode[128:124] & _0130_;
assign _0273_ = mip & _0076_;
assign _0190_ = ! _0274_;
assign _0191_ = ! _0276_;
assign _0192_ = ! _0280_;
assign _0193_ = ! _0281_;
assign _0194_ = ! _0282_;
assign _0195_ = ! _0294_;
assign _0196_ = ! _0295_;
assign _0197_ = ! _0296_;
assign _0198_ = ! _0297_;
assign _0199_ = ! _0541_;
assign _0200_ = ! _0578_;
assign _0201_ = ! _0608_;
assign _0189_ = ! _0273_;
assign _0019_ = _0190_ & _0160_;
assign _0023_ = _0191_ & _0162_;
assign _0031_ = _0192_ & _0166_;
assign _0033_ = _0193_ & _0167_;
assign _0035_ = _0194_ & _0168_;
assign _0152_ = _0195_ & _0179_;
assign _0154_ = _0196_ & _0180_;
assign _0156_ = _0197_ & _0181_;
assign _0158_ = _0198_ & _0182_;
assign _1170_ = _0199_ & _0184_;
assign _1192_ = _0200_ & _0185_;
assign _1164_ = _0201_ & _0188_;
assign _0017_ = _0189_ & _0159_;
assign _0128_ = ~ _1165_;
assign _0129_ = ~ _1167_;
assign _0575_ = _1166_ & _0129_;
assign _0576_ = _1168_ & _0128_;
assign _0577_ = _1166_ & _1168_;
assign _0859_ = _0575_ | _0576_;
assign _1190_ = _0859_ | _0577_;
assign _0098_ = ~ { _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_ };
assign _0099_ = ~ { _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_ };
assign _0100_ = ~ { _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_ };
assign _0101_ = ~ { _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_ };
assign _0102_ = ~ { _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_ };
assign _0103_ = ~ { _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_ };
assign _0104_ = ~ { _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_ };
assign _0105_ = ~ { _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_ };
assign _0106_ = ~ { _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_ };
assign _0107_ = ~ { _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_ };
assign _0122_ = ~ _1177_;
assign _0123_ = ~ _0612_;
assign _0124_ = ~ _0151_;
assign _0108_ = ~ { _1179_, _1179_, _1179_ };
assign _0109_ = ~ { _1173_, _1173_, _1173_ };
assign _0110_ = ~ { _1177_, _1177_, _1177_ };
assign _0111_ = ~ { _0612_, _0612_, _0612_ };
assign _0112_ = ~ { _1220_, _1220_, _1220_ };
assign _0113_ = ~ { _1232_, _1232_, _1232_ };
assign _0114_ = ~ { _0614_, _0614_, _0614_ };
assign _0115_ = ~ { _0151_, _0151_, _0151_ };
assign _0088_ = ~ _1175_;
assign _0089_ = ~ _1179_;
assign _0116_ = ~ _1248_;
assign _0117_ = ~ _1173_;
assign _0118_ = ~ _0153_;
assign _0090_ = ~ _1228_;
assign _0091_ = ~ _1220_;
assign _0093_ = ~ _1234_;
assign _0119_ = ~ _0616_;
assign _0120_ = ~ _0155_;
assign _0121_ = ~ _0157_;
assign _0125_ = ~ { csr_rdy, csr_rdy };
assign _0133_ = ~ activate_trap;
assign _0134_ = ~ csr_wr_en;
assign _0135_ = ~ { activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap };
assign _0136_ = ~ { csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en };
assign _0063_ = ~ _1185_;
assign _0140_ = ~ { decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131] };
assign _0704_ = { _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_ } | _0098_;
assign _0707_ = { _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_ } | _0099_;
assign _0710_ = { _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_ } | _0100_;
assign _0713_ = { _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_ } | _0101_;
assign _0716_ = { _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_ } | _0102_;
assign _0719_ = { _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_ } | _0103_;
assign _0722_ = { _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_ } | _0104_;
assign _0726_ = { _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_ } | _0105_;
assign _0729_ = { _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_ } | _0106_;
assign _0732_ = { _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_ } | _0107_;
assign _0815_ = _1178_ | _0122_;
assign _0818_ = _0613_ | _0123_;
assign _0825_ = _0152_ | _0124_;
assign _0735_ = { _1180_, _1180_, _1180_ } | _0108_;
assign _0738_ = { _1174_, _1174_, _1174_ } | _0109_;
assign _0741_ = { _1178_, _1178_, _1178_ } | _0110_;
assign _0744_ = { _0613_, _0613_, _0613_ } | _0111_;
assign _0747_ = { _1221_, _1221_, _1221_ } | _0112_;
assign _0751_ = { _1233_, _1233_, _1233_ } | _0113_;
assign _0754_ = { _0615_, _0615_, _0615_ } | _0114_;
assign _0757_ = { _0152_, _0152_, _0152_ } | _0115_;
assign _0760_ = _1176_ | _0088_;
assign _0763_ = _1180_ | _0089_;
assign _0766_ = _1249_ | _0116_;
assign _0769_ = _1174_ | _0117_;
assign _0772_ = _0154_ | _0118_;
assign _0775_ = _1229_ | _0090_;
assign _0778_ = _1221_ | _0091_;
assign _0781_ = _1235_ | _0093_;
assign _0784_ = _0617_ | _0119_;
assign _0787_ = _0156_ | _0120_;
assign _0790_ = _0158_ | _0121_;
assign _0847_ = { csr_rdy_t0, csr_rdy_t0 } | _0125_;
assign _0862_ = activate_trap_t0 | _0133_;
assign _0864_ = csr_wr_en_t0 | _0134_;
assign _0871_ = { csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0 } | _0136_;
assign _0868_ = { activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0 } | _0135_;
assign _0881_ = { decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131] } | _0140_;
assign _0705_ = { _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_ } | { _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_, _1246_ };
assign _0708_ = { _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_ } | { _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_, _1244_ };
assign _0711_ = { _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_ } | { _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_, _1179_ };
assign _0714_ = { _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_ } | { _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_, _1173_ };
assign _0717_ = { _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_ } | { _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_ };
assign _0720_ = { _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_ } | { _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_, _0612_ };
assign _0723_ = { _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_ } | { _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_ };
assign _0725_ = { _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_ } | { _1234_, _1234_, _1234_, _1234_, _1234_, _1234_, _1234_, _1234_, _1234_, _1234_, _1234_, _1234_, _1234_, _1234_, _1234_, _1234_, _1234_, _1234_, _1234_ };
assign _0727_ = { _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_ } | { _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_, _1232_ };
assign _0730_ = { _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_ } | { _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_, _0614_ };
assign _0733_ = { _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_ } | { _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_ };
assign _0816_ = _1178_ | _1177_;
assign _0819_ = _0613_ | _0612_;
assign _0826_ = _0152_ | _0151_;
assign _0736_ = { _1180_, _1180_, _1180_ } | { _1179_, _1179_, _1179_ };
assign _0739_ = { _1174_, _1174_, _1174_ } | { _1173_, _1173_, _1173_ };
assign _0742_ = { _1178_, _1178_, _1178_ } | { _1177_, _1177_, _1177_ };
assign _0745_ = { _0613_, _0613_, _0613_ } | { _0612_, _0612_, _0612_ };
assign _0748_ = { _1221_, _1221_, _1221_ } | { _1220_, _1220_, _1220_ };
assign _0750_ = { _1235_, _1235_, _1235_ } | { _1234_, _1234_, _1234_ };
assign _0752_ = { _1233_, _1233_, _1233_ } | { _1232_, _1232_, _1232_ };
assign _0755_ = { _0615_, _0615_, _0615_ } | { _0614_, _0614_, _0614_ };
assign _0758_ = { _0152_, _0152_, _0152_ } | { _0151_, _0151_, _0151_ };
assign _0761_ = _1176_ | _1175_;
assign _0764_ = _1180_ | _1179_;
assign _0767_ = _1249_ | _1248_;
assign _0770_ = _1174_ | _1173_;
assign _0773_ = _0154_ | _0153_;
assign _0776_ = _1229_ | _1228_;
assign _0779_ = _1221_ | _1220_;
assign _0782_ = _1235_ | _1234_;
assign _0785_ = _0617_ | _0616_;
assign _0788_ = _0156_ | _0155_;
assign _0791_ = _0158_ | _0157_;
assign _0863_ = activate_trap_t0 | activate_trap;
assign _0801_ = _1065_ | _1206_;
assign _0865_ = csr_wr_en_t0 | csr_wr_en;
assign _0870_ = { _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_ } | { _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_ };
assign _0874_ = { _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_, _1229_ } | { _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_, _1228_ };
assign _0869_ = { activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0 } | { activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap, activate_trap };
assign _0876_ = { _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_, _1241_ } | { _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_, _1240_ };
assign _0872_ = { csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0 } | { csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en, csr_wr_en };
assign _0861_ = return_trap_t0 | return_trap;
assign _0878_ = { return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0, return_trap_t0 } | { return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap, return_trap };
assign _0880_ = _1186_ | _1185_;
assign _0882_ = { decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131] } | { decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131] };
assign _0298_ = wr_data_t0 & _0704_;
assign _0301_ = _1015_ & _0707_;
assign _0304_ = mcycle_t0[63:45] & _0710_;
assign _0307_ = mtval_t0[31:13] & _0713_;
assign _0310_ = _1019_ & _0716_;
assign _0313_ = _1021_ & _0719_;
assign _0316_ = mepc_t0[31:13] & _0722_;
assign _0321_ = _1027_ & _0726_;
assign _0324_ = _1029_ & _0729_;
assign _0327_ = _1031_ & _0732_;
assign _0330_ = mcycle_t0[34:32] & _0735_;
assign _0333_ = mtval_t0[2:0] & _0738_;
assign _0336_ = _1035_ & _0741_;
assign _0339_ = _1037_ & _0744_;
assign _0342_ = mepc_t0[2:0] & _0747_;
assign _0347_ = _1043_ & _0751_;
assign _0350_ = _1045_ & _0754_;
assign _0353_ = _1047_ & _0757_;
assign _0356_ = minstret_t0[11] & _0760_;
assign _0359_ = _1049_ & _0763_;
assign _0362_ = mtval_t0[11] & _0766_;
assign _0365_ = _1053_ & _0769_;
assign _0368_ = _1055_ & _0772_;
assign _0371_ = mscratch_t0[11] & _0775_;
assign _0374_ = _1059_ & _0778_;
assign _0377_ = mie_t0[2] & _0781_;
assign _0380_ = _1065_ & _0784_;
assign _0383_ = _1067_ & _0787_;
assign _0386_ = _1069_ & _0790_;
assign _0389_ = minstret_t0[3] & _0760_;
assign _0392_ = _1071_ & _0763_;
assign _0395_ = mtval_t0[3] & _0766_;
assign _0398_ = _1075_ & _0769_;
assign _0401_ = _1077_ & _0772_;
assign _0404_ = mscratch_t0[3] & _0775_;
assign _0407_ = _1081_ & _0778_;
assign _0410_ = mie_t0[0] & _0781_;
assign _0415_ = _1087_ & _0784_;
assign _0418_ = _1089_ & _0787_;
assign _0421_ = _1091_ & _0790_;
assign _0424_ = mcycle_t0[38:36] & _0735_;
assign _0427_ = mtval_t0[6:4] & _0738_;
assign _0430_ = _1095_ & _0741_;
assign _0433_ = _1097_ & _0744_;
assign _0436_ = mepc_t0[6:4] & _0747_;
assign _0441_ = _1103_ & _0751_;
assign _0444_ = _1105_ & _0754_;
assign _0447_ = _1107_ & _0757_;
assign _0450_ = mcycle_t0[44] & _0763_;
assign _0453_ = mtval_t0[12] & _0769_;
assign _0456_ = _1111_ & _0815_;
assign _0459_ = _1113_ & _0818_;
assign _0462_ = mscratch_t0[12] & _0775_;
assign _0465_ = _1117_ & _0778_;
assign _0468_ = _1065_ & _0781_;
assign _0471_ = _1121_ & _0787_;
assign _0474_ = _1123_ & _0825_;
assign _0477_ = mcycle_t0[42:40] & _0735_;
assign _0480_ = mtval_t0[10:8] & _0738_;
assign _0483_ = _1127_ & _0741_;
assign _0486_ = _1129_ & _0744_;
assign _0489_ = mepc_t0[10:8] & _0747_;
assign _0494_ = _1135_ & _0751_;
assign _0497_ = _1137_ & _0754_;
assign _0500_ = _1139_ & _0757_;
assign _0503_ = minstret_t0[7] & _0760_;
assign _0506_ = _1141_ & _0763_;
assign _0509_ = mtval_t0[7] & _0766_;
assign _0512_ = _1145_ & _0769_;
assign _0515_ = _1147_ & _0772_;
assign _0518_ = mscratch_t0[7] & _0775_;
assign _0521_ = _1151_ & _0778_;
assign _0524_ = mie_t0[1] & _0781_;
assign _0529_ = _1157_ & _0784_;
assign _0532_ = _1159_ & _0787_;
assign _0535_ = _1161_ & _0790_;
assign _0538_ = _1162_ & _0847_;
assign _0582_ = _1203_ & _0864_;
assign _0585_ = _1209_ & _0862_;
assign _0587_ = _1211_ & _0864_;
assign _0590_ = _1217_ & _0871_;
assign _0593_ = _1225_ & _0871_;
assign _0596_ = _1237_ & _0871_;
assign _0601_ = return_trap_t0 & _0862_;
assign _0603_ = _1254_ & _0868_;
assign _0609_ = decode_t0[116:85] & _0881_;
assign _0299_ = _1195_ & _0705_;
assign _0302_ = _0003_ & _0708_;
assign _0305_ = minstret_t0[63:45] & _0711_;
assign _0308_ = mcycle_t0[31:13] & _0714_;
assign _0311_ = minstret_t0[31:13] & _0717_;
assign _0314_ = _1017_ & _0720_;
assign _0317_ = mcause_t0[31:13] & _0723_;
assign _0319_ = mtvec_t0[31:13] & _0725_;
assign _0322_ = mscratch_t0[31:13] & _0727_;
assign _0325_ = _1025_ & _0730_;
assign _0328_ = _1023_ & _0733_;
assign _0331_ = minstret_t0[34:32] & _0736_;
assign _0334_ = mcycle_t0[2:0] & _0739_;
assign _0337_ = minstret_t0[2:0] & _0742_;
assign _0340_ = _1033_ & _0745_;
assign _0343_ = mcause_t0[2:0] & _0748_;
assign _0345_ = { mtvec_t0[2], 2'h0 } & _0750_;
assign _0348_ = mscratch_t0[2:0] & _0752_;
assign _0351_ = _1041_ & _0755_;
assign _0354_ = _1039_ & _0758_;
assign _0357_ = mcycle_t0[43] & _0761_;
assign _0360_ = minstret_t0[43] & _0764_;
assign _0363_ = mip_t0[2] & _0767_;
assign _0366_ = mcycle_t0[11] & _0770_;
assign _0369_ = _1051_ & _0773_;
assign _0372_ = mepc_t0[11] & _0776_;
assign _0375_ = mcause_t0[11] & _0779_;
assign _0378_ = mtvec_t0[11] & _0782_;
assign _0381_ = _1063_ & _0785_;
assign _0384_ = _1061_ & _0788_;
assign _0387_ = _1057_ & _0791_;
assign _0390_ = mcycle_t0[35] & _0761_;
assign _0393_ = minstret_t0[35] & _0764_;
assign _0396_ = mip_t0[0] & _0767_;
assign _0399_ = mcycle_t0[3] & _0770_;
assign _0402_ = _1073_ & _0773_;
assign _0405_ = mepc_t0[3] & _0776_;
assign _0408_ = mcause_t0[3] & _0779_;
assign _0411_ = mtvec_t0[3] & _0782_;
assign _0413_ = mstatus_t0[0] & _0801_;
assign _0416_ = _1085_ & _0785_;
assign _0419_ = _1083_ & _0788_;
assign _0422_ = _1079_ & _0791_;
assign _0425_ = minstret_t0[38:36] & _0736_;
assign _0428_ = mcycle_t0[6:4] & _0739_;
assign _0431_ = minstret_t0[6:4] & _0742_;
assign _0434_ = _1093_ & _0745_;
assign _0437_ = mcause_t0[6:4] & _0748_;
assign _0439_ = mtvec_t0[6:4] & _0750_;
assign _0442_ = mscratch_t0[6:4] & _0752_;
assign _0445_ = _1101_ & _0755_;
assign _0448_ = _1099_ & _0758_;
assign _0451_ = minstret_t0[44] & _0764_;
assign _0454_ = mcycle_t0[12] & _0770_;
assign _0457_ = minstret_t0[12] & _0816_;
assign _0460_ = _1109_ & _0819_;
assign _0463_ = mepc_t0[12] & _0776_;
assign _0466_ = mcause_t0[12] & _0779_;
assign _0469_ = mtvec_t0[12] & _0782_;
assign _0472_ = _1119_ & _0788_;
assign _0475_ = _1115_ & _0826_;
assign _0478_ = minstret_t0[42:40] & _0736_;
assign _0481_ = mcycle_t0[10:8] & _0739_;
assign _0484_ = minstret_t0[10:8] & _0742_;
assign _0487_ = _1125_ & _0745_;
assign _0490_ = mcause_t0[10:8] & _0748_;
assign _0492_ = mtvec_t0[10:8] & _0750_;
assign _0495_ = mscratch_t0[10:8] & _0752_;
assign _0498_ = _1133_ & _0755_;
assign _0501_ = _1131_ & _0758_;
assign _0504_ = mcycle_t0[39] & _0761_;
assign _0507_ = minstret_t0[39] & _0764_;
assign _0510_ = mip_t0[1] & _0767_;
assign _0513_ = mcycle_t0[7] & _0770_;
assign _0516_ = _1143_ & _0773_;
assign _0519_ = mepc_t0[7] & _0776_;
assign _0522_ = mcause_t0[7] & _0779_;
assign _0525_ = mtvec_t0[7] & _0782_;
assign _0527_ = mstatus_t0[1] & _0801_;
assign _0530_ = _1155_ & _0785_;
assign _0533_ = _1153_ & _0788_;
assign _0536_ = _1149_ & _0791_;
assign _0580_ = mstatus_t0[0] & _0863_;
assign _1205_ = csr_wr_data_t0[7] & _0801_;
assign _0583_ = _1205_ & _0865_;
assign _1209_ = mstatus_t0[1] & _0861_;
assign _1213_ = csr_wr_data_t0[3] & _0801_;
assign _0588_ = _1213_ & _0865_;
assign _1217_ = trap_cause_t0 & _0869_;
assign _1219_ = csr_wr_data_t0 & _0870_;
assign _0591_ = _1219_ & _0872_;
assign _1225_ = { decode_t0[180:151], 2'h0 } & _0869_;
assign _1227_ = { csr_wr_data_t0[31:2], 2'h0 } & _0874_;
assign _0594_ = _1227_ & _0872_;
assign _1237_ = trap_value_t0 & _0869_;
assign _1239_ = csr_wr_data_t0 & _0876_;
assign _0597_ = _1239_ & _0872_;
assign _1254_ = mepc_t0 & _0878_;
assign _0604_ = { mtvec_t0[31:2], 2'h0 } & _0869_;
assign _0606_ = _1192_ & _0880_;
assign _0610_ = { 27'h0000000, decode_t0[136:132] } & _0882_;
assign _0706_ = _0298_ | _0299_;
assign _0709_ = _0301_ | _0302_;
assign _0712_ = _0304_ | _0305_;
assign _0715_ = _0307_ | _0308_;
assign _0718_ = _0310_ | _0311_;
assign _0721_ = _0313_ | _0314_;
assign _0724_ = _0316_ | _0317_;
assign _0728_ = _0321_ | _0322_;
assign _0731_ = _0324_ | _0325_;
assign _0734_ = _0327_ | _0328_;
assign _0737_ = _0330_ | _0331_;
assign _0740_ = _0333_ | _0334_;
assign _0743_ = _0336_ | _0337_;
assign _0746_ = _0339_ | _0340_;
assign _0749_ = _0342_ | _0343_;
assign _0753_ = _0347_ | _0348_;
assign _0756_ = _0350_ | _0351_;
assign _0759_ = _0353_ | _0354_;
assign _0762_ = _0356_ | _0357_;
assign _0765_ = _0359_ | _0360_;
assign _0768_ = _0362_ | _0363_;
assign _0771_ = _0365_ | _0366_;
assign _0774_ = _0368_ | _0369_;
assign _0777_ = _0371_ | _0372_;
assign _0780_ = _0374_ | _0375_;
assign _0783_ = _0377_ | _0378_;
assign _0786_ = _0380_ | _0381_;
assign _0789_ = _0383_ | _0384_;
assign _0792_ = _0386_ | _0387_;
assign _0793_ = _0389_ | _0390_;
assign _0794_ = _0392_ | _0393_;
assign _0795_ = _0395_ | _0396_;
assign _0796_ = _0398_ | _0399_;
assign _0797_ = _0401_ | _0402_;
assign _0798_ = _0404_ | _0405_;
assign _0799_ = _0407_ | _0408_;
assign _0800_ = _0410_ | _0411_;
assign _0802_ = _0415_ | _0416_;
assign _0803_ = _0418_ | _0419_;
assign _0804_ = _0421_ | _0422_;
assign _0805_ = _0424_ | _0425_;
assign _0806_ = _0427_ | _0428_;
assign _0807_ = _0430_ | _0431_;
assign _0808_ = _0433_ | _0434_;
assign _0809_ = _0436_ | _0437_;
assign _0810_ = _0441_ | _0442_;
assign _0811_ = _0444_ | _0445_;
assign _0812_ = _0447_ | _0448_;
assign _0813_ = _0450_ | _0451_;
assign _0814_ = _0453_ | _0454_;
assign _0817_ = _0456_ | _0457_;
assign _0820_ = _0459_ | _0460_;
assign _0821_ = _0462_ | _0463_;
assign _0822_ = _0465_ | _0466_;
assign _0823_ = _0468_ | _0469_;
assign _0824_ = _0471_ | _0472_;
assign _0827_ = _0474_ | _0475_;
assign _0828_ = _0477_ | _0478_;
assign _0829_ = _0480_ | _0481_;
assign _0830_ = _0483_ | _0484_;
assign _0831_ = _0486_ | _0487_;
assign _0832_ = _0489_ | _0490_;
assign _0833_ = _0494_ | _0495_;
assign _0834_ = _0497_ | _0498_;
assign _0835_ = _0500_ | _0501_;
assign _0836_ = _0503_ | _0504_;
assign _0837_ = _0506_ | _0507_;
assign _0838_ = _0509_ | _0510_;
assign _0839_ = _0512_ | _0513_;
assign _0840_ = _0515_ | _0516_;
assign _0841_ = _0518_ | _0519_;
assign _0842_ = _0521_ | _0522_;
assign _0843_ = _0524_ | _0525_;
assign _0844_ = _0529_ | _0530_;
assign _0845_ = _0532_ | _0533_;
assign _0846_ = _0535_ | _0536_;
assign _0866_ = _0582_ | _0583_;
assign _0867_ = _0587_ | _0588_;
assign _0873_ = _0590_ | _0591_;
assign _0875_ = _0593_ | _0594_;
assign _0877_ = _0596_ | _0597_;
assign _0879_ = _0603_ | _0604_;
assign _0883_ = _0609_ | _0610_;
assign _0901_ = wr_data ^ _1194_;
assign _0902_ = _1014_ ^ _0002_;
assign _0903_ = mcycle[63:45] ^ minstret[63:45];
assign _0904_ = mtval[31:13] ^ mcycle[31:13];
assign _0905_ = _1018_ ^ minstret[31:13];
assign _0906_ = _1020_ ^ _1016_;
assign _0907_ = mepc[31:13] ^ mcause[31:13];
assign _0908_ = _1026_ ^ mscratch[31:13];
assign _0909_ = _1028_ ^ _1024_;
assign _0910_ = _1030_ ^ _1022_;
assign _0911_ = mcycle[34:32] ^ minstret[34:32];
assign _0912_ = mtval[2:0] ^ mcycle[2:0];
assign _0913_ = _1034_ ^ minstret[2:0];
assign _0914_ = _1036_ ^ _1032_;
assign _0915_ = mepc[2:0] ^ mcause[2:0];
assign _0916_ = _1042_ ^ mscratch[2:0];
assign _0917_ = _1044_ ^ _1040_;
assign _0918_ = _1046_ ^ _1038_;
assign _0919_ = minstret[11] ^ mcycle[43];
assign _0920_ = _1048_ ^ minstret[43];
assign _0921_ = mtval[11] ^ mip[2];
assign _0922_ = _1052_ ^ mcycle[11];
assign _0923_ = _1054_ ^ _1050_;
assign _0924_ = mscratch[11] ^ mepc[11];
assign _0925_ = _1058_ ^ mcause[11];
assign _0926_ = mie[2] ^ mtvec[11];
assign _0927_ = _1064_ ^ _1062_;
assign _0928_ = _1066_ ^ _1060_;
assign _0929_ = _1068_ ^ _1056_;
assign _0930_ = minstret[3] ^ mcycle[35];
assign _0931_ = _1070_ ^ minstret[35];
assign _0932_ = mtval[3] ^ mip[0];
assign _0933_ = _1074_ ^ mcycle[3];
assign _0934_ = _1076_ ^ _1072_;
assign _0935_ = mscratch[3] ^ mepc[3];
assign _0936_ = _1080_ ^ mcause[3];
assign _0937_ = mie[0] ^ mtvec[3];
assign _0938_ = _1086_ ^ _1084_;
assign _0939_ = _1088_ ^ _1082_;
assign _0940_ = _1090_ ^ _1078_;
assign _0941_ = mcycle[38:36] ^ minstret[38:36];
assign _0942_ = mtval[6:4] ^ mcycle[6:4];
assign _0943_ = _1094_ ^ minstret[6:4];
assign _0944_ = _1096_ ^ _1092_;
assign _0945_ = mepc[6:4] ^ mcause[6:4];
assign _0946_ = _1102_ ^ mscratch[6:4];
assign _0947_ = _1104_ ^ _1100_;
assign _0948_ = _1106_ ^ _1098_;
assign _0949_ = mcycle[44] ^ minstret[44];
assign _0950_ = mtval[12] ^ mcycle[12];
assign _0951_ = _1110_ ^ minstret[12];
assign _0952_ = _1112_ ^ _1108_;
assign _0953_ = mscratch[12] ^ mepc[12];
assign _0954_ = _1116_ ^ mcause[12];
assign _0955_ = _1064_ ^ mtvec[12];
assign _0956_ = _1120_ ^ _1118_;
assign _0957_ = _1122_ ^ _1114_;
assign _0958_ = mcycle[42:40] ^ minstret[42:40];
assign _0959_ = mtval[10:8] ^ mcycle[10:8];
assign _0960_ = _1126_ ^ minstret[10:8];
assign _0961_ = _1128_ ^ _1124_;
assign _0962_ = mepc[10:8] ^ mcause[10:8];
assign _0963_ = _1134_ ^ mscratch[10:8];
assign _0964_ = _1136_ ^ _1132_;
assign _0965_ = _1138_ ^ _1130_;
assign _0966_ = minstret[7] ^ mcycle[39];
assign _0967_ = _1140_ ^ minstret[39];
assign _0968_ = mtval[7] ^ mip[1];
assign _0969_ = _1144_ ^ mcycle[7];
assign _0970_ = _1146_ ^ _1142_;
assign _0971_ = mscratch[7] ^ mepc[7];
assign _0972_ = _1150_ ^ mcause[7];
assign _0973_ = mie[1] ^ mtvec[7];
assign _0974_ = _1156_ ^ _1154_;
assign _0975_ = _1158_ ^ _1152_;
assign _0976_ = _1160_ ^ _1148_;
assign _0977_ = _0000_ ^ _0001_;
assign _0980_ = _1201_ ^ mstatus[0];
assign _0981_ = _1202_ ^ _1204_;
assign _0983_ = _1210_ ^ _1212_;
assign _0984_ = _1216_ ^ _1218_;
assign _0985_ = _1224_ ^ _1226_;
assign _0986_ = _1236_ ^ _1238_;
assign _0987_ = _1253_ ^ { mtvec[31:2], 2'h0 };
assign _0988_ = _1257_ ^ _1191_;
assign _0989_ = decode[116:85] ^ { 27'h0000000, decode[136:132] };
assign _0300_ = { _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_, _1247_ } & _0901_;
assign _0303_ = { _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_, _1245_ } & _0902_;
assign _0306_ = { _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_, _1180_ } & _0903_;
assign _0309_ = { _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_ } & _0904_;
assign _0312_ = { _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_ } & _0905_;
assign _0315_ = { _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_, _0613_ } & _0906_;
assign _0318_ = { _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_ } & _0907_;
assign _0320_ = { _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_, _1235_ } & mtvec[31:13];
assign _0323_ = { _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_, _1233_ } & _0908_;
assign _0326_ = { _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_, _0615_ } & _0909_;
assign _0329_ = { _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_ } & _0910_;
assign _0332_ = { _1180_, _1180_, _1180_ } & _0911_;
assign _0335_ = { _1174_, _1174_, _1174_ } & _0912_;
assign _0338_ = { _1178_, _1178_, _1178_ } & _0913_;
assign _0341_ = { _0613_, _0613_, _0613_ } & _0914_;
assign _0344_ = { _1221_, _1221_, _1221_ } & _0915_;
assign _0346_ = { _1235_, _1235_, _1235_ } & { mtvec[2], 2'h0 };
assign _0349_ = { _1233_, _1233_, _1233_ } & _0916_;
assign _0352_ = { _0615_, _0615_, _0615_ } & _0917_;
assign _0355_ = { _0152_, _0152_, _0152_ } & _0918_;
assign _0358_ = _1176_ & _0919_;
assign _0361_ = _1180_ & _0920_;
assign _0364_ = _1249_ & _0921_;
assign _0367_ = _1174_ & _0922_;
assign _0370_ = _0154_ & _0923_;
assign _0373_ = _1229_ & _0924_;
assign _0376_ = _1221_ & _0925_;
assign _0379_ = _1235_ & _0926_;
assign _0382_ = _0617_ & _0927_;
assign _0385_ = _0156_ & _0928_;
assign _0388_ = _0158_ & _0929_;
assign _0391_ = _1176_ & _0930_;
assign _0394_ = _1180_ & _0931_;
assign _0397_ = _1249_ & _0932_;
assign _0400_ = _1174_ & _0933_;
assign _0403_ = _0154_ & _0934_;
assign _0406_ = _1229_ & _0935_;
assign _0409_ = _1221_ & _0936_;
assign _0412_ = _1235_ & _0937_;
assign _0414_ = _1065_ & mstatus[0];
assign _0417_ = _0617_ & _0938_;
assign _0420_ = _0156_ & _0939_;
assign _0423_ = _0158_ & _0940_;
assign _0426_ = { _1180_, _1180_, _1180_ } & _0941_;
assign _0429_ = { _1174_, _1174_, _1174_ } & _0942_;
assign _0432_ = { _1178_, _1178_, _1178_ } & _0943_;
assign _0435_ = { _0613_, _0613_, _0613_ } & _0944_;
assign _0438_ = { _1221_, _1221_, _1221_ } & _0945_;
assign _0440_ = { _1235_, _1235_, _1235_ } & mtvec[6:4];
assign _0443_ = { _1233_, _1233_, _1233_ } & _0946_;
assign _0446_ = { _0615_, _0615_, _0615_ } & _0947_;
assign _0449_ = { _0152_, _0152_, _0152_ } & _0948_;
assign _0452_ = _1180_ & _0949_;
assign _0455_ = _1174_ & _0950_;
assign _0458_ = _1178_ & _0951_;
assign _0461_ = _0613_ & _0952_;
assign _0464_ = _1229_ & _0953_;
assign _0467_ = _1221_ & _0954_;
assign _0470_ = _1235_ & _0955_;
assign _0473_ = _0156_ & _0956_;
assign _0476_ = _0152_ & _0957_;
assign _0479_ = { _1180_, _1180_, _1180_ } & _0958_;
assign _0482_ = { _1174_, _1174_, _1174_ } & _0959_;
assign _0485_ = { _1178_, _1178_, _1178_ } & _0960_;
assign _0488_ = { _0613_, _0613_, _0613_ } & _0961_;
assign _0491_ = { _1221_, _1221_, _1221_ } & _0962_;
assign _0493_ = { _1235_, _1235_, _1235_ } & mtvec[10:8];
assign _0496_ = { _1233_, _1233_, _1233_ } & _0963_;
assign _0499_ = { _0615_, _0615_, _0615_ } & _0964_;
assign _0502_ = { _0152_, _0152_, _0152_ } & _0965_;
assign _0505_ = _1176_ & _0966_;
assign _0508_ = _1180_ & _0967_;
assign _0511_ = _1249_ & _0968_;
assign _0514_ = _1174_ & _0969_;
assign _0517_ = _0154_ & _0970_;
assign _0520_ = _1229_ & _0971_;
assign _0523_ = _1221_ & _0972_;
assign _0526_ = _1235_ & _0973_;
assign _0528_ = _1065_ & mstatus[1];
assign _0531_ = _0617_ & _0974_;
assign _0534_ = _0156_ & _0975_;
assign _0537_ = _0158_ & _0976_;
assign _1162_ = { _1172_, _1172_ } & _0977_;
assign _0539_ = { csr_rdy_t0, csr_rdy_t0 } & _0978_;
assign _1198_ = { mip_t0[0], mip_t0[0], mip_t0[0], mip_t0[0] } & { _0979_[3:2], _0061_ };
assign _0581_ = activate_trap_t0 & _0980_;
assign _0584_ = csr_wr_en_t0 & _0981_;
assign _0586_ = activate_trap_t0 & _0982_;
assign _0589_ = csr_wr_en_t0 & _0983_;
assign _0592_ = { csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0 } & _0984_;
assign _0595_ = { csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0 } & _0985_;
assign _0598_ = { csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0, csr_wr_en_t0 } & _0986_;
assign _0602_ = activate_trap_t0 & _0062_;
assign _0605_ = { activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0, activate_trap_t0 } & _0987_;
assign _0607_ = _1186_ & _0988_;
assign _0611_ = { decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131] } & _0989_;
assign _1015_ = _0300_ | _0706_;
assign csr_wr_data_t0 = _0303_ | _0709_;
assign _1017_ = _0306_ | _0712_;
assign _1019_ = _0309_ | _0715_;
assign _1021_ = _0312_ | _0718_;
assign _1023_ = _0315_ | _0721_;
assign _1025_ = _0318_ | _0724_;
assign _1027_ = _0320_ | _0319_;
assign _1029_ = _0323_ | _0728_;
assign _1031_ = _0326_ | _0731_;
assign csr_rd_data_t0[31:13] = _0329_ | _0734_;
assign _1033_ = _0332_ | _0737_;
assign _1035_ = _0335_ | _0740_;
assign _1037_ = _0338_ | _0743_;
assign _1039_ = _0341_ | _0746_;
assign _1041_ = _0344_ | _0749_;
assign _1043_ = _0346_ | _0345_;
assign _1045_ = _0349_ | _0753_;
assign _1047_ = _0352_ | _0756_;
assign csr_rd_data_t0[2:0] = _0355_ | _0759_;
assign _1049_ = _0358_ | _0762_;
assign _1051_ = _0361_ | _0765_;
assign _1053_ = _0364_ | _0768_;
assign _1055_ = _0367_ | _0771_;
assign _1057_ = _0370_ | _0774_;
assign _1059_ = _0373_ | _0777_;
assign _1061_ = _0376_ | _0780_;
assign _1063_ = _0379_ | _0783_;
assign _1067_ = _0382_ | _0786_;
assign _1069_ = _0385_ | _0789_;
assign csr_rd_data_t0[11] = _0388_ | _0792_;
assign _1071_ = _0391_ | _0793_;
assign _1073_ = _0394_ | _0794_;
assign _1075_ = _0397_ | _0795_;
assign _1077_ = _0400_ | _0796_;
assign _1079_ = _0403_ | _0797_;
assign _1081_ = _0406_ | _0798_;
assign _1083_ = _0409_ | _0799_;
assign _1085_ = _0412_ | _0800_;
assign _1087_ = _0414_ | _0413_;
assign _1089_ = _0417_ | _0802_;
assign _1091_ = _0420_ | _0803_;
assign csr_rd_data_t0[3] = _0423_ | _0804_;
assign _1093_ = _0426_ | _0805_;
assign _1095_ = _0429_ | _0806_;
assign _1097_ = _0432_ | _0807_;
assign _1099_ = _0435_ | _0808_;
assign _1101_ = _0438_ | _0809_;
assign _1103_ = _0440_ | _0439_;
assign _1105_ = _0443_ | _0810_;
assign _1107_ = _0446_ | _0811_;
assign csr_rd_data_t0[6:4] = _0449_ | _0812_;
assign _1109_ = _0452_ | _0813_;
assign _1111_ = _0455_ | _0814_;
assign _1113_ = _0458_ | _0817_;
assign _1115_ = _0461_ | _0820_;
assign _1117_ = _0464_ | _0821_;
assign _1119_ = _0467_ | _0822_;
assign _1121_ = _0470_ | _0823_;
assign _1123_ = _0473_ | _0824_;
assign csr_rd_data_t0[12] = _0476_ | _0827_;
assign _1125_ = _0479_ | _0828_;
assign _1127_ = _0482_ | _0829_;
assign _1129_ = _0485_ | _0830_;
assign _1131_ = _0488_ | _0831_;
assign _1133_ = _0491_ | _0832_;
assign _1135_ = _0493_ | _0492_;
assign _1137_ = _0496_ | _0833_;
assign _1139_ = _0499_ | _0834_;
assign csr_rd_data_t0[10:8] = _0502_ | _0835_;
assign _1141_ = _0505_ | _0836_;
assign _1143_ = _0508_ | _0837_;
assign _1145_ = _0511_ | _0838_;
assign _1147_ = _0514_ | _0839_;
assign _1149_ = _0517_ | _0840_;
assign _1151_ = _0520_ | _0841_;
assign _1153_ = _0523_ | _0842_;
assign _1155_ = _0526_ | _0843_;
assign _1157_ = _0528_ | _0527_;
assign _1159_ = _0531_ | _0844_;
assign _1161_ = _0534_ | _0845_;
assign csr_rd_data_t0[7] = _0537_ | _0846_;
assign next_state_t0 = _0539_ | _0538_;
assign _1203_ = _0581_ | _0580_;
assign _1208_ = _0584_ | _0866_;
assign _1211_ = _0586_ | _0585_;
assign _1215_ = _0589_ | _0867_;
assign _1223_ = _0592_ | _0873_;
assign _1231_ = _0595_ | _0875_;
assign _1243_ = _0598_ | _0877_;
assign _1252_ = _0602_ | _0601_;
assign _1256_ = _0605_ | _0879_;
assign _1259_ = _0607_ | _0606_;
assign wr_data_t0 = _0611_ | _0883_;
assign _0016_ = | mip;
assign _0018_ = | { csr_wr_en, return_trap, activate_trap };
assign _0020_ = { _1206_, csr_wr_en } != 2'h1;
assign _0022_ = | { csr_wr_en, activate_trap };
assign _0024_ = { _1228_, csr_wr_en } != 2'h1;
assign _0026_ = { _1220_, csr_wr_en } != 2'h1;
assign _0028_ = { _1240_, csr_wr_en } != 2'h1;
assign _0030_ = | { return_trap, activate_trap };
assign _0032_ = | { csr_rdy, _1185_ };
assign _0034_ = | { _1171_, _1163_, csr_rdy };
assign _0036_ = { _1171_, csr_rd_vld } != 2'h2;
assign _0038_ = { _1163_, _1181_ } != 2'h2;
assign _0040_ = & { _0016_, rstz };
assign _0042_ = & { _0018_, _0020_ };
assign _0044_ = & { _1199_, csr_wr_en };
assign _0046_ = & { _1234_, csr_wr_en };
assign _0048_ = & { _1232_, csr_wr_en, rstz };
assign _0050_ = & { _0024_, _0022_, rstz };
assign _0052_ = & { _0026_, _0022_, rstz };
assign _0054_ = & { _0028_, _0022_, rstz };
assign _0056_ = & { _0030_, rstz };
assign _0058_ = & { _0038_, _0036_, _0034_ };
assign _0060_ = | { mip[2], mip[0] };
assign _0062_ = ~ _1250_;
assign _0061_ = ~ _1196_[1:0];
assign _0092_ = ~ _1199_;
assign _0131_ = ~ csr_data;
assign _0132_ = ~ wr_data;
assign _0285_ = _1176_ & _0089_;
assign _0288_ = _1229_ & _0091_;
assign _0291_ = _1200_ & _0093_;
assign _0202_ = csr_data_t0 & _0132_;
assign _0286_ = _1180_ & _0088_;
assign _0289_ = _1221_ & _0090_;
assign _0292_ = _1235_ & _0092_;
assign _0579_ = wr_data_t0 & _0131_;
assign _0287_ = _1176_ & _1180_;
assign _0290_ = _1229_ & _1221_;
assign _0293_ = _1200_ & _1235_;
assign _0204_ = csr_data_t0 & wr_data_t0;
assign _0701_ = _0285_ | _0286_;
assign _0702_ = _0288_ | _0289_;
assign _0703_ = _0291_ | _0292_;
assign _0860_ = _0202_ | _0579_;
assign _0613_ = _0701_ | _0287_;
assign _0615_ = _0702_ | _0290_;
assign _0617_ = _0703_ | _0293_;
assign _1195_ = _0860_ | _0204_;
assign _0612_ = _1175_ | _1179_;
assign _0614_ = _1228_ | _1220_;
assign _0616_ = _1199_ | _1234_;
assign _0151_ = | { _0612_, _1240_, _1177_, _1173_ };
assign _0153_ = | { _1179_, _1177_, _1175_ };
assign _0155_ = | { _1232_, _1228_, _1220_ };
assign _0157_ = | { _1248_, _1240_, _1179_, _1177_, _1175_, _1173_ };
assign _1014_ = _1246_ ? _1194_ : wr_data;
assign csr_wr_data = _1244_ ? _0002_ : _1014_;
assign _1016_ = _1179_ ? minstret[63:45] : mcycle[63:45];
assign _1018_ = _1173_ ? mcycle[31:13] : mtval[31:13];
assign _1020_ = _1177_ ? minstret[31:13] : _1018_;
assign _1022_ = _0612_ ? _1016_ : _1020_;
assign _1024_ = _1220_ ? mcause[31:13] : mepc[31:13];
assign _1026_ = _1234_ ? mtvec[31:13] : 19'h00000;
assign _1028_ = _1232_ ? mscratch[31:13] : _1026_;
assign _1030_ = _0614_ ? _1024_ : _1028_;
assign csr_rd_data[31:13] = _0151_ ? _1022_ : _1030_;
assign _1032_ = _1179_ ? minstret[34:32] : mcycle[34:32];
assign _1034_ = _1173_ ? mcycle[2:0] : mtval[2:0];
assign _1036_ = _1177_ ? minstret[2:0] : _1034_;
assign _1038_ = _0612_ ? _1032_ : _1036_;
assign _1040_ = _1220_ ? mcause[2:0] : mepc[2:0];
assign _1042_ = _1234_ ? { mtvec[2], 2'h0 } : 3'h0;
assign _1044_ = _1232_ ? mscratch[2:0] : _1042_;
assign _1046_ = _0614_ ? _1040_ : _1044_;
assign csr_rd_data[2:0] = _0151_ ? _1038_ : _1046_;
assign _1048_ = _1175_ ? mcycle[43] : minstret[11];
assign _1050_ = _1179_ ? minstret[43] : _1048_;
assign _1052_ = _1248_ ? mip[2] : mtval[11];
assign _1054_ = _1173_ ? mcycle[11] : _1052_;
assign _1056_ = _0153_ ? _1050_ : _1054_;
assign _1058_ = _1228_ ? mepc[11] : mscratch[11];
assign _1060_ = _1220_ ? mcause[11] : _1058_;
assign _1062_ = _1234_ ? mtvec[11] : mie[2];
assign _1066_ = _0616_ ? _1062_ : _1064_;
assign _1068_ = _0155_ ? _1060_ : _1066_;
assign csr_rd_data[11] = _0157_ ? _1056_ : _1068_;
assign _1070_ = _1175_ ? mcycle[35] : minstret[3];
assign _1072_ = _1179_ ? minstret[35] : _1070_;
assign _1074_ = _1248_ ? mip[0] : mtval[3];
assign _1076_ = _1173_ ? mcycle[3] : _1074_;
assign _1078_ = _0153_ ? _1072_ : _1076_;
assign _1080_ = _1228_ ? mepc[3] : mscratch[3];
assign _1082_ = _1220_ ? mcause[3] : _1080_;
assign _1084_ = _1234_ ? mtvec[3] : mie[0];
assign _1086_ = _1206_ ? mstatus[0] : 1'h0;
assign _1088_ = _0616_ ? _1084_ : _1086_;
assign _1090_ = _0155_ ? _1082_ : _1088_;
assign csr_rd_data[3] = _0157_ ? _1078_ : _1090_;
assign _1092_ = _1179_ ? minstret[38:36] : mcycle[38:36];
assign _1094_ = _1173_ ? mcycle[6:4] : mtval[6:4];
assign _1096_ = _1177_ ? minstret[6:4] : _1094_;
assign _1098_ = _0612_ ? _1092_ : _1096_;
assign _1100_ = _1220_ ? mcause[6:4] : mepc[6:4];
assign _1102_ = _1234_ ? mtvec[6:4] : 3'h0;
assign _1104_ = _1232_ ? mscratch[6:4] : _1102_;
assign _1106_ = _0614_ ? _1100_ : _1104_;
assign csr_rd_data[6:4] = _0151_ ? _1098_ : _1106_;
assign _1108_ = _1179_ ? minstret[44] : mcycle[44];
assign _1110_ = _1173_ ? mcycle[12] : mtval[12];
assign _1112_ = _1177_ ? minstret[12] : _1110_;
assign _1114_ = _0612_ ? _1108_ : _1112_;
assign _1116_ = _1228_ ? mepc[12] : mscratch[12];
assign _1118_ = _1220_ ? mcause[12] : _1116_;
assign _1064_ = _1206_ ? 1'h1 : 1'h0;
assign _1120_ = _1234_ ? mtvec[12] : _1064_;
assign _1122_ = _0155_ ? _1118_ : _1120_;
assign csr_rd_data[12] = _0151_ ? _1114_ : _1122_;
assign _1124_ = _1179_ ? minstret[42:40] : mcycle[42:40];
assign _1126_ = _1173_ ? mcycle[10:8] : mtval[10:8];
assign _1128_ = _1177_ ? minstret[10:8] : _1126_;
assign _1130_ = _0612_ ? _1124_ : _1128_;
assign _1132_ = _1220_ ? mcause[10:8] : mepc[10:8];
assign _1134_ = _1234_ ? mtvec[10:8] : 3'h0;
assign _1136_ = _1232_ ? mscratch[10:8] : _1134_;
assign _1138_ = _0614_ ? _1132_ : _1136_;
assign csr_rd_data[10:8] = _0151_ ? _1130_ : _1138_;
assign _1140_ = _1175_ ? mcycle[39] : minstret[7];
assign _1142_ = _1179_ ? minstret[39] : _1140_;
assign _1144_ = _1248_ ? mip[1] : mtval[7];
assign _1146_ = _1173_ ? mcycle[7] : _1144_;
assign _1148_ = _0153_ ? _1142_ : _1146_;
assign _1150_ = _1228_ ? mepc[7] : mscratch[7];
assign _1152_ = _1220_ ? mcause[7] : _1150_;
assign _1154_ = _1234_ ? mtvec[7] : mie[1];
assign _1156_ = _1206_ ? mstatus[1] : 1'h0;
assign _1158_ = _0616_ ? _1154_ : _1156_;
assign _1160_ = _0155_ ? _1152_ : _1158_;
assign csr_rd_data[7] = _0157_ ? _1148_ : _1160_;
assign _0978_ = _1171_ ? _0001_ : _0000_;
assign next_state = csr_rdy ? 2'h0 : _0978_;
assign _0171_ = | { _0019_, _0021_ };
assign _0172_ = | { _1200_, csr_wr_en_t0 };
assign _0173_ = | { _1235_, csr_wr_en_t0 };
assign _0174_ = | { _1233_, csr_wr_en_t0 };
assign _0175_ = | { _0023_, _0025_ };
assign _0176_ = | { _0023_, _0027_ };
assign _0177_ = | { _0023_, _0029_ };
assign _0178_ = | { _0035_, _0037_, _0039_ };
assign _0691_ = { _0016_, rstz } | { _0017_, 1'h0 };
assign _0692_ = { _0018_, _0020_ } | { _0019_, _0021_ };
assign _0693_ = { _1199_, csr_wr_en } | { _1200_, csr_wr_en_t0 };
assign _0694_ = { _1234_, csr_wr_en } | { _1235_, csr_wr_en_t0 };
assign _0695_ = { _1232_, csr_wr_en, rstz } | { _1233_, csr_wr_en_t0, 1'h0 };
assign _0696_ = { _0024_, _0022_, rstz } | { _0025_, _0023_, 1'h0 };
assign _0697_ = { _0026_, _0022_, rstz } | { _0027_, _0023_, 1'h0 };
assign _0698_ = { _0028_, _0022_, rstz } | { _0029_, _0023_, 1'h0 };
assign _0699_ = { _0030_, rstz } | { _0031_, 1'h0 };
assign _0700_ = { _0038_, _0036_, _0034_ } | { _0039_, _0037_, _0035_ };
assign _0141_ = & _0691_;
assign _0142_ = & _0692_;
assign _0143_ = & _0693_;
assign _0144_ = & _0694_;
assign _0145_ = & _0695_;
assign _0146_ = & _0696_;
assign _0147_ = & _0697_;
assign _0148_ = & _0698_;
assign _0149_ = & _0699_;
assign _0150_ = & _0700_;
assign _0041_ = _0017_ & _0141_;
assign _0043_ = _0171_ & _0142_;
assign _0045_ = _0172_ & _0143_;
assign _0047_ = _0173_ & _0144_;
assign _0049_ = _0174_ & _0145_;
assign _0051_ = _0175_ & _0146_;
assign _0053_ = _0176_ & _0147_;
assign _0055_ = _0177_ & _0148_;
assign _0057_ = _0031_ & _0149_;
assign _0059_ = _0178_ & _0150_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME core_interrupt_t0 */
always_ff @(posedge clk)
if (!rstz) core_interrupt_t0 <= 1'h0;
else core_interrupt_t0 <= _0017_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME mip_t0 */
always_ff @(posedge clk)
if (!rstz) mip_t0 <= 3'h0;
else mip_t0 <= { _0015_, _0011_, _0007_ };
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME trap_jump_t0 */
always_ff @(posedge clk)
if (!rstz) trap_jump_t0 <= 1'h0;
else trap_jump_t0 <= _1252_;
assign _0064_ = ~ _0040_;
assign _0885_ = _0979_[2] ^ core_interrupt_cause[2];
assign _0886_ = _1197_[3] ^ core_interrupt_cause[3];
assign _0898_ = _1253_[1:0] ^ trap_handle[1:0];
assign _0631_ = _1198_[3] | core_interrupt_cause_t0[3];
assign _0679_ = _1254_[1:0] | trap_handle_t0[1:0];
assign _0629_ = _0885_ | core_interrupt_cause_t0[2];
assign _0632_ = _0886_ | _0631_;
assign _0680_ = _0898_ | _0679_;
assign _0228_ = _0040_ & _1198_[3];
assign _0264_ = { _0056_, _0056_ } & _1254_[1:0];
assign _0226_ = _0064_ & core_interrupt_cause_t0[2];
assign _0229_ = _0064_ & core_interrupt_cause_t0[3];
assign _0265_ = { _0074_, _0074_ } & trap_handle_t0[1:0];
assign _0227_ = _0629_ & _0041_;
assign _0230_ = _0632_ & _0041_;
assign _0266_ = _0680_ & { _0057_, _0057_ };
assign _0633_ = _0228_ | _0229_;
assign _0681_ = _0264_ | _0265_;
assign _0630_ = _0226_ | _0227_;
assign _0634_ = _0633_ | _0230_;
assign _0682_ = _0681_ | _0266_;
reg core_interrupt_cause_t0_reg__2_ ;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME core_interrupt_cause_t0_reg__2_  */
always_ff @(posedge clk)
if (_0060_) core_interrupt_cause_t0_reg__2_  <= 1'h0;
else core_interrupt_cause_t0_reg__2_  <= _0630_;
assign core_interrupt_cause_t0[2] = core_interrupt_cause_t0_reg__2_ ;
reg core_interrupt_cause_t0_reg__3_ ;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME core_interrupt_cause_t0_reg__3_  */
always_ff @(posedge clk)
if (mip[2]) core_interrupt_cause_t0_reg__3_  <= 1'h0;
else core_interrupt_cause_t0_reg__3_  <= _0634_;
assign core_interrupt_cause_t0[3] = core_interrupt_cause_t0_reg__3_ ;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME trap_handle_t0[1:0] */
always_ff @(posedge clk)
if (activate_trap) trap_handle_t0[1:0] <= 2'h0;
else trap_handle_t0[1:0] <= _0682_;
assign _0065_ = ~ _0042_;
assign _0066_ = ~ _0044_;
assign _0067_ = ~ _0046_;
assign _0073_ = ~ _0032_;
assign _0075_ = ~ _0058_;
assign _0884_ = _1193_ ^ csr_wr_vld;
assign _0887_ = { _1207_, _1214_ } ^ mstatus[1:0];
assign _0888_ = csr_wr_data[11] ^ mie[2];
assign _0889_ = csr_wr_data[7] ^ mie[1];
assign _0890_ = csr_wr_data[3] ^ mie[0];
assign _0891_ = csr_wr_data[31:2] ^ mtvec[31:2];
assign _0897_ = _1258_ ^ regwr_csr;
assign _0900_ = next_state ^ state;
assign _0625_ = _1188_ | csr_wr_vld_t0;
assign _0635_ = { _1208_, _1215_ } | mstatus_t0[1:0];
assign _0639_ = csr_wr_data_t0[11] | mie_t0[2];
assign _0643_ = csr_wr_data_t0[7] | mie_t0[1];
assign _0647_ = csr_wr_data_t0[3] | mie_t0[0];
assign _0651_ = csr_wr_data_t0[31:2] | mtvec_t0[31:2];
assign _0675_ = _1259_ | regwr_csr_t0;
assign _0687_ = next_state_t0 | state_t0;
assign _0626_ = _0884_ | _0625_;
assign _0636_ = _0887_ | _0635_;
assign _0640_ = _0888_ | _0639_;
assign _0644_ = _0889_ | _0643_;
assign _0648_ = _0890_ | _0647_;
assign _0652_ = _0891_ | _0651_;
assign _0676_ = _0897_ | _0675_;
assign _0688_ = _0900_ | _0687_;
assign _0223_ = _1185_ & _1188_;
assign _0231_ = { _0042_, _0042_ } & { _1208_, _1215_ };
assign _0234_ = _0044_ & csr_wr_data_t0[11];
assign _0237_ = _0044_ & csr_wr_data_t0[7];
assign _0240_ = _0044_ & csr_wr_data_t0[3];
assign _0243_ = { _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_, _0046_ } & csr_wr_data_t0[31:2];
assign _0261_ = _0032_ & _1259_;
assign _0270_ = { _0058_, _0058_ } & next_state_t0;
assign _0224_ = _0063_ & csr_wr_vld_t0;
assign _0232_ = { _0065_, _0065_ } & mstatus_t0[1:0];
assign _0235_ = _0066_ & mie_t0[2];
assign _0238_ = _0066_ & mie_t0[1];
assign _0241_ = _0066_ & mie_t0[0];
assign _0244_ = { _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_ } & mtvec_t0[31:2];
assign _0262_ = _0073_ & regwr_csr_t0;
assign _0271_ = { _0075_, _0075_ } & state_t0;
assign _0225_ = _0626_ & _1186_;
assign _0233_ = _0636_ & { _0043_, _0043_ };
assign _0236_ = _0640_ & _0045_;
assign _0239_ = _0644_ & _0045_;
assign _0242_ = _0648_ & _0045_;
assign _0245_ = _0652_ & { _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_, _0047_ };
assign _0263_ = _0676_ & _0033_;
assign _0272_ = _0688_ & { _0059_, _0059_ };
assign _0627_ = _0223_ | _0224_;
assign _0637_ = _0231_ | _0232_;
assign _0641_ = _0234_ | _0235_;
assign _0645_ = _0237_ | _0238_;
assign _0649_ = _0240_ | _0241_;
assign _0653_ = _0243_ | _0244_;
assign _0677_ = _0261_ | _0262_;
assign _0689_ = _0270_ | _0271_;
assign _0628_ = _0627_ | _0225_;
assign _0638_ = _0637_ | _0233_;
assign _0642_ = _0641_ | _0236_;
assign _0646_ = _0645_ | _0239_;
assign _0650_ = _0649_ | _0242_;
assign _0654_ = _0653_ | _0245_;
assign _0678_ = _0677_ | _0263_;
assign _0690_ = _0689_ | _0272_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME csr_wr_vld_t0 */
always_ff @(posedge clk)
if (!rstz) csr_wr_vld_t0 <= 1'h0;
else csr_wr_vld_t0 <= _0628_;
reg [1:0] _2528_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME _2528_ */
always_ff @(posedge clk)
if (!rstz) _2528_ <= 2'h0;
else _2528_ <= _0638_;
assign mstatus_t0[1:0] = _2528_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME mie_t0[2] */
always_ff @(posedge clk)
if (!rstz) mie_t0[2] <= 1'h0;
else mie_t0[2] <= _0642_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME mie_t0[1] */
always_ff @(posedge clk)
if (!rstz) mie_t0[1] <= 1'h0;
else mie_t0[1] <= _0646_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME mie_t0[0] */
always_ff @(posedge clk)
if (!rstz) mie_t0[0] <= 1'h0;
else mie_t0[0] <= _0650_;
reg [29:0] _2532_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME _2532_ */
always_ff @(posedge clk)
if (!rstz) _2532_ <= 30'h00000000;
else _2532_ <= _0654_;
assign mtvec_t0[31:2] = _2532_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME regwr_csr_t0 */
always_ff @(posedge clk)
if (!rstz) regwr_csr_t0 <= 1'h0;
else regwr_csr_t0 <= _0678_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_23175af27fd2ffc5d196  */
/* PC_TAINT_INFO STATE_NAME state_t0 */
always_ff @(posedge clk)
if (!rstz) state_t0 <= 2'h0;
else state_t0 <= _0690_;
assign _1165_ = decode[131:129] == /* src = "generated/sv2v_out.v:425.22-425.38" */ 3'h2;
assign _1167_ = decode[131:129] == /* src = "generated/sv2v_out.v:425.44-425.60" */ 3'h3;
assign _1169_ = ! /* src = "generated/sv2v_out.v:425.67-425.86" */ decode[136:132];
assign _1181_ = csr_vld && /* src = "generated/sv2v_out.v:411.9-411.29" */ decode[6];
assign _1183_ = _1163_ && /* src = "generated/sv2v_out.v:424.13-424.39" */ csr_vld;
assign _1185_ = _1183_ && /* src = "generated/sv2v_out.v:424.12-424.53" */ decode[6];
assign _1187_ = _1189_ && /* src = "generated/sv2v_out.v:425.20-425.87" */ _1169_;
assign csr_rd_vld = mcycle_rd_vld && /* src = "generated/sv2v_out.v:430.22-430.54" */ minstret_rd_vld;
assign csr_rd_en = _1171_ && /* src = "generated/sv2v_out.v:431.21-431.50" */ csr_rd_vld;
assign csr_wr_en = csr_rdy && /* src = "generated/sv2v_out.v:432.21-432.50" */ csr_wr_vld;
assign mcycle_wrenl = csr_wr_en && /* src = "generated/sv2v_out.v:558.24-558.66" */ _1173_;
assign mcycle_wrenh = csr_wr_en && /* src = "generated/sv2v_out.v:559.24-559.67" */ _1175_;
assign minstret_wrenl = csr_wr_en && /* src = "generated/sv2v_out.v:573.26-573.70" */ _1177_;
assign minstret_wrenh = csr_wr_en && /* src = "generated/sv2v_out.v:574.26-574.71" */ _1179_;
assign _1189_ = _1165_ || /* src = "generated/sv2v_out.v:425.21-425.61" */ _1167_;
assign _1191_ = | /* src = "generated/sv2v_out.v:426.17-426.34" */ decode[128:124];
assign _1193_ = ~ /* src = "generated/sv2v_out.v:425.18-425.88" */ _1187_;
assign _1194_ = csr_data | /* src = "generated/sv2v_out.v:494.39-494.57" */ wr_data;
assign { _0979_[3:2], _1196_[1:0] } = mip[1] ? /* src = "generated/sv2v_out.v:555.13-555.19|generated/sv2v_out.v:555.9-556.58" */ 4'h7 : 4'hx;
assign _1197_ = mip[0] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:553.13-553.19|generated/sv2v_out.v:553.9-556.58" */ 4'h3 : { _0979_[3:2], _1196_[1:0] };
assign _1201_ = return_trap ? /* src = "generated/sv2v_out.v:535.13-535.24|generated/sv2v_out.v:535.9-538.7" */ 1'h1 : 1'hx;
assign _1202_ = activate_trap ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:528.13-528.26|generated/sv2v_out.v:528.9-538.7" */ mstatus[0] : _1201_;
assign _1204_ = _1206_ ? /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:512.5-527.12" */ csr_wr_data[7] : 1'hx;
assign _1207_ = csr_wr_en ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:511.8-511.17|generated/sv2v_out.v:511.4-538.7" */ _1204_ : _1202_;
assign _0982_ = return_trap ? /* src = "generated/sv2v_out.v:535.13-535.24|generated/sv2v_out.v:535.9-538.7" */ mstatus[1] : 1'hx;
assign _1210_ = activate_trap ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:528.13-528.26|generated/sv2v_out.v:528.9-538.7" */ 1'h0 : _0982_;
assign _1212_ = _1206_ ? /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:512.5-527.12" */ csr_wr_data[3] : 1'hx;
assign _1214_ = csr_wr_en ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:511.8-511.17|generated/sv2v_out.v:511.4-538.7" */ _1212_ : _1210_;
assign _1216_ = activate_trap ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:528.13-528.26|generated/sv2v_out.v:528.9-538.7" */ trap_cause : 32'hxxxxxxxx;
assign _1218_ = _1220_ ? /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:512.5-527.12" */ csr_wr_data : 32'hxxxxxxxx;
assign _1222_ = csr_wr_en ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:511.8-511.17|generated/sv2v_out.v:511.4-538.7" */ _1218_ : _1216_;
assign _1224_ = activate_trap ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:528.13-528.26|generated/sv2v_out.v:528.9-538.7" */ { decode[180:151], 2'h0 } : 32'hxxxxxxxx;
assign _1226_ = _1228_ ? /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:512.5-527.12" */ { csr_wr_data[31:2], 2'h0 } : 32'hxxxxxxxx;
assign _1230_ = csr_wr_en ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:511.8-511.17|generated/sv2v_out.v:511.4-538.7" */ _1226_ : _1224_;
assign _1236_ = activate_trap ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:528.13-528.26|generated/sv2v_out.v:528.9-538.7" */ trap_value : 32'hxxxxxxxx;
assign _1238_ = _1240_ ? /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:512.5-527.12" */ csr_wr_data : 32'hxxxxxxxx;
assign _1242_ = csr_wr_en ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:511.8-511.17|generated/sv2v_out.v:511.4-538.7" */ _1238_ : _1236_;
assign _1244_ = decode[130:129] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:493.3-497.10" */ 2'h3;
assign _1246_ = decode[130:129] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:493.3-497.10" */ 2'h2;
assign _1179_ = decode[148:137] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:463.3-488.10" */ 12'hb82;
assign _1175_ = decode[148:137] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:463.3-488.10" */ 12'hb80;
assign _1177_ = decode[148:137] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:463.3-488.10" */ 12'hb02;
assign _1173_ = decode[148:137] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:463.3-488.10" */ 12'hb00;
assign _1248_ = decode[148:137] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:463.3-488.10" */ 12'h344;
assign _1240_ = decode[148:137] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:463.3-488.10" */ 12'h343;
assign _1220_ = decode[148:137] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:463.3-488.10" */ 12'h342;
assign _1228_ = decode[148:137] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:463.3-488.10" */ 12'h341;
assign _1232_ = decode[148:137] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:463.3-488.10" */ 12'h340;
assign _1234_ = decode[148:137] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:463.3-488.10" */ 12'h305;
assign _1199_ = decode[148:137] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:463.3-488.10" */ 12'h304;
assign _1206_ = decode[148:137] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:463.3-488.10" */ 12'h300;
assign _1250_ = return_trap ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:443.12-443.23|generated/sv2v_out.v:443.8-448.22" */ 1'h1 : 1'h0;
assign _1251_ = activate_trap ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:439.12-439.25|generated/sv2v_out.v:439.8-448.22" */ 1'h1 : _1250_;
assign _1253_ = return_trap ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:443.12-443.23|generated/sv2v_out.v:443.8-448.22" */ mepc : 32'hxxxxxxxx;
assign _1255_ = activate_trap ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:439.12-439.25|generated/sv2v_out.v:439.8-448.22" */ { mtvec[31:2], 2'h0 } : _1253_;
assign _1257_ = csr_rdy ? /* src = "generated/sv2v_out.v:428.12-428.25|generated/sv2v_out.v:428.8-429.22" */ 1'h0 : 1'hx;
assign _1258_ = _1185_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:424.12-424.53|generated/sv2v_out.v:424.8-429.22" */ _1191_ : _1257_;
assign _0001_ = csr_rd_vld ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:414.9-414.19|generated/sv2v_out.v:414.5-415.24" */ 2'h2 : 2'hx;
assign _0000_ = _1181_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:411.9-411.29|generated/sv2v_out.v:411.5-412.24" */ 2'h1 : 2'hx;
assign csr_rdy = state == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:409.3-417.10" */ 2'h2;
assign _1171_ = state == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:409.3-417.10" */ 2'h1;
assign _1163_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:409.3-417.10" */ state;
assign _1260_ = | /* src = "generated/sv2v_out.v:550.22-550.28" */ mip;
assign wr_data = decode[131] ? /* src = "generated/sv2v_out.v:400.20-400.89" */ { 27'h0000000, decode[136:132] } : decode[116:85];
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:563.4-572.3" */
paramodsimplif_b656ed3944a4d79ba92b  u_hpmcounter0 (
.clk(clk),
.clk_t0(clk_t0),
.count(mcycle),
.count_t0(mcycle_t0),
.count_vld(mcycle_rd_vld),
.count_vld_t0(mcycle_rd_vld_t0),
.incr(1'h1),
.incr_t0(1'h0),
.load_data(csr_wr_data),
.load_data_t0(csr_wr_data_t0),
.load_high(mcycle_wrenh),
.load_high_t0(mcycle_wrenh_t0),
.load_low(mcycle_wrenl),
.load_low_t0(mcycle_wrenl_t0),
.rstz(rstz)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:578.4-587.3" */
paramodsimplif_b656ed3944a4d79ba92b  u_hpmcounter1 (
.clk(clk),
.clk_t0(clk_t0),
.count(minstret),
.count_t0(minstret_t0),
.count_vld(minstret_rd_vld),
.count_vld_t0(minstret_rd_vld_t0),
.incr(instret),
.incr_t0(instret_t0),
.load_data(csr_wr_data),
.load_data_t0(csr_wr_data_t0),
.load_high(minstret_wrenh),
.load_high_t0(minstret_wrenh_t0),
.load_low(minstret_wrenl),
.load_low_t0(minstret_wrenl_t0),
.rstz(rstz)
);
assign _0979_[1:0] = _0061_;
assign _1196_[3:2] = _0979_[3:2];
assign core_interrupt_cause[1:0] = 2'h3;
assign core_interrupt_cause_t0[1:0] = 2'h0;
assign mstatus[3:2] = 2'h3;
assign mstatus_t0[3:2] = 2'h0;
assign mtvec[1:0] = 2'h0;
assign mtvec_t0[1:0] = 2'h0;
// Added block to randomize initial values.
`ifdef RANDOMIZE_INIT
  initial begin
    mscratch_t0 = '0;
    mepc_t0 = '0;
    mcause_t0 = '0;
    mtval_t0 = '0;
    csr_data_t0 = '0;
    trap_handle_t0[31:2] = '0;
    csr_wr_vld = '0;
    core_interrupt = '0;
    core_interrupt_cause_reg__2_ = '0;
    core_interrupt_cause_reg__3_ = '0;
    _1442_ = '0;
    mie[2] = '0;
    mie[1] = '0;
    mie[0] = '0;
    mip = '0;
    _1447_ = '0;
    mscratch = '0;
    mepc = '0;
    mcause = '0;
    mtval = '0;
    trap_jump = '0;
    csr_data = '0;
    regwr_csr = '0;
    trap_handle[1:0] = '0;
    trap_handle[31:2] = '0;
    state = '0;
    core_interrupt_t0 = '0;
    mip_t0 = '0;
    trap_jump_t0 = '0;
    core_interrupt_cause_t0_reg__2_ = '0;
    core_interrupt_cause_t0_reg__3_ = '0;
    trap_handle_t0[1:0] = '0;
    csr_wr_vld_t0 = '0;
    _2528_ = '0;
    mie_t0[2] = '0;
    mie_t0[1] = '0;
    mie_t0[0] = '0;
    _2532_ = '0;
    regwr_csr_t0 = '0;
    state_t0 = '0;
  end
`endif // RANDOMIZE_INIT
endmodule

module paramodsimplif_8a2982a34f91f245ed13 (instr, base, offset, addr, misaligned_jmp, misaligned_ldst, instr_t0, addr_t0, base_t0, misaligned_jmp_t0, misaligned_ldst_t0, offset_t0);
/* src = "generated/sv2v_out.v:1678.4-1688.29" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1678.4-1688.29" */
wire _001_;
/* src = "generated/sv2v_out.v:1678.4-1688.29" */
wire _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1678.4-1688.29" */
wire _003_;
wire [31:0] _004_;
wire [31:0] _005_;
wire [4:0] _006_;
wire [1:0] _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire [1:0] _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire [31:0] _022_;
wire [31:0] _023_;
wire _024_;
wire _025_;
wire _026_;
wire [4:0] _027_;
wire [1:0] _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire [1:0] _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire [31:0] _052_;
wire [31:0] _053_;
wire [31:0] _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire [31:0] _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire [31:0] _071_;
wire [31:0] _072_;
/* src = "generated/sv2v_out.v:1666.31-1666.59" */
wire _073_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1666.31-1666.59" */
wire _074_;
/* src = "generated/sv2v_out.v:1666.101-1666.128" */
wire _075_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1666.101-1666.128" */
wire _076_;
/* src = "generated/sv2v_out.v:1679.10-1679.39" */
wire _077_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1679.10-1679.39" */
wire _078_;
/* src = "generated/sv2v_out.v:1679.45-1679.75" */
wire _079_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1679.45-1679.75" */
wire _080_;
/* src = "generated/sv2v_out.v:1680.11-1680.41" */
wire _081_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1680.11-1680.41" */
wire _082_;
/* src = "generated/sv2v_out.v:1682.16-1682.46" */
wire _083_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1682.16-1682.46" */
wire _084_;
/* src = "generated/sv2v_out.v:1680.10-1680.66" */
wire _085_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1680.10-1680.66" */
wire _086_;
/* src = "generated/sv2v_out.v:1682.15-1682.73" */
wire _087_;
/* src = "generated/sv2v_out.v:1666.30-1666.95" */
wire _088_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1666.30-1666.95" */
wire _089_;
/* src = "generated/sv2v_out.v:1666.29-1666.129" */
wire _090_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1666.29-1666.129" */
wire _091_;
/* src = "generated/sv2v_out.v:1679.9-1679.76" */
wire _092_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1679.9-1679.76" */
wire _093_;
/* src = "generated/sv2v_out.v:1666.135-1666.153" */
wire _094_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1666.135-1666.153" */
wire _095_;
/* src = "generated/sv2v_out.v:1644.20-1644.24" */
output [31:0] addr;
wire [31:0] addr;
/* src = "generated/sv2v_out.v:1650.13-1650.21" */
wire [31:0] addr_raw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1650.13-1650.21" */
wire [31:0] addr_raw_t0;
/* cellift = 32'd1 */
output [31:0] addr_t0;
wire [31:0] addr_t0;
/* src = "generated/sv2v_out.v:1649.7-1649.12" */
wire align;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1649.7-1649.12" */
wire align_t0;
/* src = "generated/sv2v_out.v:1642.20-1642.24" */
input [31:0] base;
wire [31:0] base;
/* cellift = 32'd1 */
input [31:0] base_t0;
wire [31:0] base_t0;
/* src = "generated/sv2v_out.v:1641.20-1641.25" */
input [31:0] instr;
wire [31:0] instr;
/* cellift = 32'd1 */
input [31:0] instr_t0;
wire [31:0] instr_t0;
/* src = "generated/sv2v_out.v:1645.14-1645.28" */
output misaligned_jmp;
wire misaligned_jmp;
/* cellift = 32'd1 */
output misaligned_jmp_t0;
wire misaligned_jmp_t0;
/* src = "generated/sv2v_out.v:1646.13-1646.28" */
output misaligned_ldst;
wire misaligned_ldst;
/* cellift = 32'd1 */
output misaligned_ldst_t0;
wire misaligned_ldst_t0;
/* src = "generated/sv2v_out.v:1643.20-1643.26" */
input [31:0] offset;
wire [31:0] offset;
/* cellift = 32'd1 */
input [31:0] offset_t0;
wire [31:0] offset_t0;
assign addr_raw = base + /* src = "generated/sv2v_out.v:1657.14-1657.27" */ offset;
assign addr[0] = _009_ & /* src = "generated/sv2v_out.v:1659.13-1659.33" */ addr_raw[0];
assign _004_ = ~ base_t0;
assign _005_ = ~ offset_t0;
assign _022_ = base & _004_;
assign _023_ = offset & _005_;
assign _071_ = _022_ + _023_;
assign _052_ = base | base_t0;
assign _053_ = offset | offset_t0;
assign _072_ = _052_ + _053_;
assign _064_ = _071_ ^ _072_;
assign _054_ = _064_ | base_t0;
assign addr_raw_t0 = _054_ | offset_t0;
assign _024_ = align_t0 & addr_raw[0];
assign _025_ = addr_raw_t0[0] & _009_;
assign _026_ = align_t0 & addr_raw_t0[0];
assign _055_ = _024_ | _025_;
assign addr_t0[0] = _055_ | _026_;
assign _017_ = | instr_t0[6:2];
assign _018_ = | instr_t0[13:12];
assign _006_ = ~ instr_t0[6:2];
assign _007_ = ~ instr_t0[13:12];
assign _027_ = instr[6:2] & _006_;
assign _028_ = instr[13:12] & _007_;
assign _065_ = _027_ == { _006_[4:3], 1'h0, _006_[1:0] };
assign _066_ = _027_ == { _006_[4:3], 2'h0, _006_[0] };
assign _067_ = _027_ == { _006_[4:3], 3'h0 };
assign _068_ = _027_ == { 1'h0, _006_[3], 3'h0 };
assign _069_ = _028_ == { _007_[1], 1'h0 };
assign _070_ = _028_ == { 1'h0, _007_[0] };
assign _074_ = _065_ & _017_;
assign align_t0 = _066_ & _017_;
assign _076_ = _067_ & _017_;
assign _080_ = _068_ & _017_;
assign _082_ = _069_ & _018_;
assign _084_ = _070_ & _018_;
assign _029_ = _091_ & _094_;
assign _032_ = _082_ & _094_;
assign _035_ = _084_ & addr[0];
assign _030_ = _095_ & _090_;
assign _033_ = _095_ & _081_;
assign _036_ = addr_t0[0] & _083_;
assign _031_ = _091_ & _095_;
assign _034_ = _082_ & _095_;
assign _037_ = _084_ & addr_t0[0];
assign _056_ = _029_ | _030_;
assign _057_ = _032_ | _033_;
assign _058_ = _035_ | _036_;
assign misaligned_jmp_t0 = _056_ | _031_;
assign _086_ = _057_ | _034_;
assign _003_ = _058_ | _037_;
assign _019_ = | { addr_raw_t0[1], addr_t0[0] };
assign _014_ = ~ { addr_raw_t0[1], addr_t0[0] };
assign _047_ = { addr_raw[1], addr[0] } & _014_;
assign _020_ = ! _027_;
assign _021_ = ! _047_;
assign _078_ = _020_ & _017_;
assign _095_ = _021_ & _019_;
assign _008_ = ~ _073_;
assign _010_ = ~ _088_;
assign _012_ = ~ _077_;
assign _009_ = ~ align;
assign _011_ = ~ _075_;
assign _013_ = ~ _079_;
assign _038_ = _074_ & _009_;
assign _041_ = _089_ & _011_;
assign _044_ = _078_ & _013_;
assign _039_ = align_t0 & _008_;
assign _042_ = _076_ & _010_;
assign _045_ = _080_ & _012_;
assign _040_ = _074_ & align_t0;
assign _043_ = _089_ & _076_;
assign _046_ = _078_ & _080_;
assign _059_ = _038_ | _039_;
assign _060_ = _041_ | _042_;
assign _061_ = _044_ | _045_;
assign _089_ = _059_ | _040_;
assign _091_ = _060_ | _043_;
assign _093_ = _061_ | _046_;
assign _015_ = ~ _085_;
assign _062_ = _086_ | _015_;
assign _063_ = _093_ | _092_;
assign _048_ = _003_ & _062_;
assign _050_ = _001_ & _063_;
assign _049_ = _086_ & _016_;
assign _051_ = _093_ & _000_;
assign _001_ = _049_ | _048_;
assign misaligned_ldst_t0 = _051_ | _050_;
assign _016_ = ~ _002_;
assign _073_ = instr[6:2] == /* src = "generated/sv2v_out.v:1666.31-1666.59" */ 5'h1b;
assign align = instr[6:2] == /* src = "generated/sv2v_out.v:1666.65-1666.94" */ 5'h19;
assign _075_ = instr[6:2] == /* src = "generated/sv2v_out.v:1666.101-1666.128" */ 5'h18;
assign _077_ = ! /* src = "generated/sv2v_out.v:1679.10-1679.39" */ instr[6:2];
assign _079_ = instr[6:2] == /* src = "generated/sv2v_out.v:1679.45-1679.75" */ 5'h08;
assign _081_ = instr[13:12] == /* src = "generated/sv2v_out.v:1680.11-1680.41" */ 2'h2;
assign _083_ = instr[13:12] == /* src = "generated/sv2v_out.v:1682.16-1682.46" */ 2'h1;
assign misaligned_jmp = _090_ && /* src = "generated/sv2v_out.v:1666.28-1666.154" */ _094_;
assign _085_ = _081_ && /* src = "generated/sv2v_out.v:1680.10-1680.66" */ _094_;
assign _087_ = _083_ && /* src = "generated/sv2v_out.v:1682.15-1682.73" */ addr[0];
assign _088_ = _073_ || /* src = "generated/sv2v_out.v:1666.30-1666.95" */ align;
assign _090_ = _088_ || /* src = "generated/sv2v_out.v:1666.29-1666.129" */ _075_;
assign _092_ = _077_ || /* src = "generated/sv2v_out.v:1679.9-1679.76" */ _079_;
assign _094_ = | /* src = "generated/sv2v_out.v:1680.47-1680.65" */ { addr_raw[1], addr[0] };
assign _002_ = _087_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1682.15-1682.73|generated/sv2v_out.v:1682.11-1685.30" */ 1'h1 : 1'h0;
assign _000_ = _085_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1680.10-1680.66|generated/sv2v_out.v:1680.6-1685.30" */ 1'h1 : _002_;
assign misaligned_ldst = _092_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1679.9-1679.76|generated/sv2v_out.v:1679.5-1688.29" */ _000_ : 1'h0;
assign addr[31:1] = addr_raw[31:1];
assign addr_t0[31:1] = addr_raw_t0[31:1];
endmodule

module paramodsimplif_db7b5d87aea4226b70fe (clk, rstz, instr_addr, instr_data, instr_req, instr_ack, fetch, immediate, regrd_rs1, regrd_rs2, regrd_rs1_en, regrd_rs2_en, fetch_vld, fetch_rdy, branch_target, branch, regwr_data, regwr_sel, regwr_en, clk_t0, branch_t0
, branch_target_t0, regwr_data_t0, regwr_en_t0, regwr_sel_t0, fetch_rdy_t0, immediate_t0, instr_data_t0, regrd_rs1_t0, regrd_rs1_en_t0, regrd_rs2_t0, regrd_rs2_en_t0, fetch_t0, fetch_vld_t0, instr_ack_t0, instr_addr_t0, instr_req_t0);
/* src = "generated/sv2v_out.v:1380.2-1392.6" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1380.2-1392.6" */
wire _001_;
/* src = "generated/sv2v_out.v:1380.2-1392.6" */
wire [31:0] _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1380.2-1392.6" */
wire [31:0] _003_;
/* src = "generated/sv2v_out.v:1328.2-1351.5" */
wire [1:0] _004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1328.2-1351.5" */
wire [1:0] _005_;
/* src = "generated/sv2v_out.v:1328.2-1351.5" */
wire [1:0] _006_;
/* src = "generated/sv2v_out.v:1328.2-1351.5" */
wire [1:0] _007_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1328.2-1351.5" */
wire [1:0] _008_;
/* src = "generated/sv2v_out.v:1328.2-1351.5" */
wire [1:0] _009_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1328.2-1351.5" */
wire [1:0] _010_;
/* src = "generated/sv2v_out.v:1311.11-1311.39" */
wire [31:0] _011_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1311.11-1311.39" */
wire [31:0] _012_;
/* src = "generated/sv2v_out.v:1318.10-1318.27" */
wire [31:0] _013_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1318.10-1318.27" */
wire [31:0] _014_;
wire _015_;
/* cellift = 32'd1 */
wire _016_;
wire _017_;
/* cellift = 32'd1 */
wire _018_;
wire _019_;
/* cellift = 32'd1 */
wire _020_;
wire _021_;
/* cellift = 32'd1 */
wire _022_;
wire _023_;
/* cellift = 32'd1 */
wire _024_;
wire _025_;
/* cellift = 32'd1 */
wire _026_;
wire _027_;
/* cellift = 32'd1 */
wire _028_;
wire _029_;
wire [31:0] _030_;
wire [31:0] _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire [1:0] _036_;
wire [2:0] _037_;
wire [1:0] _038_;
wire [1:0] _039_;
wire _040_;
wire _041_;
wire [1:0] _042_;
wire [1:0] _043_;
wire [1:0] _044_;
wire _045_;
wire _046_;
wire [31:0] _047_;
wire [31:0] _048_;
wire [31:0] _049_;
wire _050_;
wire _051_;
wire [1:0] _052_;
wire [1:0] _053_;
wire [1:0] _054_;
wire [1:0] _055_;
wire [31:0] _056_;
wire _057_;
wire [31:0] _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire [31:0] _082_;
wire [31:0] _083_;
wire [31:0] _084_;
wire [31:0] _085_;
wire [31:0] _086_;
wire [31:0] _087_;
wire [31:0] _088_;
wire [31:0] _089_;
wire _090_;
wire _091_;
wire _092_;
wire [31:0] _093_;
wire [31:0] _094_;
wire [31:0] _095_;
wire [31:0] _096_;
wire [31:0] _097_;
wire [31:0] _098_;
wire [31:0] _099_;
wire [31:0] _100_;
wire [31:0] _101_;
wire [1:0] _102_;
wire [2:0] _103_;
wire [1:0] _104_;
wire [1:0] _105_;
wire _106_;
wire _107_;
wire _108_;
wire [1:0] _109_;
wire [1:0] _110_;
wire [1:0] _111_;
wire [1:0] _112_;
wire [1:0] _113_;
wire [1:0] _114_;
wire [1:0] _115_;
wire [1:0] _116_;
wire [1:0] _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire [31:0] _135_;
wire [31:0] _136_;
wire [31:0] _137_;
wire [31:0] _138_;
wire [31:0] _139_;
wire [31:0] _140_;
wire [31:0] _141_;
wire [31:0] _142_;
wire [31:0] _143_;
wire _144_;
wire _145_;
wire [1:0] _146_;
wire [1:0] _147_;
wire [1:0] _148_;
wire [1:0] _149_;
wire [1:0] _150_;
wire [1:0] _151_;
wire [1:0] _152_;
wire [1:0] _153_;
wire [1:0] _154_;
wire [31:0] _155_;
wire [31:0] _156_;
wire [31:0] _157_;
wire [31:0] _158_;
wire [31:0] _159_;
wire [31:0] _160_;
wire [31:0] _161_;
wire [31:0] _162_;
wire [31:0] _163_;
wire [31:0] _164_;
wire _165_;
wire _166_;
wire [31:0] _167_;
wire [31:0] _168_;
wire [31:0] _169_;
wire [31:0] _170_;
wire [31:0] _171_;
wire [31:0] _172_;
wire [31:0] _173_;
wire [31:0] _174_;
wire [31:0] _175_;
wire [31:0] _176_;
wire [31:0] _177_;
wire [31:0] _178_;
wire [31:0] _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire [31:0] _184_;
wire [31:0] _185_;
wire [31:0] _186_;
wire [31:0] _187_;
wire [31:0] _188_;
wire [31:0] _189_;
wire [31:0] _190_;
wire [31:0] _191_;
wire [31:0] _192_;
wire [31:0] _193_;
wire [31:0] _194_;
wire [31:0] _195_;
wire [1:0] _196_;
wire [3:0] _197_;
wire [3:0] _198_;
wire _199_;
wire [1:0] _200_;
wire [1:0] _201_;
wire [1:0] _202_;
wire [1:0] _203_;
wire [1:0] _204_;
wire [1:0] _205_;
wire [1:0] _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire [31:0] _214_;
wire [31:0] _215_;
wire [31:0] _216_;
wire [31:0] _217_;
wire [31:0] _218_;
wire [31:0] _219_;
wire [31:0] _220_;
wire [31:0] _221_;
wire [31:0] _222_;
wire [31:0] _223_;
wire _224_;
wire [1:0] _225_;
wire [1:0] _226_;
wire [1:0] _227_;
wire [1:0] _228_;
wire [1:0] _229_;
wire [31:0] _230_;
wire [31:0] _231_;
wire [31:0] _232_;
wire [31:0] _233_;
wire [31:0] _234_;
wire [31:0] _235_;
wire [31:0] _236_;
wire _237_;
wire [31:0] _238_;
wire [31:0] _239_;
wire [31:0] _240_;
wire _241_;
/* cellift = 32'd1 */
wire _242_;
wire [31:0] _243_;
wire [31:0] _244_;
wire [31:0] _245_;
wire [31:0] _246_;
wire _247_;
wire [31:0] _248_;
wire [31:0] _249_;
wire [31:0] _250_;
wire [1:0] _251_;
wire [1:0] _252_;
wire [31:0] _253_;
wire [31:0] _254_;
wire [31:0] _255_;
wire _256_;
wire [1:0] _257_;
wire [31:0] _258_;
wire [31:0] _259_;
wire [31:0] _260_;
wire [31:0] _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire [31:0] _267_;
wire [31:0] _268_;
wire [31:0] _269_;
wire [31:0] _270_;
wire [1:0] _271_;
/* cellift = 32'd1 */
wire [1:0] _272_;
wire [1:0] _273_;
/* cellift = 32'd1 */
wire [1:0] _274_;
/* src = "generated/sv2v_out.v:1317.12-1317.30" */
wire _275_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1317.12-1317.30" */
wire _276_;
/* src = "generated/sv2v_out.v:1357.14-1357.27" */
wire _277_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1357.14-1357.27" */
wire _278_;
/* src = "generated/sv2v_out.v:1357.33-1357.46" */
wire _279_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1357.33-1357.46" */
wire _280_;
/* src = "generated/sv2v_out.v:1366.13-1366.26" */
wire _281_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1366.13-1366.26" */
wire _282_;
/* src = "generated/sv2v_out.v:1357.12-1357.61" */
wire _283_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1357.12-1357.61" */
wire _284_;
/* src = "generated/sv2v_out.v:1366.12-1366.40" */
wire _285_;
/* src = "generated/sv2v_out.v:1371.12-1371.34" */
wire _286_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1371.12-1371.34" */
wire _287_;
/* src = "generated/sv2v_out.v:1378.18-1378.68" */
wire _288_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1378.18-1378.68" */
wire _289_;
/* src = "generated/sv2v_out.v:1381.7-1381.70" */
wire _290_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1381.7-1381.70" */
wire _291_;
/* src = "generated/sv2v_out.v:1357.13-1357.47" */
wire _292_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1357.13-1357.47" */
wire _293_;
/* src = "generated/sv2v_out.v:1373.20-1373.30" */
wire _294_;
/* src = "generated/sv2v_out.v:1378.58-1378.68" */
wire _295_;
wire [31:0] _296_;
/* cellift = 32'd1 */
wire [31:0] _297_;
wire [31:0] _298_;
/* cellift = 32'd1 */
wire [31:0] _299_;
wire [31:0] _300_;
/* cellift = 32'd1 */
wire [31:0] _301_;
wire [31:0] _302_;
/* cellift = 32'd1 */
wire [31:0] _303_;
wire [31:0] _304_;
/* cellift = 32'd1 */
wire [31:0] _305_;
wire [31:0] _306_;
/* cellift = 32'd1 */
wire [31:0] _307_;
wire _308_;
wire _309_;
/* cellift = 32'd1 */
wire _310_;
wire _311_;
wire _312_;
/* cellift = 32'd1 */
wire _313_;
/* unused_bits = "1" */
wire [1:0] _314_;
/* cellift = 32'd1 */
/* unused_bits = "1" */
wire [1:0] _315_;
wire [31:0] _316_;
/* cellift = 32'd1 */
wire [31:0] _317_;
wire [31:0] _318_;
/* cellift = 32'd1 */
wire [31:0] _319_;
wire [31:0] _320_;
/* cellift = 32'd1 */
wire [31:0] _321_;
wire [31:0] _322_;
/* cellift = 32'd1 */
wire [31:0] _323_;
/* src = "generated/sv2v_out.v:1378.18-1378.83" */
wire [31:0] _324_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1378.18-1378.83" */
wire [31:0] _325_;
/* src = "generated/sv2v_out.v:1292.13-1292.19" */
input branch;
wire branch;
/* cellift = 32'd1 */
input branch_t0;
wire branch_t0;
/* src = "generated/sv2v_out.v:1291.20-1291.33" */
input [31:0] branch_target;
wire [31:0] branch_target;
/* cellift = 32'd1 */
input [31:0] branch_target_t0;
wire [31:0] branch_target_t0;
/* src = "generated/sv2v_out.v:1277.13-1277.16" */
input clk;
wire clk;
/* cellift = 32'd1 */
input clk_t0;
wire clk_t0;
/* src = "generated/sv2v_out.v:1283.20-1283.25" */
output [63:0] fetch;
reg [63:0] fetch;
/* src = "generated/sv2v_out.v:1290.13-1290.22" */
input fetch_rdy;
wire fetch_rdy;
/* cellift = 32'd1 */
input fetch_rdy_t0;
wire fetch_rdy_t0;
/* cellift = 32'd1 */
output [63:0] fetch_t0;
reg [63:0] fetch_t0;
/* src = "generated/sv2v_out.v:1289.13-1289.22" */
output fetch_vld;
reg fetch_vld;
/* cellift = 32'd1 */
output fetch_vld_t0;
reg fetch_vld_t0;
/* src = "generated/sv2v_out.v:1284.21-1284.30" */
output [31:0] immediate;
wire [31:0] immediate;
/* cellift = 32'd1 */
output [31:0] immediate_t0;
wire [31:0] immediate_t0;
/* src = "generated/sv2v_out.v:1282.13-1282.22" */
input instr_ack;
wire instr_ack;
/* cellift = 32'd1 */
input instr_ack_t0;
wire instr_ack_t0;
/* src = "generated/sv2v_out.v:1279.20-1279.30" */
output [31:0] instr_addr;
wire [31:0] instr_addr;
/* cellift = 32'd1 */
output [31:0] instr_addr_t0;
wire [31:0] instr_addr_t0;
/* src = "generated/sv2v_out.v:1280.20-1280.30" */
input [31:0] instr_data;
wire [31:0] instr_data;
/* cellift = 32'd1 */
input [31:0] instr_data_t0;
wire [31:0] instr_data_t0;
/* src = "generated/sv2v_out.v:1281.14-1281.23" */
output instr_req;
wire instr_req;
/* cellift = 32'd1 */
output instr_req_t0;
wire instr_req_t0;
/* src = "generated/sv2v_out.v:1300.6-1300.15" */
wire instr_vld;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1300.6-1300.15" */
wire instr_vld_t0;
/* src = "generated/sv2v_out.v:1301.13-1301.23" */
wire [31:0] next_instr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1301.13-1301.23" */
wire [31:0] next_instr_t0;
/* src = "generated/sv2v_out.v:1303.12-1303.22" */
wire [1:0] next_state;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1303.12-1303.22" */
wire [1:0] next_state_t0;
/* src = "generated/sv2v_out.v:1296.13-1296.15" */
reg [31:0] pc /* verilator public */;
/* src = "generated/sv2v_out.v:1297.13-1297.20" */
reg [31:0] pc_last;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1297.13-1297.20" */
reg [31:0] pc_last_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1296.13-1296.15" */
reg [31:0] pc_t0 /* verilator public */;
/* src = "generated/sv2v_out.v:1299.7-1299.15" */
wire pipe_rdy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1299.7-1299.15" */
wire pipe_rdy_t0;
/* src = "generated/sv2v_out.v:1285.21-1285.30" */
output [31:0] regrd_rs1;
wire [31:0] regrd_rs1;
/* src = "generated/sv2v_out.v:1287.14-1287.26" */
output regrd_rs1_en;
wire regrd_rs1_en;
/* cellift = 32'd1 */
output regrd_rs1_en_t0;
wire regrd_rs1_en_t0;
/* cellift = 32'd1 */
output [31:0] regrd_rs1_t0;
wire [31:0] regrd_rs1_t0;
/* src = "generated/sv2v_out.v:1286.21-1286.30" */
output [31:0] regrd_rs2;
wire [31:0] regrd_rs2;
/* src = "generated/sv2v_out.v:1288.14-1288.26" */
output regrd_rs2_en;
wire regrd_rs2_en;
/* cellift = 32'd1 */
output regrd_rs2_en_t0;
wire regrd_rs2_en_t0;
/* cellift = 32'd1 */
output [31:0] regrd_rs2_t0;
wire [31:0] regrd_rs2_t0;
/* src = "generated/sv2v_out.v:1293.20-1293.30" */
input [31:0] regwr_data;
wire [31:0] regwr_data;
/* cellift = 32'd1 */
input [31:0] regwr_data_t0;
wire [31:0] regwr_data_t0;
/* src = "generated/sv2v_out.v:1295.13-1295.21" */
input regwr_en;
wire regwr_en;
/* cellift = 32'd1 */
input regwr_en_t0;
wire regwr_en_t0;
/* src = "generated/sv2v_out.v:1294.19-1294.28" */
input [4:0] regwr_sel;
wire [4:0] regwr_sel;
/* cellift = 32'd1 */
input [4:0] regwr_sel_t0;
wire [4:0] regwr_sel_t0;
/* src = "generated/sv2v_out.v:1278.13-1278.17" */
input rstz;
wire rstz;
/* src = "generated/sv2v_out.v:1298.13-1298.24" */
reg [31:0] skid_buffer;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1298.13-1298.24" */
reg [31:0] skid_buffer_t0;
/* src = "generated/sv2v_out.v:1302.12-1302.17" */
reg [1:0] state;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1302.12-1302.17" */
reg [1:0] state_t0;
assign _011_ = branch_target + /* src = "generated/sv2v_out.v:1311.11-1311.39" */ 32'd4;
assign _013_ = pc + /* src = "generated/sv2v_out.v:1318.10-1318.27" */ 32'd4;
assign _030_ = ~ branch_target_t0;
assign _031_ = ~ pc_t0;
assign _082_ = branch_target & _030_;
assign _083_ = pc & _031_;
assign _267_ = _082_ + 32'd4;
assign _269_ = _083_ + 32'd4;
assign _170_ = branch_target | branch_target_t0;
assign _171_ = pc | pc_t0;
assign _268_ = _170_ + 32'd4;
assign _270_ = _171_ + 32'd4;
assign _243_ = _267_ ^ _268_;
assign _244_ = _269_ ^ _270_;
assign _012_ = _243_ | branch_target_t0;
assign _014_ = _244_ | pc_t0;
assign _249_ = _300_ ^ fetch[63:32];
assign _250_ = _306_ ^ fetch[31:0];
assign _034_ = ~ _025_;
assign _035_ = ~ _027_;
assign _184_ = instr_data_t0 | skid_buffer_t0;
assign _188_ = _301_ | fetch_t0[63:32];
assign _192_ = _307_ | fetch_t0[31:0];
assign _185_ = _248_ | _184_;
assign _189_ = _249_ | _188_;
assign _193_ = _250_ | _192_;
assign _093_ = { _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_ } & instr_data_t0;
assign _096_ = { _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_ } & _301_;
assign _099_ = { _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_ } & _307_;
assign _094_ = { _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_ } & skid_buffer_t0;
assign _097_ = { _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_ } & fetch_t0[63:32];
assign _100_ = { _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_ } & fetch_t0[31:0];
assign _095_ = _185_ & { _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_ };
assign _098_ = _189_ & { _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_ };
assign _101_ = _193_ & { _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_ };
assign _186_ = _093_ | _094_;
assign _190_ = _096_ | _097_;
assign _194_ = _099_ | _100_;
assign _187_ = _186_ | _095_;
assign _191_ = _190_ | _098_;
assign _195_ = _194_ | _101_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_db7b5d87aea4226b70fe  */
/* PC_TAINT_INFO STATE_NAME skid_buffer_t0 */
always_ff @(posedge clk)
skid_buffer_t0 <= _187_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_db7b5d87aea4226b70fe  */
/* PC_TAINT_INFO STATE_NAME fetch_t0[63:32] */
always_ff @(posedge clk)
fetch_t0[63:32] <= _191_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_db7b5d87aea4226b70fe  */
/* PC_TAINT_INFO STATE_NAME fetch_t0[31:0] */
always_ff @(posedge clk)
fetch_t0[31:0] <= _195_;
assign _072_ = | { pipe_rdy_t0, _284_ };
assign _077_ = | next_state_t0;
assign _078_ = | state_t0;
assign _038_ = ~ { _284_, pipe_rdy_t0 };
assign _044_ = ~ next_state_t0;
assign _054_ = ~ state_t0;
assign _104_ = { _283_, pipe_rdy } & _038_;
assign _117_ = next_state & _044_;
assign _152_ = state & _054_;
assign _262_ = _104_ == { _038_[1], 1'h0 };
assign _263_ = _117_ == { 1'h0, _044_[0] };
assign _264_ = _152_ == _054_;
assign _265_ = _152_ == { _054_[1], 1'h0 };
assign _266_ = _152_ == { 1'h0, _054_[0] };
assign _020_ = _262_ & _072_;
assign _276_ = _263_ & _077_;
assign _282_ = _264_ & _078_;
assign _280_ = _265_ & _078_;
assign _278_ = _266_ & _078_;
/* src = "generated/sv2v_out.v:1321.2-1327.24" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_db7b5d87aea4226b70fe  */
/* PC_TAINT_INFO STATE_NAME state[0] */
always_ff @(posedge clk)
if (!rstz) state[0] <= 1'h0;
else state[0] <= _314_[0];
/* src = "generated/sv2v_out.v:1321.2-1327.24" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_db7b5d87aea4226b70fe  */
/* PC_TAINT_INFO STATE_NAME state[1] */
always_ff @(posedge clk)
if (_029_) state[1] <= 1'h0;
else state[1] <= next_state[1];
/* src = "generated/sv2v_out.v:1304.2-1320.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_db7b5d87aea4226b70fe  */
/* PC_TAINT_INFO STATE_NAME pc_last */
always_ff @(posedge clk)
if (!rstz) pc_last <= 32'd0;
else if (_015_) pc_last <= _318_;
/* src = "generated/sv2v_out.v:1304.2-1320.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_db7b5d87aea4226b70fe  */
/* PC_TAINT_INFO STATE_NAME pc */
always_ff @(posedge clk)
if (!rstz) pc <= 32'd2147483648;
else if (_015_) pc <= _322_;
/* src = "generated/sv2v_out.v:1352.2-1372.22" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_db7b5d87aea4226b70fe  */
/* PC_TAINT_INFO STATE_NAME fetch_vld */
always_ff @(posedge clk)
if (_029_) fetch_vld <= 1'h0;
else if (_023_) fetch_vld <= _312_;
/* src = "generated/sv2v_out.v:1352.2-1372.22" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_db7b5d87aea4226b70fe  */
/* PC_TAINT_INFO STATE_NAME skid_buffer */
always_ff @(posedge clk)
if (_025_) skid_buffer <= instr_data;
/* src = "generated/sv2v_out.v:1352.2-1372.22" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_db7b5d87aea4226b70fe  */
/* PC_TAINT_INFO STATE_NAME fetch[63:32] */
always_ff @(posedge clk)
if (_027_) fetch[63:32] <= _300_;
/* src = "generated/sv2v_out.v:1352.2-1372.22" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_db7b5d87aea4226b70fe  */
/* PC_TAINT_INFO STATE_NAME fetch[31:0] */
always_ff @(posedge clk)
if (_027_) fetch[31:0] <= _306_;
assign _118_ = fetch_vld_t0 & fetch_rdy;
assign _121_ = _293_ & _295_;
assign _124_ = _293_ & instr_ack;
assign _125_ = _284_ & pipe_rdy;
assign _128_ = _282_ & fetch_rdy;
assign _122_ = instr_ack_t0 & _292_;
assign _126_ = pipe_rdy_t0 & _283_;
assign _129_ = fetch_rdy_t0 & _281_;
assign _123_ = _293_ & instr_ack_t0;
assign _127_ = _284_ & pipe_rdy_t0;
assign _130_ = _282_ & fetch_rdy_t0;
assign _207_ = _118_ | _119_;
assign _208_ = _121_ | _122_;
assign _209_ = _124_ | _122_;
assign _210_ = _125_ | _126_;
assign _211_ = _128_ | _129_;
assign _287_ = _207_ | _120_;
assign _289_ = _208_ | _123_;
assign _284_ = _209_ | _123_;
assign _291_ = _210_ | _127_;
assign _001_ = _211_ | _130_;
assign _070_ = | { _276_, branch_t0 };
assign _071_ = | { _001_, _284_, _287_ };
assign _073_ = | { _001_, _284_ };
assign _036_ = ~ { _276_, branch_t0 };
assign _037_ = ~ { _001_, _284_, _287_ };
assign _039_ = ~ { _001_, _284_ };
assign _102_ = { _275_, branch } & _036_;
assign _103_ = { _285_, _283_, _286_ } & _037_;
assign _105_ = { _285_, _283_ } & _039_;
assign _079_ = ! _102_;
assign _080_ = ! _103_;
assign _081_ = ! _105_;
assign _016_ = _079_ & _070_;
assign _018_ = _080_ & _071_;
assign _022_ = _081_ & _073_;
assign _046_ = ~ _277_;
assign _045_ = ~ fetch_rdy;
assign _040_ = ~ _279_;
assign _131_ = fetch_vld_t0 & _045_;
assign _132_ = _278_ & _040_;
assign _119_ = fetch_rdy_t0 & fetch_vld;
assign _133_ = _280_ & _046_;
assign _120_ = fetch_vld_t0 & fetch_rdy_t0;
assign _134_ = _278_ & _280_;
assign _212_ = _131_ | _119_;
assign _213_ = _132_ | _133_;
assign pipe_rdy_t0 = _212_ | _120_;
assign _293_ = _213_ | _134_;
assign _042_ = ~ { _281_, _281_ };
assign _043_ = ~ { _241_, _241_ };
assign _049_ = ~ { _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_ };
assign _050_ = ~ pipe_rdy;
assign _051_ = ~ _283_;
assign _052_ = ~ { fetch_rdy, fetch_rdy };
assign _053_ = ~ { instr_ack, instr_ack };
assign _055_ = ~ { branch, branch };
assign _047_ = ~ { branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch };
assign _048_ = ~ { _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_ };
assign _056_ = ~ { _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_ };
assign _057_ = ~ _290_;
assign _058_ = ~ { _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_ };
assign _200_ = { _282_, _282_ } | _042_;
assign _204_ = { _242_, _242_ } | _043_;
assign _220_ = { _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_ } | _049_;
assign _224_ = _284_ | _051_;
assign _225_ = { fetch_rdy_t0, fetch_rdy_t0 } | _052_;
assign _226_ = { instr_ack_t0, instr_ack_t0 } | _053_;
assign _229_ = { branch_t0, branch_t0 } | _055_;
assign _214_ = { branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0 } | _047_;
assign _217_ = { _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_ } | _048_;
assign _234_ = { _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_ } | _056_;
assign _237_ = _291_ | _057_;
assign _238_ = { _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_ } | _058_;
assign _201_ = { _282_, _282_ } | { _281_, _281_ };
assign _203_ = { _278_, _278_ } | { _277_, _277_ };
assign _205_ = { _242_, _242_ } | { _241_, _241_ };
assign _219_ = { pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0, pipe_rdy_t0 } | { pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy, pipe_rdy };
assign _221_ = { _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_ } | { _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_ };
assign _227_ = { instr_ack_t0, instr_ack_t0 } | { instr_ack, instr_ack };
assign _230_ = { _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_ } | { _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_ };
assign _215_ = { branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0 } | { branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch, branch };
assign _218_ = { _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_ } | { _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_ };
assign _235_ = { _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_ } | { _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_, _290_ };
assign _239_ = { _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_ } | { _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_, _288_ };
assign _109_ = _008_ & _200_;
assign _114_ = _274_ & _204_;
assign _135_ = _325_ & _214_;
assign _138_ = _297_ & _220_;
assign _141_ = _303_ & _220_;
assign _144_ = _310_ & _224_;
assign _146_ = state_t0 & _225_;
assign _148_ = state_t0 & _226_;
assign _153_ = next_state_t0 & _229_;
assign _155_ = _317_ & _214_;
assign _157_ = _321_ & _214_;
assign _160_ = instr_data_t0 & _217_;
assign _162_ = _003_ & _234_;
assign _165_ = _001_ & _237_;
assign _167_ = pc_t0 & _238_;
assign _110_ = _010_ & _201_;
assign _112_ = _005_ & _203_;
assign _115_ = _272_ & _205_;
assign _297_ = pc_last_t0 & _218_;
assign _299_ = pc_last_t0 & _219_;
assign _139_ = _299_ & _221_;
assign _305_ = instr_data_t0 & _219_;
assign _142_ = _305_ & _221_;
assign _149_ = { pipe_rdy_t0, 1'h0 } & _227_;
assign _317_ = pc_t0 & _230_;
assign _136_ = branch_target_t0 & _215_;
assign _321_ = _014_ & _230_;
assign _158_ = _012_ & _215_;
assign _303_ = skid_buffer_t0 & _218_;
assign _163_ = instr_data_t0 & _235_;
assign _168_ = pc_last_t0 & _239_;
assign _202_ = _109_ | _110_;
assign _206_ = _114_ | _115_;
assign _216_ = _135_ | _136_;
assign _222_ = _138_ | _139_;
assign _223_ = _141_ | _142_;
assign _228_ = _148_ | _149_;
assign _231_ = _155_ | _136_;
assign _232_ = _157_ | _158_;
assign _233_ = _160_ | _303_;
assign _236_ = _162_ | _163_;
assign _240_ = _167_ | _168_;
assign _251_ = _007_ ^ _009_;
assign _252_ = _273_ ^ _271_;
assign _253_ = _324_ ^ branch_target;
assign _254_ = _296_ ^ _298_;
assign _255_ = _302_ ^ _304_;
assign _256_ = _309_ ^ _311_;
assign _257_ = state ^ _006_;
assign _258_ = _316_ ^ branch_target;
assign _259_ = _320_ ^ _011_;
assign _248_ = instr_data ^ skid_buffer;
assign _260_ = _002_ ^ instr_data;
assign _261_ = pc ^ pc_last;
assign _111_ = { _282_, _282_ } & _251_;
assign _113_ = { _278_, _278_ } & { _004_[1], _060_ };
assign _116_ = { _242_, _242_ } & _252_;
assign _137_ = { branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0 } & _253_;
assign _140_ = { _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_ } & _254_;
assign _143_ = { _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_ } & _255_;
assign _310_ = _001_ & _062_;
assign _145_ = _284_ & _256_;
assign _147_ = { fetch_rdy_t0, fetch_rdy_t0 } & { state[1], _061_ };
assign _150_ = { instr_ack_t0, instr_ack_t0 } & _257_;
assign _151_ = { instr_ack_t0, instr_ack_t0 } & { _059_, _006_[0] };
assign _154_ = { branch_t0, branch_t0 } & { next_state[1], _063_ };
assign _156_ = { branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0 } & _258_;
assign _159_ = { branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0, branch_t0 } & _259_;
assign _161_ = { _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_, _001_ } & _248_;
assign _164_ = { _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_, _291_ } & _260_;
assign _166_ = _291_ & _064_;
assign _169_ = { _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_, _289_ } & _261_;
assign _272_ = _111_ | _202_;
assign _274_ = _113_ | _112_;
assign next_state_t0 = _116_ | _206_;
assign instr_addr_t0 = _137_ | _216_;
assign _301_ = _140_ | _222_;
assign _307_ = _143_ | _223_;
assign _313_ = _145_ | _144_;
assign _010_ = _147_ | _146_;
assign _008_ = _150_ | _228_;
assign _005_ = _151_ | _149_;
assign _315_ = _154_ | _153_;
assign _319_ = _156_ | _231_;
assign _323_ = _159_ | _232_;
assign _003_ = _161_ | _233_;
assign next_instr_t0 = _164_ | _236_;
assign instr_vld_t0 = _166_ | _165_;
assign _325_ = _169_ | _240_;
assign _015_ = | { _275_, branch };
assign _017_ = | { _285_, _283_, _286_ };
assign _019_ = { _283_, pipe_rdy } != 2'h2;
assign _021_ = | { _285_, _283_ };
assign _066_ = ~ branch;
assign _023_ = & { _019_, _017_ };
assign _025_ = & { _050_, _066_, _283_, rstz };
assign _027_ = & { _019_, _066_, _021_, rstz };
assign _065_ = ~ rstz;
assign _029_ = | { _065_, branch };
assign _062_ = ~ _308_;
assign _064_ = ~ _000_;
assign _059_ = ~ _006_[1];
assign _060_ = ~ _004_[0];
assign _061_ = ~ state[0];
assign _063_ = ~ next_state[0];
assign _041_ = ~ _281_;
assign _106_ = _280_ & _041_;
assign _107_ = _282_ & _040_;
assign _108_ = _280_ & _282_;
assign _199_ = _106_ | _107_;
assign _242_ = _199_ | _108_;
assign _241_ = _279_ | _281_;
assign _271_ = _281_ ? _009_ : _007_;
assign _273_ = _277_ ? _004_ : 2'h1;
assign next_state = _241_ ? _271_ : _273_;
assign _074_ = | { _020_, _018_ };
assign _075_ = | { pipe_rdy_t0, _284_, branch_t0 };
assign _076_ = | { _022_, _020_, branch_t0 };
assign _196_ = { _019_, _017_ } | { _020_, _018_ };
assign _197_ = { _066_, _050_, _283_, rstz } | { branch_t0, pipe_rdy_t0, _284_, 1'h0 };
assign _198_ = { _019_, _066_, _021_, rstz } | { _020_, branch_t0, _022_, 1'h0 };
assign _067_ = & _196_;
assign _068_ = & _197_;
assign _069_ = & _198_;
assign _024_ = _074_ & _067_;
assign _026_ = _075_ & _068_;
assign _028_ = _076_ & _069_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_db7b5d87aea4226b70fe  */
/* PC_TAINT_INFO STATE_NAME state_t0[0] */
always_ff @(posedge clk)
if (!rstz) state_t0[0] <= 1'h0;
else state_t0[0] <= _315_[0];
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_db7b5d87aea4226b70fe  */
/* PC_TAINT_INFO STATE_NAME state_t0[1] */
always_ff @(posedge clk)
if (_029_) state_t0[1] <= 1'h0;
else state_t0[1] <= next_state_t0[1];
assign _032_ = ~ _015_;
assign _033_ = ~ _023_;
assign _245_ = _318_ ^ pc_last;
assign _246_ = _322_ ^ pc;
assign _247_ = _312_ ^ fetch_vld;
assign _172_ = _319_ | pc_last_t0;
assign _176_ = _323_ | pc_t0;
assign _180_ = _313_ | fetch_vld_t0;
assign _173_ = _245_ | _172_;
assign _177_ = _246_ | _176_;
assign _181_ = _247_ | _180_;
assign _084_ = { _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_ } & _319_;
assign _087_ = { _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_ } & _323_;
assign _090_ = _023_ & _313_;
assign _085_ = { _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_ } & pc_last_t0;
assign _088_ = { _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_ } & pc_t0;
assign _091_ = _033_ & fetch_vld_t0;
assign _086_ = _173_ & { _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_ };
assign _089_ = _177_ & { _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_ };
assign _092_ = _181_ & _024_;
assign _174_ = _084_ | _085_;
assign _178_ = _087_ | _088_;
assign _182_ = _090_ | _091_;
assign _175_ = _174_ | _086_;
assign _179_ = _178_ | _089_;
assign _183_ = _182_ | _092_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_db7b5d87aea4226b70fe  */
/* PC_TAINT_INFO STATE_NAME pc_last_t0 */
always_ff @(posedge clk)
if (!rstz) pc_last_t0 <= 32'd0;
else pc_last_t0 <= _175_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_db7b5d87aea4226b70fe  */
/* PC_TAINT_INFO STATE_NAME pc_t0 */
always_ff @(posedge clk)
if (!rstz) pc_t0 <= 32'd0;
else pc_t0 <= _179_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_db7b5d87aea4226b70fe  */
/* PC_TAINT_INFO STATE_NAME fetch_vld_t0 */
always_ff @(posedge clk)
if (_029_) fetch_vld_t0 <= 1'h0;
else fetch_vld_t0 <= _183_;
assign _275_ = next_state == /* src = "generated/sv2v_out.v:1317.12-1317.30" */ 2'h1;
assign _286_ = fetch_vld && /* src = "generated/sv2v_out.v:1371.12-1371.34" */ fetch_rdy;
assign _288_ = _292_ && /* src = "generated/sv2v_out.v:1378.18-1378.68" */ _295_;
assign _283_ = _292_ && /* src = "generated/sv2v_out.v:1381.8-1381.57" */ instr_ack;
assign _290_ = _283_ && /* src = "generated/sv2v_out.v:1381.7-1381.70" */ pipe_rdy;
assign _285_ = _281_ && /* src = "generated/sv2v_out.v:1385.12-1385.40" */ fetch_rdy;
assign pipe_rdy = _294_ || /* src = "generated/sv2v_out.v:1373.20-1373.43" */ fetch_rdy;
assign _292_ = _277_ || /* src = "generated/sv2v_out.v:1381.9-1381.43" */ _279_;
assign _294_ = ~ /* src = "generated/sv2v_out.v:1373.20-1373.30" */ fetch_vld;
assign _295_ = ~ /* src = "generated/sv2v_out.v:1378.58-1378.68" */ instr_ack;
assign instr_addr = branch ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1375.7-1375.27|generated/sv2v_out.v:1375.3-1378.85" */ branch_target : _324_;
assign _296_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1366.12-1366.40|generated/sv2v_out.v:1366.8-1372.22" */ pc_last : 32'hxxxxxxxx;
assign _298_ = pipe_rdy ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1358.8-1358.16|generated/sv2v_out.v:1358.4-1364.31" */ pc_last : 32'hxxxxxxxx;
assign _300_ = _283_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1357.12-1357.61|generated/sv2v_out.v:1357.8-1372.22" */ _298_ : _296_;
assign _302_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1366.12-1366.40|generated/sv2v_out.v:1366.8-1372.22" */ skid_buffer : 32'hxxxxxxxx;
assign _304_ = pipe_rdy ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1358.8-1358.16|generated/sv2v_out.v:1358.4-1364.31" */ instr_data : 32'hxxxxxxxx;
assign _306_ = _283_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1357.12-1357.61|generated/sv2v_out.v:1357.8-1372.22" */ _304_ : _302_;
assign _308_ = _286_ ? /* src = "generated/sv2v_out.v:1371.12-1371.34|generated/sv2v_out.v:1371.8-1372.22" */ 1'h0 : 1'hx;
assign _309_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1366.12-1366.40|generated/sv2v_out.v:1366.8-1372.22" */ 1'h1 : _308_;
assign _311_ = pipe_rdy ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1358.8-1358.16|generated/sv2v_out.v:1358.4-1364.31" */ 1'h1 : 1'hx;
assign _312_ = _283_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1357.12-1357.61|generated/sv2v_out.v:1357.8-1372.22" */ _311_ : _309_;
assign _009_ = fetch_rdy ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1348.9-1348.18|generated/sv2v_out.v:1348.5-1349.24" */ 2'h1 : state;
assign _007_ = instr_ack ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1342.9-1342.18|generated/sv2v_out.v:1342.5-1346.25" */ _006_ : state;
assign _006_ = pipe_rdy ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1334.10-1334.18|generated/sv2v_out.v:1334.6-1337.25" */ 2'h1 : 2'h3;
assign _004_ = instr_ack ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1333.9-1333.18|generated/sv2v_out.v:1333.5-1340.24" */ _006_ : 2'h2;
assign _281_ = state == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1330.3-1350.10" */ 2'h3;
assign _279_ = state == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1330.3-1350.10" */ 2'h2;
assign _277_ = state == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1330.3-1350.10" */ 2'h1;
assign _314_ = branch ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1324.12-1324.18|generated/sv2v_out.v:1324.8-1327.24" */ 2'h1 : next_state;
assign _316_ = _275_ ? /* src = "generated/sv2v_out.v:1317.12-1317.30|generated/sv2v_out.v:1317.8-1320.6" */ pc : 32'hxxxxxxxx;
assign _318_ = branch ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1309.12-1309.18|generated/sv2v_out.v:1309.8-1320.6" */ branch_target : _316_;
assign _320_ = _275_ ? /* src = "generated/sv2v_out.v:1317.12-1317.30|generated/sv2v_out.v:1317.8-1320.6" */ _013_ : 32'hxxxxxxxx;
assign _322_ = branch ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1309.12-1309.18|generated/sv2v_out.v:1309.8-1320.6" */ _011_ : _320_;
assign _002_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1385.12-1385.40|generated/sv2v_out.v:1385.8-1392.6" */ skid_buffer : instr_data;
assign _000_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1385.12-1385.40|generated/sv2v_out.v:1385.8-1392.6" */ 1'h1 : 1'h0;
assign next_instr = _290_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1381.7-1381.70|generated/sv2v_out.v:1381.3-1392.6" */ instr_data : _002_;
assign instr_vld = _290_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1381.7-1381.70|generated/sv2v_out.v:1381.3-1392.6" */ 1'h1 : _000_;
assign _324_ = _288_ ? /* src = "generated/sv2v_out.v:1378.18-1378.83" */ pc_last : pc;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:1393.12-1407.3" */
kronos_RF u_rf (
.clk(clk),
.clk_t0(clk_t0),
.fetch_rdy(fetch_rdy),
.fetch_rdy_t0(fetch_rdy_t0),
.immediate(immediate),
.immediate_t0(immediate_t0),
.instr_data(next_instr),
.instr_data_t0(next_instr_t0),
.instr_vld(instr_vld),
.instr_vld_t0(instr_vld_t0),
.regrd_rs1(regrd_rs1),
.regrd_rs1_en(regrd_rs1_en),
.regrd_rs1_en_t0(regrd_rs1_en_t0),
.regrd_rs1_t0(regrd_rs1_t0),
.regrd_rs2(regrd_rs2),
.regrd_rs2_en(regrd_rs2_en),
.regrd_rs2_en_t0(regrd_rs2_en_t0),
.regrd_rs2_t0(regrd_rs2_t0),
.regwr_data(regwr_data),
.regwr_data_t0(regwr_data_t0),
.regwr_en(regwr_en),
.regwr_en_t0(regwr_en_t0),
.regwr_sel(regwr_sel),
.regwr_sel_t0(regwr_sel_t0),
.rstz(rstz)
);
assign instr_req = 1'h1;
assign instr_req_t0 = 1'h0;
// Added block to randomize initial values.
`ifdef RANDOMIZE_INIT
  initial begin
    skid_buffer_t0 = '0;
    fetch_t0[63:32] = '0;
    fetch_t0[31:0] = '0;
    state[0] = '0;
    state[1] = '0;
    pc_last = '0;
    pc = '0;
    fetch_vld = '0;
    skid_buffer = '0;
    fetch[63:32] = '0;
    fetch[31:0] = '0;
    state_t0[0] = '0;
    state_t0[1] = '0;
    pc_last_t0 = '0;
    pc_t0 = '0;
    fetch_vld_t0 = '0;
  end
`endif // RANDOMIZE_INIT
endmodule

module paramodsimplif_1b215dccbb32fdcc253c (clk, rstz, instr_addr, instr_data, instr_req, instr_ack, data_addr, data_rd_data, data_wr_data, data_mask, data_wr_en, data_req, data_ack, software_interrupt, timer_interrupt, external_interrupt, clk_t0, timer_interrupt_t0, software_interrupt_t0, external_interrupt_t0, data_ack_t0
, data_addr_t0, data_mask_t0, data_rd_data_t0, data_req_t0, data_wr_data_t0, data_wr_en_t0, instr_data_t0, instr_ack_t0, instr_addr_t0, instr_req_t0);
/* src = "generated/sv2v_out.v:174.7-174.13" */
wire branch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:174.7-174.13" */
wire branch_t0;
/* src = "generated/sv2v_out.v:173.14-173.27" */
wire [31:0] branch_target;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:173.14-173.27" */
wire [31:0] branch_target_t0;
/* src = "generated/sv2v_out.v:152.13-152.16" */
input clk;
wire clk;
/* cellift = 32'd1 */
input clk_t0;
wire clk_t0;
/* src = "generated/sv2v_out.v:164.13-164.21" */
input data_ack;
wire data_ack;
/* cellift = 32'd1 */
input data_ack_t0;
wire data_ack_t0;
/* src = "generated/sv2v_out.v:158.21-158.30" */
output [31:0] data_addr;
wire [31:0] data_addr;
/* cellift = 32'd1 */
output [31:0] data_addr_t0;
wire [31:0] data_addr_t0;
/* src = "generated/sv2v_out.v:161.20-161.29" */
output [3:0] data_mask;
wire [3:0] data_mask;
/* cellift = 32'd1 */
output [3:0] data_mask_t0;
wire [3:0] data_mask_t0;
/* src = "generated/sv2v_out.v:159.20-159.32" */
input [31:0] data_rd_data;
wire [31:0] data_rd_data;
/* cellift = 32'd1 */
input [31:0] data_rd_data_t0;
wire [31:0] data_rd_data_t0;
/* src = "generated/sv2v_out.v:163.14-163.22" */
output data_req;
wire data_req;
/* cellift = 32'd1 */
output data_req_t0;
wire data_req_t0;
/* src = "generated/sv2v_out.v:160.21-160.33" */
output [31:0] data_wr_data;
wire [31:0] data_wr_data;
/* cellift = 32'd1 */
output [31:0] data_wr_data_t0;
wire [31:0] data_wr_data_t0;
/* src = "generated/sv2v_out.v:162.14-162.24" */
output data_wr_en;
wire data_wr_en;
/* cellift = 32'd1 */
output data_wr_en_t0;
wire data_wr_en_t0;
/* src = "generated/sv2v_out.v:180.15-180.21" */
wire [180:0] decode;
/* src = "generated/sv2v_out.v:184.7-184.17" */
wire decode_rdy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:184.7-184.17" */
wire decode_rdy_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:180.15-180.21" */
wire [180:0] decode_t0;
/* src = "generated/sv2v_out.v:183.7-183.17" */
wire decode_vld;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:183.7-183.17" */
wire decode_vld_t0;
/* src = "generated/sv2v_out.v:167.13-167.31" */
input external_interrupt;
wire external_interrupt;
/* cellift = 32'd1 */
input external_interrupt_t0;
wire external_interrupt_t0;
/* src = "generated/sv2v_out.v:179.14-179.19" */
wire [63:0] fetch;
/* src = "generated/sv2v_out.v:182.7-182.16" */
wire fetch_rdy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:182.7-182.16" */
wire fetch_rdy_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:179.14-179.19" */
wire [63:0] fetch_t0;
/* src = "generated/sv2v_out.v:181.7-181.16" */
wire fetch_vld;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:181.7-181.16" */
wire fetch_vld_t0;
/* src = "generated/sv2v_out.v:168.14-168.23" */
wire [31:0] immediate;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:168.14-168.23" */
wire [31:0] immediate_t0;
/* src = "generated/sv2v_out.v:157.13-157.22" */
input instr_ack;
wire instr_ack;
/* cellift = 32'd1 */
input instr_ack_t0;
wire instr_ack_t0;
/* src = "generated/sv2v_out.v:154.21-154.31" */
output [31:0] instr_addr;
wire [31:0] instr_addr;
/* cellift = 32'd1 */
output [31:0] instr_addr_t0;
wire [31:0] instr_addr_t0;
/* src = "generated/sv2v_out.v:155.20-155.30" */
input [31:0] instr_data;
wire [31:0] instr_data;
/* cellift = 32'd1 */
input [31:0] instr_data_t0;
wire [31:0] instr_data_t0;
/* src = "generated/sv2v_out.v:156.14-156.23" */
output instr_req;
wire instr_req;
/* cellift = 32'd1 */
output instr_req_t0;
wire instr_req_t0;
/* src = "generated/sv2v_out.v:169.14-169.23" */
wire [31:0] regrd_rs1;
/* src = "generated/sv2v_out.v:171.7-171.19" */
wire regrd_rs1_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:171.7-171.19" */
wire regrd_rs1_en_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:169.14-169.23" */
wire [31:0] regrd_rs1_t0;
/* src = "generated/sv2v_out.v:170.14-170.23" */
wire [31:0] regrd_rs2;
/* src = "generated/sv2v_out.v:172.7-172.19" */
wire regrd_rs2_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:172.7-172.19" */
wire regrd_rs2_en_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:170.14-170.23" */
wire [31:0] regrd_rs2_t0;
/* src = "generated/sv2v_out.v:175.14-175.24" */
wire [31:0] regwr_data;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:175.14-175.24" */
wire [31:0] regwr_data_t0;
/* src = "generated/sv2v_out.v:177.7-177.15" */
wire regwr_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:177.7-177.15" */
wire regwr_en_t0;
/* src = "generated/sv2v_out.v:185.7-185.20" */
wire regwr_pending;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:185.7-185.20" */
wire regwr_pending_t0;
/* src = "generated/sv2v_out.v:176.13-176.22" */
wire [4:0] regwr_sel;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:176.13-176.22" */
wire [4:0] regwr_sel_t0;
/* src = "generated/sv2v_out.v:153.13-153.17" */
input rstz;
wire rstz;
/* src = "generated/sv2v_out.v:165.13-165.31" */
input software_interrupt;
wire software_interrupt;
/* cellift = 32'd1 */
input software_interrupt_t0;
wire software_interrupt_t0;
/* src = "generated/sv2v_out.v:166.13-166.28" */
input timer_interrupt;
wire timer_interrupt;
/* cellift = 32'd1 */
input timer_interrupt_t0;
wire timer_interrupt_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:238.4-260.3" */
paramodsimplif_9e9afc4272f55a9beacc  u_ex (
.branch(branch),
.branch_t0(branch_t0),
.branch_target(branch_target),
.branch_target_t0(branch_target_t0),
.clk(clk),
.clk_t0(clk_t0),
.data_ack(data_ack),
.data_ack_t0(data_ack_t0),
.data_addr(data_addr),
.data_addr_t0(data_addr_t0),
.data_mask(data_mask),
.data_mask_t0(data_mask_t0),
.data_rd_data(data_rd_data),
.data_rd_data_t0(data_rd_data_t0),
.data_req(data_req),
.data_req_t0(data_req_t0),
.data_wr_data(data_wr_data),
.data_wr_data_t0(data_wr_data_t0),
.data_wr_en(data_wr_en),
.data_wr_en_t0(data_wr_en_t0),
.decode(decode),
.decode_rdy(decode_rdy),
.decode_rdy_t0(decode_rdy_t0),
.decode_t0(decode_t0),
.decode_vld(decode_vld),
.decode_vld_t0(decode_vld_t0),
.external_interrupt(external_interrupt),
.external_interrupt_t0(external_interrupt_t0),
.regwr_data(regwr_data),
.regwr_data_t0(regwr_data_t0),
.regwr_en(regwr_en),
.regwr_en_t0(regwr_en_t0),
.regwr_pending(regwr_pending),
.regwr_pending_t0(regwr_pending_t0),
.regwr_sel(regwr_sel),
.regwr_sel_t0(regwr_sel_t0),
.rstz(rstz),
.software_interrupt(software_interrupt),
.software_interrupt_t0(software_interrupt_t0),
.timer_interrupt(timer_interrupt),
.timer_interrupt_t0(timer_interrupt_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:214.4-233.3" */
paramodsimplif_62dbb6e3107130a7cf75  u_id (
.clk(clk),
.clk_t0(clk_t0),
.decode(decode),
.decode_rdy(decode_rdy),
.decode_rdy_t0(decode_rdy_t0),
.decode_t0(decode_t0),
.decode_vld(decode_vld),
.decode_vld_t0(decode_vld_t0),
.fetch(fetch),
.fetch_rdy(fetch_rdy),
.fetch_rdy_t0(fetch_rdy_t0),
.fetch_t0(fetch_t0),
.fetch_vld(fetch_vld),
.fetch_vld_t0(fetch_vld_t0),
.flush(branch),
.flush_t0(branch_t0),
.immediate(immediate),
.immediate_t0(immediate_t0),
.regrd_rs1(regrd_rs1),
.regrd_rs1_en(regrd_rs1_en),
.regrd_rs1_en_t0(regrd_rs1_en_t0),
.regrd_rs1_t0(regrd_rs1_t0),
.regrd_rs2(regrd_rs2),
.regrd_rs2_en(regrd_rs2_en),
.regrd_rs2_en_t0(regrd_rs2_en_t0),
.regrd_rs2_t0(regrd_rs2_t0),
.regwr_data(regwr_data),
.regwr_data_t0(regwr_data_t0),
.regwr_en(regwr_en),
.regwr_en_t0(regwr_en_t0),
.regwr_pending(regwr_pending),
.regwr_pending_t0(regwr_pending_t0),
.regwr_sel(regwr_sel),
.regwr_sel_t0(regwr_sel_t0),
.rstz(rstz)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:189.4-209.3" */
paramodsimplif_db7b5d87aea4226b70fe  u_if (
.branch(branch),
.branch_t0(branch_t0),
.branch_target(branch_target),
.branch_target_t0(branch_target_t0),
.clk(clk),
.clk_t0(clk_t0),
.fetch(fetch),
.fetch_rdy(fetch_rdy),
.fetch_rdy_t0(fetch_rdy_t0),
.fetch_t0(fetch_t0),
.fetch_vld(fetch_vld),
.fetch_vld_t0(fetch_vld_t0),
.immediate(immediate),
.immediate_t0(immediate_t0),
.instr_ack(instr_ack),
.instr_ack_t0(instr_ack_t0),
.instr_addr(instr_addr),
.instr_addr_t0(instr_addr_t0),
.instr_data(instr_data),
.instr_data_t0(instr_data_t0),
.instr_req(instr_req),
.instr_req_t0(instr_req_t0),
.regrd_rs1(regrd_rs1),
.regrd_rs1_en(regrd_rs1_en),
.regrd_rs1_en_t0(regrd_rs1_en_t0),
.regrd_rs1_t0(regrd_rs1_t0),
.regrd_rs2(regrd_rs2),
.regrd_rs2_en(regrd_rs2_en),
.regrd_rs2_en_t0(regrd_rs2_en_t0),
.regrd_rs2_t0(regrd_rs2_t0),
.regwr_data(regwr_data),
.regwr_data_t0(regwr_data_t0),
.regwr_en(regwr_en),
.regwr_en_t0(regwr_en_t0),
.regwr_sel(regwr_sel),
.regwr_sel_t0(regwr_sel_t0),
.rstz(rstz)
);
endmodule

module paramodsimplif_62dbb6e3107130a7cf75 (clk, rstz, flush, fetch, immediate, regrd_rs1, regrd_rs2, regrd_rs1_en, regrd_rs2_en, fetch_vld, fetch_rdy, decode, decode_vld, decode_rdy, regwr_data, regwr_sel, regwr_en, regwr_pending, clk_t0, decode_t0, decode_rdy_t0
, decode_vld_t0, regwr_data_t0, regwr_en_t0, regwr_pending_t0, regwr_sel_t0, fetch_rdy_t0, immediate_t0, regrd_rs1_t0, regrd_rs1_en_t0, regrd_rs2_t0, regrd_rs2_en_t0, fetch_t0, fetch_vld_t0, flush_t0);
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0001_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0003_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0005_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0007_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0009_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0011_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0013_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0015_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0016_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0017_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0018_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0019_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0021_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0022_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0023_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire [3:0] _0024_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire [3:0] _0025_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0026_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0027_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0028_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0029_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0030_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0031_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire [3:0] _0032_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire [3:0] _0033_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire [31:0] _0034_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire [31:0] _0035_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0036_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0037_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire [3:0] _0038_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire [3:0] _0039_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0040_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0041_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0042_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0043_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
/* unused_bits = "1" */
wire [1:0] _0044_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
/* unused_bits = "1" */
wire [1:0] _0045_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire [1:0] _0046_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire [1:0] _0047_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire [1:0] _0048_;
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0049_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1020.2-1188.5" */
wire _0050_;
wire _0051_;
/* cellift = 32'd1 */
wire _0052_;
wire _0053_;
/* cellift = 32'd1 */
wire _0054_;
wire _0055_;
wire _0056_;
wire _0057_;
wire _0058_;
/* cellift = 32'd1 */
wire _0059_;
wire _0060_;
/* cellift = 32'd1 */
wire _0061_;
wire _0062_;
wire _0063_;
/* cellift = 32'd1 */
wire _0064_;
wire _0065_;
/* cellift = 32'd1 */
wire _0066_;
wire _0067_;
/* cellift = 32'd1 */
wire _0068_;
wire _0069_;
/* cellift = 32'd1 */
wire _0070_;
wire _0071_;
wire _0072_;
wire [1:0] _0073_;
wire [2:0] _0074_;
wire [2:0] _0075_;
wire [4:0] _0076_;
wire [2:0] _0077_;
wire [5:0] _0078_;
wire [5:0] _0079_;
wire [1:0] _0080_;
wire _0081_;
wire _0082_;
wire _0083_;
wire _0084_;
wire _0085_;
wire _0086_;
wire _0087_;
wire _0088_;
wire _0089_;
wire [3:0] _0090_;
wire _0091_;
wire _0092_;
wire _0093_;
wire _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire [31:0] _0101_;
wire [31:0] _0102_;
wire [31:0] _0103_;
wire [31:0] _0104_;
wire [31:0] _0105_;
wire [3:0] _0106_;
wire [31:0] _0107_;
wire [31:0] _0108_;
wire [31:0] _0109_;
wire [1:0] _0110_;
wire [6:0] _0111_;
wire [3:0] _0112_;
wire [4:0] _0113_;
wire [4:0] _0114_;
wire [11:0] _0115_;
wire [4:0] _0116_;
wire [4:0] _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire [1:0] _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire [1:0] _0136_;
wire _0137_;
wire [1:0] _0138_;
wire _0139_;
wire _0140_;
wire [31:0] _0141_;
wire [2:0] _0142_;
wire _0143_;
wire [2:0] _0144_;
wire [3:0] _0145_;
wire [2:0] _0146_;
wire [4:0] _0147_;
wire [5:0] _0148_;
wire [4:0] _0149_;
wire [31:0] _0150_;
wire [3:0] _0151_;
wire [1:0] _0152_;
wire [31:0] _0153_;
wire [31:0] _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire [3:0] _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
/* cellift = 32'd1 */
wire _0169_;
/* cellift = 32'd1 */
wire _0170_;
/* cellift = 32'd1 */
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire _0186_;
wire _0187_;
wire _0188_;
wire _0189_;
wire _0190_;
wire _0191_;
wire _0192_;
wire _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire _0199_;
/* cellift = 32'd1 */
wire _0200_;
wire _0201_;
wire _0202_;
wire _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
wire _0221_;
wire _0222_;
wire _0223_;
wire _0224_;
wire _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire _0241_;
wire _0242_;
wire _0243_;
wire _0244_;
wire _0245_;
wire _0246_;
wire _0247_;
wire _0248_;
wire _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire [31:0] _0261_;
wire [31:0] _0262_;
wire [31:0] _0263_;
wire [31:0] _0264_;
wire [31:0] _0265_;
wire [31:0] _0266_;
wire [31:0] _0267_;
wire [31:0] _0268_;
wire [31:0] _0269_;
wire [3:0] _0270_;
wire [3:0] _0271_;
wire [3:0] _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire _0276_;
wire _0277_;
wire _0278_;
wire [31:0] _0279_;
wire [31:0] _0280_;
wire [31:0] _0281_;
wire [31:0] _0282_;
wire [31:0] _0283_;
wire [31:0] _0284_;
wire [3:0] _0285_;
wire [3:0] _0286_;
wire [3:0] _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire [1:0] _0294_;
wire [2:0] _0295_;
wire [2:0] _0296_;
wire [4:0] _0297_;
wire [2:0] _0298_;
wire [5:0] _0299_;
wire [5:0] _0300_;
wire [1:0] _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire [3:0] _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire _0324_;
wire _0325_;
wire _0326_;
wire _0327_;
wire _0328_;
wire _0329_;
wire _0330_;
wire _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire _0335_;
wire _0336_;
wire _0337_;
wire _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire _0344_;
wire _0345_;
wire _0346_;
wire _0347_;
wire _0348_;
wire _0349_;
wire _0350_;
wire _0351_;
wire _0352_;
wire _0353_;
wire _0354_;
wire _0355_;
wire _0356_;
wire _0357_;
wire _0358_;
wire [31:0] _0359_;
wire [31:0] _0360_;
wire [31:0] _0361_;
wire [31:0] _0362_;
wire [31:0] _0363_;
wire [31:0] _0364_;
wire [31:0] _0365_;
wire [31:0] _0366_;
wire [31:0] _0367_;
wire [31:0] _0368_;
wire [31:0] _0369_;
wire [31:0] _0370_;
wire [31:0] _0371_;
wire [31:0] _0372_;
wire [31:0] _0373_;
wire [31:0] _0374_;
wire [3:0] _0375_;
wire [3:0] _0376_;
wire [3:0] _0377_;
wire [3:0] _0378_;
wire [3:0] _0379_;
wire [31:0] _0380_;
wire [31:0] _0381_;
wire [31:0] _0382_;
wire [31:0] _0383_;
wire [31:0] _0384_;
wire [31:0] _0385_;
wire [31:0] _0386_;
wire [31:0] _0387_;
wire [31:0] _0388_;
wire [1:0] _0389_;
wire [6:0] _0390_;
wire [3:0] _0391_;
wire [4:0] _0392_;
wire [4:0] _0393_;
wire [11:0] _0394_;
wire [4:0] _0395_;
wire [4:0] _0396_;
wire [4:0] _0397_;
wire [4:0] _0398_;
wire _0399_;
wire _0400_;
wire _0401_;
wire _0402_;
wire _0403_;
wire _0404_;
wire _0405_;
wire _0406_;
wire _0407_;
wire _0408_;
wire _0409_;
wire _0410_;
wire _0411_;
wire _0412_;
wire _0413_;
wire _0414_;
wire _0415_;
wire _0416_;
wire _0417_;
wire _0418_;
wire _0419_;
wire _0420_;
wire _0421_;
wire _0422_;
wire _0423_;
wire _0424_;
wire _0425_;
wire _0426_;
wire _0427_;
wire _0428_;
wire _0429_;
wire _0430_;
wire _0431_;
wire _0432_;
wire _0433_;
wire _0434_;
wire _0435_;
wire _0436_;
wire _0437_;
wire _0438_;
wire _0439_;
wire _0440_;
wire _0441_;
wire _0442_;
wire _0443_;
wire _0444_;
wire _0445_;
wire _0446_;
wire _0447_;
wire _0448_;
wire _0449_;
wire _0450_;
wire _0451_;
wire _0452_;
wire _0453_;
wire _0454_;
wire _0455_;
wire _0456_;
wire _0457_;
wire _0458_;
wire _0459_;
wire _0460_;
wire _0461_;
wire _0462_;
wire _0463_;
wire _0464_;
wire _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire _0469_;
wire _0470_;
wire [1:0] _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire _0477_;
wire [1:0] _0478_;
wire [1:0] _0479_;
wire _0480_;
wire _0481_;
wire [1:0] _0482_;
wire [1:0] _0483_;
wire _0484_;
wire _0485_;
wire _0486_;
wire _0487_;
wire [31:0] _0488_;
wire [31:0] _0489_;
wire [31:0] _0490_;
wire [2:0] _0491_;
wire _0492_;
wire _0493_;
wire _0494_;
wire [2:0] _0495_;
wire [3:0] _0496_;
wire [3:0] _0497_;
wire [3:0] _0498_;
wire [2:0] _0499_;
wire [4:0] _0500_;
wire [5:0] _0501_;
wire [4:0] _0502_;
wire [31:0] _0503_;
wire [31:0] _0504_;
wire [31:0] _0505_;
wire [31:0] _0506_;
wire [31:0] _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire [3:0] _0512_;
wire [3:0] _0513_;
wire [3:0] _0514_;
wire [3:0] _0515_;
wire [3:0] _0516_;
wire [1:0] _0517_;
wire [31:0] _0518_;
wire [31:0] _0519_;
wire [31:0] _0520_;
wire [31:0] _0521_;
wire [31:0] _0522_;
wire [31:0] _0523_;
wire _0524_;
wire _0525_;
wire _0526_;
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire _0534_;
wire _0535_;
wire _0536_;
wire _0537_;
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0542_;
wire _0543_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire _0560_;
wire _0561_;
wire _0562_;
wire _0563_;
wire _0564_;
wire _0565_;
wire _0566_;
wire [31:0] _0567_;
wire [31:0] _0568_;
wire [31:0] _0569_;
wire [31:0] _0570_;
wire [31:0] _0571_;
wire [31:0] _0572_;
wire [31:0] _0573_;
wire [31:0] _0574_;
wire [31:0] _0575_;
wire [31:0] _0576_;
wire [31:0] _0577_;
wire [31:0] _0578_;
wire [3:0] _0579_;
wire [3:0] _0580_;
wire [3:0] _0581_;
wire [3:0] _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire [31:0] _0591_;
wire [31:0] _0592_;
wire [31:0] _0593_;
wire [31:0] _0594_;
wire [31:0] _0595_;
wire [31:0] _0596_;
wire [31:0] _0597_;
wire [31:0] _0598_;
wire [3:0] _0599_;
wire [3:0] _0600_;
wire [3:0] _0601_;
wire [3:0] _0602_;
wire _0603_;
wire _0604_;
wire _0605_;
wire _0606_;
wire _0607_;
wire _0608_;
wire _0609_;
wire _0610_;
wire [2:0] _0611_;
wire _0612_;
wire _0613_;
wire _0614_;
wire _0615_;
wire _0616_;
wire _0617_;
wire _0618_;
wire _0619_;
wire _0620_;
wire _0621_;
wire _0622_;
wire _0623_;
wire _0624_;
wire _0625_;
wire _0626_;
wire _0627_;
wire _0628_;
wire _0629_;
wire _0630_;
wire _0631_;
wire _0632_;
wire _0633_;
wire _0634_;
wire _0635_;
wire _0636_;
wire _0637_;
wire _0638_;
wire _0639_;
wire _0640_;
wire _0641_;
wire _0642_;
wire _0643_;
wire _0644_;
wire _0645_;
wire _0646_;
wire _0647_;
wire _0648_;
wire _0649_;
wire _0650_;
wire _0651_;
wire [31:0] _0652_;
wire [31:0] _0653_;
wire [31:0] _0654_;
wire [31:0] _0655_;
wire [31:0] _0656_;
wire [31:0] _0657_;
wire [31:0] _0658_;
wire [31:0] _0659_;
wire [31:0] _0660_;
wire [31:0] _0661_;
wire [31:0] _0662_;
wire [31:0] _0663_;
wire [31:0] _0664_;
wire [31:0] _0665_;
wire [3:0] _0666_;
wire [3:0] _0667_;
wire [3:0] _0668_;
wire [3:0] _0669_;
wire [31:0] _0670_;
wire [31:0] _0671_;
wire [31:0] _0672_;
wire [31:0] _0673_;
wire [31:0] _0674_;
wire [31:0] _0675_;
wire [31:0] _0676_;
wire [31:0] _0677_;
wire [31:0] _0678_;
wire [4:0] _0679_;
wire [4:0] _0680_;
wire _0681_;
wire _0682_;
wire _0683_;
wire _0684_;
wire _0685_;
wire _0686_;
wire _0687_;
wire _0688_;
wire _0689_;
wire _0690_;
wire _0691_;
wire _0692_;
wire _0693_;
wire _0694_;
wire _0695_;
wire _0696_;
wire _0697_;
wire _0698_;
wire _0699_;
wire _0700_;
wire _0701_;
wire _0702_;
wire _0703_;
wire _0704_;
wire _0705_;
wire _0706_;
wire _0707_;
wire [1:0] _0708_;
wire _0709_;
wire [1:0] _0710_;
wire _0711_;
wire _0712_;
wire [31:0] _0713_;
wire [31:0] _0714_;
wire [31:0] _0715_;
wire _0716_;
wire [3:0] _0717_;
wire [3:0] _0718_;
wire [3:0] _0719_;
wire [31:0] _0720_;
wire [31:0] _0721_;
wire [31:0] _0722_;
wire [31:0] _0723_;
wire _0724_;
wire [3:0] _0725_;
wire [3:0] _0726_;
wire [3:0] _0727_;
wire [3:0] _0728_;
wire [31:0] _0729_;
wire [31:0] _0730_;
wire [31:0] _0731_;
wire [31:0] _0732_;
wire [31:0] _0733_;
wire [31:0] _0734_;
wire _0735_;
/* cellift = 32'd1 */
wire _0736_;
wire _0737_;
/* cellift = 32'd1 */
wire _0738_;
wire _0739_;
/* cellift = 32'd1 */
wire _0740_;
wire _0741_;
/* cellift = 32'd1 */
wire _0742_;
wire _0743_;
/* cellift = 32'd1 */
wire _0744_;
wire _0745_;
wire _0746_;
wire _0747_;
wire _0748_;
wire _0749_;
wire _0750_;
wire _0751_;
wire _0752_;
wire _0753_;
wire _0754_;
wire [31:0] _0755_;
wire [31:0] _0756_;
wire [31:0] _0757_;
wire [3:0] _0758_;
wire _0759_;
wire _0760_;
wire [31:0] _0761_;
wire [31:0] _0762_;
wire [3:0] _0763_;
wire _0764_;
wire _0765_;
wire _0766_;
wire _0767_;
wire _0768_;
wire _0769_;
wire _0770_;
wire _0771_;
wire _0772_;
wire _0773_;
wire _0774_;
wire _0775_;
wire _0776_;
wire [31:0] _0777_;
wire [31:0] _0778_;
wire [31:0] _0779_;
wire [31:0] _0780_;
wire [3:0] _0781_;
wire [31:0] _0782_;
wire [31:0] _0783_;
wire [31:0] _0784_;
wire [31:0] _0785_;
wire [3:0] _0786_;
wire [3:0] _0787_;
wire [31:0] _0788_;
wire [31:0] _0789_;
wire _0790_;
wire _0791_;
wire _0792_;
wire _0793_;
wire _0794_;
wire _0795_;
wire _0796_;
wire _0797_;
wire _0798_;
wire _0799_;
wire _0800_;
wire _0801_;
wire _0802_;
wire _0803_;
wire _0804_;
wire _0805_;
wire _0806_;
wire _0807_;
wire _0808_;
wire _0809_;
wire _0810_;
wire _0811_;
wire _0812_;
wire _0813_;
wire _0814_;
wire _0815_;
wire _0816_;
wire _0817_;
wire _0818_;
/* cellift = 32'd1 */
wire _0819_;
wire _0820_;
/* cellift = 32'd1 */
wire _0821_;
wire _0822_;
/* cellift = 32'd1 */
wire _0823_;
wire _0824_;
/* cellift = 32'd1 */
wire _0825_;
wire _0826_;
/* cellift = 32'd1 */
wire _0827_;
wire _0828_;
/* cellift = 32'd1 */
wire _0829_;
wire _0830_;
/* cellift = 32'd1 */
wire _0831_;
wire _0832_;
/* cellift = 32'd1 */
wire _0833_;
wire _0834_;
wire _0835_;
/* cellift = 32'd1 */
wire _0836_;
wire _0837_;
/* cellift = 32'd1 */
wire _0838_;
wire [31:0] _0839_;
/* cellift = 32'd1 */
wire [31:0] _0840_;
wire [31:0] _0841_;
/* cellift = 32'd1 */
wire [31:0] _0842_;
wire [31:0] _0843_;
/* cellift = 32'd1 */
wire [31:0] _0844_;
wire [31:0] _0845_;
/* cellift = 32'd1 */
wire [31:0] _0846_;
wire [3:0] _0847_;
/* cellift = 32'd1 */
wire [3:0] _0848_;
wire [31:0] _0849_;
/* cellift = 32'd1 */
wire [31:0] _0850_;
wire [31:0] _0851_;
/* cellift = 32'd1 */
wire [31:0] _0852_;
wire [3:0] _0853_;
/* src = "generated/sv2v_out.v:1038.7-1038.37" */
wire _0854_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1038.7-1038.37" */
wire _0855_;
/* src = "generated/sv2v_out.v:1039.8-1039.38" */
wire _0856_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1039.8-1039.38" */
wire _0857_;
/* src = "generated/sv2v_out.v:1041.13-1041.43" */
wire _0858_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1041.13-1041.43" */
wire _0859_;
/* src = "generated/sv2v_out.v:1067.19-1067.35" */
wire _0860_;
/* src = "generated/sv2v_out.v:1091.10-1091.26" */
wire _0861_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1091.10-1091.26" */
wire _0862_;
/* src = "generated/sv2v_out.v:1091.32-1091.48" */
wire _0863_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1091.32-1091.48" */
wire _0864_;
/* src = "generated/sv2v_out.v:1100.11-1100.25" */
wire _0865_;
/* src = "generated/sv2v_out.v:1105.16-1105.31" */
wire _0866_;
/* src = "generated/sv2v_out.v:1147.13-1147.39" */
wire _0867_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1147.13-1147.39" */
wire _0868_;
/* src = "generated/sv2v_out.v:1147.45-1147.63" */
wire _0869_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1147.45-1147.63" */
wire _0870_;
/* src = "generated/sv2v_out.v:1147.70-1147.87" */
wire _0871_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1147.70-1147.87" */
wire _0872_;
/* src = "generated/sv2v_out.v:1150.13-1150.42" */
wire _0873_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1150.13-1150.42" */
wire _0874_;
/* src = "generated/sv2v_out.v:1163.17-1163.37" */
wire _0875_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1163.17-1163.37" */
wire _0876_;
/* src = "generated/sv2v_out.v:1167.17-1167.37" */
wire _0877_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1167.17-1167.37" */
wire _0878_;
/* src = "generated/sv2v_out.v:1171.17-1171.37" */
wire _0879_;
/* src = "generated/sv2v_out.v:1232.25-1232.53" */
wire _0880_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1232.25-1232.53" */
wire _0881_;
/* src = "generated/sv2v_out.v:1232.59-1232.89" */
wire _0882_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1232.59-1232.89" */
wire _0883_;
/* src = "generated/sv2v_out.v:1232.96-1232.126" */
wire _0884_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1232.96-1232.126" */
wire _0885_;
/* src = "generated/sv2v_out.v:1232.133-1232.160" */
wire _0886_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1232.133-1232.160" */
wire _0887_;
/* src = "generated/sv2v_out.v:1232.167-1232.194" */
wire _0888_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1232.167-1232.194" */
wire _0889_;
/* src = "generated/sv2v_out.v:1232.201-1232.229" */
wire _0890_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1232.201-1232.229" */
wire _0891_;
/* src = "generated/sv2v_out.v:1232.236-1232.265" */
wire _0892_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1232.236-1232.265" */
wire _0893_;
/* src = "generated/sv2v_out.v:1232.272-1232.301" */
wire _0894_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1232.272-1232.301" */
wire _0895_;
/* src = "generated/sv2v_out.v:1240.18-1240.47" */
wire _0896_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1240.18-1240.47" */
wire _0897_;
/* src = "generated/sv2v_out.v:1244.18-1244.46" */
wire _0898_;
/* src = "generated/sv2v_out.v:996.35-996.51" */
wire _0899_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:996.35-996.51" */
wire _0900_;
/* src = "generated/sv2v_out.v:997.35-997.51" */
wire _0901_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:997.35-997.51" */
wire _0902_;
/* src = "generated/sv2v_out.v:1147.12-1147.64" */
wire _0903_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1147.12-1147.64" */
wire _0904_;
/* src = "generated/sv2v_out.v:1147.11-1147.88" */
wire _0905_;
/* src = "generated/sv2v_out.v:1150.12-1150.67" */
wire _0906_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1150.12-1150.67" */
wire _0907_;
/* src = "generated/sv2v_out.v:1150.11-1150.91" */
wire _0908_;
/* src = "generated/sv2v_out.v:1158.11-1158.54" */
wire _0909_;
/* src = "generated/sv2v_out.v:1228.12-1228.34" */
wire _0910_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1228.12-1228.34" */
wire _0911_;
/* src = "generated/sv2v_out.v:1239.18-1239.57" */
wire _0912_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1239.18-1239.57" */
wire _0913_;
/* src = "generated/sv2v_out.v:1244.17-1244.55" */
wire _0914_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1244.17-1244.55" */
wire _0915_;
/* src = "generated/sv2v_out.v:1250.12-1250.36" */
wire _0916_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1250.12-1250.36" */
wire _0917_;
/* src = "generated/sv2v_out.v:1091.9-1091.49" */
wire _0918_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1091.9-1091.49" */
wire _0919_;
/* src = "generated/sv2v_out.v:1232.24-1232.90" */
wire _0920_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1232.24-1232.90" */
wire _0921_;
/* src = "generated/sv2v_out.v:1232.23-1232.127" */
wire _0922_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1232.23-1232.127" */
wire _0923_;
/* src = "generated/sv2v_out.v:1232.22-1232.161" */
wire _0924_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1232.22-1232.161" */
wire _0925_;
/* src = "generated/sv2v_out.v:1232.21-1232.195" */
wire _0926_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1232.21-1232.195" */
wire _0927_;
/* src = "generated/sv2v_out.v:1232.20-1232.230" */
wire _0928_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1232.20-1232.230" */
wire _0929_;
/* src = "generated/sv2v_out.v:1232.19-1232.266" */
wire _0930_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1232.19-1232.266" */
wire _0931_;
/* src = "generated/sv2v_out.v:1232.18-1232.302" */
wire _0932_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1232.18-1232.302" */
wire _0933_;
/* src = "generated/sv2v_out.v:1238.19-1238.84" */
wire _0934_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1238.19-1238.84" */
wire _0935_;
/* src = "generated/sv2v_out.v:1238.18-1238.98" */
wire _0936_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1238.18-1238.98" */
wire _0937_;
/* src = "generated/sv2v_out.v:995.48-995.150" */
wire _0938_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:995.48-995.150" */
wire _0939_;
/* src = "generated/sv2v_out.v:995.47-995.186" */
wire _0940_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:995.47-995.186" */
wire _0941_;
/* src = "generated/sv2v_out.v:995.46-995.223" */
wire _0942_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:995.46-995.223" */
wire _0943_;
/* src = "generated/sv2v_out.v:995.45-995.257" */
wire _0944_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:995.45-995.257" */
wire _0945_;
/* src = "generated/sv2v_out.v:995.22-995.39" */
wire _0946_;
/* src = "generated/sv2v_out.v:1189.42-1189.54" */
wire _0947_;
/* src = "generated/sv2v_out.v:1244.51-1244.55" */
wire _0948_;
/* src = "generated/sv2v_out.v:1252.22-1252.33" */
wire _0949_;
/* src = "generated/sv2v_out.v:1252.50-1252.56" */
wire _0950_;
/* src = "generated/sv2v_out.v:1252.22-1252.46" */
wire _0951_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1252.22-1252.46" */
wire _0952_;
wire _0953_;
wire _0954_;
/* cellift = 32'd1 */
wire _0955_;
wire [2:0] _0956_;
/* cellift = 32'd1 */
wire [2:0] _0957_;
wire [2:0] _0958_;
/* cellift = 32'd1 */
wire [2:0] _0959_;
wire _0960_;
/* cellift = 32'd1 */
wire _0961_;
wire _0962_;
/* cellift = 32'd1 */
wire _0963_;
wire _0964_;
wire _0965_;
wire _0966_;
wire _0967_;
/* cellift = 32'd1 */
wire _0968_;
wire _0969_;
/* cellift = 32'd1 */
wire _0970_;
wire _0971_;
/* cellift = 32'd1 */
wire _0972_;
/* src = "generated/sv2v_out.v:1040.12-1040.29" */
wire [3:0] _0973_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1040.12-1040.29" */
wire [3:0] _0974_;
/* src = "generated/sv2v_out.v:1042.13-1042.39" */
wire [3:0] _0975_;
/* src = "generated/sv2v_out.v:964.14-964.18" */
wire [31:0] addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:964.14-964.18" */
wire [31:0] addr_t0;
/* src = "generated/sv2v_out.v:955.12-955.17" */
wire [3:0] aluop;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:955.12-955.17" */
wire [3:0] aluop_t0;
/* src = "generated/sv2v_out.v:965.13-965.17" */
wire [31:0] base;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:965.13-965.17" */
wire [31:0] base_t0;
/* src = "generated/sv2v_out.v:957.7-957.13" */
wire branch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:957.7-957.13" */
wire branch_t0;
/* src = "generated/sv2v_out.v:925.13-925.16" */
input clk;
wire clk;
/* cellift = 32'd1 */
input clk_t0;
wire clk_t0;
/* src = "generated/sv2v_out.v:958.6-958.9" */
wire csr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:958.6-958.9" */
wire csr_t0;
/* src = "generated/sv2v_out.v:936.21-936.27" */
output [180:0] decode;
reg [180:0] decode;
/* src = "generated/sv2v_out.v:938.13-938.23" */
input decode_rdy;
wire decode_rdy;
/* cellift = 32'd1 */
input decode_rdy_t0;
wire decode_rdy_t0;
/* cellift = 32'd1 */
output [180:0] decode_t0;
reg [180:0] decode_t0;
/* src = "generated/sv2v_out.v:937.13-937.23" */
output decode_vld;
reg decode_vld;
/* cellift = 32'd1 */
output decode_vld_t0;
reg decode_vld_t0;
/* src = "generated/sv2v_out.v:928.20-928.25" */
input [63:0] fetch;
wire [63:0] fetch;
/* src = "generated/sv2v_out.v:935.14-935.23" */
output fetch_rdy;
wire fetch_rdy;
/* cellift = 32'd1 */
output fetch_rdy_t0;
wire fetch_rdy_t0;
/* cellift = 32'd1 */
input [63:0] fetch_t0;
wire [63:0] fetch_t0;
/* src = "generated/sv2v_out.v:934.13-934.22" */
input fetch_vld;
wire fetch_vld;
/* cellift = 32'd1 */
input fetch_vld_t0;
wire fetch_vld_t0;
/* src = "generated/sv2v_out.v:927.13-927.18" */
input flush;
wire flush;
/* cellift = 32'd1 */
input flush_t0;
wire flush_t0;
/* src = "generated/sv2v_out.v:961.7-961.14" */
wire illegal;
/* src = "generated/sv2v_out.v:963.7-963.21" */
wire illegal_opcode;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:963.7-963.21" */
wire illegal_opcode_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:961.7-961.14" */
wire illegal_t0;
/* src = "generated/sv2v_out.v:929.20-929.29" */
input [31:0] immediate;
wire [31:0] immediate;
/* cellift = 32'd1 */
input [31:0] immediate_t0;
wire [31:0] immediate_t0;
/* src = "generated/sv2v_out.v:962.6-962.17" */
wire instr_valid;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:962.6-962.17" */
wire instr_valid_t0;
/* src = "generated/sv2v_out.v:960.6-960.15" */
wire is_fencei;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:960.6-960.15" */
wire is_fencei_t0;
/* src = "generated/sv2v_out.v:967.7-967.21" */
wire misaligned_jmp;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:967.7-967.21" */
wire misaligned_jmp_t0;
/* src = "generated/sv2v_out.v:968.7-968.22" */
wire misaligned_ldst;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:968.7-968.22" */
wire misaligned_ldst_t0;
/* src = "generated/sv2v_out.v:966.13-966.19" */
wire [31:0] offset;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:966.13-966.19" */
wire [31:0] offset_t0;
/* src = "generated/sv2v_out.v:953.13-953.16" */
wire [31:0] op1;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:953.13-953.16" */
wire [31:0] op1_t0;
/* src = "generated/sv2v_out.v:954.13-954.16" */
wire [31:0] op2;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:954.13-954.16" */
wire [31:0] op2_t0;
/* src = "generated/sv2v_out.v:930.20-930.29" */
input [31:0] regrd_rs1;
wire [31:0] regrd_rs1;
/* src = "generated/sv2v_out.v:932.13-932.25" */
input regrd_rs1_en;
wire regrd_rs1_en;
/* cellift = 32'd1 */
input regrd_rs1_en_t0;
wire regrd_rs1_en_t0;
/* cellift = 32'd1 */
input [31:0] regrd_rs1_t0;
wire [31:0] regrd_rs1_t0;
/* src = "generated/sv2v_out.v:931.20-931.29" */
input [31:0] regrd_rs2;
wire [31:0] regrd_rs2;
/* src = "generated/sv2v_out.v:933.13-933.25" */
input regrd_rs2_en;
wire regrd_rs2_en;
/* cellift = 32'd1 */
input regrd_rs2_en_t0;
wire regrd_rs2_en_t0;
/* cellift = 32'd1 */
input [31:0] regrd_rs2_t0;
wire [31:0] regrd_rs2_t0;
/* src = "generated/sv2v_out.v:956.7-956.16" */
wire regwr_alu;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:956.7-956.16" */
wire regwr_alu_t0;
/* src = "generated/sv2v_out.v:939.20-939.30" */
input [31:0] regwr_data;
wire [31:0] regwr_data;
/* cellift = 32'd1 */
input [31:0] regwr_data_t0;
wire [31:0] regwr_data_t0;
/* src = "generated/sv2v_out.v:941.13-941.21" */
input regwr_en;
wire regwr_en;
/* cellift = 32'd1 */
input regwr_en_t0;
wire regwr_en_t0;
/* src = "generated/sv2v_out.v:942.13-942.26" */
input regwr_pending;
wire regwr_pending;
/* cellift = 32'd1 */
input regwr_pending_t0;
wire regwr_pending_t0;
/* src = "generated/sv2v_out.v:940.19-940.28" */
input [4:0] regwr_sel;
wire [4:0] regwr_sel;
/* cellift = 32'd1 */
input [4:0] regwr_sel_t0;
wire [4:0] regwr_sel_t0;
/* src = "generated/sv2v_out.v:975.14-975.22" */
wire [31:0] rs1_data;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:975.14-975.22" */
wire [31:0] rs1_data_t0;
/* src = "generated/sv2v_out.v:973.7-973.18" */
wire rs1_forward;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:973.7-973.18" */
wire rs1_forward_t0;
/* src = "generated/sv2v_out.v:976.14-976.22" */
wire [31:0] rs2_data;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:976.14-976.22" */
wire [31:0] rs2_data_t0;
/* src = "generated/sv2v_out.v:974.7-974.18" */
wire rs2_forward;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:974.7-974.18" */
wire rs2_forward_t0;
/* src = "generated/sv2v_out.v:926.13-926.17" */
input rstz;
wire rstz;
/* src = "generated/sv2v_out.v:977.7-977.12" */
wire stall;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:977.7-977.12" */
wire stall_t0;
/* src = "generated/sv2v_out.v:972.13-972.23" */
wire [31:0] store_data;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:972.13-972.23" */
wire [31:0] store_data_t0;
assign fetch_rdy = _0951_ & /* src = "generated/sv2v_out.v:1252.21-1252.56" */ _0950_;
assign rs1_forward = regwr_en & /* src = "generated/sv2v_out.v:996.23-996.52" */ _0899_;
assign rs2_forward = regwr_en & /* src = "generated/sv2v_out.v:997.23-997.52" */ _0901_;
assign _0222_ = _0952_ & _0950_;
assign _0225_ = regwr_en_t0 & _0899_;
assign _0228_ = regwr_en_t0 & _0901_;
assign _0223_ = stall_t0 & _0951_;
assign _0226_ = _0900_ & regwr_en;
assign _0229_ = _0902_ & regwr_en;
assign _0224_ = _0952_ & stall_t0;
assign _0227_ = regwr_en_t0 & _0900_;
assign _0230_ = regwr_en_t0 & _0902_;
assign _0524_ = _0222_ | _0223_;
assign _0525_ = _0225_ | _0226_;
assign _0526_ = _0228_ | _0229_;
assign fetch_rdy_t0 = _0524_ | _0224_;
assign rs1_forward_t0 = _0525_ | _0227_;
assign rs2_forward_t0 = _0526_ | _0230_;
assign _0746_ = misaligned_jmp ^ decode[1];
assign _0747_ = misaligned_ldst ^ decode[0];
assign _0748_ = illegal ^ decode[2];
assign _0749_ = _0914_ ^ decode[5];
assign _0750_ = csr ^ decode[6];
assign _0751_ = _0854_ ^ decode[11];
assign _0752_ = _0896_ ^ decode[12];
assign _0753_ = _0912_ ^ decode[13];
assign _0754_ = _0936_ ^ decode[14];
assign _0755_ = addr ^ decode[52:21];
assign _0756_ = op1 ^ decode[116:85];
assign _0757_ = op2 ^ decode[84:53];
assign _0758_ = aluop ^ decode[19:16];
assign _0759_ = _0932_ ^ decode[20];
assign _0760_ = regwr_alu ^ decode[15];
assign _0761_ = fetch[31:0] ^ decode[148:117];
assign _0762_ = fetch[63:32] ^ decode[180:149];
assign _0531_ = misaligned_jmp_t0 | decode_t0[1];
assign _0535_ = misaligned_ldst_t0 | decode_t0[0];
assign _0539_ = illegal_t0 | decode_t0[2];
assign _0543_ = _0915_ | decode_t0[5];
assign _0547_ = csr_t0 | decode_t0[6];
assign _0551_ = _0855_ | decode_t0[11];
assign _0555_ = _0897_ | decode_t0[12];
assign _0559_ = _0913_ | decode_t0[13];
assign _0563_ = _0937_ | decode_t0[14];
assign _0567_ = addr_t0 | decode_t0[52:21];
assign _0571_ = op1_t0 | decode_t0[116:85];
assign _0575_ = op2_t0 | decode_t0[84:53];
assign _0579_ = aluop_t0 | decode_t0[19:16];
assign _0583_ = _0933_ | decode_t0[20];
assign _0587_ = regwr_alu_t0 | decode_t0[15];
assign _0591_ = fetch_t0[31:0] | decode_t0[148:117];
assign _0595_ = fetch_t0[63:32] | decode_t0[180:149];
assign _0532_ = _0746_ | _0531_;
assign _0536_ = _0747_ | _0535_;
assign _0540_ = _0748_ | _0539_;
assign _0544_ = _0749_ | _0543_;
assign _0548_ = _0750_ | _0547_;
assign _0552_ = _0751_ | _0551_;
assign _0556_ = _0752_ | _0555_;
assign _0560_ = _0753_ | _0559_;
assign _0564_ = _0754_ | _0563_;
assign _0568_ = _0755_ | _0567_;
assign _0572_ = _0756_ | _0571_;
assign _0576_ = _0757_ | _0575_;
assign _0580_ = _0758_ | _0579_;
assign _0584_ = _0759_ | _0583_;
assign _0588_ = _0760_ | _0587_;
assign _0592_ = _0761_ | _0591_;
assign _0596_ = _0762_ | _0595_;
assign _0234_ = _0053_ & misaligned_jmp_t0;
assign _0237_ = _0053_ & misaligned_ldst_t0;
assign _0240_ = _0053_ & illegal_t0;
assign _0243_ = _0053_ & _0915_;
assign _0246_ = _0053_ & csr_t0;
assign _0249_ = _0053_ & _0855_;
assign _0252_ = _0053_ & _0897_;
assign _0255_ = _0053_ & _0913_;
assign _0258_ = _0053_ & _0937_;
assign _0261_ = { _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_ } & addr_t0;
assign _0264_ = { _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_ } & op1_t0;
assign _0267_ = { _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_ } & op2_t0;
assign _0270_ = { _0053_, _0053_, _0053_, _0053_ } & aluop_t0;
assign _0273_ = _0053_ & _0933_;
assign _0276_ = _0053_ & regwr_alu_t0;
assign _0279_ = { _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_ } & fetch_t0[31:0];
assign _0282_ = { _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_, _0053_ } & fetch_t0[63:32];
assign _0235_ = _0072_ & decode_t0[1];
assign _0238_ = _0072_ & decode_t0[0];
assign _0241_ = _0072_ & decode_t0[2];
assign _0244_ = _0072_ & decode_t0[5];
assign _0247_ = _0072_ & decode_t0[6];
assign _0250_ = _0072_ & decode_t0[11];
assign _0253_ = _0072_ & decode_t0[12];
assign _0256_ = _0072_ & decode_t0[13];
assign _0259_ = _0072_ & decode_t0[14];
assign _0262_ = { _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_ } & decode_t0[52:21];
assign _0265_ = { _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_ } & decode_t0[116:85];
assign _0268_ = { _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_ } & decode_t0[84:53];
assign _0271_ = { _0072_, _0072_, _0072_, _0072_ } & decode_t0[19:16];
assign _0274_ = _0072_ & decode_t0[20];
assign _0277_ = _0072_ & decode_t0[15];
assign _0280_ = { _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_ } & decode_t0[148:117];
assign _0283_ = { _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_ } & decode_t0[180:149];
assign _0236_ = _0532_ & _0054_;
assign _0239_ = _0536_ & _0054_;
assign _0242_ = _0540_ & _0054_;
assign _0245_ = _0544_ & _0054_;
assign _0248_ = _0548_ & _0054_;
assign _0251_ = _0552_ & _0054_;
assign _0254_ = _0556_ & _0054_;
assign _0257_ = _0560_ & _0054_;
assign _0260_ = _0564_ & _0054_;
assign _0263_ = _0568_ & { _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_ };
assign _0266_ = _0572_ & { _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_ };
assign _0269_ = _0576_ & { _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_ };
assign _0272_ = _0580_ & { _0054_, _0054_, _0054_, _0054_ };
assign _0275_ = _0584_ & _0054_;
assign _0278_ = _0588_ & _0054_;
assign _0281_ = _0592_ & { _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_ };
assign _0284_ = _0596_ & { _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_ };
assign _0533_ = _0234_ | _0235_;
assign _0537_ = _0237_ | _0238_;
assign _0541_ = _0240_ | _0241_;
assign _0545_ = _0243_ | _0244_;
assign _0549_ = _0246_ | _0247_;
assign _0553_ = _0249_ | _0250_;
assign _0557_ = _0252_ | _0253_;
assign _0561_ = _0255_ | _0256_;
assign _0565_ = _0258_ | _0259_;
assign _0569_ = _0261_ | _0262_;
assign _0573_ = _0264_ | _0265_;
assign _0577_ = _0267_ | _0268_;
assign _0581_ = _0270_ | _0271_;
assign _0585_ = _0273_ | _0274_;
assign _0589_ = _0276_ | _0277_;
assign _0593_ = _0279_ | _0280_;
assign _0597_ = _0282_ | _0283_;
assign _0534_ = _0533_ | _0236_;
assign _0538_ = _0537_ | _0239_;
assign _0542_ = _0541_ | _0242_;
assign _0546_ = _0545_ | _0245_;
assign _0550_ = _0549_ | _0248_;
assign _0554_ = _0553_ | _0251_;
assign _0558_ = _0557_ | _0254_;
assign _0562_ = _0561_ | _0257_;
assign _0566_ = _0565_ | _0260_;
assign _0570_ = _0569_ | _0263_;
assign _0574_ = _0573_ | _0266_;
assign _0578_ = _0577_ | _0269_;
assign _0582_ = _0581_ | _0272_;
assign _0586_ = _0585_ | _0275_;
assign _0590_ = _0589_ | _0278_;
assign _0594_ = _0593_ | _0281_;
assign _0598_ = _0597_ | _0284_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[1] */
always_ff @(posedge clk)
decode_t0[1] <= _0534_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[0] */
always_ff @(posedge clk)
decode_t0[0] <= _0538_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[2] */
always_ff @(posedge clk)
decode_t0[2] <= _0542_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[5] */
always_ff @(posedge clk)
decode_t0[5] <= _0546_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[6] */
always_ff @(posedge clk)
decode_t0[6] <= _0550_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[11] */
always_ff @(posedge clk)
decode_t0[11] <= _0554_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[12] */
always_ff @(posedge clk)
decode_t0[12] <= _0558_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[13] */
always_ff @(posedge clk)
decode_t0[13] <= _0562_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[14] */
always_ff @(posedge clk)
decode_t0[14] <= _0566_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[52:21] */
always_ff @(posedge clk)
decode_t0[52:21] <= _0570_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[116:85] */
always_ff @(posedge clk)
decode_t0[116:85] <= _0574_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[84:53] */
always_ff @(posedge clk)
decode_t0[84:53] <= _0578_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[19:16] */
always_ff @(posedge clk)
decode_t0[19:16] <= _0582_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[20] */
always_ff @(posedge clk)
decode_t0[20] <= _0586_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[15] */
always_ff @(posedge clk)
decode_t0[15] <= _0590_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[148:117] */
always_ff @(posedge clk)
decode_t0[148:117] <= _0594_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[180:149] */
always_ff @(posedge clk)
decode_t0[180:149] <= _0598_;
assign _0183_ = | fetch_t0[13:12];
assign _0188_ = | fetch_t0[31:20];
assign _0189_ = | { fetch_t0[19:15], regwr_sel_t0 };
assign _0190_ = | { fetch_t0[24:20], regwr_sel_t0 };
assign _0191_ = | fetch_t0[1:0];
assign _0197_ = | fetch_t0[6:2];
assign _0198_ = | addr_t0[1:0];
assign _0679_ = regwr_sel_t0 | fetch_t0[19:15];
assign _0680_ = regwr_sel_t0 | fetch_t0[24:20];
assign _0110_ = ~ fetch_t0[13:12];
assign _0115_ = ~ fetch_t0[31:20];
assign _0116_ = ~ _0679_;
assign _0117_ = ~ _0680_;
assign _0132_ = ~ fetch_t0[1:0];
assign _0144_ = ~ fetch_t0[14:12];
assign _0149_ = ~ fetch_t0[6:2];
assign _0152_ = ~ addr_t0[1:0];
assign _0389_ = fetch[13:12] & _0110_;
assign _0394_ = fetch[31:20] & _0115_;
assign _0395_ = regwr_sel & _0116_;
assign _0397_ = regwr_sel & _0117_;
assign _0471_ = fetch[1:0] & _0132_;
assign _0495_ = fetch[14:12] & _0144_;
assign _0502_ = fetch[6:2] & _0149_;
assign _0517_ = addr[1:0] & _0152_;
assign _0396_ = fetch[19:15] & _0116_;
assign _0398_ = fetch[24:20] & _0117_;
assign _0790_ = _0389_ == { 1'h0, _0110_[0] };
assign _0791_ = _0390_ == { 1'h0, _0111_[5], 5'h00 };
assign _0792_ = _0394_ == { 11'h000, _0115_[0] };
assign _0793_ = _0394_ == { 2'h0, _0115_[9:8], 6'h00, _0115_[1], 1'h0 };
assign _0794_ = _0394_ == { 3'h0, _0115_[8], 5'h00, _0115_[2], 1'h0, _0115_[0] };
assign _0795_ = _0395_ == _0396_;
assign _0796_ = _0397_ == _0398_;
assign _0797_ = _0471_ == _0132_;
assign _0798_ = _0495_ == { 1'h0, _0144_[1:0] };
assign _0799_ = _0495_ == { 1'h0, _0144_[1], 1'h0 };
assign _0800_ = _0495_ == { 2'h0, _0144_[0] };
assign _0801_ = _0495_ == { _0144_[2], 2'h0 };
assign _0802_ = _0495_ == { _0144_[2], 1'h0, _0144_[0] };
assign _0803_ = _0495_ == { _0144_[2:1], 1'h0 };
assign _0804_ = _0495_ == _0144_;
assign _0805_ = _0502_ == { 2'h0, _0149_[2], 1'h0, _0149_[0] };
assign _0806_ = _0502_ == { 1'h0, _0149_[3:2], 1'h0, _0149_[0] };
assign _0807_ = _0502_ == { _0149_[4:3], 3'h0 };
assign _0808_ = _0502_ == { _0149_[4:3], 1'h0, _0149_[1:0] };
assign _0809_ = _0502_ == { 1'h0, _0149_[3], 3'h0 };
assign _0810_ = _0502_ == { _0149_[4:3], 2'h0, _0149_[0] };
assign _0811_ = _0502_ == { 3'h0, _0149_[1:0] };
assign _0812_ = _0502_ == { _0149_[4:2], 2'h0 };
assign _0813_ = _0502_ == { 1'h0, _0149_[3:2], 2'h0 };
assign _0814_ = _0502_ == { 2'h0, _0149_[2], 2'h0 };
assign _0815_ = _0517_ == _0152_;
assign _0816_ = _0517_ == { _0152_[1], 1'h0 };
assign _0817_ = _0517_ == { 1'h0, _0152_[0] };
assign _0859_ = _0790_ & _0183_;
assign _0003_ = _0791_ & _0184_;
assign _0876_ = _0792_ & _0188_;
assign _0878_ = _0793_ & _0188_;
assign _0023_ = _0794_ & _0188_;
assign _0900_ = _0795_ & _0189_;
assign _0902_ = _0796_ & _0190_;
assign illegal_opcode_t0 = _0797_ & _0191_;
assign _0959_[2] = _0798_ & _0193_;
assign _0959_[1] = _0799_ & _0193_;
assign _0862_ = _0800_ & _0193_;
assign _0963_ = _0801_ & _0193_;
assign _0864_ = _0802_ & _0193_;
assign _0957_[1] = _0803_ & _0193_;
assign _0957_[2] = _0804_ & _0193_;
assign _0883_ = _0805_ & _0197_;
assign _0881_ = _0806_ & _0197_;
assign _0889_ = _0807_ & _0197_;
assign _0891_ = _0808_ & _0197_;
assign _0855_ = _0809_ & _0197_;
assign _0893_ = _0810_ & _0197_;
assign _0895_ = _0811_ & _0197_;
assign _0171_ = _0812_ & _0197_;
assign _0887_ = _0813_ & _0197_;
assign _0885_ = _0814_ & _0197_;
assign _0968_ = _0815_ & _0198_;
assign _0970_ = _0816_ & _0198_;
assign _0972_ = _0817_ & _0198_;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_vld */
always_ff @(posedge clk)
if (_0055_) decode_vld <= 1'h0;
else if (_0051_) decode_vld <= _0954_;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[1] */
always_ff @(posedge clk)
if (_0053_) decode[1] <= misaligned_jmp;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[0] */
always_ff @(posedge clk)
if (_0053_) decode[0] <= misaligned_ldst;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[2] */
always_ff @(posedge clk)
if (_0053_) decode[2] <= illegal;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[5] */
always_ff @(posedge clk)
if (_0053_) decode[5] <= _0914_;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[6] */
always_ff @(posedge clk)
if (_0053_) decode[6] <= csr;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[11] */
always_ff @(posedge clk)
if (_0053_) decode[11] <= _0854_;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[12] */
always_ff @(posedge clk)
if (_0053_) decode[12] <= _0896_;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[13] */
always_ff @(posedge clk)
if (_0053_) decode[13] <= _0912_;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[14] */
always_ff @(posedge clk)
if (_0053_) decode[14] <= _0936_;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[52:21] */
always_ff @(posedge clk)
if (_0053_) decode[52:21] <= addr;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[116:85] */
always_ff @(posedge clk)
if (_0053_) decode[116:85] <= op1;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[84:53] */
always_ff @(posedge clk)
if (_0053_) decode[84:53] <= op2;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[19:16] */
always_ff @(posedge clk)
if (_0053_) decode[19:16] <= aluop;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[20] */
always_ff @(posedge clk)
if (_0053_) decode[20] <= _0932_;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[15] */
always_ff @(posedge clk)
if (_0053_) decode[15] <= regwr_alu;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[148:117] */
always_ff @(posedge clk)
if (_0053_) decode[148:117] <= fetch[31:0];
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[180:149] */
always_ff @(posedge clk)
if (_0053_) decode[180:149] <= fetch[63:32];
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[10:7] */
always_ff @(posedge clk)
if (_0053_)
if (!_0854_) decode[10:7] <= 4'hf;
else decode[10:7] <= _0032_;
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[4] */
always_ff @(posedge clk)
if (_0053_)
if (_0056_) decode[4] <= 1'h0;
else decode[4] <= _0046_[1];
/* src = "generated/sv2v_out.v:1223.2-1251.23" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode[3] */
always_ff @(posedge clk)
if (_0053_)
if (_0057_) decode[3] <= 1'h0;
else decode[3] <= _0044_[0];
assign _0399_ = _0868_ & _0869_;
assign _0402_ = _0904_ & _0871_;
assign _0405_ = _0874_ & _0869_;
assign _0408_ = _0907_ & _0871_;
assign _0411_ = _0870_ & _0871_;
assign _0414_ = fetch_vld_t0 & fetch_rdy;
assign _0417_ = branch_t0 & _0888_;
assign _0420_ = _0171_ & _0948_;
assign _0423_ = decode_vld_t0 & decode_rdy;
assign _0426_ = _0872_ & _0944_;
assign _0400_ = _0870_ & _0867_;
assign _0403_ = _0872_ & _0903_;
assign _0406_ = _0870_ & _0873_;
assign _0409_ = _0872_ & _0906_;
assign _0412_ = _0872_ & _0869_;
assign _0415_ = fetch_rdy_t0 & fetch_vld;
assign _0418_ = _0889_ & branch;
assign _0421_ = csr_t0 & _0898_;
assign _0427_ = _0945_ & _0946_;
assign _0401_ = _0868_ & _0870_;
assign _0404_ = _0904_ & _0872_;
assign _0407_ = _0874_ & _0870_;
assign _0410_ = _0907_ & _0872_;
assign _0413_ = _0870_ & _0872_;
assign _0416_ = fetch_vld_t0 & fetch_rdy_t0;
assign _0419_ = branch_t0 & _0889_;
assign _0422_ = _0171_ & csr_t0;
assign _0428_ = _0872_ & _0945_;
assign _0681_ = _0399_ | _0400_;
assign _0682_ = _0402_ | _0403_;
assign _0683_ = _0405_ | _0406_;
assign _0684_ = _0408_ | _0409_;
assign _0685_ = _0411_ | _0412_;
assign _0686_ = _0414_ | _0415_;
assign _0687_ = _0417_ | _0418_;
assign _0688_ = _0420_ | _0421_;
assign _0689_ = _0423_ | _0424_;
assign _0690_ = _0426_ | _0427_;
assign _0904_ = _0681_ | _0401_;
assign _0009_ = _0682_ | _0404_;
assign _0907_ = _0683_ | _0407_;
assign _0011_ = _0684_ | _0410_;
assign _0170_ = _0685_ | _0413_;
assign _0911_ = _0686_ | _0416_;
assign _0913_ = _0687_ | _0419_;
assign _0915_ = _0688_ | _0422_;
assign _0917_ = _0689_ | _0425_;
assign regwr_alu_t0 = _0690_ | _0428_;
assign _0173_ = | { _0917_, _0911_ };
assign _0175_ = | { _0891_, _0883_, _0881_ };
assign _0176_ = | { _0885_, _0883_, _0881_ };
assign _0177_ = | { _0893_, _0889_, _0891_, _0897_, _0855_ };
assign _0178_ = | { _0893_, _0897_, _0855_ };
assign _0179_ = | { _0959_[2:1], _0957_[2:1], _0864_, _0862_ };
assign _0180_ = | { _0963_, _0959_[2:1], _0957_[2:1], _0862_ };
assign _0181_ = | { _0887_, _0885_ };
assign _0182_ = | { _0736_, _0887_, _0885_, _0855_ };
assign _0184_ = | fetch_t0[31:25];
assign _0185_ = | fetch_t0[31:28];
assign _0186_ = | fetch_t0[19:15];
assign _0187_ = | fetch_t0[11:7];
assign _0192_ = | { _0959_[2:1], _0862_ };
assign _0194_ = | { _0959_[1], _0862_, _0169_ };
assign _0195_ = | { _0963_, _0959_[1], _0864_, _0862_, _0169_ };
assign _0196_ = | { _0963_, _0957_[2:1], _0864_, _0862_, _0169_ };
assign _0193_ = | fetch_t0[14:12];
assign _0073_ = ~ { _0917_, _0911_ };
assign _0074_ = ~ { _0891_, _0883_, _0881_ };
assign _0075_ = ~ { _0885_, _0883_, _0881_ };
assign _0076_ = ~ { _0897_, _0893_, _0891_, _0889_, _0855_ };
assign _0077_ = ~ { _0897_, _0893_, _0855_ };
assign _0078_ = ~ { _0959_[2:1], _0957_[2:1], _0864_, _0862_ };
assign _0079_ = ~ { _0963_, _0959_[2:1], _0957_[2:1], _0862_ };
assign _0080_ = ~ { _0887_, _0885_ };
assign _0090_ = ~ { _0736_, _0887_, _0885_, _0855_ };
assign _0111_ = ~ fetch_t0[31:25];
assign _0112_ = ~ fetch_t0[31:28];
assign _0113_ = ~ fetch_t0[19:15];
assign _0114_ = ~ fetch_t0[11:7];
assign _0142_ = ~ { _0959_[2:1], _0862_ };
assign _0146_ = ~ { _0959_[1], _0862_, _0169_ };
assign _0147_ = ~ { _0963_, _0959_[1], _0864_, _0862_, _0169_ };
assign _0148_ = ~ { _0963_, _0957_[2:1], _0864_, _0862_, _0169_ };
assign _0294_ = { _0916_, _0910_ } & _0073_;
assign _0295_ = { _0890_, _0882_, _0880_ } & _0074_;
assign _0296_ = { _0884_, _0882_, _0880_ } & _0075_;
assign _0297_ = { _0896_, _0892_, _0890_, _0888_, _0854_ } & _0076_;
assign _0298_ = { _0896_, _0892_, _0854_ } & _0077_;
assign _0299_ = { _0958_[2:1], _0956_[2:1], _0863_, _0861_ } & _0078_;
assign _0300_ = { _0962_, _0958_[2:1], _0956_[2:1], _0861_ } & _0079_;
assign _0301_ = { _0886_, _0884_ } & _0080_;
assign _0317_ = { _0735_, _0886_, _0884_, _0854_ } & _0090_;
assign _0390_ = fetch[31:25] & _0111_;
assign _0391_ = fetch[31:28] & _0112_;
assign _0392_ = fetch[19:15] & _0113_;
assign _0393_ = fetch[11:7] & _0114_;
assign _0491_ = { _0958_[2:1], _0861_ } & _0142_;
assign _0499_ = { _0958_[1], _0861_, _0860_ } & _0146_;
assign _0500_ = { _0962_, _0958_[1], _0863_, _0861_, _0860_ } & _0147_;
assign _0501_ = { _0962_, _0956_[2:1], _0863_, _0861_, _0860_ } & _0148_;
assign _0201_ = ! _0294_;
assign _0202_ = ! _0295_;
assign _0203_ = ! _0296_;
assign _0204_ = ! _0297_;
assign _0205_ = ! _0298_;
assign _0206_ = ! _0299_;
assign _0207_ = ! _0300_;
assign _0208_ = ! _0301_;
assign _0209_ = ! _0317_;
assign _0210_ = ! _0389_;
assign _0211_ = ! _0390_;
assign _0212_ = ! _0391_;
assign _0213_ = ! _0392_;
assign _0215_ = ! _0394_;
assign _0214_ = ! _0393_;
assign _0216_ = ! _0491_;
assign _0217_ = ! _0499_;
assign _0218_ = ! _0500_;
assign _0219_ = ! _0501_;
assign _0220_ = ! _0495_;
assign _0221_ = ! _0502_;
assign _0052_ = _0201_ & _0173_;
assign _0059_ = _0202_ & _0175_;
assign _0061_ = _0203_ & _0176_;
assign _0064_ = _0204_ & _0177_;
assign _0068_ = _0205_ & _0178_;
assign _0027_ = _0206_ & _0179_;
assign _0070_ = _0207_ & _0180_;
assign _0066_ = _0208_ & _0181_;
assign _0200_ = _0209_ & _0182_;
assign _0857_ = _0210_ & _0183_;
assign _0005_ = _0211_ & _0184_;
assign _0868_ = _0212_ & _0185_;
assign _0870_ = _0213_ & _0186_;
assign _0874_ = _0215_ & _0188_;
assign _0872_ = _0214_ & _0187_;
assign _0961_ = _0216_ & _0192_;
assign _0041_ = _0217_ & _0194_;
assign _0037_ = _0218_ & _0195_;
assign _0029_ = _0219_ & _0196_;
assign _0169_ = _0220_ & _0193_;
assign _0897_ = _0221_ & _0197_;
assign _0118_ = ~ _0880_;
assign _0121_ = ~ _0922_;
assign _0122_ = ~ _0924_;
assign _0123_ = ~ _0926_;
assign _0125_ = ~ _0928_;
assign _0126_ = ~ _0930_;
assign _0127_ = ~ _0934_;
assign _0120_ = ~ _0920_;
assign _0129_ = ~ _0938_;
assign _0130_ = ~ _0940_;
assign _0131_ = ~ _0942_;
assign _0095_ = ~ _0863_;
assign _0119_ = ~ _0882_;
assign _0083_ = ~ _0888_;
assign _0128_ = ~ is_fencei;
assign _0124_ = ~ _0890_;
assign _0098_ = ~ _0892_;
assign _0096_ = ~ _0884_;
assign _0086_ = ~ _0886_;
assign _0429_ = _0862_ & _0095_;
assign _0432_ = _0881_ & _0119_;
assign _0435_ = _0921_ & _0096_;
assign _0438_ = _0923_ & _0086_;
assign _0441_ = _0925_ & _0083_;
assign _0444_ = _0927_ & _0124_;
assign _0447_ = _0929_ & _0098_;
assign _0450_ = _0931_ & _0081_;
assign _0453_ = _0891_ & _0098_;
assign _0456_ = _0935_ & _0128_;
assign _0459_ = _0921_ & _0124_;
assign _0462_ = _0939_ & _0098_;
assign _0465_ = _0941_ & _0096_;
assign _0468_ = _0943_ & _0086_;
assign _0430_ = _0864_ & _0093_;
assign _0433_ = _0883_ & _0118_;
assign _0436_ = _0885_ & _0120_;
assign _0439_ = _0887_ & _0121_;
assign _0442_ = _0889_ & _0122_;
assign _0445_ = _0891_ & _0123_;
assign _0448_ = _0893_ & _0125_;
assign _0451_ = _0895_ & _0126_;
assign _0454_ = _0893_ & _0124_;
assign _0457_ = is_fencei_t0 & _0127_;
assign _0460_ = _0891_ & _0120_;
assign _0463_ = _0893_ & _0129_;
assign _0466_ = _0885_ & _0130_;
assign _0469_ = _0887_ & _0131_;
assign _0431_ = _0862_ & _0864_;
assign _0434_ = _0881_ & _0883_;
assign _0437_ = _0921_ & _0885_;
assign _0440_ = _0923_ & _0887_;
assign _0443_ = _0925_ & _0889_;
assign _0446_ = _0927_ & _0891_;
assign _0449_ = _0929_ & _0893_;
assign _0452_ = _0931_ & _0895_;
assign _0455_ = _0891_ & _0893_;
assign _0458_ = _0935_ & is_fencei_t0;
assign _0461_ = _0921_ & _0891_;
assign _0464_ = _0939_ & _0893_;
assign _0467_ = _0941_ & _0885_;
assign _0470_ = _0943_ & _0887_;
assign _0691_ = _0429_ | _0430_;
assign _0692_ = _0432_ | _0433_;
assign _0693_ = _0435_ | _0436_;
assign _0694_ = _0438_ | _0439_;
assign _0695_ = _0441_ | _0442_;
assign _0696_ = _0444_ | _0445_;
assign _0697_ = _0447_ | _0448_;
assign _0698_ = _0450_ | _0451_;
assign _0699_ = _0453_ | _0454_;
assign _0700_ = _0456_ | _0457_;
assign _0701_ = _0459_ | _0460_;
assign _0702_ = _0462_ | _0463_;
assign _0703_ = _0465_ | _0466_;
assign _0704_ = _0468_ | _0469_;
assign _0919_ = _0691_ | _0431_;
assign _0921_ = _0692_ | _0434_;
assign _0923_ = _0693_ | _0437_;
assign _0925_ = _0694_ | _0440_;
assign _0927_ = _0695_ | _0443_;
assign _0929_ = _0696_ | _0446_;
assign _0931_ = _0697_ | _0449_;
assign _0933_ = _0698_ | _0452_;
assign _0935_ = _0699_ | _0455_;
assign _0937_ = _0700_ | _0458_;
assign _0939_ = _0701_ | _0461_;
assign _0941_ = _0702_ | _0464_;
assign _0943_ = _0703_ | _0467_;
assign _0945_ = _0704_ | _0470_;
assign _0091_ = ~ _0860_;
assign _0094_ = ~ _0069_;
assign _0097_ = ~ _0735_;
assign _0084_ = ~ _0896_;
assign _0099_ = ~ _0737_;
assign _0100_ = ~ _0199_;
assign _0101_ = ~ { _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_ };
assign _0102_ = ~ { _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_ };
assign _0103_ = ~ { _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_ };
assign _0104_ = ~ { _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_, _0880_ };
assign _0105_ = ~ { _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_ };
assign _0106_ = ~ { _0886_, _0886_, _0886_, _0886_ };
assign _0107_ = ~ { _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_ };
assign _0108_ = ~ { _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_ };
assign _0109_ = ~ { _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_ };
assign _0135_ = ~ _0877_;
assign _0136_ = ~ { _0877_, _0877_ };
assign _0137_ = ~ _0875_;
assign _0138_ = ~ { _0875_, _0875_ };
assign _0139_ = ~ _0873_;
assign _0140_ = ~ _0909_;
assign _0092_ = ~ _0062_;
assign _0141_ = ~ { _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_ };
assign _0093_ = ~ _0861_;
assign _0143_ = ~ _0865_;
assign _0145_ = ~ { _0918_, _0918_, _0918_, _0918_ };
assign _0150_ = ~ { _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_ };
assign _0081_ = ~ _0894_;
assign _0082_ = ~ _0898_;
assign _0151_ = ~ { _0856_, _0856_, _0856_, _0856_ };
assign _0153_ = ~ { rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward };
assign _0154_ = ~ { rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward };
assign _0622_ = _0070_ | _0094_;
assign _0625_ = _0864_ | _0095_;
assign _0631_ = _0885_ | _0096_;
assign _0634_ = _0887_ | _0086_;
assign _0637_ = _0736_ | _0097_;
assign _0640_ = _0897_ | _0084_;
assign _0643_ = _0893_ | _0098_;
assign _0646_ = _0738_ | _0099_;
assign _0649_ = _0200_ | _0100_;
assign _0652_ = { _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_ } | _0101_;
assign _0656_ = { _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_ } | _0102_;
assign _0659_ = { _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_ } | _0103_;
assign _0662_ = { _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_ } | _0104_;
assign _0663_ = { _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_ } | _0105_;
assign _0667_ = { _0887_, _0887_, _0887_, _0887_ } | _0106_;
assign _0670_ = { _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_ } | _0107_;
assign _0673_ = { _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_ } | _0108_;
assign _0676_ = { _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_ } | _0109_;
assign _0707_ = _0878_ | _0135_;
assign _0708_ = { _0878_, _0878_ } | _0136_;
assign _0709_ = _0876_ | _0137_;
assign _0710_ = { _0876_, _0876_ } | _0138_;
assign _0711_ = _0874_ | _0139_;
assign _0618_ = _0027_ | _0092_;
assign _0713_ = { _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_ } | _0141_;
assign _0619_ = _0862_ | _0093_;
assign _0716_ = _0005_ | _0143_;
assign _0717_ = { _0919_, _0919_, _0919_, _0919_ } | _0145_;
assign _0721_ = { _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_ } | _0150_;
assign _0628_ = _0171_ | _0082_;
assign _0726_ = { _0857_, _0857_, _0857_, _0857_ } | _0151_;
assign _0729_ = { rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0 } | _0153_;
assign _0732_ = { rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0 } | _0154_;
assign _0617_ = _0169_ | _0860_;
assign _0623_ = _0070_ | _0069_;
assign _0626_ = _0864_ | _0863_;
assign _0632_ = _0885_ | _0884_;
assign _0635_ = _0887_ | _0886_;
assign _0638_ = _0736_ | _0735_;
assign _0641_ = _0897_ | _0896_;
assign _0644_ = _0893_ | _0892_;
assign _0647_ = _0738_ | _0737_;
assign _0650_ = _0200_ | _0199_;
assign _0653_ = { _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_ } | { _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_, _0886_ };
assign _0655_ = { _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_ } | { _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_, _0854_ };
assign _0657_ = { _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_ } | { _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_, _0739_ };
assign _0660_ = { _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_ } | { _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_, _0898_ };
assign _0664_ = { _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_ } | { _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_, _0741_ };
assign _0666_ = { _0885_, _0885_, _0885_, _0885_ } | { _0884_, _0884_, _0884_, _0884_ };
assign _0668_ = { _0887_, _0887_, _0887_, _0887_ } | { _0886_, _0886_, _0886_, _0886_ };
assign _0671_ = { _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_ } | { _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_, _0967_ };
assign _0674_ = { _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_ } | { _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_, _0971_ };
assign _0677_ = { _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_ } | { _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_, _0743_ };
assign _0712_ = _0170_ | _0909_;
assign _0714_ = { _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_ } | { _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_, _0960_ };
assign _0620_ = _0862_ | _0861_;
assign _0718_ = { _0919_, _0919_, _0919_, _0919_ } | { _0918_, _0918_, _0918_, _0918_ };
assign _0720_ = { _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_ } | { _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_, _0063_ };
assign _0722_ = { _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_ } | { _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_, _0067_ };
assign _0724_ = _0895_ | _0894_;
assign _0629_ = _0171_ | _0898_;
assign _0725_ = { _0859_, _0859_, _0859_, _0859_ } | { _0858_, _0858_, _0858_, _0858_ };
assign _0727_ = { _0857_, _0857_, _0857_, _0857_ } | { _0856_, _0856_, _0856_, _0856_ };
assign _0730_ = { rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0 } | { rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward, rs1_forward };
assign _0733_ = { rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0 } | { rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward, rs2_forward };
assign _0320_ = _0819_ & _0618_;
assign _0324_ = _0821_ & _0619_;
assign _0327_ = _0001_ & _0622_;
assign _0332_ = _0823_ & _0625_;
assign _0335_ = _0007_ & _0628_;
assign _0338_ = _0041_ & _0631_;
assign _0341_ = _0827_ & _0634_;
assign _0344_ = _0829_ & _0637_;
assign _0347_ = _0029_ & _0640_;
assign _0350_ = _0059_ & _0643_;
assign _0353_ = _0836_ & _0646_;
assign _0356_ = _0838_ & _0649_;
assign _0359_ = immediate_t0 & _0652_;
assign _0364_ = _0842_ & _0656_;
assign _0367_ = rs1_data_t0 & _0659_;
assign _0370_ = fetch_t0[63:32] & _0662_;
assign _0372_ = _0846_ & _0663_;
assign _0377_ = _0848_ & _0667_;
assign _0380_ = { rs2_data_t0[15:0], rs2_data_t0[31:16] } & _0670_;
assign _0383_ = rs2_data_t0 & _0673_;
assign _0386_ = _0852_ & _0676_;
assign _0476_ = _0023_ & _0707_;
assign _0478_ = { _0023_, _0023_ } & _0708_;
assign _0480_ = _0021_ & _0709_;
assign _0482_ = _0047_ & _0710_;
assign _0484_ = _0019_ & _0711_;
assign _0488_ = fetch_t0[63:32] & _0713_;
assign _0493_ = _0003_ & _0716_;
assign _0496_ = { 1'h0, fetch_t0[14:12] } & _0717_;
assign _0505_ = fetch_t0[63:32] & _0721_;
assign _0514_ = _0039_ & _0726_;
assign _0518_ = regrd_rs1_t0 & _0729_;
assign _0521_ = regrd_rs2_t0 & _0732_;
assign _0318_ = _0015_ & _0617_;
assign _0322_ = _0009_ & _0617_;
assign _0328_ = _0005_ & _0623_;
assign _0330_ = _0005_ & _0620_;
assign _0333_ = _0001_ & _0626_;
assign _0336_ = _0013_ & _0629_;
assign _0339_ = _0043_ & _0632_;
assign _0342_ = _0050_ & _0635_;
assign _0345_ = _0825_ & _0638_;
assign _0348_ = _0037_ & _0641_;
assign _0351_ = _0169_ & _0644_;
assign _0354_ = _0833_ & _0647_;
assign _0357_ = _0831_ & _0650_;
assign _0360_ = rs2_data_t0 & _0653_;
assign _0362_ = store_data_t0 & _0655_;
assign _0365_ = _0840_ & _0657_;
assign _0368_ = _0035_ & _0660_;
assign _0373_ = _0844_ & _0664_;
assign _0375_ = _0025_ & _0666_;
assign _0378_ = { fetch_t0[30], fetch_t0[14:12] } & _0668_;
assign _0381_ = { rs2_data_t0[7:0], rs2_data_t0[31:8] } & _0671_;
assign _0384_ = { rs2_data_t0[23:0], rs2_data_t0[31:24] } & _0674_;
assign _0387_ = _0850_ & _0677_;
assign _0486_ = _0017_ & _0712_;
assign _0489_ = rs1_data_t0 & _0714_;
assign _0325_ = _0011_ & _0620_;
assign _0497_ = { fetch_t0[30], fetch_t0[14:12] } & _0718_;
assign _0503_ = immediate_t0 & _0720_;
assign _0506_ = rs1_data_t0 & _0722_;
assign _0508_ = _0031_ & _0724_;
assign _0510_ = _0027_ & _0629_;
assign _0512_ = { addr_t0[1], addr_t0[1], addr_t0[1], addr_t0[1] } & _0725_;
assign _0515_ = _0974_ & _0727_;
assign _0519_ = regwr_data_t0 & _0730_;
assign _0522_ = regwr_data_t0 & _0733_;
assign _0621_ = _0324_ | _0325_;
assign _0624_ = _0327_ | _0328_;
assign _0627_ = _0332_ | _0333_;
assign _0630_ = _0335_ | _0336_;
assign _0633_ = _0338_ | _0339_;
assign _0636_ = _0341_ | _0342_;
assign _0639_ = _0344_ | _0345_;
assign _0642_ = _0347_ | _0348_;
assign _0645_ = _0350_ | _0351_;
assign _0648_ = _0353_ | _0354_;
assign _0651_ = _0356_ | _0357_;
assign _0654_ = _0359_ | _0360_;
assign _0658_ = _0364_ | _0365_;
assign _0661_ = _0367_ | _0368_;
assign _0665_ = _0372_ | _0373_;
assign _0669_ = _0377_ | _0378_;
assign _0672_ = _0380_ | _0381_;
assign _0675_ = _0383_ | _0384_;
assign _0678_ = _0386_ | _0387_;
assign _0715_ = _0488_ | _0489_;
assign _0719_ = _0496_ | _0497_;
assign _0723_ = _0505_ | _0506_;
assign _0728_ = _0514_ | _0515_;
assign _0731_ = _0518_ | _0519_;
assign _0734_ = _0521_ | _0522_;
assign _0766_ = _0820_ ^ _0010_;
assign _0767_ = _0000_ ^ _0004_;
assign _0768_ = _0822_ ^ _0000_;
assign _0769_ = _0006_ ^ _0012_;
assign _0770_ = _0040_ ^ _0042_;
assign _0771_ = _0826_ ^ _0049_;
assign _0772_ = _0828_ ^ _0824_;
assign _0773_ = _0028_ ^ _0036_;
assign _0774_ = _0834_ ^ _0860_;
assign _0775_ = _0835_ ^ _0832_;
assign _0776_ = _0837_ ^ _0830_;
assign _0777_ = immediate ^ rs2_data;
assign _0778_ = _0841_ ^ _0839_;
assign _0779_ = rs1_data ^ _0034_;
assign _0780_ = _0845_ ^ _0843_;
assign _0781_ = _0847_ ^ { fetch[30], fetch[14:12] };
assign _0782_ = { rs2_data[15:0], rs2_data[31:16] } ^ { rs2_data[7:0], rs2_data[31:8] };
assign _0783_ = rs2_data ^ { rs2_data[23:0], rs2_data[31:24] };
assign _0784_ = _0851_ ^ _0849_;
assign _0785_ = fetch[63:32] ^ rs1_data;
assign _0786_ = { 1'h0, fetch[14:12] } ^ { fetch[30], fetch[14:12] };
assign _0787_ = _0038_ ^ _0973_;
assign _0788_ = regrd_rs1 ^ regwr_data;
assign _0789_ = regrd_rs2 ^ regwr_data;
assign _0319_ = _0169_ & _0014_;
assign _0321_ = _0027_ & _0161_;
assign _0323_ = _0169_ & _0008_;
assign _0326_ = _0862_ & _0766_;
assign _0329_ = _0070_ & _0767_;
assign _0331_ = _0862_ & _0156_;
assign _0334_ = _0864_ & _0768_;
assign _0337_ = _0171_ & _0769_;
assign _0340_ = _0885_ & _0770_;
assign _0343_ = _0887_ & _0771_;
assign _0346_ = _0736_ & _0772_;
assign _0349_ = _0897_ & _0773_;
assign _0352_ = _0893_ & _0774_;
assign _0355_ = _0738_ & _0775_;
assign _0358_ = _0200_ & _0776_;
assign _0361_ = { _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_, _0887_ } & _0777_;
assign _0363_ = { _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_, _0855_ } & { store_data[31:3], _0162_, store_data[1:0] };
assign _0366_ = { _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_, _0740_ } & _0778_;
assign _0369_ = { _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_, _0171_ } & _0779_;
assign _0371_ = { _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_, _0881_ } & fetch[63:32];
assign _0374_ = { _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_, _0742_ } & _0780_;
assign _0376_ = { _0885_, _0885_, _0885_, _0885_ } & _0024_;
assign _0379_ = { _0887_, _0887_, _0887_, _0887_ } & _0781_;
assign _0382_ = { _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_, _0968_ } & _0782_;
assign _0385_ = { _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_, _0972_ } & _0783_;
assign _0388_ = { _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_, _0744_ } & _0784_;
assign _0955_ = _0911_ & _0155_;
assign _0477_ = _0878_ & _0158_;
assign _0479_ = { _0878_, _0878_ } & { _0164_, _0048_[0] };
assign _0481_ = _0876_ & _0159_;
assign _0483_ = { _0876_, _0876_ } & { _0046_[1], _0165_ };
assign _0485_ = _0874_ & _0160_;
assign _0487_ = _0170_ & _0016_;
assign _0490_ = { _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_, _0961_ } & _0785_;
assign _0492_ = _0862_ & _0010_;
assign _0494_ = _0005_ & _0157_;
assign _0498_ = { _0919_, _0919_, _0919_, _0919_ } & _0786_;
assign _0504_ = { _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_, _0064_ } & { immediate[31:3], _0166_, immediate[1:0] };
assign _0507_ = { _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_, _0068_ } & _0785_;
assign _0509_ = _0895_ & _0030_;
assign _0511_ = _0171_ & _0026_;
assign _0513_ = { _0859_, _0859_, _0859_, _0859_ } & _0163_;
assign _0516_ = { _0857_, _0857_, _0857_, _0857_ } & _0787_;
assign _0520_ = { rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0, rs1_forward_t0 } & _0788_;
assign _0523_ = { rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0, rs2_forward_t0 } & _0789_;
assign _0819_ = _0319_ | _0318_;
assign _0013_ = _0321_ | _0320_;
assign _0821_ = _0323_ | _0322_;
assign _0007_ = _0326_ | _0621_;
assign _0050_ = _0329_ | _0624_;
assign _0823_ = _0331_ | _0330_;
assign _0043_ = _0334_ | _0627_;
assign _0825_ = _0337_ | _0630_;
assign _0827_ = _0340_ | _0633_;
assign _0829_ = _0343_ | _0636_;
assign _0831_ = _0346_ | _0639_;
assign _0833_ = _0349_ | _0642_;
assign _0836_ = _0352_ | _0645_;
assign _0838_ = _0355_ | _0648_;
assign instr_valid_t0 = _0358_ | _0651_;
assign _0840_ = _0361_ | _0654_;
assign _0842_ = _0363_ | _0362_;
assign op2_t0 = _0366_ | _0658_;
assign _0844_ = _0369_ | _0661_;
assign _0846_ = _0371_ | _0370_;
assign op1_t0 = _0374_ | _0665_;
assign _0848_ = _0376_ | _0375_;
assign aluop_t0 = _0379_ | _0669_;
assign _0850_ = _0382_ | _0672_;
assign _0852_ = _0385_ | _0675_;
assign store_data_t0 = _0388_ | _0678_;
assign _0021_ = _0477_ | _0476_;
assign _0047_ = _0479_ | _0478_;
assign _0019_ = _0481_ | _0480_;
assign _0045_ = _0483_ | _0482_;
assign _0017_ = _0485_ | _0484_;
assign _0015_ = _0487_ | _0486_;
assign _0035_ = _0490_ | _0715_;
assign _0031_ = _0492_ | _0325_;
assign _0001_ = _0494_ | _0493_;
assign _0025_ = _0498_ | _0719_;
assign offset_t0 = _0504_ | _0503_;
assign base_t0 = _0507_ | _0723_;
assign is_fencei_t0 = _0509_ | _0508_;
assign csr_t0 = _0511_ | _0510_;
assign _0039_ = _0513_ | _0512_;
assign _0033_ = _0516_ | _0728_;
assign rs1_data_t0 = _0520_ | _0731_;
assign rs2_data_t0 = _0523_ | _0734_;
assign _0051_ = | { _0916_, _0910_ };
assign _0168_ = ~ flush;
assign _0053_ = & { _0910_, _0168_, rstz };
assign _0167_ = ~ rstz;
assign _0055_ = | { _0167_, flush };
assign _0056_ = | { _0140_, _0091_, _0082_, _0875_, _0873_ };
assign _0057_ = | { _0140_, _0091_, _0082_, _0873_ };
assign _0155_ = ~ _0953_;
assign _0156_ = ~ _0004_;
assign _0157_ = ~ _0002_;
assign _0158_ = ~ _0022_;
assign _0159_ = ~ _0020_;
assign _0160_ = ~ _0018_;
assign _0161_ = ~ _0818_;
assign _0162_ = ~ store_data[2];
assign _0163_ = ~ _0975_;
assign _0164_ = ~ _0048_[1];
assign _0165_ = ~ _0046_[0];
assign _0166_ = ~ immediate[2];
assign _0058_ = | { _0890_, _0882_, _0880_ };
assign _0060_ = | { _0884_, _0882_, _0880_ };
assign _0063_ = | { _0896_, _0892_, _0890_, _0888_, _0854_ };
assign _0067_ = | { _0896_, _0892_, _0854_ };
assign _0062_ = | { _0958_[2:1], _0956_[2:1], _0863_, _0861_ };
assign _0069_ = | { _0962_, _0958_[2:1], _0956_[2:1], _0861_ };
assign _0085_ = ~ _0060_;
assign _0087_ = ~ _0065_;
assign _0088_ = ~ _0969_;
assign _0089_ = ~ _0967_;
assign _0133_ = ~ illegal_opcode;
assign _0134_ = ~ decode_rdy;
assign _0302_ = _0895_ & _0082_;
assign _0305_ = _0889_ & _0084_;
assign _0308_ = _0061_ & _0086_;
assign _0311_ = _0066_ & _0082_;
assign _0314_ = _0970_ & _0089_;
assign _0472_ = instr_valid_t0 & _0133_;
assign _0475_ = decode_vld_t0 & _0134_;
assign _0303_ = _0171_ & _0081_;
assign _0306_ = _0897_ & _0083_;
assign _0309_ = _0887_ & _0085_;
assign _0312_ = _0171_ & _0087_;
assign _0315_ = _0968_ & _0088_;
assign _0473_ = illegal_opcode_t0 & instr_valid;
assign _0424_ = decode_rdy_t0 & decode_vld;
assign _0304_ = _0895_ & _0171_;
assign _0307_ = _0889_ & _0897_;
assign _0310_ = _0061_ & _0887_;
assign _0313_ = _0066_ & _0171_;
assign _0316_ = _0970_ & _0968_;
assign _0474_ = instr_valid_t0 & illegal_opcode_t0;
assign _0425_ = decode_vld_t0 & decode_rdy_t0;
assign _0612_ = _0302_ | _0303_;
assign _0613_ = _0305_ | _0306_;
assign _0614_ = _0308_ | _0309_;
assign _0615_ = _0311_ | _0312_;
assign _0616_ = _0314_ | _0315_;
assign _0705_ = _0472_ | _0473_;
assign _0706_ = _0475_ | _0424_;
assign _0736_ = _0612_ | _0304_;
assign _0738_ = _0613_ | _0307_;
assign _0740_ = _0614_ | _0310_;
assign _0742_ = _0615_ | _0313_;
assign _0744_ = _0616_ | _0316_;
assign illegal_t0 = _0705_ | _0474_;
assign _0952_ = _0706_ | _0425_;
assign _0065_ = | { _0886_, _0884_ };
assign _0735_ = _0894_ | _0898_;
assign _0737_ = _0888_ | _0896_;
assign _0739_ = _0060_ | _0886_;
assign _0741_ = _0065_ | _0898_;
assign _0743_ = _0969_ | _0967_;
assign _0199_ = | { _0735_, _0886_, _0884_, _0854_ };
assign _0818_ = _0860_ ? _0014_ : 1'h0;
assign _0012_ = _0062_ ? 1'h1 : _0818_;
assign _0820_ = _0860_ ? _0008_ : 1'h0;
assign _0006_ = _0861_ ? _0010_ : _0820_;
assign _0049_ = _0069_ ? _0004_ : _0000_;
assign _0822_ = _0861_ ? _0004_ : 1'h1;
assign _0042_ = _0863_ ? _0000_ : _0822_;
assign _0824_ = _0898_ ? _0012_ : _0006_;
assign _0826_ = _0884_ ? _0042_ : _0040_;
assign _0828_ = _0886_ ? _0049_ : _0826_;
assign _0830_ = _0735_ ? _0824_ : _0828_;
assign _0832_ = _0896_ ? _0036_ : _0028_;
assign _0834_ = _0058_ ? 1'h1 : 1'h0;
assign _0835_ = _0892_ ? _0860_ : _0834_;
assign _0837_ = _0737_ ? _0832_ : _0835_;
assign instr_valid = _0199_ ? _0830_ : _0837_;
assign _0839_ = _0886_ ? rs2_data : immediate;
assign _0841_ = _0854_ ? store_data : 32'd4;
assign op2 = _0739_ ? _0839_ : _0841_;
assign _0843_ = _0898_ ? _0034_ : rs1_data;
assign _0845_ = _0880_ ? 32'd0 : fetch[63:32];
assign op1 = _0741_ ? _0843_ : _0845_;
assign _0847_ = _0884_ ? _0024_ : 4'h0;
assign aluop = _0886_ ? { fetch[30], fetch[14:12] } : _0847_;
assign _0849_ = _0967_ ? { rs2_data[7:0], rs2_data[31:8] } : { rs2_data[15:0], rs2_data[31:16] };
assign _0851_ = _0971_ ? { rs2_data[23:0], rs2_data[31:24] } : rs2_data;
assign store_data = _0743_ ? _0849_ : _0851_;
assign _0174_ = | { _0911_, flush_t0 };
assign _0611_ = { _0910_, _0168_, rstz } | { _0911_, flush_t0, 1'h0 };
assign _0172_ = & _0611_;
assign _0054_ = _0174_ & _0172_;
assign _0072_ = ~ _0053_;
assign _0763_ = _0032_ ^ decode[10:7];
assign _0764_ = _0046_[1] ^ decode[4];
assign _0765_ = _0044_[0] ^ decode[3];
assign _0599_ = _0033_ | decode_t0[10:7];
assign _0603_ = _0047_[1] | decode_t0[4];
assign _0607_ = _0045_[0] | decode_t0[3];
assign _0600_ = _0763_ | _0599_;
assign _0604_ = _0764_ | _0603_;
assign _0608_ = _0765_ | _0607_;
assign _0285_ = { _0053_, _0053_, _0053_, _0053_ } & _0033_;
assign _0288_ = _0053_ & _0047_[1];
assign _0291_ = _0053_ & _0045_[0];
assign _0286_ = { _0072_, _0072_, _0072_, _0072_ } & decode_t0[10:7];
assign _0289_ = _0072_ & decode_t0[4];
assign _0292_ = _0072_ & decode_t0[3];
assign _0287_ = _0600_ & { _0054_, _0054_, _0054_, _0054_ };
assign _0290_ = _0604_ & _0054_;
assign _0293_ = _0608_ & _0054_;
assign _0601_ = _0285_ | _0286_;
assign _0605_ = _0288_ | _0289_;
assign _0609_ = _0291_ | _0292_;
assign _0602_ = _0601_ | _0287_;
assign _0606_ = _0605_ | _0290_;
assign _0610_ = _0609_ | _0293_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[10:7] */
always_ff @(posedge clk)
if (!_0854_) decode_t0[10:7] <= 4'h0;
else decode_t0[10:7] <= _0602_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[4] */
always_ff @(posedge clk)
if (_0056_) decode_t0[4] <= 1'h0;
else decode_t0[4] <= _0606_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_t0[3] */
always_ff @(posedge clk)
if (_0057_) decode_t0[3] <= 1'h0;
else decode_t0[3] <= _0610_;
assign _0071_ = ~ _0051_;
assign _0745_ = _0954_ ^ decode_vld;
assign _0527_ = _0955_ | decode_vld_t0;
assign _0528_ = _0745_ | _0527_;
assign _0231_ = _0051_ & _0955_;
assign _0232_ = _0071_ & decode_vld_t0;
assign _0233_ = _0528_ & _0052_;
assign _0529_ = _0231_ | _0232_;
assign _0530_ = _0529_ | _0233_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_62dbb6e3107130a7cf75  */
/* PC_TAINT_INFO STATE_NAME decode_vld_t0 */
always_ff @(posedge clk)
if (_0055_) decode_vld_t0 <= 1'h0;
else decode_vld_t0 <= _0530_;
assign _0853_ = 4'h0 << addr[1:0];
assign _0974_ = { _0198_, _0198_, _0198_, _0198_ } | _0853_;
assign _0856_ = ! /* src = "generated/sv2v_out.v:1039.8-1039.38" */ fetch[13:12];
assign _0858_ = fetch[13:12] == /* src = "generated/sv2v_out.v:1041.13-1041.43" */ 2'h1;
assign _0866_ = fetch[31:25] == /* src = "generated/sv2v_out.v:1134.16-1134.31" */ 7'h20;
assign _0865_ = ! /* src = "generated/sv2v_out.v:1140.11-1140.25" */ fetch[31:25];
assign _0867_ = ! /* src = "generated/sv2v_out.v:1147.13-1147.39" */ fetch[31:28];
assign _0869_ = ! /* src = "generated/sv2v_out.v:1158.12-1158.30" */ fetch[19:15];
assign _0871_ = ! /* src = "generated/sv2v_out.v:1158.36-1158.53" */ fetch[11:7];
assign _0873_ = ! /* src = "generated/sv2v_out.v:1159.12-1159.32" */ fetch[31:20];
assign _0875_ = fetch[31:20] == /* src = "generated/sv2v_out.v:1163.17-1163.37" */ 12'h001;
assign _0877_ = fetch[31:20] == /* src = "generated/sv2v_out.v:1167.17-1167.37" */ 12'h302;
assign _0879_ = fetch[31:20] == /* src = "generated/sv2v_out.v:1171.17-1171.37" */ 12'h105;
assign _0899_ = regwr_sel == /* src = "generated/sv2v_out.v:996.35-996.51" */ fetch[19:15];
assign _0901_ = regwr_sel == /* src = "generated/sv2v_out.v:997.35-997.51" */ fetch[24:20];
assign _0903_ = _0867_ && /* src = "generated/sv2v_out.v:1147.12-1147.64" */ _0869_;
assign _0905_ = _0903_ && /* src = "generated/sv2v_out.v:1147.11-1147.88" */ _0871_;
assign _0906_ = _0873_ && /* src = "generated/sv2v_out.v:1150.12-1150.67" */ _0869_;
assign _0908_ = _0906_ && /* src = "generated/sv2v_out.v:1150.11-1150.91" */ _0871_;
assign _0909_ = _0869_ && /* src = "generated/sv2v_out.v:1158.11-1158.54" */ _0871_;
assign _0910_ = fetch_vld && /* src = "generated/sv2v_out.v:1228.12-1228.34" */ fetch_rdy;
assign _0912_ = branch && /* src = "generated/sv2v_out.v:1239.18-1239.57" */ _0888_;
assign _0914_ = _0898_ && /* src = "generated/sv2v_out.v:1244.17-1244.55" */ _0948_;
assign _0916_ = decode_vld && /* src = "generated/sv2v_out.v:1250.12-1250.36" */ decode_rdy;
assign regwr_alu = _0946_ && /* src = "generated/sv2v_out.v:995.21-995.258" */ _0944_;
assign _0918_ = _0861_ || /* src = "generated/sv2v_out.v:1091.9-1091.49" */ _0863_;
assign _0920_ = _0880_ || /* src = "generated/sv2v_out.v:1232.24-1232.90" */ _0882_;
assign _0922_ = _0920_ || /* src = "generated/sv2v_out.v:1232.23-1232.127" */ _0884_;
assign _0924_ = _0922_ || /* src = "generated/sv2v_out.v:1232.22-1232.161" */ _0886_;
assign _0926_ = _0924_ || /* src = "generated/sv2v_out.v:1232.21-1232.195" */ _0888_;
assign _0928_ = _0926_ || /* src = "generated/sv2v_out.v:1232.20-1232.230" */ _0890_;
assign _0930_ = _0928_ || /* src = "generated/sv2v_out.v:1232.19-1232.266" */ _0892_;
assign _0932_ = _0930_ || /* src = "generated/sv2v_out.v:1232.18-1232.302" */ _0894_;
assign _0934_ = _0890_ || /* src = "generated/sv2v_out.v:1238.19-1238.84" */ _0892_;
assign _0936_ = _0934_ || /* src = "generated/sv2v_out.v:1238.18-1238.98" */ is_fencei;
assign _0938_ = _0920_ || /* src = "generated/sv2v_out.v:995.48-995.150" */ _0890_;
assign _0940_ = _0938_ || /* src = "generated/sv2v_out.v:995.47-995.186" */ _0892_;
assign _0942_ = _0940_ || /* src = "generated/sv2v_out.v:995.46-995.223" */ _0884_;
assign _0944_ = _0942_ || /* src = "generated/sv2v_out.v:995.45-995.257" */ _0886_;
assign illegal_opcode = fetch[1:0] != /* src = "generated/sv2v_out.v:988.26-988.46" */ 2'h3;
assign _0946_ = | /* src = "generated/sv2v_out.v:995.22-995.39" */ fetch[11:7];
assign _0947_ = ~ /* src = "generated/sv2v_out.v:1189.42-1189.54" */ instr_valid;
assign _0948_ = ~ /* src = "generated/sv2v_out.v:1244.51-1244.55" */ csr;
assign _0949_ = ~ /* src = "generated/sv2v_out.v:1252.22-1252.33" */ decode_vld;
assign _0950_ = ~ /* src = "generated/sv2v_out.v:1252.50-1252.56" */ stall;
assign illegal = _0947_ | /* src = "generated/sv2v_out.v:1189.42-1189.71" */ illegal_opcode;
assign _0951_ = _0949_ | /* src = "generated/sv2v_out.v:1252.22-1252.46" */ decode_rdy;
assign _0953_ = _0916_ ? /* src = "generated/sv2v_out.v:1250.12-1250.36|generated/sv2v_out.v:1250.8-1251.23" */ 1'h0 : 1'hx;
assign _0954_ = _0910_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1228.12-1228.34|generated/sv2v_out.v:1228.8-1251.23" */ 1'h1 : _0953_;
assign _0022_ = _0879_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1171.17-1171.37|generated/sv2v_out.v:1171.13-1174.11" */ 1'h1 : 1'h0;
assign _0048_ = _0879_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1171.17-1171.37|generated/sv2v_out.v:1171.13-1174.11" */ 2'h3 : 2'h0;
assign _0020_ = _0877_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1167.17-1167.37|generated/sv2v_out.v:1167.13-1174.11" */ 1'h1 : _0022_;
assign _0046_ = _0877_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1167.17-1167.37|generated/sv2v_out.v:1167.13-1174.11" */ 2'h2 : _0048_;
assign _0018_ = _0875_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1163.17-1163.37|generated/sv2v_out.v:1163.13-1174.11" */ 1'h1 : _0020_;
assign _0044_ = _0875_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1163.17-1163.37|generated/sv2v_out.v:1163.13-1174.11" */ 2'h1 : _0046_;
assign _0016_ = _0873_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1159.12-1159.32|generated/sv2v_out.v:1159.8-1174.11" */ 1'h1 : _0018_;
assign _0014_ = _0909_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1158.11-1158.54|generated/sv2v_out.v:1158.7-1174.11" */ _0016_ : 1'h0;
assign _0026_ = _0062_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1156.5-1184.12" */ 1'h1 : 1'h0;
assign _0034_ = _0960_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1156.5-1184.12" */ rs1_data : fetch[63:32];
assign _0960_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1156.5-1184.12" */ { _0958_[2:1], _0861_ };
assign _0010_ = _0908_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1150.11-1150.91|generated/sv2v_out.v:1150.7-1153.10" */ 1'h1 : 1'h0;
assign _0008_ = _0905_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1147.11-1147.88|generated/sv2v_out.v:1147.7-1148.27" */ 1'h1 : 1'h0;
assign _0030_ = _0861_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1145.5-1154.12" */ _0010_ : 1'h0;
assign _0002_ = _0866_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1105.16-1105.31|generated/sv2v_out.v:1105.12-1106.27" */ 1'h1 : 1'h0;
assign _0000_ = _0865_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1103.11-1103.25|generated/sv2v_out.v:1103.7-1106.27" */ 1'h1 : _0002_;
assign _0004_ = _0865_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1100.11-1100.25|generated/sv2v_out.v:1100.7-1101.27" */ 1'h1 : 1'h0;
assign _0958_[2] = fetch[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1097.5-1107.12" */ 3'h3;
assign _0024_ = _0918_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1091.9-1091.49|generated/sv2v_out.v:1091.5-1094.29" */ { fetch[30], fetch[14:12] } : { 1'h0, fetch[14:12] };
assign _0040_ = _0964_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1086.5-1088.12" */ 1'h1 : 1'h0;
assign _0964_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1086.5-1088.12" */ { _0958_[1], _0861_, _0860_ };
assign _0036_ = _0965_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1078.5-1080.12" */ 1'h1 : 1'h0;
assign _0965_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1078.5-1080.12" */ { _0962_, _0958_[1], _0863_, _0861_, _0860_ };
assign _0958_[1] = fetch[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1078.5-1080.12" */ 3'h2;
assign _0028_ = _0966_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1071.5-1073.12" */ 1'h1 : 1'h0;
assign _0966_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1071.5-1073.12" */ { _0962_, _0956_[2:1], _0863_, _0861_, _0860_ };
assign _0860_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1071.5-1073.12" */ fetch[14:12];
assign _0861_ = fetch[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1071.5-1073.12" */ 3'h1;
assign _0962_ = fetch[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1071.5-1073.12" */ 3'h4;
assign _0863_ = fetch[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1071.5-1073.12" */ 3'h5;
assign _0956_[1] = fetch[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1071.5-1073.12" */ 3'h6;
assign _0956_[2] = fetch[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1071.5-1073.12" */ 3'h7;
assign _0882_ = fetch[6:2] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1048.3-1187.10" */ 5'h05;
assign _0880_ = fetch[6:2] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1048.3-1187.10" */ 5'h0d;
assign offset = _0063_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1048.3-1187.10" */ immediate : 32'd4;
assign _0888_ = fetch[6:2] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1048.3-1187.10" */ 5'h18;
assign _0890_ = fetch[6:2] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1048.3-1187.10" */ 5'h1b;
assign base = _0067_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1048.3-1187.10" */ rs1_data : fetch[63:32];
assign _0854_ = fetch[6:2] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1048.3-1187.10" */ 5'h08;
assign _0896_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1048.3-1187.10" */ fetch[6:2];
assign _0892_ = fetch[6:2] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1048.3-1187.10" */ 5'h19;
assign is_fencei = _0894_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1048.3-1187.10" */ _0030_ : 1'h0;
assign _0894_ = fetch[6:2] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1048.3-1187.10" */ 5'h03;
assign csr = _0898_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1048.3-1187.10" */ _0026_ : 1'h0;
assign _0898_ = fetch[6:2] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1048.3-1187.10" */ 5'h1c;
assign _0886_ = fetch[6:2] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1048.3-1187.10" */ 5'h0c;
assign _0884_ = fetch[6:2] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1048.3-1187.10" */ 5'h04;
assign _0038_ = _0858_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1041.13-1041.43|generated/sv2v_out.v:1041.9-1044.17" */ _0975_ : 4'hf;
assign _0032_ = _0856_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1039.8-1039.38|generated/sv2v_out.v:1039.4-1044.17" */ _0973_ : _0038_;
assign _0967_ = addr[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1032.3-1037.10" */ 2'h3;
assign _0969_ = addr[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1032.3-1037.10" */ 2'h2;
assign _0971_ = addr[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1032.3-1037.10" */ 2'h1;
assign _0973_ = 4'h1 << /* src = "generated/sv2v_out.v:1040.12-1040.29" */ addr[1:0];
assign _0975_ = addr[1] ? /* src = "generated/sv2v_out.v:1042.13-1042.39" */ 4'hc : 4'h3;
assign rs1_data = rs1_forward ? /* src = "generated/sv2v_out.v:998.21-998.57" */ regwr_data : regrd_rs1;
assign rs2_data = rs2_forward ? /* src = "generated/sv2v_out.v:999.21-999.57" */ regwr_data : regrd_rs2;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:1193.4-1200.3" */
paramodsimplif_8a2982a34f91f245ed13  u_agu (
.addr(addr),
.addr_t0(addr_t0),
.base(base),
.base_t0(base_t0),
.instr(fetch[31:0]),
.instr_t0(fetch_t0[31:0]),
.misaligned_jmp(misaligned_jmp),
.misaligned_jmp_t0(misaligned_jmp_t0),
.misaligned_ldst(misaligned_ldst),
.misaligned_ldst_t0(misaligned_ldst_t0),
.offset(offset),
.offset_t0(offset_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:1201.16-1206.3" */
kronos_branch u_branch (
.branch(branch),
.branch_t0(branch_t0),
.op(fetch[14:12]),
.op_t0(fetch_t0[14:12]),
.rs1(rs1_data),
.rs1_t0(rs1_data_t0),
.rs2(rs2_data),
.rs2_t0(rs2_data_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:1207.13-1222.3" */
kronos_hcu u_hcu (
.clk(clk),
.clk_t0(clk_t0),
.decode_rdy(decode_rdy),
.decode_rdy_t0(decode_rdy_t0),
.decode_vld(decode_vld),
.decode_vld_t0(decode_vld_t0),
.fetch_rdy(fetch_rdy),
.fetch_rdy_t0(fetch_rdy_t0),
.fetch_vld(fetch_vld),
.fetch_vld_t0(fetch_vld_t0),
.flush(flush),
.flush_t0(flush_t0),
.instr(fetch[31:0]),
.instr_t0(fetch_t0[31:0]),
.regrd_rs1_en(regrd_rs1_en),
.regrd_rs1_en_t0(regrd_rs1_en_t0),
.regrd_rs2_en(regrd_rs2_en),
.regrd_rs2_en_t0(regrd_rs2_en_t0),
.regwr_en(regwr_en),
.regwr_en_t0(regwr_en_t0),
.regwr_pending(regwr_pending),
.regwr_pending_t0(regwr_pending_t0),
.regwr_sel(regwr_sel),
.regwr_sel_t0(regwr_sel_t0),
.rstz(rstz),
.stall(stall),
.stall_t0(stall_t0)
);
assign _0956_[0] = _0863_;
assign _0957_[0] = _0864_;
assign _0958_[0] = _0861_;
assign _0959_[0] = _0862_;
// Added block to randomize initial values.
`ifdef RANDOMIZE_INIT
  initial begin
    decode_t0[1] = '0;
    decode_t0[0] = '0;
    decode_t0[2] = '0;
    decode_t0[5] = '0;
    decode_t0[6] = '0;
    decode_t0[11] = '0;
    decode_t0[12] = '0;
    decode_t0[13] = '0;
    decode_t0[14] = '0;
    decode_t0[52:21] = '0;
    decode_t0[116:85] = '0;
    decode_t0[84:53] = '0;
    decode_t0[19:16] = '0;
    decode_t0[20] = '0;
    decode_t0[15] = '0;
    decode_t0[148:117] = '0;
    decode_t0[180:149] = '0;
    decode_vld = '0;
    decode[1] = '0;
    decode[0] = '0;
    decode[2] = '0;
    decode[5] = '0;
    decode[6] = '0;
    decode[11] = '0;
    decode[12] = '0;
    decode[13] = '0;
    decode[14] = '0;
    decode[52:21] = '0;
    decode[116:85] = '0;
    decode[84:53] = '0;
    decode[19:16] = '0;
    decode[20] = '0;
    decode[15] = '0;
    decode[148:117] = '0;
    decode[180:149] = '0;
    decode[10:7] = '0;
    decode[4] = '0;
    decode[3] = '0;
    decode_t0[10:7] = '0;
    decode_t0[4] = '0;
    decode_t0[3] = '0;
    decode_vld_t0 = '0;
  end
`endif // RANDOMIZE_INIT
endmodule

module paramodsimplif_b656ed3944a4d79ba92b (clk, rstz, incr, load_data, load_low, load_high, count, count_vld, clk_t0, incr_t0, load_data_t0, load_high_t0, load_low_t0, count_t0, count_vld_t0);
/* src = "generated/sv2v_out.v:300.19-300.35" */
wire [31:0] _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:300.19-300.35" */
wire [31:0] _001_;
/* src = "generated/sv2v_out.v:304.20-304.37" */
wire [31:0] _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:304.20-304.37" */
wire [31:0] _003_;
wire _004_;
/* cellift = 32'd1 */
wire _005_;
wire _006_;
/* cellift = 32'd1 */
wire _007_;
wire _008_;
/* cellift = 32'd1 */
wire _009_;
wire _010_;
/* cellift = 32'd1 */
wire _011_;
wire _012_;
/* cellift = 32'd1 */
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire [31:0] _018_;
wire [31:0] _019_;
wire _020_;
wire _021_;
wire [2:0] _022_;
wire [1:0] _023_;
wire [1:0] _024_;
wire [31:0] _025_;
wire [31:0] _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire [31:0] _037_;
wire [31:0] _038_;
wire [31:0] _039_;
wire [31:0] _040_;
wire [31:0] _041_;
wire [31:0] _042_;
wire [31:0] _043_;
wire [31:0] _044_;
wire [2:0] _045_;
wire [1:0] _046_;
wire [1:0] _047_;
wire [31:0] _048_;
wire [31:0] _049_;
wire [31:0] _050_;
wire [31:0] _051_;
wire [31:0] _052_;
wire [31:0] _053_;
wire [31:0] _054_;
wire [31:0] _055_;
wire [31:0] _056_;
wire [31:0] _057_;
wire [31:0] _058_;
wire [31:0] _059_;
wire [31:0] _060_;
wire [31:0] _061_;
wire [31:0] _062_;
wire [31:0] _063_;
wire [1:0] _064_;
wire [1:0] _065_;
wire [31:0] _066_;
wire [31:0] _067_;
wire [31:0] _068_;
wire [31:0] _069_;
wire [31:0] _070_;
wire [31:0] _071_;
wire [31:0] _072_;
wire [31:0] _073_;
wire [31:0] _074_;
wire [31:0] _075_;
wire [31:0] _076_;
wire [31:0] _077_;
wire [31:0] _078_;
wire [31:0] _079_;
wire _080_;
wire _081_;
wire [31:0] _082_;
wire [31:0] _083_;
wire [31:0] _084_;
wire [31:0] _085_;
/* src = "generated/sv2v_out.v:301.19-301.44" */
wire _086_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:301.19-301.44" */
wire _087_;
wire [31:0] _088_;
/* cellift = 32'd1 */
wire [31:0] _089_;
wire [31:0] _090_;
/* cellift = 32'd1 */
wire [31:0] _091_;
wire [31:0] _092_;
/* cellift = 32'd1 */
wire [31:0] _093_;
wire [31:0] _094_;
/* cellift = 32'd1 */
wire [31:0] _095_;
wire [31:0] _096_;
/* cellift = 32'd1 */
wire [31:0] _097_;
/* src = "generated/sv2v_out.v:275.13-275.16" */
input clk;
wire clk;
/* cellift = 32'd1 */
input clk_t0;
wire clk_t0;
/* src = "generated/sv2v_out.v:281.21-281.26" */
output [63:0] count;
wire [63:0] count;
/* src = "generated/sv2v_out.v:284.13-284.23" */
reg [31:0] count_high;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:284.13-284.23" */
reg [31:0] count_high_t0;
/* src = "generated/sv2v_out.v:283.13-283.22" */
reg [31:0] count_low;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:283.13-283.22" */
reg [31:0] count_low_t0;
/* cellift = 32'd1 */
output [63:0] count_t0;
wire [63:0] count_t0;
/* src = "generated/sv2v_out.v:282.14-282.23" */
output count_vld;
wire count_vld;
/* cellift = 32'd1 */
output count_vld_t0;
reg count_vld_t0;
/* src = "generated/sv2v_out.v:277.13-277.17" */
input incr;
wire incr;
/* src = "generated/sv2v_out.v:285.6-285.15" */
reg incr_high;
/* cellift = 32'd1 */
input incr_t0;
wire incr_t0;
/* src = "generated/sv2v_out.v:278.20-278.29" */
input [31:0] load_data;
wire [31:0] load_data;
/* cellift = 32'd1 */
input [31:0] load_data_t0;
wire [31:0] load_data_t0;
/* src = "generated/sv2v_out.v:280.13-280.22" */
input load_high;
wire load_high;
/* cellift = 32'd1 */
input load_high_t0;
wire load_high_t0;
/* src = "generated/sv2v_out.v:279.13-279.21" */
input load_low;
wire load_low;
/* cellift = 32'd1 */
input load_low_t0;
wire load_low_t0;
/* src = "generated/sv2v_out.v:276.13-276.17" */
input rstz;
wire rstz;
assign _000_ = count_low + /* src = "generated/sv2v_out.v:300.19-300.35" */ 1'h1;
assign _002_ = count_high + /* src = "generated/sv2v_out.v:304.20-304.37" */ 1'h1;
assign _019_ = ~ count_high_t0;
assign _038_ = count_high & _019_;
assign _082_ = _037_ + 32'd1;
assign _084_ = _038_ + 32'd1;
assign _054_ = count_low | count_low_t0;
assign _055_ = count_high | count_high_t0;
assign _083_ = _054_ + 32'd1;
assign _085_ = _055_ + 32'd1;
assign _074_ = _082_ ^ _083_;
assign _075_ = _084_ ^ _085_;
assign _001_ = _074_ | count_low_t0;
assign _003_ = _075_ | count_high_t0;
assign _030_ = | { load_low_t0, load_high_t0 };
assign _034_ = | count_low_t0;
assign _023_ = ~ { load_high_t0, load_low_t0 };
assign _018_ = ~ count_low_t0;
assign _046_ = { load_high, load_low } & _023_;
assign _037_ = count_low & _018_;
assign _080_ = _046_ == { _023_[1], 1'h0 };
assign _081_ = _037_ == _018_;
assign _007_ = _080_ & _030_;
assign _087_ = _081_ & _034_;
/* src = "generated/sv2v_out.v:286.2-306.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_b656ed3944a4d79ba92b  */
/* PC_TAINT_INFO STATE_NAME count_low */
always_ff @(posedge clk)
if (!rstz) count_low <= 32'd0;
else if (_010_) count_low <= _096_;
/* src = "generated/sv2v_out.v:286.2-306.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_b656ed3944a4d79ba92b  */
/* PC_TAINT_INFO STATE_NAME count_high */
always_ff @(posedge clk)
if (!rstz) count_high <= 32'd0;
else if (_012_) count_high <= _090_;
/* src = "generated/sv2v_out.v:286.2-306.6" */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_b656ed3944a4d79ba92b  */
/* PC_TAINT_INFO STATE_NAME incr_high */
always_ff @(posedge clk)
if (_014_) incr_high <= 1'h0;
else incr_high <= _086_;
assign _031_ = | { count_vld_t0, load_high_t0 };
assign _029_ = | { load_low_t0, load_high_t0, incr_t0 };
assign _022_ = ~ { load_high_t0, load_low_t0, incr_t0 };
assign _024_ = ~ { count_vld_t0, load_high_t0 };
assign _045_ = { load_high, load_low, incr } & _022_;
assign _047_ = { incr_high, load_high } & _024_;
assign _035_ = ! _045_;
assign _036_ = ! _047_;
assign _005_ = _035_ & _029_;
assign _009_ = _036_ & _031_;
assign _025_ = ~ { load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high };
assign _026_ = ~ { load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low };
assign _067_ = { load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0 } | _025_;
assign _071_ = { load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0 } | _026_;
assign _066_ = { count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0, count_vld_t0 } | { incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high, incr_high };
assign _068_ = { load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0 } | { load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high, load_high };
assign _070_ = { incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0, incr_t0 } | { incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr, incr };
assign _072_ = { load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0 } | { load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low, load_low };
assign _048_ = _089_ & _067_;
assign _095_ = _093_ & _067_;
assign _051_ = _095_ & _071_;
assign _089_ = _003_ & _066_;
assign _049_ = load_data_t0 & _068_;
assign _093_ = _001_ & _070_;
assign _052_ = load_data_t0 & _072_;
assign _069_ = _048_ | _049_;
assign _073_ = _051_ | _052_;
assign _078_ = _088_ ^ load_data;
assign _079_ = _094_ ^ load_data;
assign _050_ = { load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0, load_high_t0 } & _078_;
assign _053_ = { load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0, load_low_t0 } & _079_;
assign _091_ = _050_ | _069_;
assign _097_ = _053_ | _073_;
assign _004_ = | { load_high, load_low, incr };
assign _006_ = { load_high, load_low } != 2'h2;
assign _008_ = | { incr_high, load_high };
assign _015_ = ~ load_low;
assign _010_ = & { _004_, _006_ };
assign _012_ = & { _008_, _015_ };
assign _016_ = ~ incr;
assign _017_ = ~ rstz;
assign _014_ = | { _017_, _016_, load_high, load_low };
assign _032_ = | { _005_, _007_ };
assign _033_ = | { _009_, load_low_t0 };
assign _064_ = { _004_, _006_ } | { _005_, _007_ };
assign _065_ = { _008_, _015_ } | { _009_, load_low_t0 };
assign _027_ = & _064_;
assign _028_ = & _065_;
assign _011_ = _032_ & _027_;
assign _013_ = _033_ & _028_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_b656ed3944a4d79ba92b  */
/* PC_TAINT_INFO STATE_NAME count_vld_t0 */
always_ff @(posedge clk)
if (_014_) count_vld_t0 <= 1'h0;
else count_vld_t0 <= _087_;
assign _020_ = ~ _010_;
assign _021_ = ~ _012_;
assign _076_ = _096_ ^ count_low;
assign _077_ = _090_ ^ count_high;
assign _056_ = _097_ | count_low_t0;
assign _060_ = _091_ | count_high_t0;
assign _057_ = _076_ | _056_;
assign _061_ = _077_ | _060_;
assign _039_ = { _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_ } & _097_;
assign _042_ = { _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_, _012_ } & _091_;
assign _040_ = { _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_ } & count_low_t0;
assign _043_ = { _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_, _021_ } & count_high_t0;
assign _041_ = _057_ & { _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_ };
assign _044_ = _061_ & { _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_, _013_ };
assign _058_ = _039_ | _040_;
assign _062_ = _042_ | _043_;
assign _059_ = _058_ | _041_;
assign _063_ = _062_ | _044_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_b656ed3944a4d79ba92b  */
/* PC_TAINT_INFO STATE_NAME count_low_t0 */
always_ff @(posedge clk)
if (!rstz) count_low_t0 <= 32'd0;
else count_low_t0 <= _059_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME paramodsimplif_b656ed3944a4d79ba92b  */
/* PC_TAINT_INFO STATE_NAME count_high_t0 */
always_ff @(posedge clk)
if (!rstz) count_high_t0 <= 32'd0;
else count_high_t0 <= _063_;
assign _086_ = count_low == /* src = "generated/sv2v_out.v:301.19-301.44" */ 32'd4294967295;
assign count_vld = ~ /* src = "generated/sv2v_out.v:311.24-311.34" */ incr_high;
assign _088_ = incr_high ? /* src = "generated/sv2v_out.v:303.9-303.18|generated/sv2v_out.v:303.5-304.38" */ _002_ : 32'hxxxxxxxx;
assign _090_ = load_high ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:296.13-296.22|generated/sv2v_out.v:296.9-305.7" */ load_data : _088_;
assign _092_ = incr ? /* src = "generated/sv2v_out.v:299.9-299.13|generated/sv2v_out.v:299.5-302.8" */ _000_ : 32'hxxxxxxxx;
assign _094_ = load_high ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:296.13-296.22|generated/sv2v_out.v:296.9-305.7" */ 32'hxxxxxxxx : _092_;
assign _096_ = load_low ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:294.8-294.16|generated/sv2v_out.v:294.4-305.7" */ load_data : _094_;
assign count = { count_high, count_low };
assign count_t0 = { count_high_t0, count_low_t0 };
// Added block to randomize initial values.
`ifdef RANDOMIZE_INIT
  initial begin
    count_low = '0;
    count_high = '0;
    incr_high = '0;
    count_vld_t0 = '0;
    count_low_t0 = '0;
    count_high_t0 = '0;
  end
`endif // RANDOMIZE_INIT
endmodule

module kronos_RF(clk, rstz, instr_data, instr_vld, fetch_rdy, immediate, regrd_rs1, regrd_rs2, regrd_rs1_en, regrd_rs2_en, regwr_data, regwr_sel, regwr_en, clk_t0, regwr_data_t0, regwr_en_t0, regwr_sel_t0, instr_vld_t0, fetch_rdy_t0, immediate_t0, instr_data_t0
, regrd_rs1_t0, regrd_rs1_en_t0, regrd_rs2_t0, regrd_rs2_en_t0);
/* src = "generated/sv2v_out.v:1627.2-1629.33" */
wire [4:0] _0000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1627.2-1629.33" */
wire [4:0] _0001_;
/* src = "generated/sv2v_out.v:1627.2-1629.33" */
wire [31:0] _0002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1627.2-1629.33" */
wire [31:0] _0003_;
/* src = "generated/sv2v_out.v:1627.2-1629.33" */
wire [31:0] _0004_;
/* src = "generated/sv2v_out.v:1549.2-1587.5" */
wire _0005_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1549.2-1587.5" */
wire _0006_;
/* src = "generated/sv2v_out.v:1549.2-1587.5" */
wire [3:0] _0007_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1549.2-1587.5" */
wire [3:0] _0008_;
/* src = "generated/sv2v_out.v:1549.2-1587.5" */
wire _0009_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1549.2-1587.5" */
wire _0010_;
/* src = "generated/sv2v_out.v:1549.2-1587.5" */
wire _0011_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1549.2-1587.5" */
wire _0012_;
wire _0013_;
/* cellift = 32'd1 */
wire _0014_;
wire _0015_;
/* cellift = 32'd1 */
wire _0016_;
wire _0017_;
/* cellift = 32'd1 */
wire _0018_;
wire _0019_;
/* cellift = 32'd1 */
wire _0020_;
wire _0021_;
/* cellift = 32'd1 */
wire _0022_;
wire _0023_;
/* cellift = 32'd1 */
wire _0024_;
wire _0025_;
/* cellift = 32'd1 */
wire _0026_;
wire _0027_;
/* cellift = 32'd1 */
wire _0028_;
wire _0029_;
/* cellift = 32'd1 */
wire _0030_;
wire [1:0] _0031_;
wire [2:0] _0032_;
wire [2:0] _0033_;
wire [2:0] _0034_;
wire [4:0] _0035_;
wire [2:0] _0036_;
wire [4:0] _0037_;
wire [4:0] _0038_;
wire [4:0] _0039_;
wire [4:0] _0040_;
wire [4:0] _0041_;
wire [4:0] _0042_;
wire _0043_;
wire _0044_;
wire _0045_;
wire _0046_;
wire _0047_;
wire _0048_;
wire _0049_;
wire _0050_;
wire _0051_;
wire _0052_;
wire _0053_;
wire _0054_;
wire _0055_;
wire _0056_;
wire _0057_;
wire _0058_;
wire _0059_;
wire _0060_;
wire _0061_;
wire _0062_;
wire _0063_;
wire _0064_;
wire _0065_;
wire [31:0] _0066_;
wire [31:0] _0067_;
wire [31:0] _0068_;
wire [31:0] _0069_;
wire [31:0] _0070_;
wire [31:0] _0071_;
wire [31:0] _0072_;
wire [31:0] _0073_;
wire [31:0] _0074_;
wire [31:0] _0075_;
wire _0076_;
wire [31:0] _0077_;
wire [31:0] _0078_;
wire [31:0] _0079_;
wire [31:0] _0080_;
wire [31:0] _0081_;
wire [11:0] _0082_;
wire [7:0] _0083_;
wire [3:0] _0084_;
wire _0085_;
wire _0086_;
wire _0087_;
wire _0088_;
wire _0089_;
wire _0090_;
wire _0091_;
wire _0092_;
wire _0093_;
wire _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire _0109_;
wire _0110_;
wire _0111_;
wire _0112_;
wire _0113_;
wire _0114_;
wire _0115_;
wire _0116_;
wire _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire _0139_;
wire _0140_;
wire _0141_;
wire _0142_;
wire _0143_;
wire _0144_;
wire _0145_;
wire _0146_;
wire _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
wire _0152_;
wire _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire _0186_;
wire _0187_;
wire _0188_;
wire _0189_;
wire _0190_;
wire _0191_;
wire _0192_;
wire _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire _0199_;
wire _0200_;
wire _0201_;
wire _0202_;
wire _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
wire _0221_;
wire _0222_;
wire _0223_;
wire _0224_;
wire _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire _0241_;
wire _0242_;
wire _0243_;
wire _0244_;
wire [1:0] _0245_;
wire [2:0] _0246_;
wire [2:0] _0247_;
wire [2:0] _0248_;
wire [4:0] _0249_;
wire [2:0] _0250_;
wire [4:0] _0251_;
wire [4:0] _0252_;
wire [4:0] _0253_;
wire [4:0] _0254_;
wire [4:0] _0255_;
wire [4:0] _0256_;
wire [4:0] _0257_;
wire [4:0] _0258_;
wire [4:0] _0259_;
wire [4:0] _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire _0271_;
wire _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire _0276_;
wire _0277_;
wire _0278_;
wire _0279_;
wire _0280_;
wire _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire _0285_;
wire _0286_;
wire _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire _0294_;
wire _0295_;
wire _0296_;
wire _0297_;
wire _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire [31:0] _0324_;
wire [31:0] _0325_;
wire [31:0] _0326_;
wire [31:0] _0327_;
wire [31:0] _0328_;
wire [31:0] _0329_;
wire [31:0] _0330_;
wire [31:0] _0331_;
wire [31:0] _0332_;
wire [31:0] _0333_;
wire [31:0] _0334_;
wire [31:0] _0335_;
wire [31:0] _0336_;
wire [31:0] _0337_;
wire [31:0] _0338_;
wire [31:0] _0339_;
wire [31:0] _0340_;
wire [31:0] _0341_;
wire [31:0] _0342_;
wire [31:0] _0343_;
wire [31:0] _0344_;
wire [31:0] _0345_;
wire [31:0] _0346_;
wire [31:0] _0347_;
wire [31:0] _0348_;
wire [31:0] _0349_;
wire [31:0] _0350_;
wire [31:0] _0351_;
wire [31:0] _0352_;
wire [31:0] _0353_;
wire [31:0] _0354_;
wire [31:0] _0355_;
wire [31:0] _0356_;
wire [31:0] _0357_;
wire [31:0] _0358_;
wire [31:0] _0359_;
wire [31:0] _0360_;
wire [31:0] _0361_;
wire [31:0] _0362_;
wire [31:0] _0363_;
wire [31:0] _0364_;
wire [31:0] _0365_;
wire [31:0] _0366_;
wire [31:0] _0367_;
wire [31:0] _0368_;
wire [31:0] _0369_;
wire [31:0] _0370_;
wire [31:0] _0371_;
wire [31:0] _0372_;
wire [31:0] _0373_;
wire [31:0] _0374_;
wire [31:0] _0375_;
wire [31:0] _0376_;
wire [31:0] _0377_;
wire [31:0] _0378_;
wire [31:0] _0379_;
wire [31:0] _0380_;
wire [31:0] _0381_;
wire [31:0] _0382_;
wire [31:0] _0383_;
wire [31:0] _0384_;
wire [31:0] _0385_;
wire [31:0] _0386_;
wire [31:0] _0387_;
wire [31:0] _0388_;
wire [31:0] _0389_;
wire [31:0] _0390_;
wire [31:0] _0391_;
wire [31:0] _0392_;
wire [31:0] _0393_;
wire [31:0] _0394_;
wire [31:0] _0395_;
wire [31:0] _0396_;
wire [31:0] _0397_;
wire [31:0] _0398_;
wire [31:0] _0399_;
wire [31:0] _0400_;
wire [31:0] _0401_;
wire [31:0] _0402_;
wire [31:0] _0403_;
wire [31:0] _0404_;
wire [31:0] _0405_;
wire [31:0] _0406_;
wire [31:0] _0407_;
wire [31:0] _0408_;
wire [31:0] _0409_;
wire [31:0] _0410_;
wire [31:0] _0411_;
wire [31:0] _0412_;
wire [31:0] _0413_;
wire [31:0] _0414_;
wire [31:0] _0415_;
wire [31:0] _0416_;
wire [31:0] _0417_;
wire [31:0] _0418_;
wire [31:0] _0419_;
wire [31:0] _0420_;
wire [31:0] _0421_;
wire [31:0] _0422_;
wire [31:0] _0423_;
wire [31:0] _0424_;
wire [31:0] _0425_;
wire [31:0] _0426_;
wire [31:0] _0427_;
wire [31:0] _0428_;
wire [31:0] _0429_;
wire [31:0] _0430_;
wire [31:0] _0431_;
wire [31:0] _0432_;
wire [31:0] _0433_;
wire [31:0] _0434_;
wire [31:0] _0435_;
wire [31:0] _0436_;
wire [31:0] _0437_;
wire [31:0] _0438_;
wire [31:0] _0439_;
wire [31:0] _0440_;
wire [31:0] _0441_;
wire [31:0] _0442_;
wire [31:0] _0443_;
wire [31:0] _0444_;
wire [31:0] _0445_;
wire [31:0] _0446_;
wire [31:0] _0447_;
wire [31:0] _0448_;
wire [31:0] _0449_;
wire [31:0] _0450_;
wire [31:0] _0451_;
wire [31:0] _0452_;
wire [31:0] _0453_;
wire [31:0] _0454_;
wire [31:0] _0455_;
wire [31:0] _0456_;
wire [31:0] _0457_;
wire [31:0] _0458_;
wire [31:0] _0459_;
wire [31:0] _0460_;
wire [31:0] _0461_;
wire [31:0] _0462_;
wire [31:0] _0463_;
wire [31:0] _0464_;
wire [31:0] _0465_;
wire [31:0] _0466_;
wire [31:0] _0467_;
wire [31:0] _0468_;
wire [31:0] _0469_;
wire [31:0] _0470_;
wire [31:0] _0471_;
wire [31:0] _0472_;
wire [31:0] _0473_;
wire [31:0] _0474_;
wire [31:0] _0475_;
wire [31:0] _0476_;
wire [31:0] _0477_;
wire [31:0] _0478_;
wire [31:0] _0479_;
wire [31:0] _0480_;
wire [31:0] _0481_;
wire [31:0] _0482_;
wire [31:0] _0483_;
wire [31:0] _0484_;
wire [31:0] _0485_;
wire [31:0] _0486_;
wire [31:0] _0487_;
wire [31:0] _0488_;
wire [31:0] _0489_;
wire [31:0] _0490_;
wire [31:0] _0491_;
wire [31:0] _0492_;
wire [31:0] _0493_;
wire [31:0] _0494_;
wire [31:0] _0495_;
wire [31:0] _0496_;
wire [31:0] _0497_;
wire [31:0] _0498_;
wire [31:0] _0499_;
wire [31:0] _0500_;
wire [31:0] _0501_;
wire [31:0] _0502_;
wire [31:0] _0503_;
wire [31:0] _0504_;
wire [31:0] _0505_;
wire [31:0] _0506_;
wire [31:0] _0507_;
wire [31:0] _0508_;
wire [31:0] _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0517_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
wire _0525_;
wire _0526_;
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire _0534_;
wire _0535_;
wire _0536_;
wire _0537_;
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0542_;
wire _0543_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire _0560_;
wire _0561_;
wire _0562_;
wire _0563_;
wire _0564_;
wire _0565_;
wire _0566_;
wire _0567_;
wire _0568_;
wire _0569_;
wire _0570_;
wire _0571_;
wire _0572_;
wire _0573_;
wire _0574_;
wire _0575_;
wire _0576_;
wire _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire _0596_;
wire _0597_;
wire _0598_;
wire _0599_;
wire _0600_;
wire _0601_;
wire _0602_;
wire _0603_;
wire _0604_;
wire _0605_;
wire _0606_;
wire [31:0] _0607_;
wire [31:0] _0608_;
wire [31:0] _0609_;
wire [31:0] _0610_;
wire [31:0] _0611_;
wire [31:0] _0612_;
wire [31:0] _0613_;
wire [31:0] _0614_;
wire [31:0] _0615_;
wire [31:0] _0616_;
wire [31:0] _0617_;
wire [31:0] _0618_;
wire [31:0] _0619_;
wire [31:0] _0620_;
wire [31:0] _0621_;
wire [31:0] _0622_;
wire [11:0] _0623_;
wire [11:0] _0624_;
wire [11:0] _0625_;
wire [7:0] _0626_;
wire [7:0] _0627_;
wire [7:0] _0628_;
wire _0629_;
wire _0630_;
wire _0631_;
wire _0632_;
wire _0633_;
wire _0634_;
wire [3:0] _0635_;
wire [3:0] _0636_;
wire [3:0] _0637_;
wire _0638_;
wire _0639_;
wire _0640_;
wire _0641_;
wire _0642_;
wire _0643_;
/* cellift = 32'd1 */
wire _0644_;
wire _0645_;
/* cellift = 32'd1 */
wire _0646_;
wire _0647_;
/* cellift = 32'd1 */
wire _0648_;
wire _0649_;
/* cellift = 32'd1 */
wire _0650_;
wire _0651_;
/* cellift = 32'd1 */
wire _0652_;
wire _0653_;
/* cellift = 32'd1 */
wire _0654_;
wire _0655_;
/* cellift = 32'd1 */
wire _0656_;
wire _0657_;
/* cellift = 32'd1 */
wire _0658_;
wire _0659_;
/* cellift = 32'd1 */
wire _0660_;
wire _0661_;
/* cellift = 32'd1 */
wire _0662_;
wire _0663_;
/* cellift = 32'd1 */
wire _0664_;
wire _0665_;
/* cellift = 32'd1 */
wire _0666_;
wire _0667_;
/* cellift = 32'd1 */
wire _0668_;
wire _0669_;
/* cellift = 32'd1 */
wire _0670_;
wire _0671_;
/* cellift = 32'd1 */
wire _0672_;
wire _0673_;
/* cellift = 32'd1 */
wire _0674_;
wire _0675_;
/* cellift = 32'd1 */
wire _0676_;
wire _0677_;
/* cellift = 32'd1 */
wire _0678_;
wire _0679_;
/* cellift = 32'd1 */
wire _0680_;
wire _0681_;
/* cellift = 32'd1 */
wire _0682_;
wire _0683_;
/* cellift = 32'd1 */
wire _0684_;
wire _0685_;
/* cellift = 32'd1 */
wire _0686_;
wire _0687_;
/* cellift = 32'd1 */
wire _0688_;
wire _0689_;
/* cellift = 32'd1 */
wire _0690_;
wire _0691_;
/* cellift = 32'd1 */
wire _0692_;
wire _0693_;
/* cellift = 32'd1 */
wire _0694_;
wire _0695_;
/* cellift = 32'd1 */
wire _0696_;
wire _0697_;
/* cellift = 32'd1 */
wire _0698_;
wire _0699_;
/* cellift = 32'd1 */
wire _0700_;
wire _0701_;
/* cellift = 32'd1 */
wire _0702_;
wire _0703_;
/* cellift = 32'd1 */
wire _0704_;
wire _0705_;
/* cellift = 32'd1 */
wire _0706_;
wire _0707_;
/* cellift = 32'd1 */
wire _0708_;
wire _0709_;
/* cellift = 32'd1 */
wire _0710_;
wire _0711_;
/* cellift = 32'd1 */
wire _0712_;
wire _0713_;
/* cellift = 32'd1 */
wire _0714_;
wire _0715_;
/* cellift = 32'd1 */
wire _0716_;
wire _0717_;
/* cellift = 32'd1 */
wire _0718_;
wire _0719_;
/* cellift = 32'd1 */
wire _0720_;
wire _0721_;
/* cellift = 32'd1 */
wire _0722_;
wire _0723_;
/* cellift = 32'd1 */
wire _0724_;
wire _0725_;
/* cellift = 32'd1 */
wire _0726_;
wire _0727_;
/* cellift = 32'd1 */
wire _0728_;
wire _0729_;
/* cellift = 32'd1 */
wire _0730_;
wire _0731_;
/* cellift = 32'd1 */
wire _0732_;
wire _0733_;
/* cellift = 32'd1 */
wire _0734_;
wire _0735_;
/* cellift = 32'd1 */
wire _0736_;
wire _0737_;
/* cellift = 32'd1 */
wire _0738_;
wire [31:0] _0739_;
wire [31:0] _0740_;
wire [31:0] _0741_;
wire [31:0] _0742_;
wire [31:0] _0743_;
wire [31:0] _0744_;
wire _0745_;
wire _0746_;
wire _0747_;
wire _0748_;
wire _0749_;
wire _0750_;
wire _0751_;
wire _0752_;
wire _0753_;
wire [4:0] _0754_;
wire [4:0] _0755_;
wire [4:0] _0756_;
wire [4:0] _0757_;
wire [4:0] _0758_;
wire [4:0] _0759_;
wire [10:0] _0760_;
wire [10:0] _0761_;
wire [10:0] _0762_;
wire [20:0] _0763_;
wire [20:0] _0764_;
wire [20:0] _0765_;
wire [31:0] _0766_;
wire [31:0] _0767_;
wire [31:0] _0768_;
wire [31:0] _0769_;
wire [31:0] _0770_;
wire [31:0] _0771_;
wire [31:0] _0772_;
wire [31:0] _0773_;
wire [31:0] _0774_;
wire [31:0] _0775_;
wire [31:0] _0776_;
wire [31:0] _0777_;
wire [31:0] _0778_;
wire [31:0] _0779_;
wire [31:0] _0780_;
wire [31:0] _0781_;
wire [31:0] _0782_;
wire [31:0] _0783_;
wire [31:0] _0784_;
wire [31:0] _0785_;
wire [31:0] _0786_;
wire [31:0] _0787_;
wire [31:0] _0788_;
wire [31:0] _0789_;
wire [31:0] _0790_;
wire [31:0] _0791_;
wire [31:0] _0792_;
wire [31:0] _0793_;
wire [31:0] _0794_;
wire [31:0] _0795_;
wire [31:0] _0796_;
wire [31:0] _0797_;
wire [31:0] _0798_;
wire [31:0] _0799_;
wire [31:0] _0800_;
wire [31:0] _0801_;
wire [31:0] _0802_;
wire [31:0] _0803_;
wire [31:0] _0804_;
wire [31:0] _0805_;
wire [31:0] _0806_;
wire [31:0] _0807_;
wire [31:0] _0808_;
wire [31:0] _0809_;
wire [31:0] _0810_;
wire [31:0] _0811_;
wire [31:0] _0812_;
wire [31:0] _0813_;
wire [31:0] _0814_;
wire [31:0] _0815_;
wire [31:0] _0816_;
wire [31:0] _0817_;
wire [31:0] _0818_;
wire [31:0] _0819_;
wire [31:0] _0820_;
wire [31:0] _0821_;
wire [31:0] _0822_;
wire [31:0] _0823_;
wire [31:0] _0824_;
wire [31:0] _0825_;
wire [31:0] _0826_;
wire [31:0] _0827_;
wire [31:0] _0828_;
wire [31:0] _0829_;
wire [31:0] _0830_;
wire [31:0] _0831_;
wire [31:0] _0832_;
wire [31:0] _0833_;
wire [31:0] _0834_;
wire [31:0] _0835_;
wire [31:0] _0836_;
wire [31:0] _0837_;
wire [31:0] _0838_;
wire [31:0] _0839_;
wire [31:0] _0840_;
wire [31:0] _0841_;
wire [31:0] _0842_;
wire [31:0] _0843_;
wire [31:0] _0844_;
wire [31:0] _0845_;
wire [31:0] _0846_;
wire [31:0] _0847_;
wire [31:0] _0848_;
wire [31:0] _0849_;
wire [31:0] _0850_;
wire [31:0] _0851_;
wire [31:0] _0852_;
wire [31:0] _0853_;
wire [31:0] _0854_;
wire [31:0] _0855_;
wire [31:0] _0856_;
wire [31:0] _0857_;
wire [31:0] _0858_;
wire [31:0] _0859_;
wire [31:0] _0860_;
wire [31:0] _0861_;
wire _0862_;
wire _0863_;
wire _0864_;
wire _0865_;
wire _0866_;
wire _0867_;
wire _0868_;
wire _0869_;
wire _0870_;
wire _0871_;
wire _0872_;
wire _0873_;
wire _0874_;
wire _0875_;
wire _0876_;
wire _0877_;
wire _0878_;
wire _0879_;
wire _0880_;
wire _0881_;
wire _0882_;
wire _0883_;
wire _0884_;
wire _0885_;
wire _0886_;
wire _0887_;
wire _0888_;
wire _0889_;
wire _0890_;
wire _0891_;
wire _0892_;
wire _0893_;
wire _0894_;
wire _0895_;
wire _0896_;
wire _0897_;
wire _0898_;
wire _0899_;
wire _0900_;
wire _0901_;
wire _0902_;
wire _0903_;
wire _0904_;
wire _0905_;
wire _0906_;
wire _0907_;
wire _0908_;
wire _0909_;
wire _0910_;
wire _0911_;
wire _0912_;
wire _0913_;
wire _0914_;
wire _0915_;
wire _0916_;
wire _0917_;
wire _0918_;
wire _0919_;
wire _0920_;
wire _0921_;
wire [2:0] _0922_;
wire [2:0] _0923_;
wire [1:0] _0924_;
wire [1:0] _0925_;
wire [4:0] _0926_;
wire [4:0] _0927_;
wire [4:0] _0928_;
wire [4:0] _0929_;
wire _0930_;
wire _0931_;
wire _0932_;
wire _0933_;
wire _0934_;
wire _0935_;
wire _0936_;
wire _0937_;
wire _0938_;
wire _0939_;
wire _0940_;
wire _0941_;
wire _0942_;
wire _0943_;
wire _0944_;
wire _0945_;
wire _0946_;
wire _0947_;
wire _0948_;
wire _0949_;
wire _0950_;
wire [31:0] _0951_;
wire [31:0] _0952_;
wire [31:0] _0953_;
wire [31:0] _0954_;
wire [31:0] _0955_;
wire [31:0] _0956_;
wire [31:0] _0957_;
wire [31:0] _0958_;
wire [31:0] _0959_;
wire [31:0] _0960_;
wire [31:0] _0961_;
wire [31:0] _0962_;
wire [31:0] _0963_;
wire [31:0] _0964_;
wire [31:0] _0965_;
wire [31:0] _0966_;
wire [31:0] _0967_;
wire [31:0] _0968_;
wire [31:0] _0969_;
wire [31:0] _0970_;
wire [31:0] _0971_;
wire [31:0] _0972_;
wire [31:0] _0973_;
wire [31:0] _0974_;
wire [31:0] _0975_;
wire [31:0] _0976_;
wire [31:0] _0977_;
wire [31:0] _0978_;
wire [31:0] _0979_;
wire [31:0] _0980_;
wire [31:0] _0981_;
wire [31:0] _0982_;
wire [31:0] _0983_;
wire [31:0] _0984_;
wire [31:0] _0985_;
wire [31:0] _0986_;
wire [31:0] _0987_;
wire [31:0] _0988_;
wire [31:0] _0989_;
wire [31:0] _0990_;
wire [31:0] _0991_;
wire [31:0] _0992_;
wire [31:0] _0993_;
wire [31:0] _0994_;
wire [31:0] _0995_;
wire [31:0] _0996_;
wire [31:0] _0997_;
wire [31:0] _0998_;
wire [31:0] _0999_;
wire [31:0] _1000_;
wire [31:0] _1001_;
wire [31:0] _1002_;
wire [31:0] _1003_;
wire [31:0] _1004_;
wire [31:0] _1005_;
wire [31:0] _1006_;
wire [31:0] _1007_;
wire [31:0] _1008_;
wire [31:0] _1009_;
wire [31:0] _1010_;
wire [31:0] _1011_;
wire [31:0] _1012_;
wire [31:0] _1013_;
wire [31:0] _1014_;
wire [31:0] _1015_;
wire [31:0] _1016_;
wire [31:0] _1017_;
wire [31:0] _1018_;
wire [31:0] _1019_;
wire [31:0] _1020_;
wire [31:0] _1021_;
wire [31:0] _1022_;
wire [31:0] _1023_;
wire [31:0] _1024_;
wire [31:0] _1025_;
wire [31:0] _1026_;
wire [31:0] _1027_;
wire [31:0] _1028_;
wire [31:0] _1029_;
wire [31:0] _1030_;
wire [31:0] _1031_;
wire [31:0] _1032_;
wire _1033_;
wire _1034_;
wire _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire _1046_;
wire _1047_;
wire _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1052_;
wire _1053_;
wire _1054_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire _1061_;
wire _1062_;
wire _1063_;
wire _1064_;
wire _1065_;
wire [31:0] _1066_;
wire [4:0] _1067_;
wire [31:0] _1068_;
wire [31:0] _1069_;
wire [31:0] _1070_;
wire [31:0] _1071_;
wire [31:0] _1072_;
wire [31:0] _1073_;
wire [31:0] _1074_;
wire [31:0] _1075_;
wire [31:0] _1076_;
wire [31:0] _1077_;
wire [31:0] _1078_;
wire [31:0] _1079_;
wire [31:0] _1080_;
wire [31:0] _1081_;
wire [31:0] _1082_;
wire [11:0] _1083_;
wire [11:0] _1084_;
wire [11:0] _1085_;
wire [7:0] _1086_;
wire [7:0] _1087_;
wire [7:0] _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire [3:0] _1095_;
wire [3:0] _1096_;
wire [3:0] _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire [31:0] _1102_;
wire [31:0] _1103_;
wire [31:0] _1104_;
wire [31:0] _1105_;
wire [31:0] _1106_;
wire [31:0] _1107_;
wire [31:0] _1108_;
wire [31:0] _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire [4:0] _1122_;
wire [4:0] _1123_;
wire [4:0] _1124_;
wire [4:0] _1125_;
wire [4:0] _1126_;
wire [4:0] _1127_;
wire [4:0] _1128_;
wire [4:0] _1129_;
wire [10:0] _1130_;
wire [10:0] _1131_;
wire [10:0] _1132_;
wire [10:0] _1133_;
wire [20:0] _1134_;
wire [20:0] _1135_;
wire [20:0] _1136_;
wire [20:0] _1137_;
wire [31:0] _1138_;
wire [31:0] _1139_;
wire [31:0] _1140_;
wire [31:0] _1141_;
wire [31:0] _1142_;
wire [31:0] _1143_;
wire [31:0] _1144_;
wire [31:0] _1145_;
wire [31:0] _1146_;
wire [31:0] _1147_;
wire [31:0] _1148_;
wire [31:0] _1149_;
wire [31:0] _1150_;
wire [31:0] _1151_;
wire [31:0] _1152_;
wire [31:0] _1153_;
wire [31:0] _1154_;
wire [31:0] _1155_;
wire [31:0] _1156_;
wire [31:0] _1157_;
wire [31:0] _1158_;
wire [31:0] _1159_;
wire [31:0] _1160_;
wire [31:0] _1161_;
wire [31:0] _1162_;
wire [31:0] _1163_;
wire [31:0] _1164_;
wire [31:0] _1165_;
wire [31:0] _1166_;
wire [31:0] _1167_;
wire [31:0] _1168_;
wire [31:0] _1169_;
wire [31:0] _1170_;
wire [31:0] _1171_;
wire [31:0] _1172_;
wire [31:0] _1173_;
wire [31:0] _1174_;
wire [31:0] _1175_;
wire [31:0] _1176_;
wire [31:0] _1177_;
wire [31:0] _1178_;
wire [31:0] _1179_;
wire [31:0] _1180_;
wire [31:0] _1181_;
wire [31:0] _1182_;
wire [31:0] _1183_;
wire [31:0] _1184_;
wire [31:0] _1185_;
wire [31:0] _1186_;
wire [31:0] _1187_;
wire [31:0] _1188_;
wire [31:0] _1189_;
wire [31:0] _1190_;
wire [31:0] _1191_;
wire [31:0] _1192_;
wire [31:0] _1193_;
wire [31:0] _1194_;
wire [31:0] _1195_;
wire [31:0] _1196_;
wire [31:0] _1197_;
wire [31:0] _1198_;
wire [31:0] _1199_;
wire [31:0] _1200_;
wire [31:0] _1201_;
wire [31:0] _1202_;
wire [31:0] _1203_;
wire [31:0] _1204_;
wire [31:0] _1205_;
wire [31:0] _1206_;
wire [31:0] _1207_;
wire [31:0] _1208_;
wire [31:0] _1209_;
wire [31:0] _1210_;
wire [31:0] _1211_;
wire [31:0] _1212_;
wire [31:0] _1213_;
wire [31:0] _1214_;
wire [31:0] _1215_;
wire [31:0] _1216_;
wire [31:0] _1217_;
wire [31:0] _1218_;
wire [31:0] _1219_;
wire [31:0] _1220_;
wire [31:0] _1221_;
wire [31:0] _1222_;
wire [31:0] _1223_;
wire [31:0] _1224_;
wire [31:0] _1225_;
wire [31:0] _1226_;
wire [31:0] _1227_;
wire [31:0] _1228_;
wire [31:0] _1229_;
wire [31:0] _1230_;
wire [31:0] _1231_;
wire [31:0] _1232_;
wire [31:0] _1233_;
wire [31:0] _1234_;
wire [31:0] _1235_;
wire [31:0] _1236_;
wire [31:0] _1237_;
wire [31:0] _1238_;
wire [31:0] _1239_;
wire [31:0] _1240_;
wire [31:0] _1241_;
wire [31:0] _1242_;
wire [31:0] _1243_;
wire [31:0] _1244_;
wire [31:0] _1245_;
wire [31:0] _1246_;
wire [31:0] _1247_;
wire [31:0] _1248_;
wire [31:0] _1249_;
wire [31:0] _1250_;
wire [31:0] _1251_;
wire [31:0] _1252_;
wire [31:0] _1253_;
wire [31:0] _1254_;
wire [31:0] _1255_;
wire [31:0] _1256_;
wire [31:0] _1257_;
wire [31:0] _1258_;
wire [31:0] _1259_;
wire [31:0] _1260_;
wire [31:0] _1261_;
wire [31:0] _1262_;
wire [31:0] _1263_;
wire [31:0] _1264_;
wire [31:0] _1265_;
wire _1266_;
wire _1267_;
wire _1268_;
wire _1269_;
wire _1270_;
wire _1271_;
wire _1272_;
wire _1273_;
wire _1274_;
wire _1275_;
wire _1276_;
wire [31:0] _1277_;
wire [31:0] _1278_;
wire [31:0] _1279_;
wire [31:0] _1280_;
wire [31:0] _1281_;
wire [31:0] _1282_;
wire [31:0] _1283_;
wire [31:0] _1284_;
wire [31:0] _1285_;
wire [31:0] _1286_;
wire [31:0] _1287_;
wire [31:0] _1288_;
wire [31:0] _1289_;
wire [31:0] _1290_;
wire [31:0] _1291_;
wire [31:0] _1292_;
wire [31:0] _1293_;
wire [31:0] _1294_;
wire [31:0] _1295_;
wire [31:0] _1296_;
wire [31:0] _1297_;
wire [31:0] _1298_;
wire [31:0] _1299_;
wire [31:0] _1300_;
wire [31:0] _1301_;
wire [31:0] _1302_;
wire [31:0] _1303_;
wire [31:0] _1304_;
wire [31:0] _1305_;
wire [31:0] _1306_;
wire [31:0] _1307_;
wire [31:0] _1308_;
wire [31:0] _1309_;
wire [31:0] _1310_;
wire [31:0] _1311_;
wire [31:0] _1312_;
wire [31:0] _1313_;
wire [31:0] _1314_;
wire [31:0] _1315_;
wire [31:0] _1316_;
wire [31:0] _1317_;
wire [31:0] _1318_;
wire [31:0] _1319_;
wire [31:0] _1320_;
wire [31:0] _1321_;
wire [31:0] _1322_;
wire [31:0] _1323_;
wire [31:0] _1324_;
wire [31:0] _1325_;
wire [31:0] _1326_;
wire [31:0] _1327_;
wire [31:0] _1328_;
wire [11:0] _1329_;
wire [7:0] _1330_;
wire _1331_;
wire _1332_;
wire [3:0] _1333_;
wire _1334_;
wire [31:0] _1335_;
wire [31:0] _1336_;
wire _1337_;
wire _1338_;
wire _1339_;
wire [4:0] _1340_;
wire [4:0] _1341_;
wire [10:0] _1342_;
wire [20:0] _1343_;
wire [31:0] _1344_;
wire [31:0] _1345_;
wire [31:0] _1346_;
wire [31:0] _1347_;
wire [31:0] _1348_;
wire [31:0] _1349_;
wire [31:0] _1350_;
wire [31:0] _1351_;
wire [31:0] _1352_;
wire [31:0] _1353_;
wire [31:0] _1354_;
wire [31:0] _1355_;
wire [31:0] _1356_;
wire [31:0] _1357_;
wire [31:0] _1358_;
wire [31:0] _1359_;
wire [31:0] _1360_;
wire [31:0] _1361_;
wire [31:0] _1362_;
wire [31:0] _1363_;
wire [31:0] _1364_;
wire [31:0] _1365_;
wire [31:0] _1366_;
wire [31:0] _1367_;
wire [31:0] _1368_;
wire [31:0] _1369_;
wire [31:0] _1370_;
wire [31:0] _1371_;
wire [31:0] _1372_;
wire [31:0] _1373_;
wire [31:0] _1374_;
wire [31:0] _1375_;
wire _1376_;
wire _1377_;
wire _1378_;
wire _1379_;
wire _1380_;
wire _1381_;
wire _1382_;
wire _1383_;
wire _1384_;
wire _1385_;
wire _1386_;
wire _1387_;
wire _1388_;
wire _1389_;
wire _1390_;
wire _1391_;
wire _1392_;
wire _1393_;
wire _1394_;
wire _1395_;
wire _1396_;
wire _1397_;
wire _1398_;
wire _1399_;
/* src = "generated/sv2v_out.v:1550.16-1550.46" */
wire _1400_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1550.16-1550.46" */
wire _1401_;
/* src = "generated/sv2v_out.v:1550.52-1550.81" */
wire _1402_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1550.52-1550.81" */
wire _1403_;
/* src = "generated/sv2v_out.v:1550.88-1550.117" */
wire _1404_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1550.88-1550.117" */
wire _1405_;
/* src = "generated/sv2v_out.v:1554.15-1554.43" */
wire _1406_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1554.15-1554.43" */
wire _1407_;
/* src = "generated/sv2v_out.v:1554.49-1554.79" */
wire _1408_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1554.49-1554.79" */
wire _1409_;
/* src = "generated/sv2v_out.v:1590.22-1590.50" */
wire _1410_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1590.22-1590.50" */
wire _1411_;
/* src = "generated/sv2v_out.v:1590.58-1590.74" */
wire _1412_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1590.58-1590.74" */
wire _1413_;
/* src = "generated/sv2v_out.v:1590.80-1590.96" */
wire _1414_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1590.80-1590.96" */
wire _1415_;
/* src = "generated/sv2v_out.v:1590.103-1590.119" */
wire _1416_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1590.103-1590.119" */
wire _1417_;
/* src = "generated/sv2v_out.v:1592.69-1592.96" */
wire _1418_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1592.69-1592.96" */
wire _1419_;
/* src = "generated/sv2v_out.v:1601.8-1601.16" */
wire _1420_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1601.8-1601.16" */
wire _1421_;
/* src = "generated/sv2v_out.v:1603.26-1603.42" */
wire _1422_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1603.26-1603.42" */
wire _1423_;
/* src = "generated/sv2v_out.v:1607.8-1607.16" */
wire _1424_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1607.8-1607.16" */
wire _1425_;
/* src = "generated/sv2v_out.v:1609.26-1609.42" */
wire _1426_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1609.26-1609.42" */
wire _1427_;
/* src = "generated/sv2v_out.v:1619.8-1619.28" */
wire _1428_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1619.8-1619.28" */
wire _1429_;
/* src = "generated/sv2v_out.v:1621.8-1621.28" */
wire _1430_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1621.8-1621.28" */
wire _1431_;
/* src = "generated/sv2v_out.v:1598.12-1598.34" */
wire _1432_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1598.12-1598.34" */
wire _1433_;
/* src = "generated/sv2v_out.v:1603.13-1603.43" */
wire _1434_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1603.13-1603.43" */
wire _1435_;
/* src = "generated/sv2v_out.v:1609.13-1609.43" */
wire _1436_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1609.13-1609.43" */
wire _1437_;
/* src = "generated/sv2v_out.v:1618.12-1618.31" */
wire _1438_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1618.12-1618.31" */
wire _1439_;
/* src = "generated/sv2v_out.v:1624.12-1624.32" */
wire _1440_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1624.12-1624.32" */
wire _1441_;
/* src = "generated/sv2v_out.v:1550.15-1550.82" */
wire _1442_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1550.15-1550.82" */
wire _1443_;
/* src = "generated/sv2v_out.v:1563.12-1563.32" */
wire _1444_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1563.12-1563.32" */
wire _1445_;
/* src = "generated/sv2v_out.v:1579.7-1579.27" */
wire _1446_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1579.7-1579.27" */
wire _1447_;
/* src = "generated/sv2v_out.v:1590.57-1590.97" */
wire _1448_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1590.57-1590.97" */
wire _1449_;
/* src = "generated/sv2v_out.v:1590.56-1590.120" */
wire _1450_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1590.56-1590.120" */
wire _1451_;
/* src = "generated/sv2v_out.v:1592.32-1592.97" */
wire _1452_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1592.32-1592.97" */
wire _1453_;
/* src = "generated/sv2v_out.v:1592.31-1592.133" */
wire _1454_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1592.31-1592.133" */
wire _1455_;
/* src = "generated/sv2v_out.v:1592.30-1592.167" */
wire _1456_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1592.30-1592.167" */
wire _1457_;
/* src = "generated/sv2v_out.v:1592.29-1592.203" */
wire _1458_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1592.29-1592.203" */
wire _1459_;
/* src = "generated/sv2v_out.v:1592.28-1592.240" */
wire _1460_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1592.28-1592.240" */
wire _1461_;
/* src = "generated/sv2v_out.v:1593.28-1593.90" */
wire _1462_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1593.28-1593.90" */
wire _1463_;
wire [31:0] _1464_;
/* cellift = 32'd1 */
wire [31:0] _1465_;
wire [31:0] _1466_;
/* cellift = 32'd1 */
wire [31:0] _1467_;
wire [31:0] _1468_;
/* cellift = 32'd1 */
wire [31:0] _1469_;
wire [31:0] _1470_;
/* cellift = 32'd1 */
wire [31:0] _1471_;
wire [31:0] _1472_;
/* cellift = 32'd1 */
wire [31:0] _1473_;
wire [31:0] _1474_;
/* cellift = 32'd1 */
wire [31:0] _1475_;
wire [31:0] _1476_;
/* cellift = 32'd1 */
wire [31:0] _1477_;
wire [31:0] _1478_;
/* cellift = 32'd1 */
wire [31:0] _1479_;
wire [31:0] _1480_;
/* cellift = 32'd1 */
wire [31:0] _1481_;
wire [31:0] _1482_;
/* cellift = 32'd1 */
wire [31:0] _1483_;
wire [31:0] _1484_;
/* cellift = 32'd1 */
wire [31:0] _1485_;
wire [31:0] _1486_;
/* cellift = 32'd1 */
wire [31:0] _1487_;
wire [31:0] _1488_;
/* cellift = 32'd1 */
wire [31:0] _1489_;
wire [31:0] _1490_;
/* cellift = 32'd1 */
wire [31:0] _1491_;
wire [31:0] _1492_;
/* cellift = 32'd1 */
wire [31:0] _1493_;
wire [31:0] _1494_;
/* cellift = 32'd1 */
wire [31:0] _1495_;
wire [31:0] _1496_;
/* cellift = 32'd1 */
wire [31:0] _1497_;
wire [31:0] _1498_;
/* cellift = 32'd1 */
wire [31:0] _1499_;
wire [31:0] _1500_;
/* cellift = 32'd1 */
wire [31:0] _1501_;
wire [31:0] _1502_;
/* cellift = 32'd1 */
wire [31:0] _1503_;
wire [31:0] _1504_;
/* cellift = 32'd1 */
wire [31:0] _1505_;
wire [31:0] _1506_;
/* cellift = 32'd1 */
wire [31:0] _1507_;
wire [31:0] _1508_;
/* cellift = 32'd1 */
wire [31:0] _1509_;
wire [31:0] _1510_;
/* cellift = 32'd1 */
wire [31:0] _1511_;
wire [31:0] _1512_;
/* cellift = 32'd1 */
wire [31:0] _1513_;
wire [31:0] _1514_;
/* cellift = 32'd1 */
wire [31:0] _1515_;
wire [31:0] _1516_;
/* cellift = 32'd1 */
wire [31:0] _1517_;
wire [31:0] _1518_;
/* cellift = 32'd1 */
wire [31:0] _1519_;
wire [31:0] _1520_;
/* cellift = 32'd1 */
wire [31:0] _1521_;
wire [31:0] _1522_;
/* cellift = 32'd1 */
wire [31:0] _1523_;
wire [31:0] _1524_;
/* cellift = 32'd1 */
wire [31:0] _1525_;
wire [31:0] _1526_;
/* cellift = 32'd1 */
wire [31:0] _1527_;
wire [31:0] _1528_;
/* cellift = 32'd1 */
wire [31:0] _1529_;
wire [31:0] _1530_;
/* cellift = 32'd1 */
wire [31:0] _1531_;
wire [31:0] _1532_;
/* cellift = 32'd1 */
wire [31:0] _1533_;
wire [31:0] _1534_;
/* cellift = 32'd1 */
wire [31:0] _1535_;
wire [31:0] _1536_;
/* cellift = 32'd1 */
wire [31:0] _1537_;
wire [31:0] _1538_;
/* cellift = 32'd1 */
wire [31:0] _1539_;
wire [31:0] _1540_;
/* cellift = 32'd1 */
wire [31:0] _1541_;
wire [31:0] _1542_;
/* cellift = 32'd1 */
wire [31:0] _1543_;
wire [31:0] _1544_;
/* cellift = 32'd1 */
wire [31:0] _1545_;
wire [31:0] _1546_;
/* cellift = 32'd1 */
wire [31:0] _1547_;
wire [31:0] _1548_;
/* cellift = 32'd1 */
wire [31:0] _1549_;
wire [31:0] _1550_;
/* cellift = 32'd1 */
wire [31:0] _1551_;
wire [31:0] _1552_;
/* cellift = 32'd1 */
wire [31:0] _1553_;
wire [31:0] _1554_;
/* cellift = 32'd1 */
wire [31:0] _1555_;
wire [31:0] _1556_;
/* cellift = 32'd1 */
wire [31:0] _1557_;
wire [31:0] _1558_;
/* cellift = 32'd1 */
wire [31:0] _1559_;
wire [31:0] _1560_;
/* cellift = 32'd1 */
wire [31:0] _1561_;
wire [31:0] _1562_;
/* cellift = 32'd1 */
wire [31:0] _1563_;
wire [31:0] _1564_;
/* cellift = 32'd1 */
wire [31:0] _1565_;
wire [31:0] _1566_;
/* cellift = 32'd1 */
wire [31:0] _1567_;
wire [31:0] _1568_;
/* cellift = 32'd1 */
wire [31:0] _1569_;
wire [31:0] _1570_;
/* cellift = 32'd1 */
wire [31:0] _1571_;
wire [31:0] _1572_;
/* cellift = 32'd1 */
wire [31:0] _1573_;
wire [31:0] _1574_;
/* cellift = 32'd1 */
wire [31:0] _1575_;
wire [31:0] _1576_;
/* cellift = 32'd1 */
wire [31:0] _1577_;
wire [31:0] _1578_;
/* cellift = 32'd1 */
wire [31:0] _1579_;
wire [31:0] _1580_;
/* cellift = 32'd1 */
wire [31:0] _1581_;
wire [31:0] _1582_;
/* cellift = 32'd1 */
wire [31:0] _1583_;
wire _1584_;
/* cellift = 32'd1 */
wire _1585_;
wire _1586_;
/* cellift = 32'd1 */
wire _1587_;
wire _1588_;
/* cellift = 32'd1 */
wire _1589_;
wire _1590_;
/* cellift = 32'd1 */
wire _1591_;
wire _1592_;
/* cellift = 32'd1 */
wire _1593_;
wire _1594_;
/* cellift = 32'd1 */
wire _1595_;
wire _1596_;
/* cellift = 32'd1 */
wire _1597_;
wire _1598_;
/* cellift = 32'd1 */
wire _1599_;
wire _1600_;
/* cellift = 32'd1 */
wire _1601_;
wire _1602_;
/* cellift = 32'd1 */
wire _1603_;
wire _1604_;
/* cellift = 32'd1 */
wire _1605_;
wire _1606_;
/* cellift = 32'd1 */
wire _1607_;
wire _1608_;
/* cellift = 32'd1 */
wire _1609_;
wire _1610_;
/* cellift = 32'd1 */
wire _1611_;
wire _1612_;
/* cellift = 32'd1 */
wire _1613_;
wire _1614_;
/* cellift = 32'd1 */
wire _1615_;
wire _1616_;
/* cellift = 32'd1 */
wire _1617_;
wire _1618_;
/* cellift = 32'd1 */
wire _1619_;
wire _1620_;
/* cellift = 32'd1 */
wire _1621_;
wire _1622_;
/* cellift = 32'd1 */
wire _1623_;
wire _1624_;
/* cellift = 32'd1 */
wire _1625_;
wire _1626_;
/* cellift = 32'd1 */
wire _1627_;
wire _1628_;
/* cellift = 32'd1 */
wire _1629_;
wire _1630_;
/* cellift = 32'd1 */
wire _1631_;
wire _1632_;
/* cellift = 32'd1 */
wire _1633_;
wire _1634_;
/* cellift = 32'd1 */
wire _1635_;
wire _1636_;
/* cellift = 32'd1 */
wire _1637_;
wire _1638_;
/* cellift = 32'd1 */
wire _1639_;
wire _1640_;
/* cellift = 32'd1 */
wire _1641_;
wire _1642_;
/* cellift = 32'd1 */
wire _1643_;
wire _1644_;
/* cellift = 32'd1 */
wire _1645_;
wire _1646_;
/* cellift = 32'd1 */
wire _1647_;
/* src = "generated/sv2v_out.v:1606.18-1606.21" */
wire [31:0] _1648_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1606.18-1606.21" */
wire [31:0] _1649_;
/* src = "generated/sv2v_out.v:1612.18-1612.21" */
wire [31:0] _1650_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1612.18-1612.21" */
wire [31:0] _1651_;
/* src = "generated/sv2v_out.v:1626.21-1626.29" */
wire _1652_;
wire _1653_;
wire _1654_;
wire _1655_;
/* cellift = 32'd1 */
wire _1656_;
wire [31:0] _1657_;
/* cellift = 32'd1 */
wire [31:0] _1658_;
wire [31:0] _1659_;
/* cellift = 32'd1 */
wire [31:0] _1660_;
/* cellift = 32'd1 */
wire [31:0] _1661_;
wire [31:0] _1662_;
/* cellift = 32'd1 */
wire [31:0] _1663_;
wire [31:0] _1664_;
/* cellift = 32'd1 */
wire [31:0] _1665_;
wire [31:0] _1666_;
/* cellift = 32'd1 */
wire [31:0] _1667_;
wire [31:0] _1668_;
/* cellift = 32'd1 */
wire [31:0] _1669_;
/* cellift = 32'd1 */
wire [31:0] _1670_;
wire [31:0] _1671_;
/* cellift = 32'd1 */
wire [31:0] _1672_;
wire [31:0] _1673_;
/* cellift = 32'd1 */
wire [31:0] _1674_;
/* src = "generated/sv2v_out.v:1519.6-1519.10" */
wire ImmA;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1519.6-1519.10" */
wire ImmA_t0;
/* src = "generated/sv2v_out.v:1523.12-1523.16" */
wire [7:0] ImmE;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1523.12-1523.16" */
wire [7:0] ImmE_t0;
/* src = "generated/sv2v_out.v:1524.13-1524.17" */
wire [11:0] ImmF;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1524.13-1524.17" */
wire [11:0] ImmF_t0;
reg [31:0] REG__0_ ;
/* cellift = 32'd1 */
reg [31:0] REG__0__t0 ;
reg [31:0] REG__10_ ;
/* cellift = 32'd1 */
reg [31:0] REG__10__t0 ;
reg [31:0] REG__11_ ;
/* cellift = 32'd1 */
reg [31:0] REG__11__t0 ;
reg [31:0] REG__12_ ;
/* cellift = 32'd1 */
reg [31:0] REG__12__t0 ;
reg [31:0] REG__13_ ;
/* cellift = 32'd1 */
reg [31:0] REG__13__t0 ;
reg [31:0] REG__14_ ;
/* cellift = 32'd1 */
reg [31:0] REG__14__t0 ;
reg [31:0] REG__15_ ;
/* cellift = 32'd1 */
reg [31:0] REG__15__t0 ;
reg [31:0] REG__16_ ;
/* cellift = 32'd1 */
reg [31:0] REG__16__t0 ;
reg [31:0] REG__17_ ;
/* cellift = 32'd1 */
reg [31:0] REG__17__t0 ;
reg [31:0] REG__18_ ;
/* cellift = 32'd1 */
reg [31:0] REG__18__t0 ;
reg [31:0] REG__19_ ;
/* cellift = 32'd1 */
reg [31:0] REG__19__t0 ;
reg [31:0] REG__1_ ;
/* cellift = 32'd1 */
reg [31:0] REG__1__t0 ;
reg [31:0] REG__20_ ;
/* cellift = 32'd1 */
reg [31:0] REG__20__t0 ;
reg [31:0] REG__21_ ;
/* cellift = 32'd1 */
reg [31:0] REG__21__t0 ;
reg [31:0] REG__22_ ;
/* cellift = 32'd1 */
reg [31:0] REG__22__t0 ;
reg [31:0] REG__23_ ;
/* cellift = 32'd1 */
reg [31:0] REG__23__t0 ;
reg [31:0] REG__24_ ;
/* cellift = 32'd1 */
reg [31:0] REG__24__t0 ;
reg [31:0] REG__25_ ;
/* cellift = 32'd1 */
reg [31:0] REG__25__t0 ;
reg [31:0] REG__26_ ;
/* cellift = 32'd1 */
reg [31:0] REG__26__t0 ;
reg [31:0] REG__27_ ;
/* cellift = 32'd1 */
reg [31:0] REG__27__t0 ;
reg [31:0] REG__28_ ;
/* cellift = 32'd1 */
reg [31:0] REG__28__t0 ;
reg [31:0] REG__29_ ;
/* cellift = 32'd1 */
reg [31:0] REG__29__t0 ;
reg [31:0] REG__2_ ;
/* cellift = 32'd1 */
reg [31:0] REG__2__t0 ;
reg [31:0] REG__30_ ;
/* cellift = 32'd1 */
reg [31:0] REG__30__t0 ;
reg [31:0] REG__31_ ;
/* cellift = 32'd1 */
reg [31:0] REG__31__t0 ;
reg [31:0] REG__3_ ;
/* cellift = 32'd1 */
reg [31:0] REG__3__t0 ;
reg [31:0] REG__4_ ;
/* cellift = 32'd1 */
reg [31:0] REG__4__t0 ;
reg [31:0] REG__5_ ;
/* cellift = 32'd1 */
reg [31:0] REG__5__t0 ;
reg [31:0] REG__6_ ;
/* cellift = 32'd1 */
reg [31:0] REG__6__t0 ;
reg [31:0] REG__7_ ;
/* cellift = 32'd1 */
reg [31:0] REG__7__t0 ;
reg [31:0] REG__8_ ;
/* cellift = 32'd1 */
reg [31:0] REG__8__t0 ;
reg [31:0] REG__9_ ;
/* cellift = 32'd1 */
reg [31:0] REG__9__t0 ;
/* src = "generated/sv2v_out.v:1497.13-1497.16" */
input clk;
wire clk;
/* cellift = 32'd1 */
input clk_t0;
wire clk_t0;
/* src = "generated/sv2v_out.v:1532.7-1532.16" */
wire csr_regrd;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1532.7-1532.16" */
wire csr_regrd_t0;
/* src = "generated/sv2v_out.v:1501.13-1501.22" */
input fetch_rdy;
wire fetch_rdy;
/* cellift = 32'd1 */
input fetch_rdy_t0;
wire fetch_rdy_t0;
/* src = "generated/sv2v_out.v:1530.6-1530.14" */
wire format_B;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1530.6-1530.14" */
wire format_B_t0;
/* src = "generated/sv2v_out.v:1527.6-1527.14" */
wire format_I;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1527.6-1527.14" */
wire format_I_t0;
/* src = "generated/sv2v_out.v:1528.6-1528.14" */
wire format_J;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1528.6-1528.14" */
wire format_J_t0;
/* src = "generated/sv2v_out.v:1529.6-1529.14" */
wire format_S;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1529.6-1529.14" */
wire format_S_t0;
/* src = "generated/sv2v_out.v:1531.6-1531.14" */
wire format_U;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1531.6-1531.14" */
wire format_U_t0;
/* src = "generated/sv2v_out.v:1502.20-1502.29" */
output [31:0] immediate;
wire [31:0] immediate;
/* cellift = 32'd1 */
output [31:0] immediate_t0;
wire [31:0] immediate_t0;
/* src = "generated/sv2v_out.v:1499.20-1499.30" */
input [31:0] instr_data;
wire [31:0] instr_data;
/* cellift = 32'd1 */
input [31:0] instr_data_t0;
wire [31:0] instr_data_t0;
/* src = "generated/sv2v_out.v:1511.7-1511.16" */
wire instr_rdy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1511.7-1511.16" */
wire instr_rdy_t0;
/* src = "generated/sv2v_out.v:1500.13-1500.22" */
input instr_vld;
wire instr_vld;
/* cellift = 32'd1 */
input instr_vld_t0;
wire instr_vld_t0;
/* src = "generated/sv2v_out.v:1533.7-1533.22" */
wire is_regrd_rs1_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1533.7-1533.22" */
wire is_regrd_rs1_en_t0;
/* src = "generated/sv2v_out.v:1534.7-1534.22" */
wire is_regrd_rs2_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1534.7-1534.22" */
wire is_regrd_rs2_en_t0;
/* src = "generated/sv2v_out.v:1512.12-1512.19" */
reg [4:0] reg_rs1;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1512.12-1512.19" */
reg [4:0] reg_rs1_t0;
/* src = "generated/sv2v_out.v:1513.12-1513.19" */
reg [4:0] reg_rs2;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1513.12-1513.19" */
reg [4:0] reg_rs2_t0;
/* src = "generated/sv2v_out.v:1510.6-1510.13" */
reg reg_vld;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1510.6-1510.13" */
reg reg_vld_t0;
/* src = "generated/sv2v_out.v:1503.20-1503.29" */
output [31:0] regrd_rs1;
reg [31:0] regrd_rs1;
/* src = "generated/sv2v_out.v:1505.13-1505.25" */
output regrd_rs1_en;
reg regrd_rs1_en;
/* cellift = 32'd1 */
output regrd_rs1_en_t0;
reg regrd_rs1_en_t0;
/* cellift = 32'd1 */
output [31:0] regrd_rs1_t0;
reg [31:0] regrd_rs1_t0;
/* src = "generated/sv2v_out.v:1504.20-1504.29" */
output [31:0] regrd_rs2;
reg [31:0] regrd_rs2;
/* src = "generated/sv2v_out.v:1506.13-1506.25" */
output regrd_rs2_en;
reg regrd_rs2_en;
/* cellift = 32'd1 */
output regrd_rs2_en_t0;
reg regrd_rs2_en_t0;
/* cellift = 32'd1 */
output [31:0] regrd_rs2_t0;
reg [31:0] regrd_rs2_t0;
/* src = "generated/sv2v_out.v:1507.20-1507.30" */
input [31:0] regwr_data;
wire [31:0] regwr_data;
/* cellift = 32'd1 */
input [31:0] regwr_data_t0;
wire [31:0] regwr_data_t0;
/* src = "generated/sv2v_out.v:1509.13-1509.21" */
input regwr_en;
wire regwr_en;
/* cellift = 32'd1 */
input regwr_en_t0;
wire regwr_en_t0;
/* src = "generated/sv2v_out.v:1508.19-1508.28" */
input [4:0] regwr_sel;
wire [4:0] regwr_sel;
/* cellift = 32'd1 */
input [4:0] regwr_sel_t0;
wire [4:0] regwr_sel_t0;
/* src = "generated/sv2v_out.v:1498.13-1498.17" */
input rstz;
wire rstz;
assign _0147_ = _0652_ & _0663_;
assign _0150_ = _0656_ & _0663_;
assign _0153_ = _0660_ & _0663_;
assign _0156_ = _0001_[3] & _1399_;
assign _0162_ = _0644_ & _0675_;
assign _0165_ = _0652_ & _0675_;
assign _0168_ = _0656_ & _0675_;
assign _0171_ = _0660_ & _0675_;
assign _0159_ = _0001_[2] & _0673_;
assign _0175_ = _0644_ & _0685_;
assign _0178_ = _0652_ & _0685_;
assign _0181_ = _0656_ & _0685_;
assign _0184_ = _0660_ & _0685_;
assign _0192_ = _0644_ & _0697_;
assign _0195_ = _0652_ & _0697_;
assign _0198_ = _0656_ & _0697_;
assign _0201_ = _0660_ & _0697_;
assign _0189_ = _0001_[2] & _0695_;
assign _0205_ = _0644_ & _0707_;
assign _0208_ = _0652_ & _0707_;
assign _0211_ = _0656_ & _0707_;
assign _0214_ = _0660_ & _0707_;
assign _0187_ = _0001_[3] & _0000_[4];
assign _0220_ = _0644_ & _0719_;
assign _0223_ = _0652_ & _0719_;
assign _0226_ = _0656_ & _0719_;
assign _0229_ = _0660_ & _0719_;
assign _0217_ = _0001_[2] & _0717_;
assign _0233_ = _0644_ & _0729_;
assign _0236_ = _0652_ & _0729_;
assign _0239_ = _0656_ & _0729_;
assign _0242_ = _0660_ & _0729_;
assign _0510_ = _0650_ & _0004_[31];
assign _0513_ = _0682_ & _0004_[31];
assign _0516_ = _0684_ & _0004_[31];
assign _0519_ = _0688_ & _0004_[31];
assign _0522_ = _0690_ & _0004_[31];
assign _0525_ = _0692_ & _0004_[31];
assign _0528_ = _0694_ & _0004_[31];
assign _0531_ = _0700_ & _0004_[31];
assign _0534_ = _0702_ & _0004_[31];
assign _0537_ = _0704_ & _0004_[31];
assign _0540_ = _0706_ & _0004_[31];
assign _0543_ = _0654_ & _0004_[31];
assign _0546_ = _0710_ & _0004_[31];
assign _0549_ = _0712_ & _0004_[31];
assign _0552_ = _0714_ & _0004_[31];
assign _0555_ = _0716_ & _0004_[31];
assign _0558_ = _0722_ & _0004_[31];
assign _0561_ = _0724_ & _0004_[31];
assign _0564_ = _0726_ & _0004_[31];
assign _0567_ = _0728_ & _0004_[31];
assign _0570_ = _0732_ & _0004_[31];
assign _0573_ = _0734_ & _0004_[31];
assign _0576_ = _0658_ & _0004_[31];
assign _0579_ = _0736_ & _0004_[31];
assign _0582_ = _0738_ & _0004_[31];
assign _0585_ = _0662_ & _0004_[31];
assign _0588_ = _0666_ & _0004_[31];
assign _0591_ = _0668_ & _0004_[31];
assign _0594_ = _0670_ & _0004_[31];
assign _0597_ = _0672_ & _0004_[31];
assign _0600_ = _0678_ & _0004_[31];
assign _0603_ = _0680_ & _0004_[31];
assign _0868_ = _0644_ & _0647_;
assign _0862_ = _0001_[0] & _1396_;
assign _0872_ = _0652_ & _0647_;
assign _0876_ = _0656_ & _0647_;
assign _0875_ = _0001_[0] & _0000_[1];
assign _0879_ = _0660_ & _0647_;
assign _0865_ = _0001_[2] & _0645_;
assign _0883_ = _0644_ & _0663_;
assign _0148_ = _0664_ & _0651_;
assign _0151_ = _0664_ & _0655_;
assign _0154_ = _0664_ & _0659_;
assign _0160_ = _0674_ & _1397_;
assign _0163_ = _0676_ & _0643_;
assign _0166_ = _0676_ & _0651_;
assign _0169_ = _0676_ & _0655_;
assign _0172_ = _0676_ & _0659_;
assign _0174_ = _0674_ & _0000_[2];
assign _0176_ = _0686_ & _0643_;
assign _0179_ = _0686_ & _0651_;
assign _0182_ = _0686_ & _0655_;
assign _0185_ = _0686_ & _0659_;
assign _0188_ = _0001_[4] & _1398_;
assign _0190_ = _0696_ & _1397_;
assign _0193_ = _0698_ & _0643_;
assign _0196_ = _0698_ & _0651_;
assign _0199_ = _0698_ & _0655_;
assign _0202_ = _0698_ & _0659_;
assign _0204_ = _0696_ & _0000_[2];
assign _0206_ = _0708_ & _0643_;
assign _0209_ = _0708_ & _0651_;
assign _0212_ = _0708_ & _0655_;
assign _0215_ = _0708_ & _0659_;
assign _0157_ = _0001_[4] & _0000_[3];
assign _0218_ = _0718_ & _1397_;
assign _0221_ = _0720_ & _0643_;
assign _0224_ = _0720_ & _0651_;
assign _0227_ = _0720_ & _0655_;
assign _0230_ = _0720_ & _0659_;
assign _0232_ = _0718_ & _0000_[2];
assign _0234_ = _0730_ & _0643_;
assign _0237_ = _0730_ & _0651_;
assign _0240_ = _0730_ & _0655_;
assign _0243_ = _0730_ & _0659_;
assign _0511_ = regwr_en_t0 & _0649_;
assign _0514_ = regwr_en_t0 & _0681_;
assign _0517_ = regwr_en_t0 & _0683_;
assign _0520_ = regwr_en_t0 & _0687_;
assign _0523_ = regwr_en_t0 & _0689_;
assign _0526_ = regwr_en_t0 & _0691_;
assign _0529_ = regwr_en_t0 & _0693_;
assign _0532_ = regwr_en_t0 & _0699_;
assign _0535_ = regwr_en_t0 & _0701_;
assign _0538_ = regwr_en_t0 & _0703_;
assign _0541_ = regwr_en_t0 & _0705_;
assign _0544_ = regwr_en_t0 & _0653_;
assign _0547_ = regwr_en_t0 & _0709_;
assign _0550_ = regwr_en_t0 & _0711_;
assign _0553_ = regwr_en_t0 & _0713_;
assign _0556_ = regwr_en_t0 & _0715_;
assign _0559_ = regwr_en_t0 & _0721_;
assign _0562_ = regwr_en_t0 & _0723_;
assign _0565_ = regwr_en_t0 & _0725_;
assign _0568_ = regwr_en_t0 & _0727_;
assign _0571_ = regwr_en_t0 & _0731_;
assign _0574_ = regwr_en_t0 & _0733_;
assign _0577_ = regwr_en_t0 & _0657_;
assign _0580_ = regwr_en_t0 & _0735_;
assign _0583_ = regwr_en_t0 & _0737_;
assign _0586_ = regwr_en_t0 & _0661_;
assign _0589_ = regwr_en_t0 & _0665_;
assign _0592_ = regwr_en_t0 & _0667_;
assign _0595_ = regwr_en_t0 & _0669_;
assign _0598_ = regwr_en_t0 & _0671_;
assign _0601_ = regwr_en_t0 & _0677_;
assign _0604_ = regwr_en_t0 & _0679_;
assign _0866_ = _0646_ & _1397_;
assign _0869_ = _0648_ & _0643_;
assign _0873_ = _0648_ & _0651_;
assign _0863_ = _0001_[1] & _1395_;
assign _0877_ = _0648_ & _0655_;
assign _0871_ = _0001_[1] & _0000_[0];
assign _0880_ = _0648_ & _0659_;
assign _0882_ = _0646_ & _0000_[2];
assign _0884_ = _0664_ & _0643_;
assign _0146_ = _0644_ & _0664_;
assign _0149_ = _0652_ & _0664_;
assign _0152_ = _0656_ & _0664_;
assign _0155_ = _0660_ & _0664_;
assign _0164_ = _0644_ & _0676_;
assign _0167_ = _0652_ & _0676_;
assign _0170_ = _0656_ & _0676_;
assign _0173_ = _0660_ & _0676_;
assign _0161_ = _0001_[2] & _0674_;
assign _0177_ = _0644_ & _0686_;
assign _0180_ = _0652_ & _0686_;
assign _0183_ = _0656_ & _0686_;
assign _0186_ = _0660_ & _0686_;
assign _0194_ = _0644_ & _0698_;
assign _0197_ = _0652_ & _0698_;
assign _0200_ = _0656_ & _0698_;
assign _0203_ = _0660_ & _0698_;
assign _0191_ = _0001_[2] & _0696_;
assign _0207_ = _0644_ & _0708_;
assign _0210_ = _0652_ & _0708_;
assign _0213_ = _0656_ & _0708_;
assign _0216_ = _0660_ & _0708_;
assign _0158_ = _0001_[3] & _0001_[4];
assign _0222_ = _0644_ & _0720_;
assign _0225_ = _0652_ & _0720_;
assign _0228_ = _0656_ & _0720_;
assign _0231_ = _0660_ & _0720_;
assign _0219_ = _0001_[2] & _0718_;
assign _0235_ = _0644_ & _0730_;
assign _0238_ = _0652_ & _0730_;
assign _0241_ = _0656_ & _0730_;
assign _0244_ = _0660_ & _0730_;
assign _0512_ = _0650_ & regwr_en_t0;
assign _0515_ = _0682_ & regwr_en_t0;
assign _0518_ = _0684_ & regwr_en_t0;
assign _0521_ = _0688_ & regwr_en_t0;
assign _0524_ = _0690_ & regwr_en_t0;
assign _0527_ = _0692_ & regwr_en_t0;
assign _0530_ = _0694_ & regwr_en_t0;
assign _0533_ = _0700_ & regwr_en_t0;
assign _0536_ = _0702_ & regwr_en_t0;
assign _0539_ = _0704_ & regwr_en_t0;
assign _0542_ = _0706_ & regwr_en_t0;
assign _0545_ = _0654_ & regwr_en_t0;
assign _0548_ = _0710_ & regwr_en_t0;
assign _0551_ = _0712_ & regwr_en_t0;
assign _0554_ = _0714_ & regwr_en_t0;
assign _0557_ = _0716_ & regwr_en_t0;
assign _0560_ = _0722_ & regwr_en_t0;
assign _0563_ = _0724_ & regwr_en_t0;
assign _0566_ = _0726_ & regwr_en_t0;
assign _0569_ = _0728_ & regwr_en_t0;
assign _0572_ = _0732_ & regwr_en_t0;
assign _0575_ = _0734_ & regwr_en_t0;
assign _0578_ = _0658_ & regwr_en_t0;
assign _0581_ = _0736_ & regwr_en_t0;
assign _0584_ = _0738_ & regwr_en_t0;
assign _0587_ = _0662_ & regwr_en_t0;
assign _0590_ = _0666_ & regwr_en_t0;
assign _0593_ = _0668_ & regwr_en_t0;
assign _0596_ = _0670_ & regwr_en_t0;
assign _0599_ = _0672_ & regwr_en_t0;
assign _0602_ = _0678_ & regwr_en_t0;
assign _0605_ = _0680_ & regwr_en_t0;
assign _0870_ = _0644_ & _0648_;
assign _0874_ = _0652_ & _0648_;
assign _0878_ = _0656_ & _0648_;
assign _0864_ = _0001_[0] & _0001_[1];
assign _0881_ = _0660_ & _0648_;
assign _0867_ = _0001_[2] & _0646_;
assign _0885_ = _0883_ | _0884_;
assign _0886_ = _0147_ | _0148_;
assign _0887_ = _0150_ | _0151_;
assign _0888_ = _0153_ | _0154_;
assign _0889_ = _0156_ | _0157_;
assign _0890_ = _0159_ | _0160_;
assign _0891_ = _0162_ | _0163_;
assign _0892_ = _0165_ | _0166_;
assign _0893_ = _0168_ | _0169_;
assign _0894_ = _0171_ | _0172_;
assign _0895_ = _0159_ | _0174_;
assign _0896_ = _0175_ | _0176_;
assign _0897_ = _0178_ | _0179_;
assign _0898_ = _0181_ | _0182_;
assign _0899_ = _0184_ | _0185_;
assign _0900_ = _0187_ | _0188_;
assign _0901_ = _0189_ | _0190_;
assign _0902_ = _0192_ | _0193_;
assign _0903_ = _0195_ | _0196_;
assign _0904_ = _0198_ | _0199_;
assign _0905_ = _0201_ | _0202_;
assign _0906_ = _0189_ | _0204_;
assign _0907_ = _0205_ | _0206_;
assign _0908_ = _0208_ | _0209_;
assign _0909_ = _0211_ | _0212_;
assign _0910_ = _0214_ | _0215_;
assign _0911_ = _0187_ | _0157_;
assign _0912_ = _0217_ | _0218_;
assign _0913_ = _0220_ | _0221_;
assign _0914_ = _0223_ | _0224_;
assign _0915_ = _0226_ | _0227_;
assign _0916_ = _0229_ | _0230_;
assign _0917_ = _0217_ | _0232_;
assign _0918_ = _0233_ | _0234_;
assign _0919_ = _0236_ | _0237_;
assign _0920_ = _0239_ | _0240_;
assign _0921_ = _0242_ | _0243_;
assign _1033_ = _0510_ | _0511_;
assign _1034_ = _0513_ | _0514_;
assign _1035_ = _0516_ | _0517_;
assign _1036_ = _0519_ | _0520_;
assign _1037_ = _0522_ | _0523_;
assign _1038_ = _0525_ | _0526_;
assign _1039_ = _0528_ | _0529_;
assign _1040_ = _0531_ | _0532_;
assign _1041_ = _0534_ | _0535_;
assign _1042_ = _0537_ | _0538_;
assign _1043_ = _0540_ | _0541_;
assign _1044_ = _0543_ | _0544_;
assign _1045_ = _0546_ | _0547_;
assign _1046_ = _0549_ | _0550_;
assign _1047_ = _0552_ | _0553_;
assign _1048_ = _0555_ | _0556_;
assign _1049_ = _0558_ | _0559_;
assign _1050_ = _0561_ | _0562_;
assign _1051_ = _0564_ | _0565_;
assign _1052_ = _0567_ | _0568_;
assign _1053_ = _0570_ | _0571_;
assign _1054_ = _0573_ | _0574_;
assign _1055_ = _0576_ | _0577_;
assign _1056_ = _0579_ | _0580_;
assign _1057_ = _0582_ | _0583_;
assign _1058_ = _0585_ | _0586_;
assign _1059_ = _0588_ | _0589_;
assign _1060_ = _0591_ | _0592_;
assign _1061_ = _0594_ | _0595_;
assign _1062_ = _0597_ | _0598_;
assign _1063_ = _0600_ | _0601_;
assign _1064_ = _0603_ | _0604_;
assign _1266_ = _0862_ | _0863_;
assign _1267_ = _0156_ | _0188_;
assign _1268_ = _0865_ | _0866_;
assign _1269_ = _0868_ | _0869_;
assign _1270_ = _0862_ | _0871_;
assign _1271_ = _0872_ | _0873_;
assign _1272_ = _0875_ | _0863_;
assign _1273_ = _0876_ | _0877_;
assign _1274_ = _0875_ | _0871_;
assign _1275_ = _0879_ | _0880_;
assign _1276_ = _0865_ | _0882_;
assign _0666_ = _0885_ | _0146_;
assign _0668_ = _0886_ | _0149_;
assign _0670_ = _0887_ | _0152_;
assign _0672_ = _0888_ | _0155_;
assign _0674_ = _0889_ | _0158_;
assign _0676_ = _0890_ | _0161_;
assign _0678_ = _0891_ | _0164_;
assign _0680_ = _0892_ | _0167_;
assign _0682_ = _0893_ | _0170_;
assign _0684_ = _0894_ | _0173_;
assign _0686_ = _0895_ | _0161_;
assign _0688_ = _0896_ | _0177_;
assign _0690_ = _0897_ | _0180_;
assign _0692_ = _0898_ | _0183_;
assign _0694_ = _0899_ | _0186_;
assign _0696_ = _0900_ | _0158_;
assign _0698_ = _0901_ | _0191_;
assign _0700_ = _0902_ | _0194_;
assign _0702_ = _0903_ | _0197_;
assign _0704_ = _0904_ | _0200_;
assign _0706_ = _0905_ | _0203_;
assign _0708_ = _0906_ | _0191_;
assign _0710_ = _0907_ | _0207_;
assign _0712_ = _0908_ | _0210_;
assign _0714_ = _0909_ | _0213_;
assign _0716_ = _0910_ | _0216_;
assign _0718_ = _0911_ | _0158_;
assign _0720_ = _0912_ | _0219_;
assign _0722_ = _0913_ | _0222_;
assign _0724_ = _0914_ | _0225_;
assign _0726_ = _0915_ | _0228_;
assign _0728_ = _0916_ | _0231_;
assign _0730_ = _0917_ | _0219_;
assign _0732_ = _0918_ | _0235_;
assign _0734_ = _0919_ | _0238_;
assign _0736_ = _0920_ | _0241_;
assign _0738_ = _0921_ | _0244_;
assign _1585_ = _1033_ | _0512_;
assign _1587_ = _1034_ | _0515_;
assign _1589_ = _1035_ | _0518_;
assign _1591_ = _1036_ | _0521_;
assign _1593_ = _1037_ | _0524_;
assign _1595_ = _1038_ | _0527_;
assign _1597_ = _1039_ | _0530_;
assign _1599_ = _1040_ | _0533_;
assign _1601_ = _1041_ | _0536_;
assign _1603_ = _1042_ | _0539_;
assign _1605_ = _1043_ | _0542_;
assign _1607_ = _1044_ | _0545_;
assign _1609_ = _1045_ | _0548_;
assign _1611_ = _1046_ | _0551_;
assign _1613_ = _1047_ | _0554_;
assign _1615_ = _1048_ | _0557_;
assign _1617_ = _1049_ | _0560_;
assign _1619_ = _1050_ | _0563_;
assign _1621_ = _1051_ | _0566_;
assign _1623_ = _1052_ | _0569_;
assign _1625_ = _1053_ | _0572_;
assign _1627_ = _1054_ | _0575_;
assign _1629_ = _1055_ | _0578_;
assign _1631_ = _1056_ | _0581_;
assign _1633_ = _1057_ | _0584_;
assign _1635_ = _1058_ | _0587_;
assign _1637_ = _1059_ | _0590_;
assign _1639_ = _1060_ | _0593_;
assign _1641_ = _1061_ | _0596_;
assign _1643_ = _1062_ | _0599_;
assign _1645_ = _1063_ | _0602_;
assign _1647_ = _1064_ | _0605_;
assign _0644_ = _1266_ | _0864_;
assign _0646_ = _1267_ | _0158_;
assign _0648_ = _1268_ | _0867_;
assign _0650_ = _1269_ | _0870_;
assign _0652_ = _1270_ | _0864_;
assign _0654_ = _1271_ | _0874_;
assign _0656_ = _1272_ | _0864_;
assign _0658_ = _1273_ | _0878_;
assign _0660_ = _1274_ | _0864_;
assign _0662_ = _1275_ | _0881_;
assign _0664_ = _1276_ | _0867_;
assign _1335_ = _1673_ ^ regrd_rs1;
assign _1336_ = _1664_ ^ regrd_rs2;
assign _1337_ = is_regrd_rs1_en ^ regrd_rs1_en;
assign _1338_ = is_regrd_rs2_en ^ regrd_rs2_en;
assign _1340_ = instr_data[19:15] ^ reg_rs1;
assign _1341_ = instr_data[24:20] ^ reg_rs2;
assign _1343_ = { ImmF, ImmE, ImmA } ^ { immediate[31:12], immediate[0] };
assign _1344_ = _0002_ ^ REG__9_ ;
assign _1345_ = _0002_ ^ REG__8_ ;
assign _1346_ = _0002_ ^ REG__7_ ;
assign _1347_ = _0002_ ^ REG__6_ ;
assign _1348_ = _0002_ ^ REG__5_ ;
assign _1349_ = _0002_ ^ REG__4_ ;
assign _1350_ = _0002_ ^ REG__3_ ;
assign _1351_ = _0002_ ^ REG__31_ ;
assign _1352_ = _0002_ ^ REG__30_ ;
assign _1353_ = _0002_ ^ REG__2_ ;
assign _1354_ = _0002_ ^ REG__29_ ;
assign _1355_ = _0002_ ^ REG__28_ ;
assign _1356_ = _0002_ ^ REG__27_ ;
assign _1357_ = _0002_ ^ REG__26_ ;
assign _1358_ = _0002_ ^ REG__25_ ;
assign _1359_ = _0002_ ^ REG__24_ ;
assign _1360_ = _0002_ ^ REG__23_ ;
assign _1361_ = _0002_ ^ REG__22_ ;
assign _1362_ = _0002_ ^ REG__21_ ;
assign _1363_ = _0002_ ^ REG__20_ ;
assign _1364_ = _0002_ ^ REG__1_ ;
assign _1365_ = _0002_ ^ REG__19_ ;
assign _1366_ = _0002_ ^ REG__18_ ;
assign _1367_ = _0002_ ^ REG__17_ ;
assign _1368_ = _0002_ ^ REG__16_ ;
assign _1369_ = _0002_ ^ REG__15_ ;
assign _1370_ = _0002_ ^ REG__14_ ;
assign _1371_ = _0002_ ^ REG__13_ ;
assign _1372_ = _0002_ ^ REG__12_ ;
assign _1373_ = _0002_ ^ REG__11_ ;
assign _1374_ = _0002_ ^ REG__10_ ;
assign _1375_ = _0002_ ^ REG__0_ ;
assign _0086_ = ~ _0023_;
assign _0087_ = ~ _0025_;
assign _0088_ = ~ _0027_;
assign _0090_ = ~ _1646_;
assign _0091_ = ~ _1644_;
assign _0092_ = ~ _1642_;
assign _0093_ = ~ _1640_;
assign _0094_ = ~ _1638_;
assign _0095_ = ~ _1636_;
assign _0096_ = ~ _1634_;
assign _0097_ = ~ _1632_;
assign _0098_ = ~ _1630_;
assign _0099_ = ~ _1628_;
assign _0100_ = ~ _1626_;
assign _0101_ = ~ _1624_;
assign _0102_ = ~ _1622_;
assign _0103_ = ~ _1620_;
assign _0104_ = ~ _1618_;
assign _0105_ = ~ _1616_;
assign _0106_ = ~ _1614_;
assign _0107_ = ~ _1612_;
assign _0108_ = ~ _1610_;
assign _0109_ = ~ _1608_;
assign _0110_ = ~ _1606_;
assign _0111_ = ~ _1604_;
assign _0112_ = ~ _1602_;
assign _0113_ = ~ _1600_;
assign _0114_ = ~ _1598_;
assign _0115_ = ~ _1596_;
assign _0116_ = ~ _1594_;
assign _0117_ = ~ _1592_;
assign _0118_ = ~ _1590_;
assign _0119_ = ~ _1588_;
assign _0120_ = ~ _1586_;
assign _0121_ = ~ _1584_;
assign _1102_ = _1674_ | regrd_rs1_t0;
assign _1106_ = _1665_ | regrd_rs2_t0;
assign _1110_ = is_regrd_rs1_en_t0 | regrd_rs1_en_t0;
assign _1114_ = is_regrd_rs2_en_t0 | regrd_rs2_en_t0;
assign _1122_ = instr_data_t0[19:15] | reg_rs1_t0;
assign _1126_ = instr_data_t0[24:20] | reg_rs2_t0;
assign _1134_ = { ImmF_t0, ImmE_t0, ImmA_t0 } | { immediate_t0[31:12], immediate_t0[0] };
assign _1138_ = _0003_ | REG__9__t0 ;
assign _1142_ = _0003_ | REG__8__t0 ;
assign _1146_ = _0003_ | REG__7__t0 ;
assign _1150_ = _0003_ | REG__6__t0 ;
assign _1154_ = _0003_ | REG__5__t0 ;
assign _1158_ = _0003_ | REG__4__t0 ;
assign _1162_ = _0003_ | REG__3__t0 ;
assign _1166_ = _0003_ | REG__31__t0 ;
assign _1170_ = _0003_ | REG__30__t0 ;
assign _1174_ = _0003_ | REG__2__t0 ;
assign _1178_ = _0003_ | REG__29__t0 ;
assign _1182_ = _0003_ | REG__28__t0 ;
assign _1186_ = _0003_ | REG__27__t0 ;
assign _1190_ = _0003_ | REG__26__t0 ;
assign _1194_ = _0003_ | REG__25__t0 ;
assign _1198_ = _0003_ | REG__24__t0 ;
assign _1202_ = _0003_ | REG__23__t0 ;
assign _1206_ = _0003_ | REG__22__t0 ;
assign _1210_ = _0003_ | REG__21__t0 ;
assign _1214_ = _0003_ | REG__20__t0 ;
assign _1218_ = _0003_ | REG__1__t0 ;
assign _1222_ = _0003_ | REG__19__t0 ;
assign _1226_ = _0003_ | REG__18__t0 ;
assign _1230_ = _0003_ | REG__17__t0 ;
assign _1234_ = _0003_ | REG__16__t0 ;
assign _1238_ = _0003_ | REG__15__t0 ;
assign _1242_ = _0003_ | REG__14__t0 ;
assign _1246_ = _0003_ | REG__13__t0 ;
assign _1250_ = _0003_ | REG__12__t0 ;
assign _1254_ = _0003_ | REG__11__t0 ;
assign _1258_ = _0003_ | REG__10__t0 ;
assign _1262_ = _0003_ | REG__0__t0 ;
assign _1103_ = _1335_ | _1102_;
assign _1107_ = _1336_ | _1106_;
assign _1111_ = _1337_ | _1110_;
assign _1115_ = _1338_ | _1114_;
assign _1123_ = _1340_ | _1122_;
assign _1127_ = _1341_ | _1126_;
assign _1135_ = _1343_ | _1134_;
assign _1139_ = _1344_ | _1138_;
assign _1143_ = _1345_ | _1142_;
assign _1147_ = _1346_ | _1146_;
assign _1151_ = _1347_ | _1150_;
assign _1155_ = _1348_ | _1154_;
assign _1159_ = _1349_ | _1158_;
assign _1163_ = _1350_ | _1162_;
assign _1167_ = _1351_ | _1166_;
assign _1171_ = _1352_ | _1170_;
assign _1175_ = _1353_ | _1174_;
assign _1179_ = _1354_ | _1178_;
assign _1183_ = _1355_ | _1182_;
assign _1187_ = _1356_ | _1186_;
assign _1191_ = _1357_ | _1190_;
assign _1195_ = _1358_ | _1194_;
assign _1199_ = _1359_ | _1198_;
assign _1203_ = _1360_ | _1202_;
assign _1207_ = _1361_ | _1206_;
assign _1211_ = _1362_ | _1210_;
assign _1215_ = _1363_ | _1214_;
assign _1219_ = _1364_ | _1218_;
assign _1223_ = _1365_ | _1222_;
assign _1227_ = _1366_ | _1226_;
assign _1231_ = _1367_ | _1230_;
assign _1235_ = _1368_ | _1234_;
assign _1239_ = _1369_ | _1238_;
assign _1243_ = _1370_ | _1242_;
assign _1247_ = _1371_ | _1246_;
assign _1251_ = _1372_ | _1250_;
assign _1255_ = _1373_ | _1254_;
assign _1259_ = _1374_ | _1258_;
assign _1263_ = _1375_ | _1262_;
assign _0739_ = { _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_ } & _1674_;
assign _0742_ = { _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_ } & _1665_;
assign _0745_ = _0027_ & is_regrd_rs1_en_t0;
assign _0748_ = _0027_ & is_regrd_rs2_en_t0;
assign _0754_ = { _0027_, _0027_, _0027_, _0027_, _0027_ } & instr_data_t0[19:15];
assign _0757_ = { _0027_, _0027_, _0027_, _0027_, _0027_ } & instr_data_t0[24:20];
assign _0763_ = { _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_ } & { ImmF_t0, ImmE_t0, ImmA_t0 };
assign _0766_ = { _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_, _1646_ } & _0003_;
assign _0769_ = { _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_, _1644_ } & _0003_;
assign _0772_ = { _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_ } & _0003_;
assign _0775_ = { _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_ } & _0003_;
assign _0778_ = { _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_, _1638_ } & _0003_;
assign _0781_ = { _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_, _1636_ } & _0003_;
assign _0784_ = { _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_ } & _0003_;
assign _0787_ = { _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_ } & _0003_;
assign _0790_ = { _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_ } & _0003_;
assign _0793_ = { _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_ } & _0003_;
assign _0796_ = { _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_, _1626_ } & _0003_;
assign _0799_ = { _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_, _1624_ } & _0003_;
assign _0802_ = { _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_, _1622_ } & _0003_;
assign _0805_ = { _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_, _1620_ } & _0003_;
assign _0808_ = { _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_, _1618_ } & _0003_;
assign _0811_ = { _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_, _1616_ } & _0003_;
assign _0814_ = { _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_, _1614_ } & _0003_;
assign _0817_ = { _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_, _1612_ } & _0003_;
assign _0820_ = { _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_, _1610_ } & _0003_;
assign _0823_ = { _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_, _1608_ } & _0003_;
assign _0826_ = { _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_, _1606_ } & _0003_;
assign _0829_ = { _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_, _1604_ } & _0003_;
assign _0832_ = { _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_, _1602_ } & _0003_;
assign _0835_ = { _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_, _1600_ } & _0003_;
assign _0838_ = { _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_, _1598_ } & _0003_;
assign _0841_ = { _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_, _1596_ } & _0003_;
assign _0844_ = { _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_, _1594_ } & _0003_;
assign _0847_ = { _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_, _1592_ } & _0003_;
assign _0850_ = { _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_, _1590_ } & _0003_;
assign _0853_ = { _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_, _1588_ } & _0003_;
assign _0856_ = { _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_, _1586_ } & _0003_;
assign _0859_ = { _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_, _1584_ } & _0003_;
assign _0740_ = { _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_, _0086_ } & regrd_rs1_t0;
assign _0743_ = { _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_, _0087_ } & regrd_rs2_t0;
assign _0746_ = _0088_ & regrd_rs1_en_t0;
assign _0749_ = _0088_ & regrd_rs2_en_t0;
assign _0755_ = { _0088_, _0088_, _0088_, _0088_, _0088_ } & reg_rs1_t0;
assign _0758_ = { _0088_, _0088_, _0088_, _0088_, _0088_ } & reg_rs2_t0;
assign _0764_ = { _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_ } & { immediate_t0[31:12], immediate_t0[0] };
assign _0767_ = { _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_, _0090_ } & REG__9__t0 ;
assign _0770_ = { _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_, _0091_ } & REG__8__t0 ;
assign _0773_ = { _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_, _0092_ } & REG__7__t0 ;
assign _0776_ = { _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_, _0093_ } & REG__6__t0 ;
assign _0779_ = { _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_ } & REG__5__t0 ;
assign _0782_ = { _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_ } & REG__4__t0 ;
assign _0785_ = { _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_ } & REG__3__t0 ;
assign _0788_ = { _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_ } & REG__31__t0 ;
assign _0791_ = { _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_ } & REG__30__t0 ;
assign _0794_ = { _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_ } & REG__2__t0 ;
assign _0797_ = { _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_ } & REG__29__t0 ;
assign _0800_ = { _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_ } & REG__28__t0 ;
assign _0803_ = { _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_ } & REG__27__t0 ;
assign _0806_ = { _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_ } & REG__26__t0 ;
assign _0809_ = { _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_ } & REG__25__t0 ;
assign _0812_ = { _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_ } & REG__24__t0 ;
assign _0815_ = { _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_ } & REG__23__t0 ;
assign _0818_ = { _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_ } & REG__22__t0 ;
assign _0821_ = { _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_ } & REG__21__t0 ;
assign _0824_ = { _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_ } & REG__20__t0 ;
assign _0827_ = { _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_ } & REG__1__t0 ;
assign _0830_ = { _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_ } & REG__19__t0 ;
assign _0833_ = { _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_ } & REG__18__t0 ;
assign _0836_ = { _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_ } & REG__17__t0 ;
assign _0839_ = { _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_ } & REG__16__t0 ;
assign _0842_ = { _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_ } & REG__15__t0 ;
assign _0845_ = { _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_ } & REG__14__t0 ;
assign _0848_ = { _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_ } & REG__13__t0 ;
assign _0851_ = { _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_ } & REG__12__t0 ;
assign _0854_ = { _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_ } & REG__11__t0 ;
assign _0857_ = { _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_ } & REG__10__t0 ;
assign _0860_ = { _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_ } & REG__0__t0 ;
assign _0741_ = _1103_ & { _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_ };
assign _0744_ = _1107_ & { _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_ };
assign _0747_ = _1111_ & _0028_;
assign _0750_ = _1115_ & _0028_;
assign _0756_ = _1123_ & { _0028_, _0028_, _0028_, _0028_, _0028_ };
assign _0759_ = _1127_ & { _0028_, _0028_, _0028_, _0028_, _0028_ };
assign _0765_ = _1135_ & { _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_ };
assign _0768_ = _1139_ & { _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_, _1647_ };
assign _0771_ = _1143_ & { _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_, _1645_ };
assign _0774_ = _1147_ & { _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_ };
assign _0777_ = _1151_ & { _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_ };
assign _0780_ = _1155_ & { _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_, _1639_ };
assign _0783_ = _1159_ & { _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_ };
assign _0786_ = _1163_ & { _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_ };
assign _0789_ = _1167_ & { _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_, _1633_ };
assign _0792_ = _1171_ & { _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_ };
assign _0795_ = _1175_ & { _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_ };
assign _0798_ = _1179_ & { _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_, _1627_ };
assign _0801_ = _1183_ & { _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_, _1625_ };
assign _0804_ = _1187_ & { _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_, _1623_ };
assign _0807_ = _1191_ & { _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_, _1621_ };
assign _0810_ = _1195_ & { _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_, _1619_ };
assign _0813_ = _1199_ & { _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_, _1617_ };
assign _0816_ = _1203_ & { _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_, _1615_ };
assign _0819_ = _1207_ & { _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_, _1613_ };
assign _0822_ = _1211_ & { _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_, _1611_ };
assign _0825_ = _1215_ & { _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_, _1609_ };
assign _0828_ = _1219_ & { _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_, _1607_ };
assign _0831_ = _1223_ & { _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_, _1605_ };
assign _0834_ = _1227_ & { _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_, _1603_ };
assign _0837_ = _1231_ & { _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_, _1601_ };
assign _0840_ = _1235_ & { _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_, _1599_ };
assign _0843_ = _1239_ & { _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_, _1597_ };
assign _0846_ = _1243_ & { _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_, _1595_ };
assign _0849_ = _1247_ & { _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_, _1593_ };
assign _0852_ = _1251_ & { _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_, _1591_ };
assign _0855_ = _1255_ & { _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_, _1589_ };
assign _0858_ = _1259_ & { _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_, _1587_ };
assign _0861_ = _1263_ & { _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_, _1585_ };
assign _1104_ = _0739_ | _0740_;
assign _1108_ = _0742_ | _0743_;
assign _1112_ = _0745_ | _0746_;
assign _1116_ = _0748_ | _0749_;
assign _1124_ = _0754_ | _0755_;
assign _1128_ = _0757_ | _0758_;
assign _1136_ = _0763_ | _0764_;
assign _1140_ = _0766_ | _0767_;
assign _1144_ = _0769_ | _0770_;
assign _1148_ = _0772_ | _0773_;
assign _1152_ = _0775_ | _0776_;
assign _1156_ = _0778_ | _0779_;
assign _1160_ = _0781_ | _0782_;
assign _1164_ = _0784_ | _0785_;
assign _1168_ = _0787_ | _0788_;
assign _1172_ = _0790_ | _0791_;
assign _1176_ = _0793_ | _0794_;
assign _1180_ = _0796_ | _0797_;
assign _1184_ = _0799_ | _0800_;
assign _1188_ = _0802_ | _0803_;
assign _1192_ = _0805_ | _0806_;
assign _1196_ = _0808_ | _0809_;
assign _1200_ = _0811_ | _0812_;
assign _1204_ = _0814_ | _0815_;
assign _1208_ = _0817_ | _0818_;
assign _1212_ = _0820_ | _0821_;
assign _1216_ = _0823_ | _0824_;
assign _1220_ = _0826_ | _0827_;
assign _1224_ = _0829_ | _0830_;
assign _1228_ = _0832_ | _0833_;
assign _1232_ = _0835_ | _0836_;
assign _1236_ = _0838_ | _0839_;
assign _1240_ = _0841_ | _0842_;
assign _1244_ = _0844_ | _0845_;
assign _1248_ = _0847_ | _0848_;
assign _1252_ = _0850_ | _0851_;
assign _1256_ = _0853_ | _0854_;
assign _1260_ = _0856_ | _0857_;
assign _1264_ = _0859_ | _0860_;
assign _1105_ = _1104_ | _0741_;
assign _1109_ = _1108_ | _0744_;
assign _1113_ = _1112_ | _0747_;
assign _1117_ = _1116_ | _0750_;
assign _1125_ = _1124_ | _0756_;
assign _1129_ = _1128_ | _0759_;
assign _1137_ = _1136_ | _0765_;
assign _1141_ = _1140_ | _0768_;
assign _1145_ = _1144_ | _0771_;
assign _1149_ = _1148_ | _0774_;
assign _1153_ = _1152_ | _0777_;
assign _1157_ = _1156_ | _0780_;
assign _1161_ = _1160_ | _0783_;
assign _1165_ = _1164_ | _0786_;
assign _1169_ = _1168_ | _0789_;
assign _1173_ = _1172_ | _0792_;
assign _1177_ = _1176_ | _0795_;
assign _1181_ = _1180_ | _0798_;
assign _1185_ = _1184_ | _0801_;
assign _1189_ = _1188_ | _0804_;
assign _1193_ = _1192_ | _0807_;
assign _1197_ = _1196_ | _0810_;
assign _1201_ = _1200_ | _0813_;
assign _1205_ = _1204_ | _0816_;
assign _1209_ = _1208_ | _0819_;
assign _1213_ = _1212_ | _0822_;
assign _1217_ = _1216_ | _0825_;
assign _1221_ = _1220_ | _0828_;
assign _1225_ = _1224_ | _0831_;
assign _1229_ = _1228_ | _0834_;
assign _1233_ = _1232_ | _0837_;
assign _1237_ = _1236_ | _0840_;
assign _1241_ = _1240_ | _0843_;
assign _1245_ = _1244_ | _0846_;
assign _1249_ = _1248_ | _0849_;
assign _1253_ = _1252_ | _0852_;
assign _1257_ = _1256_ | _0855_;
assign _1261_ = _1260_ | _0858_;
assign _1265_ = _1264_ | _0861_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME regrd_rs1_t0 */
always_ff @(posedge clk)
regrd_rs1_t0 <= _1105_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME regrd_rs2_t0 */
always_ff @(posedge clk)
regrd_rs2_t0 <= _1109_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME regrd_rs1_en_t0 */
always_ff @(posedge clk)
regrd_rs1_en_t0 <= _1113_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME regrd_rs2_en_t0 */
always_ff @(posedge clk)
regrd_rs2_en_t0 <= _1117_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME reg_rs1_t0 */
always_ff @(posedge clk)
reg_rs1_t0 <= _1125_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME reg_rs2_t0 */
always_ff @(posedge clk)
reg_rs2_t0 <= _1129_;
reg [20:0] _2406_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME _2406_ */
always_ff @(posedge clk)
_2406_ <= _1137_;
assign { immediate_t0[31:12], immediate_t0[0] } = _2406_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__9__t0  */
always_ff @(posedge clk)
REG__9__t0  <= _1141_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__8__t0  */
always_ff @(posedge clk)
REG__8__t0  <= _1145_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__7__t0  */
always_ff @(posedge clk)
REG__7__t0  <= _1149_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__6__t0  */
always_ff @(posedge clk)
REG__6__t0  <= _1153_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__5__t0  */
always_ff @(posedge clk)
REG__5__t0  <= _1157_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__4__t0  */
always_ff @(posedge clk)
REG__4__t0  <= _1161_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__3__t0  */
always_ff @(posedge clk)
REG__3__t0  <= _1165_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__31__t0  */
always_ff @(posedge clk)
REG__31__t0  <= _1169_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__30__t0  */
always_ff @(posedge clk)
REG__30__t0  <= _1173_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__2__t0  */
always_ff @(posedge clk)
REG__2__t0  <= _1177_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__29__t0  */
always_ff @(posedge clk)
REG__29__t0  <= _1181_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__28__t0  */
always_ff @(posedge clk)
REG__28__t0  <= _1185_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__27__t0  */
always_ff @(posedge clk)
REG__27__t0  <= _1189_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__26__t0  */
always_ff @(posedge clk)
REG__26__t0  <= _1193_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__25__t0  */
always_ff @(posedge clk)
REG__25__t0  <= _1197_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__24__t0  */
always_ff @(posedge clk)
REG__24__t0  <= _1201_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__23__t0  */
always_ff @(posedge clk)
REG__23__t0  <= _1205_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__22__t0  */
always_ff @(posedge clk)
REG__22__t0  <= _1209_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__21__t0  */
always_ff @(posedge clk)
REG__21__t0  <= _1213_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__20__t0  */
always_ff @(posedge clk)
REG__20__t0  <= _1217_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__1__t0  */
always_ff @(posedge clk)
REG__1__t0  <= _1221_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__19__t0  */
always_ff @(posedge clk)
REG__19__t0  <= _1225_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__18__t0  */
always_ff @(posedge clk)
REG__18__t0  <= _1229_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__17__t0  */
always_ff @(posedge clk)
REG__17__t0  <= _1233_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__16__t0  */
always_ff @(posedge clk)
REG__16__t0  <= _1237_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__15__t0  */
always_ff @(posedge clk)
REG__15__t0  <= _1241_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__14__t0  */
always_ff @(posedge clk)
REG__14__t0  <= _1245_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__13__t0  */
always_ff @(posedge clk)
REG__13__t0  <= _1249_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__12__t0  */
always_ff @(posedge clk)
REG__12__t0  <= _1253_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__11__t0  */
always_ff @(posedge clk)
REG__11__t0  <= _1257_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__10__t0  */
always_ff @(posedge clk)
REG__10__t0  <= _1261_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__0__t0  */
always_ff @(posedge clk)
REG__0__t0  <= _1265_;
assign _0127_ = | { _1429_, _1439_, _1433_ };
assign _0128_ = | { _1431_, _1439_, _1433_ };
assign _0126_ = | { _1439_, _1433_ };
assign _0134_ = | instr_data_t0[14:12];
assign _0133_ = | instr_data_t0[6:2];
assign _0136_ = | { instr_data_t0[19:15], regwr_sel_t0 };
assign _0138_ = | { instr_data_t0[24:20], regwr_sel_t0 };
assign _0139_ = | { reg_rs1_t0, regwr_sel_t0 };
assign _0140_ = | { reg_rs2_t0, regwr_sel_t0 };
assign _0926_ = instr_data_t0[19:15] | regwr_sel_t0;
assign _0927_ = instr_data_t0[24:20] | regwr_sel_t0;
assign _0928_ = reg_rs1_t0 | regwr_sel_t0;
assign _0929_ = reg_rs2_t0 | regwr_sel_t0;
assign _0032_ = ~ { _1429_, _1439_, _1433_ };
assign _0033_ = ~ { _1431_, _1439_, _1433_ };
assign _0031_ = ~ { _1439_, _1433_ };
assign _0036_ = ~ instr_data_t0[14:12];
assign _0035_ = ~ instr_data_t0[6:2];
assign _0038_ = ~ _0926_;
assign _0040_ = ~ _0927_;
assign _0041_ = ~ _0928_;
assign _0042_ = ~ _0929_;
assign _0246_ = { _1428_, _1438_, _1432_ } & _0032_;
assign _0247_ = { _1430_, _1438_, _1432_ } & _0033_;
assign _0245_ = { _1438_, _1432_ } & _0031_;
assign _0250_ = instr_data[14:12] & _0036_;
assign _0249_ = instr_data[6:2] & _0035_;
assign _0252_ = instr_data[19:15] & _0038_;
assign _0255_ = instr_data[24:20] & _0040_;
assign _0257_ = reg_rs1 & _0041_;
assign _0259_ = reg_rs2 & _0042_;
assign _0253_ = regwr_sel & _0038_;
assign _0256_ = regwr_sel & _0040_;
assign _0258_ = regwr_sel & _0041_;
assign _0260_ = regwr_sel & _0042_;
assign _1376_ = _0246_ == { 1'h0, _0032_[1], 1'h0 };
assign _1377_ = _0247_ == { 1'h0, _0033_[1], 1'h0 };
assign _1378_ = _0245_ == { _0031_[1], 1'h0 };
assign _1379_ = _0249_ == { _0035_[4:3], 1'h0, _0035_[1:0] };
assign _1380_ = _0249_ == { 1'h0, _0035_[3:2], 1'h0, _0035_[0] };
assign _1381_ = _0249_ == { 2'h0, _0035_[2], 1'h0, _0035_[0] };
assign _1382_ = _0249_ == { _0035_[4:2], 2'h0 };
assign _1383_ = _0250_ == { 2'h0, _0036_[0] };
assign _1384_ = _0250_ == { 1'h0, _0036_[1], 1'h0 };
assign _1385_ = _0250_ == { 1'h0, _0036_[1:0] };
assign _1386_ = _0249_ == { 2'h0, _0035_[2], 2'h0 };
assign _1387_ = _0249_ == { _0035_[4:3], 2'h0, _0035_[0] };
assign _1388_ = _0249_ == { 1'h0, _0035_[3:2], 2'h0 };
assign _1389_ = _0249_ == { _0035_[4:3], 3'h0 };
assign _1390_ = _0249_ == { 1'h0, _0035_[3], 3'h0 };
assign _1391_ = _0252_ == _0253_;
assign _1392_ = _0255_ == _0256_;
assign _1393_ = _0257_ == _0258_;
assign _1394_ = _0259_ == _0260_;
assign _0016_ = _1376_ & _0127_;
assign _0018_ = _1377_ & _0128_;
assign _0022_ = _1378_ & _0126_;
assign format_J_t0 = _1379_ & _0133_;
assign _1407_ = _1380_ & _0133_;
assign _1409_ = _1381_ & _0133_;
assign _1411_ = _1382_ & _0133_;
assign _1413_ = _1383_ & _0134_;
assign _1415_ = _1384_ & _0134_;
assign _1417_ = _1385_ & _0134_;
assign _1401_ = _1386_ & _0133_;
assign _1403_ = _1387_ & _0133_;
assign _1419_ = _1388_ & _0133_;
assign format_B_t0 = _1389_ & _0133_;
assign format_S_t0 = _1390_ & _0133_;
assign _1423_ = _1391_ & _0136_;
assign _1427_ = _1392_ & _0138_;
assign _1429_ = _1393_ & _0139_;
assign _1431_ = _1394_ & _0140_;
/* src = "generated/sv2v_out.v:1595.2-1625.20" */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME regrd_rs1 */
always_ff @(posedge clk)
if (_0023_) regrd_rs1 <= _1673_;
/* src = "generated/sv2v_out.v:1595.2-1625.20" */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME regrd_rs2 */
always_ff @(posedge clk)
if (_0025_) regrd_rs2 <= _1664_;
/* src = "generated/sv2v_out.v:1595.2-1625.20" */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME regrd_rs1_en */
always_ff @(posedge clk)
if (_0027_) regrd_rs1_en <= is_regrd_rs1_en;
/* src = "generated/sv2v_out.v:1595.2-1625.20" */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME regrd_rs2_en */
always_ff @(posedge clk)
if (_0027_) regrd_rs2_en <= is_regrd_rs2_en;
/* src = "generated/sv2v_out.v:1595.2-1625.20" */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME reg_vld */
always_ff @(posedge clk)
if (!rstz) reg_vld <= 1'h0;
else if (_0029_) reg_vld <= _1655_;
/* src = "generated/sv2v_out.v:1595.2-1625.20" */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME reg_rs1 */
always_ff @(posedge clk)
if (_0027_) reg_rs1 <= instr_data[19:15];
/* src = "generated/sv2v_out.v:1595.2-1625.20" */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME reg_rs2 */
always_ff @(posedge clk)
if (_0027_) reg_rs2 <= instr_data[24:20];
reg [10:0] _2519_;
/* src = "generated/sv2v_out.v:1595.2-1625.20" */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME _2519_ */
always_ff @(posedge clk)
if (_0027_)
if (format_U) _2519_ <= 11'h000;
else _2519_ <= { _0009_, instr_data[30:25], _0007_ };
assign immediate[11:1] = _2519_;
reg [20:0] _2520_;
/* src = "generated/sv2v_out.v:1595.2-1625.20" */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME _2520_ */
always_ff @(posedge clk)
if (_0027_) _2520_ <= { ImmF, ImmE, ImmA };
assign { immediate[31:12], immediate[0] } = _2520_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__9_  */
always_ff @(posedge clk)
if (_1646_) REG__9_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__8_  */
always_ff @(posedge clk)
if (_1644_) REG__8_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__7_  */
always_ff @(posedge clk)
if (_1642_) REG__7_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__6_  */
always_ff @(posedge clk)
if (_1640_) REG__6_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__5_  */
always_ff @(posedge clk)
if (_1638_) REG__5_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__4_  */
always_ff @(posedge clk)
if (_1636_) REG__4_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__3_  */
always_ff @(posedge clk)
if (_1634_) REG__3_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__31_  */
always_ff @(posedge clk)
if (_1632_) REG__31_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__30_  */
always_ff @(posedge clk)
if (_1630_) REG__30_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__2_  */
always_ff @(posedge clk)
if (_1628_) REG__2_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__29_  */
always_ff @(posedge clk)
if (_1626_) REG__29_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__28_  */
always_ff @(posedge clk)
if (_1624_) REG__28_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__27_  */
always_ff @(posedge clk)
if (_1622_) REG__27_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__26_  */
always_ff @(posedge clk)
if (_1620_) REG__26_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__25_  */
always_ff @(posedge clk)
if (_1618_) REG__25_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__24_  */
always_ff @(posedge clk)
if (_1616_) REG__24_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__23_  */
always_ff @(posedge clk)
if (_1614_) REG__23_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__22_  */
always_ff @(posedge clk)
if (_1612_) REG__22_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__21_  */
always_ff @(posedge clk)
if (_1610_) REG__21_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__20_  */
always_ff @(posedge clk)
if (_1608_) REG__20_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__1_  */
always_ff @(posedge clk)
if (_1606_) REG__1_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__19_  */
always_ff @(posedge clk)
if (_1604_) REG__19_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__18_  */
always_ff @(posedge clk)
if (_1602_) REG__18_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__17_  */
always_ff @(posedge clk)
if (_1600_) REG__17_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__16_  */
always_ff @(posedge clk)
if (_1598_) REG__16_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__15_  */
always_ff @(posedge clk)
if (_1596_) REG__15_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__14_  */
always_ff @(posedge clk)
if (_1594_) REG__14_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__13_  */
always_ff @(posedge clk)
if (_1592_) REG__13_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__12_  */
always_ff @(posedge clk)
if (_1590_) REG__12_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__11_  */
always_ff @(posedge clk)
if (_1588_) REG__11_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__10_  */
always_ff @(posedge clk)
if (_1586_) REG__10_  <= _0002_;
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME REG__0_  */
always_ff @(posedge clk)
if (_1584_) REG__0_  <= _0002_;
assign _0261_ = _1411_ & _1450_;
assign _0264_ = instr_vld_t0 & instr_rdy;
assign _0267_ = regwr_en_t0 & _1422_;
assign _0270_ = regwr_en_t0 & _1426_;
assign _0273_ = reg_vld_t0 & regwr_en;
assign _0276_ = reg_vld_t0 & fetch_rdy;
assign _0262_ = _1451_ & _1410_;
assign _0265_ = instr_rdy_t0 & instr_vld;
assign _0268_ = _1423_ & regwr_en;
assign _0271_ = _1427_ & regwr_en;
assign _0274_ = regwr_en_t0 & reg_vld;
assign _0263_ = _1411_ & _1451_;
assign _0266_ = instr_vld_t0 & instr_rdy_t0;
assign _0269_ = regwr_en_t0 & _1423_;
assign _0272_ = regwr_en_t0 & _1427_;
assign _0275_ = reg_vld_t0 & regwr_en_t0;
assign _0930_ = _0261_ | _0262_;
assign _0931_ = _0264_ | _0265_;
assign _0932_ = _0267_ | _0268_;
assign _0933_ = _0270_ | _0271_;
assign _0934_ = _0273_ | _0274_;
assign _0935_ = _0276_ | _0277_;
assign csr_regrd_t0 = _0930_ | _0263_;
assign _1433_ = _0931_ | _0266_;
assign _1435_ = _0932_ | _0269_;
assign _1437_ = _0933_ | _0272_;
assign _1439_ = _0934_ | _0275_;
assign _1441_ = _0935_ | _0278_;
assign _0129_ = | { _1441_, _1439_, _1433_ };
assign _0135_ = | instr_data_t0[19:15];
assign _0137_ = | instr_data_t0[24:20];
assign _0034_ = ~ { _1441_, _1439_, _1433_ };
assign _0037_ = ~ instr_data_t0[19:15];
assign _0039_ = ~ instr_data_t0[24:20];
assign _0248_ = { _1440_, _1438_, _1432_ } & _0034_;
assign _0251_ = instr_data[19:15] & _0037_;
assign _0254_ = instr_data[24:20] & _0039_;
assign _0141_ = ! _0245_;
assign _0142_ = ! _0248_;
assign _0143_ = ! _0249_;
assign _0144_ = ! _0251_;
assign _0145_ = ! _0254_;
assign _0014_ = _0141_ & _0126_;
assign _0020_ = _0142_ & _0129_;
assign _1405_ = _0143_ & _0133_;
assign _1421_ = _0144_ & _0135_;
assign _1425_ = _0145_ & _0137_;
assign _0045_ = ~ _1442_;
assign _0047_ = ~ _1406_;
assign _0051_ = ~ format_U;
assign _0052_ = ~ _1412_;
assign _0054_ = ~ _1448_;
assign _0043_ = ~ _1400_;
assign _0057_ = ~ _1452_;
assign _0058_ = ~ _1454_;
assign _0060_ = ~ _1456_;
assign _0061_ = ~ _1458_;
assign _0063_ = ~ _1460_;
assign _0056_ = ~ _1418_;
assign _0065_ = ~ _1462_;
assign _0048_ = ~ _1408_;
assign _0050_ = ~ format_J;
assign _0053_ = ~ _1414_;
assign _0055_ = ~ _1416_;
assign _0044_ = ~ _1402_;
assign _0046_ = ~ _1404_;
assign _0064_ = ~ csr_regrd;
assign _0059_ = ~ format_B;
assign _0279_ = _1401_ & _0044_;
assign _0282_ = _1443_ & _0046_;
assign _0285_ = _1407_ & _0048_;
assign _0288_ = format_I_t0 & _0050_;
assign _0291_ = format_U_t0 & _0050_;
assign _0294_ = _1413_ & _0053_;
assign _0297_ = _1449_ & _0055_;
assign _0300_ = _1401_ & _0056_;
assign _0303_ = _1453_ & _0044_;
assign _0306_ = _1455_ & _0059_;
assign _0309_ = _1457_ & _0046_;
assign _0312_ = _1459_ & _0062_;
assign _0315_ = _1461_ & _0064_;
assign _0318_ = _1419_ & _0059_;
assign _0321_ = _1463_ & _0062_;
assign _0280_ = _1403_ & _0043_;
assign _0283_ = _1405_ & _0045_;
assign _0286_ = _1409_ & _0047_;
assign _0289_ = format_J_t0 & _0049_;
assign _0292_ = format_J_t0 & _0051_;
assign _0295_ = _1415_ & _0052_;
assign _0298_ = _1417_ & _0054_;
assign _0301_ = _1419_ & _0043_;
assign _0304_ = _1403_ & _0057_;
assign _0307_ = format_B_t0 & _0058_;
assign _0310_ = _1405_ & _0060_;
assign _0313_ = format_S_t0 & _0061_;
assign _0316_ = csr_regrd_t0 & _0063_;
assign _0319_ = format_B_t0 & _0056_;
assign _0322_ = format_S_t0 & _0065_;
assign _0281_ = _1401_ & _1403_;
assign _0284_ = _1443_ & _1405_;
assign _0287_ = _1407_ & _1409_;
assign _0290_ = format_I_t0 & format_J_t0;
assign _0293_ = format_U_t0 & format_J_t0;
assign _0296_ = _1413_ & _1415_;
assign _0299_ = _1449_ & _1417_;
assign _0302_ = _1401_ & _1419_;
assign _0305_ = _1453_ & _1403_;
assign _0308_ = _1455_ & format_B_t0;
assign _0311_ = _1457_ & _1405_;
assign _0314_ = _1459_ & format_S_t0;
assign _0317_ = _1461_ & csr_regrd_t0;
assign _0320_ = _1419_ & format_B_t0;
assign _0323_ = _1463_ & format_S_t0;
assign _0936_ = _0279_ | _0280_;
assign _0937_ = _0282_ | _0283_;
assign _0938_ = _0285_ | _0286_;
assign _0939_ = _0288_ | _0289_;
assign _0940_ = _0291_ | _0292_;
assign _0941_ = _0294_ | _0295_;
assign _0942_ = _0297_ | _0298_;
assign _0943_ = _0300_ | _0301_;
assign _0944_ = _0303_ | _0304_;
assign _0945_ = _0306_ | _0307_;
assign _0946_ = _0309_ | _0310_;
assign _0947_ = _0312_ | _0313_;
assign _0948_ = _0315_ | _0316_;
assign _0949_ = _0318_ | _0319_;
assign _0950_ = _0321_ | _0322_;
assign _1443_ = _0936_ | _0281_;
assign format_I_t0 = _0937_ | _0284_;
assign format_U_t0 = _0938_ | _0287_;
assign _1445_ = _0939_ | _0290_;
assign _1447_ = _0940_ | _0293_;
assign _1449_ = _0941_ | _0296_;
assign _1451_ = _0942_ | _0299_;
assign _1453_ = _0943_ | _0302_;
assign _1455_ = _0944_ | _0305_;
assign _1457_ = _0945_ | _0308_;
assign _1459_ = _0946_ | _0311_;
assign _1461_ = _0947_ | _0314_;
assign is_regrd_rs1_en_t0 = _0948_ | _0317_;
assign _1463_ = _0949_ | _0320_;
assign is_regrd_rs2_en_t0 = _0950_ | _0323_;
assign _1395_ = ~ _0000_[0];
assign _1396_ = ~ _0000_[1];
assign _1397_ = ~ _0000_[2];
assign _1398_ = ~ _0000_[3];
assign _1399_ = ~ _0000_[4];
assign _0643_ = _1395_ & _1396_;
assign _0645_ = _1398_ & _1399_;
assign _0647_ = _1397_ & _0645_;
assign _0649_ = _0643_ & _0647_;
assign _0651_ = _0000_[0] & _1396_;
assign _0653_ = _0651_ & _0647_;
assign _0655_ = _1395_ & _0000_[1];
assign _0657_ = _0655_ & _0647_;
assign _0659_ = _0000_[0] & _0000_[1];
assign _0661_ = _0659_ & _0647_;
assign _0663_ = _0000_[2] & _0645_;
assign _0665_ = _0643_ & _0663_;
assign _0667_ = _0651_ & _0663_;
assign _0669_ = _0655_ & _0663_;
assign _0671_ = _0659_ & _0663_;
assign _0673_ = _0000_[3] & _1399_;
assign _0675_ = _1397_ & _0673_;
assign _0677_ = _0643_ & _0675_;
assign _0679_ = _0651_ & _0675_;
assign _0681_ = _0655_ & _0675_;
assign _0683_ = _0659_ & _0675_;
assign _0685_ = _0000_[2] & _0673_;
assign _0687_ = _0643_ & _0685_;
assign _0689_ = _0651_ & _0685_;
assign _0691_ = _0655_ & _0685_;
assign _0693_ = _0659_ & _0685_;
assign _0695_ = _1398_ & _0000_[4];
assign _0697_ = _1397_ & _0695_;
assign _0699_ = _0643_ & _0697_;
assign _0701_ = _0651_ & _0697_;
assign _0703_ = _0655_ & _0697_;
assign _0705_ = _0659_ & _0697_;
assign _0707_ = _0000_[2] & _0695_;
assign _0709_ = _0643_ & _0707_;
assign _0711_ = _0651_ & _0707_;
assign _0713_ = _0655_ & _0707_;
assign _0715_ = _0659_ & _0707_;
assign _0717_ = _0000_[3] & _0000_[4];
assign _0719_ = _1397_ & _0717_;
assign _0721_ = _0643_ & _0719_;
assign _0723_ = _0651_ & _0719_;
assign _0725_ = _0655_ & _0719_;
assign _0727_ = _0659_ & _0719_;
assign _0729_ = _0000_[2] & _0717_;
assign _0731_ = _0643_ & _0729_;
assign _0733_ = _0651_ & _0729_;
assign _0735_ = _0655_ & _0729_;
assign _0737_ = _0659_ & _0729_;
assign _0066_ = ~ { instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24] };
assign _0067_ = ~ { instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23] };
assign _0068_ = ~ { instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22] };
assign _0069_ = ~ { instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21] };
assign _0070_ = ~ { instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20] };
assign _0071_ = ~ { instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19] };
assign _0072_ = ~ { instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18] };
assign _0073_ = ~ { instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17] };
assign _0074_ = ~ { instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16] };
assign _0075_ = ~ { instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15] };
assign _0077_ = ~ { _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_ };
assign _0078_ = ~ { _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_ };
assign _0079_ = ~ { _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_ };
assign _0080_ = ~ { _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_ };
assign _0081_ = ~ { _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_ };
assign _0082_ = ~ { format_U, format_U, format_U, format_U, format_U, format_U, format_U, format_U, format_U, format_U, format_U, format_U };
assign _0083_ = ~ { _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_ };
assign _0084_ = ~ { _1444_, _1444_, _1444_, _1444_ };
assign _0062_ = ~ format_S;
assign _0049_ = ~ format_I;
assign _0951_ = { instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24] } | _0066_;
assign _0954_ = { instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23] } | _0067_;
assign _0958_ = { instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22] } | _0068_;
assign _0964_ = { instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21] } | _0069_;
assign _0974_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } | _0070_;
assign _0992_ = { instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19] } | _0071_;
assign _0995_ = { instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18] } | _0072_;
assign _0999_ = { instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17] } | _0073_;
assign _1005_ = { instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16] } | _0074_;
assign _1015_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } | _0075_;
assign _1070_ = { _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_ } | _0077_;
assign _1073_ = { _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_ } | _0078_;
assign _1074_ = { _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_ } | _0079_;
assign _1078_ = { _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_ } | _0080_;
assign _1081_ = { _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_ } | _0081_;
assign _1083_ = { format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0 } | _0082_;
assign _1086_ = { _1447_, _1447_, _1447_, _1447_, _1447_, _1447_, _1447_, _1447_ } | _0083_;
assign _1089_ = format_J_t0 | _0050_;
assign _1092_ = format_B_t0 | _0059_;
assign _1095_ = { _1445_, _1445_, _1445_, _1445_ } | _0084_;
assign _1099_ = format_I_t0 | _0049_;
assign _0952_ = { instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24] } | { instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24], instr_data[24] };
assign _0955_ = { instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23] } | { instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23], instr_data[23] };
assign _0959_ = { instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22] } | { instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22], instr_data[22] };
assign _0965_ = { instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21] } | { instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21], instr_data[21] };
assign _0975_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } | { instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20], instr_data[20] };
assign _0993_ = { instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19] } | { instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19], instr_data[19] };
assign _0996_ = { instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18] } | { instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18], instr_data[18] };
assign _1000_ = { instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17] } | { instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17], instr_data[17] };
assign _1006_ = { instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16] } | { instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16], instr_data[16] };
assign _1016_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } | { instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15], instr_data[15] };
assign _1066_ = { regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0 } | { regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en, regwr_en };
assign _1067_ = { regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0, regwr_en_t0 } | { regwr_en, regwr_en, regwr_en, regwr_en, regwr_en };
assign _1068_ = { _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_ } | { _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_, _1430_ };
assign _1071_ = { _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_ } | { _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_, _1436_ };
assign _1075_ = { _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_ } | { _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_ };
assign _1077_ = { _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_, _1429_ } | { _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_ };
assign _1069_ = { _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_, _1439_ } | { _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_ };
assign _1079_ = { _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_ } | { _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_ };
assign _1084_ = { format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0 } | { format_U, format_U, format_U, format_U, format_U, format_U, format_U, format_U, format_U, format_U, format_U, format_U };
assign _1087_ = { _1447_, _1447_, _1447_, _1447_, _1447_, _1447_, _1447_, _1447_ } | { _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_ };
assign _1090_ = format_J_t0 | format_J;
assign _1093_ = format_B_t0 | format_B;
assign _1096_ = { _1445_, _1445_, _1445_, _1445_ } | { _1444_, _1444_, _1444_, _1444_ };
assign _1098_ = format_S_t0 | format_S;
assign _1100_ = format_I_t0 | format_I;
assign _0324_ = _1465_ & _0951_;
assign _0327_ = _1469_ & _0954_;
assign _0330_ = _1473_ & _0954_;
assign _0333_ = _1477_ & _0958_;
assign _0336_ = _1481_ & _0958_;
assign _0339_ = _1485_ & _0958_;
assign _0342_ = _1489_ & _0958_;
assign _0345_ = _1493_ & _0964_;
assign _0348_ = _1497_ & _0964_;
assign _0351_ = _1501_ & _0964_;
assign _0354_ = _1505_ & _0964_;
assign _0357_ = _1509_ & _0964_;
assign _0360_ = _1513_ & _0964_;
assign _0363_ = _1517_ & _0964_;
assign _0366_ = _1521_ & _0964_;
assign _0369_ = REG__0__t0  & _0974_;
assign _0372_ = REG__20__t0  & _0974_;
assign _0375_ = REG__22__t0  & _0974_;
assign _0378_ = REG__24__t0  & _0974_;
assign _0381_ = REG__26__t0  & _0974_;
assign _0384_ = REG__28__t0  & _0974_;
assign _0387_ = REG__30__t0  & _0974_;
assign _0390_ = REG__2__t0  & _0974_;
assign _0393_ = REG__4__t0  & _0974_;
assign _0396_ = REG__6__t0  & _0974_;
assign _0399_ = REG__8__t0  & _0974_;
assign _0402_ = REG__10__t0  & _0974_;
assign _0405_ = REG__12__t0  & _0974_;
assign _0408_ = REG__14__t0  & _0974_;
assign _0411_ = REG__16__t0  & _0974_;
assign _0414_ = REG__18__t0  & _0974_;
assign _0417_ = _1525_ & _0992_;
assign _0420_ = _1529_ & _0995_;
assign _0423_ = _1533_ & _0995_;
assign _0426_ = _1537_ & _0999_;
assign _0429_ = _1541_ & _0999_;
assign _0432_ = _1545_ & _0999_;
assign _0435_ = _1549_ & _0999_;
assign _0438_ = _1553_ & _1005_;
assign _0441_ = _1557_ & _1005_;
assign _0444_ = _1561_ & _1005_;
assign _0447_ = _1565_ & _1005_;
assign _0450_ = _1569_ & _1005_;
assign _0453_ = _1573_ & _1005_;
assign _0456_ = _1577_ & _1005_;
assign _0459_ = _1581_ & _1005_;
assign _0462_ = REG__0__t0  & _1015_;
assign _0465_ = REG__20__t0  & _1015_;
assign _0468_ = REG__22__t0  & _1015_;
assign _0471_ = REG__24__t0  & _1015_;
assign _0474_ = REG__26__t0  & _1015_;
assign _0477_ = REG__28__t0  & _1015_;
assign _0480_ = REG__30__t0  & _1015_;
assign _0483_ = REG__2__t0  & _1015_;
assign _0486_ = REG__4__t0  & _1015_;
assign _0489_ = REG__6__t0  & _1015_;
assign _0492_ = REG__8__t0  & _1015_;
assign _0495_ = REG__10__t0  & _1015_;
assign _0498_ = REG__12__t0  & _1015_;
assign _0501_ = REG__14__t0  & _1015_;
assign _0504_ = REG__16__t0  & _1015_;
assign _0507_ = REG__18__t0  & _1015_;
assign _0607_ = _1651_ & _1070_;
assign _0610_ = _1661_ & _1073_;
assign _0612_ = _1660_ & _1074_;
assign _0615_ = _1649_ & _1078_;
assign _0618_ = _1670_ & _1081_;
assign _0620_ = _1669_ & _1074_;
assign _0623_ = { instr_data_t0[31], instr_data_t0[31], instr_data_t0[31], instr_data_t0[31], instr_data_t0[31], instr_data_t0[31], instr_data_t0[31], instr_data_t0[31], instr_data_t0[31], instr_data_t0[31], instr_data_t0[31], instr_data_t0[31] } & _1083_;
assign _0626_ = { instr_data_t0[31], instr_data_t0[31], instr_data_t0[31], instr_data_t0[31], instr_data_t0[31], instr_data_t0[31], instr_data_t0[31], instr_data_t0[31] } & _1086_;
assign _0629_ = instr_data_t0[31] & _1089_;
assign _0632_ = _0012_ & _1092_;
assign _0635_ = instr_data_t0[11:8] & _1095_;
assign _0640_ = _0006_ & _1099_;
assign _0325_ = _1467_ & _0952_;
assign _0328_ = _1471_ & _0955_;
assign _0331_ = _1475_ & _0955_;
assign _0334_ = _1479_ & _0959_;
assign _0337_ = _1483_ & _0959_;
assign _0340_ = _1487_ & _0959_;
assign _0343_ = _1491_ & _0959_;
assign _0346_ = _1495_ & _0965_;
assign _0349_ = _1499_ & _0965_;
assign _0352_ = _1503_ & _0965_;
assign _0355_ = _1507_ & _0965_;
assign _0358_ = _1511_ & _0965_;
assign _0361_ = _1515_ & _0965_;
assign _0364_ = _1519_ & _0965_;
assign _0367_ = _1523_ & _0965_;
assign _0370_ = REG__1__t0  & _0975_;
assign _0373_ = REG__21__t0  & _0975_;
assign _0376_ = REG__23__t0  & _0975_;
assign _0379_ = REG__25__t0  & _0975_;
assign _0382_ = REG__27__t0  & _0975_;
assign _0385_ = REG__29__t0  & _0975_;
assign _0388_ = REG__31__t0  & _0975_;
assign _0391_ = REG__3__t0  & _0975_;
assign _0394_ = REG__5__t0  & _0975_;
assign _0397_ = REG__7__t0  & _0975_;
assign _0400_ = REG__9__t0  & _0975_;
assign _0403_ = REG__11__t0  & _0975_;
assign _0406_ = REG__13__t0  & _0975_;
assign _0409_ = REG__15__t0  & _0975_;
assign _0412_ = REG__17__t0  & _0975_;
assign _0415_ = REG__19__t0  & _0975_;
assign _0418_ = _1527_ & _0993_;
assign _0421_ = _1531_ & _0996_;
assign _0424_ = _1535_ & _0996_;
assign _0427_ = _1539_ & _1000_;
assign _0430_ = _1543_ & _1000_;
assign _0433_ = _1547_ & _1000_;
assign _0436_ = _1551_ & _1000_;
assign _0439_ = _1555_ & _1006_;
assign _0442_ = _1559_ & _1006_;
assign _0445_ = _1563_ & _1006_;
assign _0448_ = _1567_ & _1006_;
assign _0451_ = _1571_ & _1006_;
assign _0454_ = _1575_ & _1006_;
assign _0457_ = _1579_ & _1006_;
assign _0460_ = _1583_ & _1006_;
assign _0463_ = REG__1__t0  & _1016_;
assign _0466_ = REG__21__t0  & _1016_;
assign _0469_ = REG__23__t0  & _1016_;
assign _0472_ = REG__25__t0  & _1016_;
assign _0475_ = REG__27__t0  & _1016_;
assign _0478_ = REG__29__t0  & _1016_;
assign _0481_ = REG__31__t0  & _1016_;
assign _0484_ = REG__3__t0  & _1016_;
assign _0487_ = REG__5__t0  & _1016_;
assign _0490_ = REG__7__t0  & _1016_;
assign _0493_ = REG__9__t0  & _1016_;
assign _0496_ = REG__11__t0  & _1016_;
assign _0499_ = REG__13__t0  & _1016_;
assign _0502_ = REG__15__t0  & _1016_;
assign _0505_ = REG__17__t0  & _1016_;
assign _0508_ = REG__19__t0  & _1016_;
assign _0003_ = regwr_data_t0 & _1066_;
assign _0001_ = regwr_sel_t0 & _1067_;
assign _1658_ = regwr_data_t0 & _1068_;
assign _1660_ = _1658_ & _1069_;
assign _0608_ = regwr_data_t0 & _1071_;
assign _0613_ = _1663_ & _1075_;
assign _1667_ = regwr_data_t0 & _1077_;
assign _1669_ = _1667_ & _1069_;
assign _0616_ = regwr_data_t0 & _1079_;
assign _0621_ = _1672_ & _1075_;
assign _0624_ = instr_data_t0[31:20] & _1084_;
assign _0627_ = instr_data_t0[19:12] & _1087_;
assign _0630_ = instr_data_t0[20] & _1090_;
assign _0633_ = instr_data_t0[7] & _1093_;
assign _0636_ = instr_data_t0[24:21] & _1096_;
assign _0638_ = instr_data_t0[7] & _1098_;
assign _0641_ = instr_data_t0[20] & _1100_;
assign _0953_ = _0324_ | _0325_;
assign _0956_ = _0327_ | _0328_;
assign _0957_ = _0330_ | _0331_;
assign _0960_ = _0333_ | _0334_;
assign _0961_ = _0336_ | _0337_;
assign _0962_ = _0339_ | _0340_;
assign _0963_ = _0342_ | _0343_;
assign _0966_ = _0345_ | _0346_;
assign _0967_ = _0348_ | _0349_;
assign _0968_ = _0351_ | _0352_;
assign _0969_ = _0354_ | _0355_;
assign _0970_ = _0357_ | _0358_;
assign _0971_ = _0360_ | _0361_;
assign _0972_ = _0363_ | _0364_;
assign _0973_ = _0366_ | _0367_;
assign _0976_ = _0369_ | _0370_;
assign _0977_ = _0372_ | _0373_;
assign _0978_ = _0375_ | _0376_;
assign _0979_ = _0378_ | _0379_;
assign _0980_ = _0381_ | _0382_;
assign _0981_ = _0384_ | _0385_;
assign _0982_ = _0387_ | _0388_;
assign _0983_ = _0390_ | _0391_;
assign _0984_ = _0393_ | _0394_;
assign _0985_ = _0396_ | _0397_;
assign _0986_ = _0399_ | _0400_;
assign _0987_ = _0402_ | _0403_;
assign _0988_ = _0405_ | _0406_;
assign _0989_ = _0408_ | _0409_;
assign _0990_ = _0411_ | _0412_;
assign _0991_ = _0414_ | _0415_;
assign _0994_ = _0417_ | _0418_;
assign _0997_ = _0420_ | _0421_;
assign _0998_ = _0423_ | _0424_;
assign _1001_ = _0426_ | _0427_;
assign _1002_ = _0429_ | _0430_;
assign _1003_ = _0432_ | _0433_;
assign _1004_ = _0435_ | _0436_;
assign _1007_ = _0438_ | _0439_;
assign _1008_ = _0441_ | _0442_;
assign _1009_ = _0444_ | _0445_;
assign _1010_ = _0447_ | _0448_;
assign _1011_ = _0450_ | _0451_;
assign _1012_ = _0453_ | _0454_;
assign _1013_ = _0456_ | _0457_;
assign _1014_ = _0459_ | _0460_;
assign _1017_ = _0462_ | _0463_;
assign _1018_ = _0465_ | _0466_;
assign _1019_ = _0468_ | _0469_;
assign _1020_ = _0471_ | _0472_;
assign _1021_ = _0474_ | _0475_;
assign _1022_ = _0477_ | _0478_;
assign _1023_ = _0480_ | _0481_;
assign _1024_ = _0483_ | _0484_;
assign _1025_ = _0486_ | _0487_;
assign _1026_ = _0489_ | _0490_;
assign _1027_ = _0492_ | _0493_;
assign _1028_ = _0495_ | _0496_;
assign _1029_ = _0498_ | _0499_;
assign _1030_ = _0501_ | _0502_;
assign _1031_ = _0504_ | _0505_;
assign _1032_ = _0507_ | _0508_;
assign _1072_ = _0607_ | _0608_;
assign _1076_ = _0612_ | _0613_;
assign _1080_ = _0615_ | _0616_;
assign _1082_ = _0620_ | _0621_;
assign _1085_ = _0623_ | _0624_;
assign _1088_ = _0626_ | _0627_;
assign _1091_ = _0629_ | _0630_;
assign _1094_ = _0632_ | _0633_;
assign _1097_ = _0635_ | _0636_;
assign _1101_ = _0640_ | _0641_;
assign _1277_ = _1464_ ^ _1466_;
assign _1278_ = _1468_ ^ _1470_;
assign _1279_ = _1472_ ^ _1474_;
assign _1280_ = _1476_ ^ _1478_;
assign _1281_ = _1480_ ^ _1482_;
assign _1282_ = _1484_ ^ _1486_;
assign _1283_ = _1488_ ^ _1490_;
assign _1284_ = _1492_ ^ _1494_;
assign _1285_ = _1496_ ^ _1498_;
assign _1286_ = _1500_ ^ _1502_;
assign _1287_ = _1504_ ^ _1506_;
assign _1288_ = _1508_ ^ _1510_;
assign _1289_ = _1512_ ^ _1514_;
assign _1290_ = _1516_ ^ _1518_;
assign _1291_ = _1520_ ^ _1522_;
assign _1308_ = _1524_ ^ _1526_;
assign _1309_ = _1528_ ^ _1530_;
assign _1310_ = _1532_ ^ _1534_;
assign _1311_ = _1536_ ^ _1538_;
assign _1312_ = _1540_ ^ _1542_;
assign _1313_ = _1544_ ^ _1546_;
assign _1314_ = _1548_ ^ _1550_;
assign _1315_ = _1552_ ^ _1554_;
assign _1316_ = _1556_ ^ _1558_;
assign _1317_ = _1560_ ^ _1562_;
assign _1318_ = _1564_ ^ _1566_;
assign _1319_ = _1568_ ^ _1570_;
assign _1320_ = _1572_ ^ _1574_;
assign _1321_ = _1576_ ^ _1578_;
assign _1322_ = _1580_ ^ _1582_;
assign _1292_ = REG__0_  ^ REG__1_ ;
assign _1293_ = REG__20_  ^ REG__21_ ;
assign _1294_ = REG__22_  ^ REG__23_ ;
assign _1295_ = REG__24_  ^ REG__25_ ;
assign _1296_ = REG__26_  ^ REG__27_ ;
assign _1297_ = REG__28_  ^ REG__29_ ;
assign _1298_ = REG__30_  ^ REG__31_ ;
assign _1299_ = REG__2_  ^ REG__3_ ;
assign _1300_ = REG__4_  ^ REG__5_ ;
assign _1301_ = REG__6_  ^ REG__7_ ;
assign _1302_ = REG__8_  ^ REG__9_ ;
assign _1303_ = REG__10_  ^ REG__11_ ;
assign _1304_ = REG__12_  ^ REG__13_ ;
assign _1305_ = REG__14_  ^ REG__15_ ;
assign _1306_ = REG__16_  ^ REG__17_ ;
assign _1307_ = REG__18_  ^ REG__19_ ;
assign _1323_ = _1650_ ^ regwr_data;
assign _1325_ = _1659_ ^ _1662_;
assign _1326_ = _1648_ ^ regwr_data;
assign _1328_ = _1668_ ^ _1671_;
assign _1329_ = { instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31] } ^ instr_data[31:20];
assign _1330_ = { instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31] } ^ instr_data[19:12];
assign _1331_ = instr_data[31] ^ instr_data[20];
assign _1332_ = _0011_ ^ instr_data[7];
assign _1333_ = instr_data[11:8] ^ instr_data[24:21];
assign _1334_ = _0005_ ^ instr_data[20];
assign _0326_ = { instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24], instr_data_t0[24] } & _1277_;
assign _0329_ = { instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23] } & _1278_;
assign _0332_ = { instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23], instr_data_t0[23] } & _1279_;
assign _0335_ = { instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22] } & _1280_;
assign _0338_ = { instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22] } & _1281_;
assign _0341_ = { instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22] } & _1282_;
assign _0344_ = { instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22], instr_data_t0[22] } & _1283_;
assign _0347_ = { instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21] } & _1284_;
assign _0350_ = { instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21] } & _1285_;
assign _0353_ = { instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21] } & _1286_;
assign _0356_ = { instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21] } & _1287_;
assign _0359_ = { instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21] } & _1288_;
assign _0362_ = { instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21] } & _1289_;
assign _0365_ = { instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21] } & _1290_;
assign _0368_ = { instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21], instr_data_t0[21] } & _1291_;
assign _0371_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } & _1292_;
assign _0374_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } & _1293_;
assign _0377_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } & _1294_;
assign _0380_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } & _1295_;
assign _0383_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } & _1296_;
assign _0386_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } & _1297_;
assign _0389_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } & _1298_;
assign _0392_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } & _1299_;
assign _0395_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } & _1300_;
assign _0398_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } & _1301_;
assign _0401_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } & _1302_;
assign _0404_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } & _1303_;
assign _0407_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } & _1304_;
assign _0410_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } & _1305_;
assign _0413_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } & _1306_;
assign _0416_ = { instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20], instr_data_t0[20] } & _1307_;
assign _0419_ = { instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19], instr_data_t0[19] } & _1308_;
assign _0422_ = { instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18] } & _1309_;
assign _0425_ = { instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18], instr_data_t0[18] } & _1310_;
assign _0428_ = { instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17] } & _1311_;
assign _0431_ = { instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17] } & _1312_;
assign _0434_ = { instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17] } & _1313_;
assign _0437_ = { instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17], instr_data_t0[17] } & _1314_;
assign _0440_ = { instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16] } & _1315_;
assign _0443_ = { instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16] } & _1316_;
assign _0446_ = { instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16] } & _1317_;
assign _0449_ = { instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16] } & _1318_;
assign _0452_ = { instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16] } & _1319_;
assign _0455_ = { instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16] } & _1320_;
assign _0458_ = { instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16] } & _1321_;
assign _0461_ = { instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16], instr_data_t0[16] } & _1322_;
assign _0464_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } & _1292_;
assign _0467_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } & _1293_;
assign _0470_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } & _1294_;
assign _0473_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } & _1295_;
assign _0476_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } & _1296_;
assign _0479_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } & _1297_;
assign _0482_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } & _1298_;
assign _0485_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } & _1299_;
assign _0488_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } & _1300_;
assign _0491_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } & _1301_;
assign _0494_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } & _1302_;
assign _0497_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } & _1303_;
assign _0500_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } & _1304_;
assign _0503_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } & _1305_;
assign _0506_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } & _1306_;
assign _0509_ = { instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15], instr_data_t0[15] } & _1307_;
assign _1656_ = _1433_ & _0085_;
assign _0609_ = { _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_ } & _1323_;
assign _0611_ = { _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_, _1425_ } & _1324_;
assign _0614_ = { _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_ } & _1325_;
assign _0617_ = { _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_, _1435_ } & _1326_;
assign _0619_ = { _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_, _1421_ } & _1327_;
assign _0622_ = { _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_ } & _1328_;
assign _0625_ = { format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0, format_U_t0 } & _1329_;
assign _0628_ = { _1447_, _1447_, _1447_, _1447_, _1447_, _1447_, _1447_, _1447_ } & _1330_;
assign _0631_ = format_J_t0 & _1331_;
assign _0634_ = format_B_t0 & _1332_;
assign _0637_ = { _1445_, _1445_, _1445_, _1445_ } & _1333_;
assign _0639_ = format_S_t0 & instr_data[7];
assign _0642_ = format_I_t0 & _1334_;
assign _1651_ = _0326_ | _0953_;
assign _1465_ = _0329_ | _0956_;
assign _1467_ = _0332_ | _0957_;
assign _1469_ = _0335_ | _0960_;
assign _1471_ = _0338_ | _0961_;
assign _1473_ = _0341_ | _0962_;
assign _1475_ = _0344_ | _0963_;
assign _1477_ = _0347_ | _0966_;
assign _1479_ = _0350_ | _0967_;
assign _1481_ = _0353_ | _0968_;
assign _1483_ = _0356_ | _0969_;
assign _1485_ = _0359_ | _0970_;
assign _1487_ = _0362_ | _0971_;
assign _1489_ = _0365_ | _0972_;
assign _1491_ = _0368_ | _0973_;
assign _1493_ = _0371_ | _0976_;
assign _1513_ = _0374_ | _0977_;
assign _1515_ = _0377_ | _0978_;
assign _1517_ = _0380_ | _0979_;
assign _1519_ = _0383_ | _0980_;
assign _1521_ = _0386_ | _0981_;
assign _1523_ = _0389_ | _0982_;
assign _1495_ = _0392_ | _0983_;
assign _1497_ = _0395_ | _0984_;
assign _1499_ = _0398_ | _0985_;
assign _1501_ = _0401_ | _0986_;
assign _1503_ = _0404_ | _0987_;
assign _1505_ = _0407_ | _0988_;
assign _1507_ = _0410_ | _0989_;
assign _1509_ = _0413_ | _0990_;
assign _1511_ = _0416_ | _0991_;
assign _1649_ = _0419_ | _0994_;
assign _1525_ = _0422_ | _0997_;
assign _1527_ = _0425_ | _0998_;
assign _1529_ = _0428_ | _1001_;
assign _1531_ = _0431_ | _1002_;
assign _1533_ = _0434_ | _1003_;
assign _1535_ = _0437_ | _1004_;
assign _1537_ = _0440_ | _1007_;
assign _1539_ = _0443_ | _1008_;
assign _1541_ = _0446_ | _1009_;
assign _1543_ = _0449_ | _1010_;
assign _1545_ = _0452_ | _1011_;
assign _1547_ = _0455_ | _1012_;
assign _1549_ = _0458_ | _1013_;
assign _1551_ = _0461_ | _1014_;
assign _1553_ = _0464_ | _1017_;
assign _1573_ = _0467_ | _1018_;
assign _1575_ = _0470_ | _1019_;
assign _1577_ = _0473_ | _1020_;
assign _1579_ = _0476_ | _1021_;
assign _1581_ = _0479_ | _1022_;
assign _1583_ = _0482_ | _1023_;
assign _1555_ = _0485_ | _1024_;
assign _1557_ = _0488_ | _1025_;
assign _1559_ = _0491_ | _1026_;
assign _1561_ = _0494_ | _1027_;
assign _1563_ = _0497_ | _1028_;
assign _1565_ = _0500_ | _1029_;
assign _1567_ = _0503_ | _1030_;
assign _1569_ = _0506_ | _1031_;
assign _1571_ = _0509_ | _1032_;
assign _1661_ = _0609_ | _1072_;
assign _1663_ = _0611_ | _0610_;
assign _1665_ = _0614_ | _1076_;
assign _1670_ = _0617_ | _1080_;
assign _1672_ = _0619_ | _0618_;
assign _1674_ = _0622_ | _1082_;
assign ImmF_t0 = _0625_ | _1085_;
assign ImmE_t0 = _0628_ | _1088_;
assign _0012_ = _0631_ | _1091_;
assign _0010_ = _0634_ | _1094_;
assign _0008_ = _0637_ | _1097_;
assign _0006_ = _0639_ | _0638_;
assign ImmA_t0 = _0642_ | _1101_;
assign _0013_ = | { _1438_, _1432_ };
assign _0015_ = { _1428_, _1438_, _1432_ } != 3'h2;
assign _0017_ = { _1430_, _1438_, _1432_ } != 3'h2;
assign _0019_ = | { _1440_, _1438_, _1432_ };
assign _0021_ = { _1438_, _1432_ } != 2'h2;
assign _0023_ = & { _0015_, _0013_, rstz };
assign _0025_ = & { _0013_, _0017_, rstz };
assign _0027_ = & { _1432_, rstz };
assign _0029_ = & { _0019_, _0021_ };
assign _0085_ = ~ _1654_;
assign _0076_ = ~ fetch_rdy;
assign _0606_ = reg_vld_t0 & _0076_;
assign _0277_ = fetch_rdy_t0 & reg_vld;
assign _0278_ = reg_vld_t0 & fetch_rdy_t0;
assign _1065_ = _0606_ | _0277_;
assign instr_rdy_t0 = _1065_ | _0278_;
assign _0130_ = | { _0016_, _0014_ };
assign _0131_ = | { _0018_, _0014_ };
assign _0132_ = | { _0022_, _0020_ };
assign _0922_ = { _0015_, _0013_, rstz } | { _0016_, _0014_, 1'h0 };
assign _0923_ = { _0013_, _0017_, rstz } | { _0014_, _0018_, 1'h0 };
assign _0924_ = { _1432_, rstz } | { _1433_, 1'h0 };
assign _0925_ = { _0019_, _0021_ } | { _0020_, _0022_ };
assign _0122_ = & _0922_;
assign _0123_ = & _0923_;
assign _0124_ = & _0924_;
assign _0125_ = & _0925_;
assign _0024_ = _0130_ & _0122_;
assign _0026_ = _0131_ & _0123_;
assign _0028_ = _1433_ & _0124_;
assign _0030_ = _0132_ & _0125_;
assign _1342_ = { _0009_, instr_data[30:25], _0007_ } ^ immediate[11:1];
assign _1130_ = { _0010_, instr_data_t0[30:25], _0008_ } | immediate_t0[11:1];
assign _1131_ = _1342_ | _1130_;
assign _0760_ = { _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_ } & { _0010_, instr_data_t0[30:25], _0008_ };
assign _0761_ = { _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_, _0088_ } & immediate_t0[11:1];
assign _0762_ = _1131_ & { _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_ };
assign _1132_ = _0760_ | _0761_;
assign _1133_ = _1132_ | _0762_;
reg [10:0] _3286_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME _3286_ */
always_ff @(posedge clk)
if (format_U) _3286_ <= 11'h000;
else _3286_ <= _1133_;
assign immediate_t0[11:1] = _3286_;
assign _0089_ = ~ _0029_;
assign _1339_ = _1655_ ^ reg_vld;
assign _1118_ = _1656_ | reg_vld_t0;
assign _1119_ = _1339_ | _1118_;
assign _0751_ = _0029_ & _1656_;
assign _0752_ = _0089_ & reg_vld_t0;
assign _0753_ = _1119_ & _0030_;
assign _1120_ = _0751_ | _0752_;
assign _1121_ = _1120_ | _0753_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_RF */
/* PC_TAINT_INFO STATE_NAME reg_vld_t0 */
always_ff @(posedge clk)
if (!rstz) reg_vld_t0 <= 1'h0;
else reg_vld_t0 <= _1121_;
assign format_J = instr_data[6:2] == /* src = "generated/sv2v_out.v:1551.14-1551.42" */ 5'h1b;
assign _1406_ = instr_data[6:2] == /* src = "generated/sv2v_out.v:1554.15-1554.43" */ 5'h0d;
assign _1408_ = instr_data[6:2] == /* src = "generated/sv2v_out.v:1554.49-1554.79" */ 5'h05;
assign _1410_ = instr_data[6:2] == /* src = "generated/sv2v_out.v:1590.22-1590.50" */ 5'h1c;
assign _1412_ = instr_data[14:12] == /* src = "generated/sv2v_out.v:1590.58-1590.74" */ 3'h1;
assign _1414_ = instr_data[14:12] == /* src = "generated/sv2v_out.v:1590.80-1590.96" */ 3'h2;
assign _1416_ = instr_data[14:12] == /* src = "generated/sv2v_out.v:1590.103-1590.119" */ 3'h3;
assign _1400_ = instr_data[6:2] == /* src = "generated/sv2v_out.v:1592.33-1592.63" */ 5'h04;
assign _1402_ = instr_data[6:2] == /* src = "generated/sv2v_out.v:1592.103-1592.132" */ 5'h19;
assign _1404_ = ! /* src = "generated/sv2v_out.v:1592.173-1592.202" */ instr_data[6:2];
assign _1418_ = instr_data[6:2] == /* src = "generated/sv2v_out.v:1593.29-1593.56" */ 5'h0c;
assign format_B = instr_data[6:2] == /* src = "generated/sv2v_out.v:1593.62-1593.89" */ 5'h18;
assign format_S = instr_data[6:2] == /* src = "generated/sv2v_out.v:1593.96-1593.126" */ 5'h08;
assign _1420_ = ! /* src = "generated/sv2v_out.v:1601.8-1601.16" */ instr_data[19:15];
assign _1422_ = instr_data[19:15] == /* src = "generated/sv2v_out.v:1603.26-1603.42" */ regwr_sel;
assign _1424_ = ! /* src = "generated/sv2v_out.v:1607.8-1607.16" */ instr_data[24:20];
assign _1426_ = instr_data[24:20] == /* src = "generated/sv2v_out.v:1609.26-1609.42" */ regwr_sel;
assign _1428_ = reg_rs1 == /* src = "generated/sv2v_out.v:1619.8-1619.28" */ regwr_sel;
assign _1430_ = reg_rs2 == /* src = "generated/sv2v_out.v:1621.8-1621.28" */ regwr_sel;
assign csr_regrd = _1410_ && /* src = "generated/sv2v_out.v:1590.21-1590.121" */ _1450_;
assign _1432_ = instr_vld && /* src = "generated/sv2v_out.v:1598.12-1598.34" */ instr_rdy;
assign _1434_ = regwr_en && /* src = "generated/sv2v_out.v:1603.13-1603.43" */ _1422_;
assign _1436_ = regwr_en && /* src = "generated/sv2v_out.v:1609.13-1609.43" */ _1426_;
assign _1438_ = reg_vld && /* src = "generated/sv2v_out.v:1618.12-1618.31" */ regwr_en;
assign _1440_ = reg_vld && /* src = "generated/sv2v_out.v:1624.12-1624.32" */ fetch_rdy;
assign _1442_ = _1400_ || /* src = "generated/sv2v_out.v:1550.15-1550.82" */ _1402_;
assign format_I = _1442_ || /* src = "generated/sv2v_out.v:1550.14-1550.118" */ _1404_;
assign format_U = _1406_ || /* src = "generated/sv2v_out.v:1554.14-1554.80" */ _1408_;
assign _1444_ = format_I || /* src = "generated/sv2v_out.v:1563.12-1563.32" */ format_J;
assign _1446_ = format_U || /* src = "generated/sv2v_out.v:1579.7-1579.27" */ format_J;
assign _1448_ = _1412_ || /* src = "generated/sv2v_out.v:1590.57-1590.97" */ _1414_;
assign _1450_ = _1448_ || /* src = "generated/sv2v_out.v:1590.56-1590.120" */ _1416_;
assign _1452_ = _1400_ || /* src = "generated/sv2v_out.v:1592.32-1592.97" */ _1418_;
assign _1454_ = _1452_ || /* src = "generated/sv2v_out.v:1592.31-1592.133" */ _1402_;
assign _1456_ = _1454_ || /* src = "generated/sv2v_out.v:1592.30-1592.167" */ format_B;
assign _1458_ = _1456_ || /* src = "generated/sv2v_out.v:1592.29-1592.203" */ _1404_;
assign _1460_ = _1458_ || /* src = "generated/sv2v_out.v:1592.28-1592.240" */ format_S;
assign is_regrd_rs1_en = _1460_ || /* src = "generated/sv2v_out.v:1592.27-1592.254" */ csr_regrd;
assign _1462_ = _1418_ || /* src = "generated/sv2v_out.v:1593.28-1593.90" */ format_B;
assign is_regrd_rs2_en = _1462_ || /* src = "generated/sv2v_out.v:1593.27-1593.127" */ format_S;
assign _1650_ = instr_data[24] ? _1466_ : _1464_;
assign _1464_ = instr_data[23] ? _1470_ : _1468_;
assign _1466_ = instr_data[23] ? _1474_ : _1472_;
assign _1468_ = instr_data[22] ? _1478_ : _1476_;
assign _1470_ = instr_data[22] ? _1482_ : _1480_;
assign _1472_ = instr_data[22] ? _1486_ : _1484_;
assign _1474_ = instr_data[22] ? _1490_ : _1488_;
assign _1476_ = instr_data[21] ? _1494_ : _1492_;
assign _1478_ = instr_data[21] ? _1498_ : _1496_;
assign _1480_ = instr_data[21] ? _1502_ : _1500_;
assign _1482_ = instr_data[21] ? _1506_ : _1504_;
assign _1484_ = instr_data[21] ? _1510_ : _1508_;
assign _1486_ = instr_data[21] ? _1514_ : _1512_;
assign _1488_ = instr_data[21] ? _1518_ : _1516_;
assign _1490_ = instr_data[21] ? _1522_ : _1520_;
assign _1492_ = instr_data[20] ? REG__1_  : REG__0_ ;
assign _1512_ = instr_data[20] ? REG__21_  : REG__20_ ;
assign _1514_ = instr_data[20] ? REG__23_  : REG__22_ ;
assign _1516_ = instr_data[20] ? REG__25_  : REG__24_ ;
assign _1518_ = instr_data[20] ? REG__27_  : REG__26_ ;
assign _1520_ = instr_data[20] ? REG__29_  : REG__28_ ;
assign _1522_ = instr_data[20] ? REG__31_  : REG__30_ ;
assign _1494_ = instr_data[20] ? REG__3_  : REG__2_ ;
assign _1496_ = instr_data[20] ? REG__5_  : REG__4_ ;
assign _1498_ = instr_data[20] ? REG__7_  : REG__6_ ;
assign _1500_ = instr_data[20] ? REG__9_  : REG__8_ ;
assign _1502_ = instr_data[20] ? REG__11_  : REG__10_ ;
assign _1504_ = instr_data[20] ? REG__13_  : REG__12_ ;
assign _1506_ = instr_data[20] ? REG__15_  : REG__14_ ;
assign _1508_ = instr_data[20] ? REG__17_  : REG__16_ ;
assign _1510_ = instr_data[20] ? REG__19_  : REG__18_ ;
assign _1648_ = instr_data[19] ? _1526_ : _1524_;
assign _1524_ = instr_data[18] ? _1530_ : _1528_;
assign _1526_ = instr_data[18] ? _1534_ : _1532_;
assign _1528_ = instr_data[17] ? _1538_ : _1536_;
assign _1530_ = instr_data[17] ? _1542_ : _1540_;
assign _1532_ = instr_data[17] ? _1546_ : _1544_;
assign _1534_ = instr_data[17] ? _1550_ : _1548_;
assign _1536_ = instr_data[16] ? _1554_ : _1552_;
assign _1538_ = instr_data[16] ? _1558_ : _1556_;
assign _1540_ = instr_data[16] ? _1562_ : _1560_;
assign _1542_ = instr_data[16] ? _1566_ : _1564_;
assign _1544_ = instr_data[16] ? _1570_ : _1568_;
assign _1546_ = instr_data[16] ? _1574_ : _1572_;
assign _1548_ = instr_data[16] ? _1578_ : _1576_;
assign _1550_ = instr_data[16] ? _1582_ : _1580_;
assign _1552_ = instr_data[15] ? REG__1_  : REG__0_ ;
assign _1572_ = instr_data[15] ? REG__21_  : REG__20_ ;
assign _1574_ = instr_data[15] ? REG__23_  : REG__22_ ;
assign _1576_ = instr_data[15] ? REG__25_  : REG__24_ ;
assign _1578_ = instr_data[15] ? REG__27_  : REG__26_ ;
assign _1580_ = instr_data[15] ? REG__29_  : REG__28_ ;
assign _1582_ = instr_data[15] ? REG__31_  : REG__30_ ;
assign _1554_ = instr_data[15] ? REG__3_  : REG__2_ ;
assign _1556_ = instr_data[15] ? REG__5_  : REG__4_ ;
assign _1558_ = instr_data[15] ? REG__7_  : REG__6_ ;
assign _1560_ = instr_data[15] ? REG__9_  : REG__8_ ;
assign _1562_ = instr_data[15] ? REG__11_  : REG__10_ ;
assign _1564_ = instr_data[15] ? REG__13_  : REG__12_ ;
assign _1566_ = instr_data[15] ? REG__15_  : REG__14_ ;
assign _1568_ = instr_data[15] ? REG__17_  : REG__16_ ;
assign _1570_ = instr_data[15] ? REG__19_  : REG__18_ ;
assign _1584_ = _0649_ & _0004_[31];
assign _1586_ = _0681_ & _0004_[31];
assign _1588_ = _0683_ & _0004_[31];
assign _1590_ = _0687_ & _0004_[31];
assign _1592_ = _0689_ & _0004_[31];
assign _1594_ = _0691_ & _0004_[31];
assign _1596_ = _0693_ & _0004_[31];
assign _1598_ = _0699_ & _0004_[31];
assign _1600_ = _0701_ & _0004_[31];
assign _1602_ = _0703_ & _0004_[31];
assign _1604_ = _0705_ & _0004_[31];
assign _1606_ = _0653_ & _0004_[31];
assign _1608_ = _0709_ & _0004_[31];
assign _1610_ = _0711_ & _0004_[31];
assign _1612_ = _0713_ & _0004_[31];
assign _1614_ = _0715_ & _0004_[31];
assign _1616_ = _0721_ & _0004_[31];
assign _1618_ = _0723_ & _0004_[31];
assign _1620_ = _0725_ & _0004_[31];
assign _1622_ = _0727_ & _0004_[31];
assign _1624_ = _0731_ & _0004_[31];
assign _1626_ = _0733_ & _0004_[31];
assign _1628_ = _0657_ & _0004_[31];
assign _1630_ = _0735_ & _0004_[31];
assign _1632_ = _0737_ & _0004_[31];
assign _1634_ = _0661_ & _0004_[31];
assign _1636_ = _0665_ & _0004_[31];
assign _1638_ = _0667_ & _0004_[31];
assign _1640_ = _0669_ & _0004_[31];
assign _1642_ = _0671_ & _0004_[31];
assign _1644_ = _0677_ & _0004_[31];
assign _1646_ = _0679_ & _0004_[31];
assign _1652_ = ~ /* src = "generated/sv2v_out.v:1626.21-1626.29" */ reg_vld;
assign instr_rdy = _1652_ | /* src = "generated/sv2v_out.v:1626.21-1626.41" */ fetch_rdy;
assign _0004_[31] = regwr_en ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1628.7-1628.15|generated/sv2v_out.v:1628.3-1629.33" */ 1'h1 : 1'h0;
assign _0002_ = regwr_en ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1628.7-1628.15|generated/sv2v_out.v:1628.3-1629.33" */ regwr_data : 32'hxxxxxxxx;
assign _0000_ = regwr_en ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1628.7-1628.15|generated/sv2v_out.v:1628.3-1629.33" */ regwr_sel : 5'hxx;
assign _1653_ = _1440_ ? /* src = "generated/sv2v_out.v:1624.12-1624.32|generated/sv2v_out.v:1624.8-1625.20" */ 1'h0 : 1'hx;
assign _1654_ = _1438_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1618.12-1618.31|generated/sv2v_out.v:1618.8-1625.20" */ 1'hx : _1653_;
assign _1655_ = _1432_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1598.12-1598.34|generated/sv2v_out.v:1598.8-1625.20" */ 1'h1 : _1654_;
assign _1657_ = _1430_ ? /* src = "generated/sv2v_out.v:1621.8-1621.28|generated/sv2v_out.v:1621.4-1622.29" */ regwr_data : 32'hxxxxxxxx;
assign _1659_ = _1438_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1618.12-1618.31|generated/sv2v_out.v:1618.8-1625.20" */ _1657_ : 32'hxxxxxxxx;
assign _1324_ = _1436_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1609.13-1609.43|generated/sv2v_out.v:1609.9-1612.27" */ regwr_data : _1650_;
assign _1662_ = _1424_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1607.8-1607.16|generated/sv2v_out.v:1607.4-1612.27" */ 32'd0 : _1324_;
assign _1664_ = _1432_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1598.12-1598.34|generated/sv2v_out.v:1598.8-1625.20" */ _1662_ : _1659_;
assign _1666_ = _1428_ ? /* src = "generated/sv2v_out.v:1619.8-1619.28|generated/sv2v_out.v:1619.4-1620.29" */ regwr_data : 32'hxxxxxxxx;
assign _1668_ = _1438_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1618.12-1618.31|generated/sv2v_out.v:1618.8-1625.20" */ _1666_ : 32'hxxxxxxxx;
assign _1327_ = _1434_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1603.13-1603.43|generated/sv2v_out.v:1603.9-1606.27" */ regwr_data : _1648_;
assign _1671_ = _1420_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1601.8-1601.16|generated/sv2v_out.v:1601.4-1606.27" */ 32'd0 : _1327_;
assign _1673_ = _1432_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1598.12-1598.34|generated/sv2v_out.v:1598.8-1625.20" */ _1671_ : _1668_;
assign ImmF = format_U ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1583.7-1583.15|generated/sv2v_out.v:1583.3-1586.23" */ instr_data[31:20] : { instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31] };
assign ImmE = _1446_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1579.7-1579.27|generated/sv2v_out.v:1579.3-1582.22" */ instr_data[19:12] : { instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31], instr_data[31] };
assign _0011_ = format_J ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1575.12-1575.20|generated/sv2v_out.v:1575.8-1578.16" */ instr_data[20] : instr_data[31];
assign _0009_ = format_B ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1573.12-1573.20|generated/sv2v_out.v:1573.8-1578.16" */ instr_data[7] : _0011_;
assign _0007_ = _1444_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1563.12-1563.32|generated/sv2v_out.v:1563.8-1566.20" */ instr_data[24:21] : instr_data[11:8];
assign _0005_ = format_S ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1557.12-1557.20|generated/sv2v_out.v:1557.8-1560.16" */ instr_data[7] : 1'h0;
assign ImmA = format_I ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1555.7-1555.15|generated/sv2v_out.v:1555.3-1560.16" */ instr_data[20] : _0005_;
assign _0004_[30:0] = { _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31], _0004_[31] };
// Added block to randomize initial values.
`ifdef RANDOMIZE_INIT
  initial begin
    regrd_rs1_t0 = '0;
    regrd_rs2_t0 = '0;
    regrd_rs1_en_t0 = '0;
    regrd_rs2_en_t0 = '0;
    reg_rs1_t0 = '0;
    reg_rs2_t0 = '0;
    _2406_ = '0;
    REG__9__t0 = '0;
    REG__8__t0 = '0;
    REG__7__t0 = '0;
    REG__6__t0 = '0;
    REG__5__t0 = '0;
    REG__4__t0 = '0;
    REG__3__t0 = '0;
    REG__31__t0 = '0;
    REG__30__t0 = '0;
    REG__2__t0 = '0;
    REG__29__t0 = '0;
    REG__28__t0 = '0;
    REG__27__t0 = '0;
    REG__26__t0 = '0;
    REG__25__t0 = '0;
    REG__24__t0 = '0;
    REG__23__t0 = '0;
    REG__22__t0 = '0;
    REG__21__t0 = '0;
    REG__20__t0 = '0;
    REG__1__t0 = '0;
    REG__19__t0 = '0;
    REG__18__t0 = '0;
    REG__17__t0 = '0;
    REG__16__t0 = '0;
    REG__15__t0 = '0;
    REG__14__t0 = '0;
    REG__13__t0 = '0;
    REG__12__t0 = '0;
    REG__11__t0 = '0;
    REG__10__t0 = '0;
    REG__0__t0 = '0;
    regrd_rs1 = '0;
    regrd_rs2 = '0;
    regrd_rs1_en = '0;
    regrd_rs2_en = '0;
    reg_vld = '0;
    reg_rs1 = '0;
    reg_rs2 = '0;
    _2519_ = '0;
    _2520_ = '0;
    REG__9_ = '0;
    REG__8_ = '0;
    REG__7_ = '0;
    REG__6_ = '0;
    REG__5_ = '0;
    REG__4_ = '0;
    REG__3_ = '0;
    REG__31_ = '0;
    REG__30_ = '0;
    REG__2_ = '0;
    REG__29_ = '0;
    REG__28_ = '0;
    REG__27_ = '0;
    REG__26_ = '0;
    REG__25_ = '0;
    REG__24_ = '0;
    REG__23_ = '0;
    REG__22_ = '0;
    REG__21_ = '0;
    REG__20_ = '0;
    REG__1_ = '0;
    REG__19_ = '0;
    REG__18_ = '0;
    REG__17_ = '0;
    REG__16_ = '0;
    REG__15_ = '0;
    REG__14_ = '0;
    REG__13_ = '0;
    REG__12_ = '0;
    REG__11_ = '0;
    REG__10_ = '0;
    REG__0_ = '0;
    _3286_ = '0;
    reg_vld_t0 = '0;
  end
`endif // RANDOMIZE_INIT
endmodule

module kronos_alu(op1, op2, aluop, result, aluop_t0, op1_t0, op2_t0, result_t0);
/* src = "generated/sv2v_out.v:52.22-52.55" */
wire [32:0] _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:52.22-52.55" */
wire [32:0] _001_;
wire _002_;
/* cellift = 32'd1 */
wire _003_;
wire [32:0] _004_;
wire [32:0] _005_;
wire [32:0] _006_;
wire [32:0] _007_;
wire [1:0] _008_;
wire [4:0] _009_;
wire [31:0] _010_;
wire [31:0] _011_;
wire [31:0] _012_;
wire [31:0] _013_;
wire [31:0] _014_;
wire _015_;
wire _016_;
wire _017_;
wire [31:0] _018_;
wire [31:0] _019_;
wire [2:0] _020_;
wire [3:0] _021_;
wire [1:0] _022_;
wire [1:0] _023_;
wire [31:0] _024_;
wire _025_;
wire [31:0] _026_;
wire [31:0] _027_;
wire [31:0] _028_;
wire [31:0] _029_;
wire [31:0] _030_;
wire [31:0] _031_;
wire _032_;
/* cellift = 32'd1 */
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire [32:0] _045_;
wire [32:0] _046_;
wire [32:0] _047_;
wire [32:0] _048_;
wire [31:0] _049_;
wire [31:0] _050_;
wire [31:0] _051_;
wire _052_;
wire _053_;
wire _054_;
wire [1:0] _055_;
wire [4:0] _056_;
wire [31:0] _057_;
wire [31:0] _058_;
wire [31:0] _059_;
wire [31:0] _060_;
wire [31:0] _061_;
wire [31:0] _062_;
wire [31:0] _063_;
wire [31:0] _064_;
wire [31:0] _065_;
wire [31:0] _066_;
wire [31:0] _067_;
wire [31:0] _068_;
wire [31:0] _069_;
wire [31:0] _070_;
wire [31:0] _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire [31:0] _078_;
wire [31:0] _079_;
wire [2:0] _080_;
wire [3:0] _081_;
wire [1:0] _082_;
wire [1:0] _083_;
wire [31:0] _084_;
wire [31:0] _085_;
wire [31:0] _086_;
wire _087_;
wire _088_;
wire _089_;
wire [31:0] _090_;
wire [31:0] _091_;
wire [31:0] _092_;
wire [31:0] _093_;
wire [31:0] _094_;
wire [31:0] _095_;
wire [31:0] _096_;
wire [31:0] _097_;
wire [31:0] _098_;
wire [31:0] _099_;
wire [31:0] _100_;
wire [31:0] _101_;
wire [31:0] _102_;
wire [31:0] _103_;
wire [31:0] _104_;
wire [31:0] _105_;
wire [31:0] _106_;
wire [31:0] _107_;
wire [31:0] _108_;
wire [31:0] _109_;
wire [31:0] _110_;
wire [32:0] _111_;
wire [32:0] _112_;
wire [32:0] _113_;
wire [32:0] _114_;
wire [32:0] _115_;
wire [32:0] _116_;
wire [31:0] _117_;
wire _118_;
wire [31:0] _119_;
wire [31:0] _120_;
wire [31:0] _121_;
wire [31:0] _122_;
wire [31:0] _123_;
wire [31:0] _124_;
wire [31:0] _125_;
wire [31:0] _126_;
wire [31:0] _127_;
wire [31:0] _128_;
wire [31:0] _129_;
wire [31:0] _130_;
wire [31:0] _131_;
wire [31:0] _132_;
wire [31:0] _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire [31:0] _138_;
wire [31:0] _139_;
wire [31:0] _140_;
wire [31:0] _141_;
wire _142_;
wire _143_;
wire _144_;
wire [31:0] _145_;
wire [31:0] _146_;
wire [31:0] _147_;
wire [31:0] _148_;
wire [31:0] _149_;
wire [31:0] _150_;
wire [31:0] _151_;
wire [31:0] _152_;
wire [31:0] _153_;
wire [31:0] _154_;
wire [31:0] _155_;
wire [31:0] _156_;
wire [31:0] _157_;
wire [31:0] _158_;
wire [31:0] _159_;
wire [31:0] _160_;
wire [31:0] _161_;
wire [31:0] _162_;
wire [31:0] _163_;
wire [32:0] _164_;
wire [32:0] _165_;
wire [31:0] _166_;
wire [31:0] _167_;
wire [31:0] _168_;
wire [31:0] _169_;
wire [31:0] _170_;
wire _171_;
wire [31:0] _172_;
wire _173_;
wire [31:0] _174_;
wire [31:0] _175_;
wire [31:0] _176_;
wire [31:0] _177_;
wire [31:0] _178_;
wire [31:0] _179_;
wire [31:0] _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire [32:0] _191_;
wire [32:0] _192_;
wire [32:0] _193_;
wire [32:0] _194_;
wire [31:0] _195_;
/* cellift = 32'd1 */
wire [31:0] _196_;
wire [31:0] _197_;
/* cellift = 32'd1 */
wire [31:0] _198_;
wire [31:0] _199_;
/* cellift = 32'd1 */
wire [31:0] _200_;
wire [31:0] _201_;
/* cellift = 32'd1 */
wire [31:0] _202_;
wire _203_;
/* cellift = 32'd1 */
wire _204_;
wire [2:0] _205_;
/* cellift = 32'd1 */
wire [2:0] _206_;
wire _207_;
/* cellift = 32'd1 */
wire _208_;
wire _209_;
/* cellift = 32'd1 */
wire _210_;
wire _211_;
/* cellift = 32'd1 */
wire _212_;
wire _213_;
/* cellift = 32'd1 */
wire _214_;
wire [1:0] _215_;
/* cellift = 32'd1 */
wire [1:0] _216_;
wire _217_;
/* cellift = 32'd1 */
wire _218_;
wire _219_;
/* cellift = 32'd1 */
wire _220_;
wire _221_;
wire _222_;
/* cellift = 32'd1 */
wire _223_;
/* src = "generated/sv2v_out.v:34.6-34.12" */
wire R_sign;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:34.6-34.12" */
wire R_sign_t0;
/* src = "generated/sv2v_out.v:30.13-30.20" */
wire [31:0] adder_B;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:30.13-30.20" */
wire [31:0] adder_B_t0;
/* src = "generated/sv2v_out.v:9.19-9.24" */
input [3:0] aluop;
wire [3:0] aluop;
/* cellift = 32'd1 */
input [3:0] aluop_t0;
wire [3:0] aluop_t0;
/* src = "generated/sv2v_out.v:21.7-21.10" */
wire cin;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21.7-21.10" */
wire cin_t0;
/* src = "generated/sv2v_out.v:31.6-31.10" */
wire cout;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:31.6-31.10" */
wire cout_t0;
/* src = "generated/sv2v_out.v:38.14-38.18" */
wire [31:0] data;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:38.14-38.18" */
wire [31:0] data_t0;
/* src = "generated/sv2v_out.v:7.20-7.23" */
input [31:0] op1;
wire [31:0] op1;
/* cellift = 32'd1 */
input [31:0] op1_t0;
wire [31:0] op1_t0;
/* src = "generated/sv2v_out.v:8.20-8.23" */
input [31:0] op2;
wire [31:0] op2;
/* cellift = 32'd1 */
input [31:0] op2_t0;
wire [31:0] op2_t0;
/* src = "generated/sv2v_out.v:41.14-41.16" */
wire [31:0] p0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:41.14-41.16" */
wire [31:0] p0_t0;
/* src = "generated/sv2v_out.v:42.14-42.16" */
wire [31:0] p1;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:42.14-42.16" */
wire [31:0] p1_t0;
/* src = "generated/sv2v_out.v:43.14-43.16" */
wire [31:0] p2;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:43.14-43.16" */
wire [31:0] p2_t0;
/* src = "generated/sv2v_out.v:44.14-44.16" */
wire [31:0] p3;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:44.14-44.16" */
wire [31:0] p3_t0;
/* src = "generated/sv2v_out.v:45.14-45.16" */
wire [31:0] p4;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:45.14-45.16" */
wire [31:0] p4_t0;
/* src = "generated/sv2v_out.v:24.13-24.20" */
wire [31:0] r_adder;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:24.13-24.20" */
wire [31:0] r_adder_t0;
/* src = "generated/sv2v_out.v:25.13-25.18" */
wire [31:0] r_and;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25.13-25.18" */
wire [31:0] r_and_t0;
/* src = "generated/sv2v_out.v:37.6-37.12" */
wire r_comp;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:37.6-37.12" */
wire r_comp_t0;
/* src = "generated/sv2v_out.v:35.6-35.10" */
wire r_lt;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:35.6-35.10" */
wire r_lt_t0;
/* src = "generated/sv2v_out.v:36.6-36.11" */
wire r_ltu;
/* src = "generated/sv2v_out.v:26.13-26.17" */
wire [31:0] r_or;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26.13-26.17" */
wire [31:0] r_or_t0;
/* src = "generated/sv2v_out.v:28.14-28.21" */
wire [31:0] r_shift;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:28.14-28.21" */
wire [31:0] r_shift_t0;
/* src = "generated/sv2v_out.v:27.13-27.18" */
wire [31:0] r_xor;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:27.13-27.18" */
wire [31:0] r_xor_t0;
/* src = "generated/sv2v_out.v:10.20-10.26" */
output [31:0] result;
wire [31:0] result;
/* cellift = 32'd1 */
output [31:0] result_t0;
wire [31:0] result_t0;
/* src = "generated/sv2v_out.v:40.7-40.15" */
wire shift_in;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:40.7-40.15" */
wire shift_in_t0;
assign _000_ = { 1'h0, op1 } + /* src = "generated/sv2v_out.v:52.22-52.55" */ { 1'h0, adder_B };
assign { cout, R_sign, r_adder[30:0] } = _000_ + /* src = "generated/sv2v_out.v:52.21-52.62" */ cin;
assign r_and = op1 & /* src = "generated/sv2v_out.v:55.11-55.20" */ op2;
assign shift_in = cin & /* src = "generated/sv2v_out.v:73.20-73.33" */ op1[31];
assign _004_ = ~ { 1'h0, op1_t0 };
assign _006_ = ~ _001_;
assign _005_ = ~ { 1'h0, adder_B_t0 };
assign _007_ = ~ { 32'h00000000, cin_t0 };
assign _045_ = { 1'h0, op1 } & _004_;
assign _047_ = _000_ & _006_;
assign _046_ = { 1'h0, adder_B } & _005_;
assign _048_ = { 32'h00000000, cin } & _007_;
assign _191_ = _045_ + _046_;
assign _193_ = _047_ + _048_;
assign _111_ = { 1'h0, op1 } | { 1'h0, op1_t0 };
assign _114_ = _000_ | _001_;
assign _112_ = { 1'h0, adder_B } | { 1'h0, adder_B_t0 };
assign _115_ = { 32'h00000000, cin } | { 32'h00000000, cin_t0 };
assign _192_ = _111_ + _112_;
assign _194_ = _114_ + _115_;
assign _164_ = _191_ ^ _192_;
assign _165_ = _193_ ^ _194_;
assign _113_ = _164_ | { 1'h0, op1_t0 };
assign _116_ = _165_ | _001_;
assign _001_ = _113_ | { 1'h0, adder_B_t0 };
assign { cout_t0, R_sign_t0, r_adder_t0[30:0] } = _116_ | { 32'h00000000, cin_t0 };
assign _049_ = op1_t0 & op2;
assign _052_ = cin_t0 & op1[31];
assign _050_ = op2_t0 & op1;
assign _053_ = op1_t0[31] & cin;
assign _054_ = cin_t0 & op1_t0[31];
assign _117_ = _049_ | _050_;
assign _118_ = _052_ | _053_;
assign r_and_t0 = _117_ | _051_;
assign shift_in_t0 = _118_ | _054_;
assign _037_ = | aluop_t0;
assign _021_ = ~ aluop_t0;
assign _081_ = aluop & _021_;
assign _181_ = _081_ == { 3'h0, _021_[0] };
assign _182_ = _081_ == { 1'h0, _021_[2], 1'h0, _021_[0] };
assign _183_ = _081_ == { _021_[3:2], 1'h0, _021_[0] };
assign _184_ = _081_ == { 1'h0, _021_[2:0] };
assign _185_ = _081_ == { 1'h0, _021_[2:1], 1'h0 };
assign _186_ = _081_ == { 1'h0, _021_[2], 2'h0 };
assign _187_ = _081_ == { 2'h0, _021_[1], 1'h0 };
assign _188_ = _081_ == { 2'h0, _021_[1:0] };
assign _189_ = _083_ == _023_;
assign _190_ = _083_ == { _023_[1], 1'h0 };
assign _206_[0] = _181_ & _037_;
assign _206_[1] = _182_ & _037_;
assign _206_[2] = _183_ & _037_;
assign _210_ = _184_ & _037_;
assign _212_ = _185_ & _037_;
assign _214_ = _186_ & _037_;
assign _216_[0] = _187_ & _037_;
assign _216_[1] = _188_ & _037_;
assign _220_ = _189_ & _039_;
assign _204_ = _190_ & _039_;
assign _034_ = | { _223_, _220_ };
assign _035_ = | { _212_, _210_, _206_ };
assign _036_ = | _206_;
assign _038_ = | _216_;
assign _039_ = | { op2_t0[31], op1_t0[31] };
assign _008_ = ~ { _223_, _220_ };
assign _009_ = ~ { _212_, _210_, _206_ };
assign _020_ = ~ _206_;
assign _022_ = ~ _216_;
assign _023_ = ~ { op1_t0[31], op2_t0[31] };
assign _055_ = { _222_, _219_ } & _008_;
assign _056_ = { _211_, _209_, _205_ } & _009_;
assign _080_ = _205_ & _020_;
assign _082_ = _215_ & _022_;
assign _083_ = { op1[31], op2[31] } & _023_;
assign _040_ = ! _055_;
assign _041_ = ! _056_;
assign _042_ = ! _080_;
assign _043_ = ! _082_;
assign _044_ = ! _083_;
assign _003_ = _040_ & _034_;
assign _033_ = _041_ & _035_;
assign _208_ = _042_ & _036_;
assign _218_ = _043_ & _038_;
assign _223_ = _044_ & _039_;
assign _016_ = ~ aluop[3];
assign _017_ = ~ aluop[1];
assign _075_ = aluop_t0[3] & _017_;
assign _076_ = aluop_t0[1] & _016_;
assign _077_ = aluop_t0[3] & aluop_t0[1];
assign _137_ = _075_ | _076_;
assign cin_t0 = _137_ | _077_;
assign _010_ = ~ { _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_ };
assign _011_ = ~ { _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_ };
assign _012_ = ~ { _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_ };
assign _013_ = ~ { _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_ };
assign _014_ = ~ { _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_ };
assign _015_ = ~ _002_;
assign _024_ = ~ { cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin };
assign _025_ = ~ aluop[0];
assign _026_ = ~ { aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2] };
assign _027_ = ~ { op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0] };
assign _028_ = ~ { op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1] };
assign _029_ = ~ { op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2] };
assign _030_ = ~ { op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3] };
assign _031_ = ~ { op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4] };
assign _119_ = { _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_ } | _010_;
assign _122_ = { _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_ } | _011_;
assign _125_ = { _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_ } | _012_;
assign _128_ = { _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_ } | _013_;
assign _131_ = { _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_ } | _014_;
assign _134_ = _003_ | _015_;
assign _139_ = { cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0 } | _024_;
assign _142_ = aluop_t0[0] | _025_;
assign _145_ = { aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2] } | _026_;
assign _148_ = { op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0] } | _027_;
assign _151_ = { op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1] } | _028_;
assign _154_ = { op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2] } | _029_;
assign _157_ = { op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3] } | _030_;
assign _160_ = { op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4] } | _031_;
assign _120_ = { _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_ } | { _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_, _209_ };
assign _123_ = { _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_ } | { _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_, _207_ };
assign _126_ = { _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_ } | { _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_, _217_ };
assign _129_ = { _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_ } | { _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_ };
assign _132_ = { _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_ } | { _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_ };
assign _135_ = _003_ | _002_;
assign _140_ = { cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0 } | { cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin, cin };
assign _143_ = aluop_t0[0] | aluop[0];
assign _146_ = { aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2] } | { aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2], aluop[2] };
assign _149_ = { op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0] } | { op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0], op2[0] };
assign _152_ = { op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1] } | { op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1], op2[1] };
assign _155_ = { op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2] } | { op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2], op2[2] };
assign _158_ = { op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3] } | { op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3], op2[3] };
assign _161_ = { op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4] } | { op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4], op2[4] };
assign _057_ = r_or_t0 & _119_;
assign _060_ = _196_ & _122_;
assign _063_ = { R_sign_t0, r_adder_t0[30:0] } & _125_;
assign _066_ = _200_ & _128_;
assign _069_ = _202_ & _131_;
assign _072_ = _204_ & _134_;
assign _084_ = op2_t0 & _139_;
assign _087_ = r_lt_t0 & _142_;
assign _090_ = { op1_t0[0], op1_t0[1], op1_t0[2], op1_t0[3], op1_t0[4], op1_t0[5], op1_t0[6], op1_t0[7], op1_t0[8], op1_t0[9], op1_t0[10], op1_t0[11], op1_t0[12], op1_t0[13], op1_t0[14], op1_t0[15], op1_t0[16], op1_t0[17], op1_t0[18], op1_t0[19], op1_t0[20], op1_t0[21], op1_t0[22], op1_t0[23], op1_t0[24], op1_t0[25], op1_t0[26], op1_t0[27], op1_t0[28], op1_t0[29], op1_t0[30], op1_t0[31] } & _145_;
assign _093_ = data_t0 & _148_;
assign _096_ = p0_t0 & _151_;
assign _099_ = p1_t0 & _154_;
assign _102_ = p2_t0 & _157_;
assign _105_ = p3_t0 & _160_;
assign _108_ = { p4_t0[0], p4_t0[1], p4_t0[2], p4_t0[3], p4_t0[4], p4_t0[5], p4_t0[6], p4_t0[7], p4_t0[8], p4_t0[9], p4_t0[10], p4_t0[11], p4_t0[12], p4_t0[13], p4_t0[14], p4_t0[15], p4_t0[16], p4_t0[17], p4_t0[18], p4_t0[19], p4_t0[20], p4_t0[21], p4_t0[22], p4_t0[23], p4_t0[24], p4_t0[25], p4_t0[26], p4_t0[27], p4_t0[28], p4_t0[29], p4_t0[30], p4_t0[31] } & _145_;
assign _058_ = r_and_t0 & _120_;
assign _061_ = r_shift_t0 & _123_;
assign _064_ = { 31'h00000000, r_comp_t0 } & _126_;
assign _067_ = r_xor_t0 & _129_;
assign _070_ = _198_ & _132_;
assign _073_ = R_sign_t0 & _135_;
assign _085_ = op2_t0 & _140_;
assign _088_ = cout_t0 & _143_;
assign _091_ = op1_t0 & _146_;
assign _094_ = { shift_in_t0, data_t0[31:1] } & _149_;
assign _097_ = { shift_in_t0, shift_in_t0, p0_t0[31:2] } & _152_;
assign _100_ = { shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, p1_t0[31:4] } & _155_;
assign _103_ = { shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, p2_t0[31:8] } & _158_;
assign _106_ = { shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, shift_in_t0, p3_t0[31:16] } & _161_;
assign _109_ = p4_t0 & _146_;
assign _121_ = _057_ | _058_;
assign _124_ = _060_ | _061_;
assign _127_ = _063_ | _064_;
assign _130_ = _066_ | _067_;
assign _133_ = _069_ | _070_;
assign _136_ = _072_ | _073_;
assign _141_ = _084_ | _085_;
assign _144_ = _087_ | _088_;
assign _147_ = _090_ | _091_;
assign _150_ = _093_ | _094_;
assign _153_ = _096_ | _097_;
assign _156_ = _099_ | _100_;
assign _159_ = _102_ | _103_;
assign _162_ = _105_ | _106_;
assign _163_ = _108_ | _109_;
assign _166_ = r_or ^ r_and;
assign _167_ = _195_ ^ r_shift;
assign _168_ = { R_sign, r_adder[30:0] } ^ { 31'h00000000, r_comp };
assign _169_ = _199_ ^ r_xor;
assign _170_ = _201_ ^ _197_;
assign _171_ = _203_ ^ R_sign;
assign _172_ = op2 ^ _019_;
assign _173_ = r_lt ^ r_ltu;
assign _174_ = { op1[0], op1[1], op1[2], op1[3], op1[4], op1[5], op1[6], op1[7], op1[8], op1[9], op1[10], op1[11], op1[12], op1[13], op1[14], op1[15], op1[16], op1[17], op1[18], op1[19], op1[20], op1[21], op1[22], op1[23], op1[24], op1[25], op1[26], op1[27], op1[28], op1[29], op1[30], op1[31] } ^ op1;
assign _175_ = data ^ { shift_in, data[31:1] };
assign _176_ = p0 ^ { shift_in, shift_in, p0[31:2] };
assign _177_ = p1 ^ { shift_in, shift_in, shift_in, shift_in, p1[31:4] };
assign _178_ = p2 ^ { shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, p2[31:8] };
assign _179_ = p3 ^ { shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, p3[31:16] };
assign _180_ = { p4[0], p4[1], p4[2], p4[3], p4[4], p4[5], p4[6], p4[7], p4[8], p4[9], p4[10], p4[11], p4[12], p4[13], p4[14], p4[15], p4[16], p4[17], p4[18], p4[19], p4[20], p4[21], p4[22], p4[23], p4[24], p4[25], p4[26], p4[27], p4[28], p4[29], p4[30], p4[31] } ^ p4;
assign _059_ = { _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_, _210_ } & _166_;
assign _062_ = { _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_, _208_ } & _167_;
assign _065_ = { _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_, _218_ } & _168_;
assign _068_ = { _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_, _214_ } & _169_;
assign _071_ = { _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_ } & _170_;
assign _074_ = _003_ & _171_;
assign _086_ = { cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0, cin_t0 } & _172_;
assign _089_ = aluop_t0[0] & _173_;
assign _092_ = { aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2] } & _174_;
assign _095_ = { op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0], op2_t0[0] } & _175_;
assign _098_ = { op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1], op2_t0[1] } & _176_;
assign _101_ = { op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2], op2_t0[2] } & _177_;
assign _104_ = { op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3], op2_t0[3] } & _178_;
assign _107_ = { op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4], op2_t0[4] } & _179_;
assign _110_ = { aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2], aluop_t0[2] } & _180_;
assign _196_ = _059_ | _121_;
assign _198_ = _062_ | _124_;
assign _200_ = _065_ | _127_;
assign _202_ = _068_ | _130_;
assign result_t0 = _071_ | _133_;
assign r_lt_t0 = _074_ | _136_;
assign adder_B_t0 = _086_ | _141_;
assign r_comp_t0 = _089_ | _144_;
assign data_t0 = _092_ | _147_;
assign p0_t0 = _095_ | _150_;
assign p1_t0 = _098_ | _153_;
assign p2_t0 = _101_ | _156_;
assign p3_t0 = _104_ | _159_;
assign p4_t0 = _107_ | _162_;
assign r_shift_t0 = _110_ | _163_;
assign _002_ = | { _222_, _219_ };
assign _018_ = ~ op1;
assign _019_ = ~ op2;
assign _078_ = op1_t0 & _019_;
assign _079_ = op2_t0 & _018_;
assign _051_ = op1_t0 & op2_t0;
assign _138_ = _078_ | _079_;
assign r_or_t0 = _138_ | _051_;
assign _032_ = | { _211_, _209_, _205_ };
assign _195_ = _209_ ? r_and : r_or;
assign _197_ = _207_ ? r_shift : _195_;
assign _199_ = _217_ ? { 31'h00000000, r_comp } : { R_sign, r_adder[30:0] };
assign _201_ = _213_ ? r_xor : _199_;
assign result = _032_ ? _197_ : _201_;
assign _203_ = _221_ ? 1'h1 : 1'h0;
assign r_lt = _002_ ? R_sign : _203_;
assign r_xor_t0 = op1_t0 | op2_t0;
assign cin = aluop[3] || /* src = "generated/sv2v_out.v:46.15-46.35" */ aluop[1];
assign r_ltu = ~ /* src = "generated/sv2v_out.v:69.11-69.16" */ cout;
assign r_or = op1 | /* src = "generated/sv2v_out.v:56.10-56.19" */ op2;
assign _207_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:90.3-97.10" */ _205_;
assign _205_[0] = aluop == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:90.3-97.10" */ 4'h1;
assign _205_[1] = aluop == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:90.3-97.10" */ 4'h5;
assign _205_[2] = aluop == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:90.3-97.10" */ 4'hd;
assign _209_ = aluop == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:90.3-97.10" */ 4'h7;
assign _211_ = aluop == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:90.3-97.10" */ 4'h6;
assign _213_ = aluop == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:90.3-97.10" */ 4'h4;
assign _217_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:90.3-97.10" */ _215_;
assign _215_[0] = aluop == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:90.3-97.10" */ 4'h2;
assign _215_[1] = aluop == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:90.3-97.10" */ 4'h3;
assign _219_ = { op1[31], op2[31] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:63.3-68.10" */ 2'h3;
assign _221_ = { op1[31], op2[31] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:63.3-68.10" */ 2'h2;
assign _222_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:63.3-68.10" */ { op1[31], op2[31] };
assign adder_B = cin ? /* src = "generated/sv2v_out.v:51.14-51.30" */ _019_ : op2;
assign r_comp = aluop[0] ? /* src = "generated/sv2v_out.v:70.13-70.31" */ r_ltu : r_lt;
assign data = aluop[2] ? /* src = "generated/sv2v_out.v:72.17-72.46" */ op1 : { op1[0], op1[1], op1[2], op1[3], op1[4], op1[5], op1[6], op1[7], op1[8], op1[9], op1[10], op1[11], op1[12], op1[13], op1[14], op1[15], op1[16], op1[17], op1[18], op1[19], op1[20], op1[21], op1[22], op1[23], op1[24], op1[25], op1[26], op1[27], op1[28], op1[29], op1[30], op1[31] };
assign p0 = op2[0] ? /* src = "generated/sv2v_out.v:75.15-75.55" */ { shift_in, data[31:1] } : data;
assign p1 = op2[1] ? /* src = "generated/sv2v_out.v:76.15-76.57" */ { shift_in, shift_in, p0[31:2] } : p0;
assign p2 = op2[2] ? /* src = "generated/sv2v_out.v:77.15-77.57" */ { shift_in, shift_in, shift_in, shift_in, p1[31:4] } : p1;
assign p3 = op2[3] ? /* src = "generated/sv2v_out.v:78.15-78.57" */ { shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, p2[31:8] } : p2;
assign p4 = op2[4] ? /* src = "generated/sv2v_out.v:79.15-79.59" */ { shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, shift_in, p3[31:16] } : p3;
assign r_shift = aluop[2] ? /* src = "generated/sv2v_out.v:80.20-80.47" */ p4 : { p4[0], p4[1], p4[2], p4[3], p4[4], p4[5], p4[6], p4[7], p4[8], p4[9], p4[10], p4[11], p4[12], p4[13], p4[14], p4[15], p4[16], p4[17], p4[18], p4[19], p4[20], p4[21], p4[22], p4[23], p4[24], p4[25], p4[26], p4[27], p4[28], p4[29], p4[30], p4[31] };
assign r_xor = op1 ^ /* src = "generated/sv2v_out.v:57.11-57.20" */ op2;
assign r_adder[31] = R_sign;
assign r_adder_t0[31] = R_sign_t0;
endmodule

module kronos_branch(op, rs1, rs2, branch, branch_t0, op_t0, rs1_t0, rs2_t0);
wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire [31:0] _008_;
wire [30:0] _009_;
wire _010_;
wire [30:0] _011_;
wire _012_;
wire [1:0] _013_;
wire [2:0] _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire [31:0] _033_;
wire [31:0] _034_;
wire _035_;
wire _036_;
wire [30:0] _037_;
wire [30:0] _038_;
wire [1:0] _039_;
wire [2:0] _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire [31:0] _054_;
wire _055_;
wire _056_;
wire [30:0] _057_;
wire [30:0] _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
/* cellift = 32'd1 */
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
/* cellift = 32'd1 */
wire _073_;
wire _074_;
/* cellift = 32'd1 */
wire _075_;
/* src = "generated/sv2v_out.v:114.21-114.30" */
wire _076_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:114.21-114.30" */
wire _077_;
/* src = "generated/sv2v_out.v:114.33-114.60" */
wire _078_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:114.33-114.60" */
wire _079_;
/* src = "generated/sv2v_out.v:122.31-122.34" */
wire _080_;
/* src = "generated/sv2v_out.v:123.50-123.53" */
wire _081_;
wire [1:0] _082_;
/* cellift = 32'd1 */
wire [1:0] _083_;
wire _084_;
/* cellift = 32'd1 */
wire _085_;
wire _086_;
/* cellift = 32'd1 */
wire _087_;
wire _088_;
/* cellift = 32'd1 */
wire _089_;
/* src = "generated/sv2v_out.v:108.13-108.19" */
output branch;
wire branch;
/* cellift = 32'd1 */
output branch_t0;
wire branch_t0;
/* src = "generated/sv2v_out.v:110.7-110.9" */
wire eq;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:110.7-110.9" */
wire eq_t0;
/* src = "generated/sv2v_out.v:111.7-111.9" */
wire lt;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:111.7-111.9" */
wire lt_t0;
/* src = "generated/sv2v_out.v:105.19-105.21" */
input [2:0] op;
wire [2:0] op;
/* cellift = 32'd1 */
input [2:0] op_t0;
wire [2:0] op_t0;
/* src = "generated/sv2v_out.v:106.20-106.23" */
input [31:0] rs1;
wire [31:0] rs1;
/* cellift = 32'd1 */
input [31:0] rs1_t0;
wire [31:0] rs1_t0;
/* src = "generated/sv2v_out.v:107.20-107.23" */
input [31:0] rs2;
wire [31:0] rs2;
/* cellift = 32'd1 */
input [31:0] rs2_t0;
wire [31:0] rs2_t0;
assign _016_ = | { rs2_t0, rs1_t0 };
assign _018_ = | op_t0;
assign _054_ = rs1_t0 | rs2_t0;
assign _008_ = ~ _054_;
assign _033_ = rs1 & _008_;
assign _040_ = op & _014_;
assign _034_ = rs2 & _008_;
assign _068_ = _033_ == _034_;
assign _069_ = _040_ == { _014_[2], 1'h0, _014_[0] };
assign _070_ = _040_ == _014_;
assign _071_ = _040_ == { 2'h0, _014_[0] };
assign eq_t0 = _068_ & _016_;
assign _083_[0] = _069_ & _018_;
assign _083_[1] = _070_ & _018_;
assign _087_ = _071_ & _018_;
assign _017_ = | _083_;
assign _013_ = ~ _083_;
assign _014_ = ~ op_t0;
assign _039_ = _082_ & _013_;
assign _019_ = ! _039_;
assign _020_ = ! _040_;
assign _085_ = _019_ & _017_;
assign _089_ = _020_ & _018_;
assign _000_ = { _035_, _037_ } < { _056_, _058_ };
assign _001_ = $signed({ _055_, _037_ }) < $signed({ _036_, _058_ });
assign _002_ = { _055_, _057_ } < { _036_, _038_ };
assign _003_ = $signed({ _035_, _057_ }) < $signed({ _056_, _038_ });
assign _077_ = _000_ ^ _002_;
assign _079_ = _001_ ^ _003_;
assign _009_ = ~ rs1_t0[30:0];
assign _010_ = ~ rs1_t0[31];
assign _011_ = ~ rs2_t0[30:0];
assign _012_ = ~ rs2_t0[31];
assign _055_ = rs1[31] | rs1_t0[31];
assign _056_ = rs2[31] | rs2_t0[31];
assign _035_ = rs1[31] & _010_;
assign _036_ = rs2[31] & _012_;
assign _037_ = rs1[30:0] & _009_;
assign _038_ = rs2[30:0] & _011_;
assign _057_ = rs1[30:0] | rs1_t0[30:0];
assign _058_ = rs2[30:0] | rs2_t0[30:0];
assign _005_ = ~ _084_;
assign _006_ = ~ _088_;
assign _007_ = ~ _062_;
assign _015_ = ~ op[1];
assign _045_ = _085_ | _005_;
assign _048_ = _089_ | _006_;
assign _051_ = _063_ | _007_;
assign _059_ = op_t0[1] | _015_;
assign _046_ = _085_ | _084_;
assign _049_ = _089_ | _088_;
assign _052_ = _063_ | _062_;
assign _060_ = op_t0[1] | op[1];
assign _024_ = eq_t0 & _045_;
assign _027_ = lt_t0 & _048_;
assign _030_ = _075_ & _051_;
assign _041_ = _079_ & _059_;
assign _025_ = lt_t0 & _046_;
assign _028_ = eq_t0 & _049_;
assign _031_ = _073_ & _052_;
assign _042_ = _077_ & _060_;
assign _047_ = _024_ | _025_;
assign _050_ = _027_ | _028_;
assign _053_ = _030_ | _031_;
assign _061_ = _041_ | _042_;
assign _064_ = _080_ ^ _081_;
assign _065_ = lt ^ eq;
assign _066_ = _074_ ^ _072_;
assign _067_ = _078_ ^ _076_;
assign _026_ = _085_ & _064_;
assign _029_ = _089_ & _065_;
assign _032_ = _063_ & _066_;
assign _043_ = op_t0[1] & _067_;
assign _073_ = _026_ | _047_;
assign _075_ = _029_ | _050_;
assign branch_t0 = _032_ | _053_;
assign lt_t0 = _043_ | _061_;
assign _004_ = ~ _086_;
assign _021_ = _087_ & _005_;
assign _022_ = _085_ & _004_;
assign _023_ = _087_ & _085_;
assign _044_ = _021_ | _022_;
assign _063_ = _044_ | _023_;
assign _062_ = _086_ | _084_;
assign _072_ = _084_ ? _081_ : _080_;
assign _074_ = _088_ ? eq : lt;
assign branch = _062_ ? _072_ : _074_;
assign eq = rs1 == /* src = "generated/sv2v_out.v:113.14-113.24" */ rs2;
assign _076_ = rs1 < /* src = "generated/sv2v_out.v:114.21-114.30" */ rs2;
assign _078_ = $signed(rs1) < /* src = "generated/sv2v_out.v:114.33-114.60" */ $signed(rs2);
assign _080_ = ~ /* src = "generated/sv2v_out.v:122.31-122.34" */ eq;
assign _081_ = ~ /* src = "generated/sv2v_out.v:123.50-123.53" */ lt;
assign _084_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:120.3-125.10" */ _082_;
assign _082_[0] = op == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:120.3-125.10" */ 3'h5;
assign _082_[1] = op == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:120.3-125.10" */ 3'h7;
assign _086_ = op == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:120.3-125.10" */ 3'h1;
assign _088_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:120.3-125.10" */ op;
assign lt = op[1] ? /* src = "generated/sv2v_out.v:114.15-114.60" */ _076_ : _078_;
endmodule

module kronos_hcu(clk, rstz, flush, instr, regrd_rs1_en, regrd_rs2_en, fetch_vld, fetch_rdy, decode_vld, decode_rdy, regwr_sel, regwr_en, regwr_pending, stall, clk_t0, decode_rdy_t0, decode_vld_t0, regwr_en_t0, regwr_pending_t0, regwr_sel_t0, fetch_rdy_t0
, regrd_rs1_en_t0, regrd_rs2_en_t0, fetch_vld_t0, flush_t0, instr_t0, stall_t0);
/* src = "generated/sv2v_out.v:895.23-895.51" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:895.23-895.51" */
wire _001_;
/* src = "generated/sv2v_out.v:896.23-896.51" */
wire _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:896.23-896.51" */
wire _003_;
/* src = "generated/sv2v_out.v:897.47-897.85" */
wire _004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:897.47-897.85" */
wire _005_;
wire _006_;
wire [4:0] _007_;
wire [4:0] _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire [4:0] _031_;
wire [4:0] _032_;
wire [4:0] _033_;
wire [4:0] _034_;
wire [4:0] _035_;
wire [4:0] _036_;
wire [4:0] _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire [4:0] _053_;
wire [4:0] _054_;
wire [4:0] _055_;
wire [4:0] _056_;
wire [4:0] _057_;
wire [4:0] _058_;
wire _059_;
wire _060_;
wire _061_;
wire [4:0] _062_;
wire _063_;
wire _064_;
/* src = "generated/sv2v_out.v:895.56-895.68" */
wire _065_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:895.56-895.68" */
wire _066_;
/* src = "generated/sv2v_out.v:896.56-896.68" */
wire _067_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:896.56-896.68" */
wire _068_;
/* src = "generated/sv2v_out.v:897.60-897.84" */
wire _069_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:897.60-897.84" */
wire _070_;
/* src = "generated/sv2v_out.v:899.7-899.29" */
wire _071_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:899.7-899.29" */
wire _072_;
/* src = "generated/sv2v_out.v:897.58-897.85" */
wire _073_;
/* src = "generated/sv2v_out.v:897.45-897.86" */
wire _074_;
/* src = "generated/sv2v_out.v:897.18-897.41" */
wire _075_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:897.18-897.41" */
wire _076_;
/* src = "generated/sv2v_out.v:856.13-856.16" */
input clk;
wire clk;
/* cellift = 32'd1 */
input clk_t0;
wire clk_t0;
/* src = "generated/sv2v_out.v:865.13-865.23" */
input decode_rdy;
wire decode_rdy;
/* cellift = 32'd1 */
input decode_rdy_t0;
wire decode_rdy_t0;
/* src = "generated/sv2v_out.v:864.13-864.23" */
input decode_vld;
wire decode_vld;
/* cellift = 32'd1 */
input decode_vld_t0;
wire decode_vld_t0;
/* src = "generated/sv2v_out.v:863.13-863.22" */
input fetch_rdy;
wire fetch_rdy;
/* cellift = 32'd1 */
input fetch_rdy_t0;
wire fetch_rdy_t0;
/* src = "generated/sv2v_out.v:862.13-862.22" */
input fetch_vld;
wire fetch_vld;
/* cellift = 32'd1 */
input fetch_vld_t0;
wire fetch_vld_t0;
/* src = "generated/sv2v_out.v:858.13-858.18" */
input flush;
wire flush;
/* cellift = 32'd1 */
input flush_t0;
wire flush_t0;
/* src = "generated/sv2v_out.v:859.20-859.25" */
input [31:0] instr;
wire [31:0] instr;
/* cellift = 32'd1 */
input [31:0] instr_t0;
wire [31:0] instr_t0;
/* src = "generated/sv2v_out.v:860.13-860.25" */
input regrd_rs1_en;
wire regrd_rs1_en;
/* cellift = 32'd1 */
input regrd_rs1_en_t0;
wire regrd_rs1_en_t0;
/* src = "generated/sv2v_out.v:861.13-861.25" */
input regrd_rs2_en;
wire regrd_rs2_en;
/* cellift = 32'd1 */
input regrd_rs2_en_t0;
wire regrd_rs2_en_t0;
/* src = "generated/sv2v_out.v:867.13-867.21" */
input regwr_en;
wire regwr_en;
/* cellift = 32'd1 */
input regwr_en_t0;
wire regwr_en_t0;
/* src = "generated/sv2v_out.v:868.13-868.26" */
input regwr_pending;
wire regwr_pending;
/* cellift = 32'd1 */
input regwr_pending_t0;
wire regwr_pending_t0;
/* src = "generated/sv2v_out.v:866.19-866.28" */
input [4:0] regwr_sel;
wire [4:0] regwr_sel;
/* cellift = 32'd1 */
input [4:0] regwr_sel_t0;
wire [4:0] regwr_sel_t0;
/* src = "generated/sv2v_out.v:879.12-879.17" */
reg [4:0] rpend;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:879.12-879.17" */
reg [4:0] rpend_t0;
/* src = "generated/sv2v_out.v:877.7-877.17" */
wire rs1_hazard;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:877.7-877.17" */
wire rs1_hazard_t0;
/* src = "generated/sv2v_out.v:878.7-878.17" */
wire rs2_hazard;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:878.7-878.17" */
wire rs2_hazard_t0;
/* src = "generated/sv2v_out.v:857.13-857.17" */
input rstz;
wire rstz;
/* src = "generated/sv2v_out.v:869.14-869.19" */
output stall;
wire stall;
/* cellift = 32'd1 */
output stall_t0;
wire stall_t0;
assign _000_ = regrd_rs1_en & /* src = "generated/sv2v_out.v:895.23-895.51" */ regwr_pending;
assign rs1_hazard = _000_ & /* src = "generated/sv2v_out.v:895.22-895.69" */ _065_;
assign _002_ = regrd_rs2_en & /* src = "generated/sv2v_out.v:896.23-896.51" */ regwr_pending;
assign rs2_hazard = _002_ & /* src = "generated/sv2v_out.v:896.22-896.69" */ _067_;
assign _004_ = regwr_en & /* src = "generated/sv2v_out.v:897.47-897.85" */ _073_;
assign stall = _075_ & /* src = "generated/sv2v_out.v:897.17-897.86" */ _074_;
assign _013_ = regrd_rs1_en_t0 & regwr_pending;
assign _016_ = _001_ & _065_;
assign _019_ = regrd_rs2_en_t0 & regwr_pending;
assign _022_ = _003_ & _067_;
assign _025_ = regwr_en_t0 & _073_;
assign _028_ = _076_ & _074_;
assign _014_ = regwr_pending_t0 & regrd_rs1_en;
assign _017_ = _066_ & _000_;
assign _020_ = regwr_pending_t0 & regrd_rs2_en;
assign _023_ = _068_ & _002_;
assign _026_ = _070_ & regwr_en;
assign _029_ = _005_ & _075_;
assign _015_ = regrd_rs1_en_t0 & regwr_pending_t0;
assign _018_ = _001_ & _066_;
assign _021_ = regrd_rs2_en_t0 & regwr_pending_t0;
assign _024_ = _003_ & _068_;
assign _027_ = regwr_en_t0 & _070_;
assign _030_ = _076_ & _005_;
assign _047_ = _013_ | _014_;
assign _048_ = _016_ | _017_;
assign _049_ = _019_ | _020_;
assign _050_ = _022_ | _023_;
assign _051_ = _025_ | _026_;
assign _052_ = _028_ | _029_;
assign _001_ = _047_ | _015_;
assign rs1_hazard_t0 = _048_ | _018_;
assign _003_ = _049_ | _021_;
assign rs2_hazard_t0 = _050_ | _024_;
assign _005_ = _051_ | _027_;
assign stall_t0 = _052_ | _030_;
assign _062_ = instr[11:7] ^ rpend;
assign _006_ = ~ _071_;
assign _053_ = instr_t0[11:7] | rpend_t0;
assign _054_ = _062_ | _053_;
assign _031_ = { _071_, _071_, _071_, _071_, _071_ } & instr_t0[11:7];
assign _032_ = { _006_, _006_, _006_, _006_, _006_ } & rpend_t0;
assign _033_ = _054_ & { _072_, _072_, _072_, _072_, _072_ };
assign _055_ = _031_ | _032_;
assign _056_ = _055_ | _033_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_hcu */
/* PC_TAINT_INFO STATE_NAME rpend_t0 */
always_ff @(posedge clk)
rpend_t0 <= _056_;
assign _011_ = | { rpend_t0, instr_t0[19:15] };
assign _012_ = | { rpend_t0, instr_t0[24:20] };
assign _057_ = rpend_t0 | instr_t0[19:15];
assign _058_ = rpend_t0 | instr_t0[24:20];
assign _007_ = ~ _057_;
assign _008_ = ~ _058_;
assign _034_ = rpend & _007_;
assign _036_ = rpend & _008_;
assign _035_ = instr[19:15] & _007_;
assign _037_ = instr[24:20] & _008_;
assign _063_ = _034_ == _035_;
assign _064_ = _036_ == _037_;
assign _066_ = _063_ & _011_;
assign _068_ = _064_ & _012_;
/* src = "generated/sv2v_out.v:898.2-900.16" */
/* PC_TAINT_INFO MODULE_NAME kronos_hcu */
/* PC_TAINT_INFO STATE_NAME rpend */
always_ff @(posedge clk)
if (_071_) rpend <= instr[11:7];
assign _038_ = decode_vld_t0 & decode_rdy;
assign _041_ = fetch_vld_t0 & fetch_rdy;
assign _039_ = decode_rdy_t0 & decode_vld;
assign _042_ = fetch_rdy_t0 & fetch_vld;
assign _040_ = decode_vld_t0 & decode_rdy_t0;
assign _043_ = fetch_vld_t0 & fetch_rdy_t0;
assign _059_ = _038_ | _039_;
assign _060_ = _041_ | _042_;
assign _070_ = _059_ | _040_;
assign _072_ = _060_ | _043_;
assign _009_ = ~ rs1_hazard;
assign _010_ = ~ rs2_hazard;
assign _044_ = rs1_hazard_t0 & _010_;
assign _045_ = rs2_hazard_t0 & _009_;
assign _046_ = rs1_hazard_t0 & rs2_hazard_t0;
assign _061_ = _044_ | _045_;
assign _076_ = _061_ | _046_;
assign _065_ = rpend == /* src = "generated/sv2v_out.v:895.56-895.68" */ instr[19:15];
assign _067_ = rpend == /* src = "generated/sv2v_out.v:896.56-896.68" */ instr[24:20];
assign _069_ = decode_vld && /* src = "generated/sv2v_out.v:897.60-897.84" */ decode_rdy;
assign _071_ = fetch_vld && /* src = "generated/sv2v_out.v:899.7-899.29" */ fetch_rdy;
assign _073_ = ~ /* src = "generated/sv2v_out.v:897.58-897.85" */ _069_;
assign _074_ = ~ /* src = "generated/sv2v_out.v:897.45-897.86" */ _004_;
assign _075_ = rs1_hazard | /* src = "generated/sv2v_out.v:897.18-897.41" */ rs2_hazard;
// Added block to randomize initial values.
`ifdef RANDOMIZE_INIT
  initial begin
    rpend_t0 = '0;
    rpend = '0;
  end
`endif // RANDOMIZE_INIT
endmodule

module kronos_lsu(decode, lsu_vld, lsu_rdy, load_data, regwr_lsu, data_addr, data_rd_data, data_wr_data, data_mask, data_wr_en, data_req, data_ack, load_data_t0, decode_t0, data_ack_t0, data_addr_t0, data_mask_t0, data_rd_data_t0, data_req_t0, data_wr_data_t0, data_wr_en_t0
, lsu_rdy_t0, lsu_vld_t0, regwr_lsu_t0);
/* src = "generated/sv2v_out.v:1474.2-1480.26" */
wire [31:0] _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1474.2-1480.26" */
wire [31:0] _001_;
wire _002_;
wire _003_;
wire [31:0] _004_;
wire [31:0] _005_;
wire [31:0] _006_;
wire [1:0] _007_;
wire [4:0] _008_;
wire _009_;
wire _010_;
wire [31:0] _011_;
wire [31:0] _012_;
wire [31:0] _013_;
wire [1:0] _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire [31:0] _023_;
wire [31:0] _024_;
wire [31:0] _025_;
wire [31:0] _026_;
wire [31:0] _027_;
wire [31:0] _028_;
wire [31:0] _029_;
wire [31:0] _030_;
wire [31:0] _031_;
wire [1:0] _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire [4:0] _048_;
wire _049_;
wire _050_;
wire _051_;
wire [31:0] _052_;
wire [31:0] _053_;
wire [31:0] _054_;
wire [31:0] _055_;
wire [31:0] _056_;
wire [31:0] _057_;
wire [31:0] _058_;
wire [31:0] _059_;
wire [31:0] _060_;
wire [31:0] _061_;
wire [31:0] _062_;
wire [31:0] _063_;
wire [1:0] _064_;
wire _065_;
/* cellift = 32'd1 */
wire _066_;
wire _067_;
wire [31:0] _068_;
wire [31:0] _069_;
wire [31:0] _070_;
wire [31:0] _071_;
wire [31:0] _072_;
wire [31:0] _073_;
wire [31:0] _074_;
wire [31:0] _075_;
wire [31:0] _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire [31:0] _083_;
wire [31:0] _084_;
wire [31:0] _085_;
wire [31:0] _086_;
wire [31:0] _087_;
wire [31:0] _088_;
wire [31:0] _089_;
wire [31:0] _090_;
wire [31:0] _091_;
wire [31:0] _092_;
wire [31:0] _093_;
wire [31:0] _094_;
wire [31:0] _095_;
wire [31:0] _096_;
wire [31:0] _097_;
wire [31:0] _098_;
wire [31:0] _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire [31:0] _104_;
/* cellift = 32'd1 */
wire [31:0] _105_;
wire [31:0] _106_;
/* cellift = 32'd1 */
wire [31:0] _107_;
/* src = "generated/sv2v_out.v:1475.7-1475.37" */
wire _108_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1475.7-1475.37" */
wire _109_;
/* src = "generated/sv2v_out.v:1477.12-1477.42" */
wire _110_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1477.12-1477.42" */
wire _111_;
/* src = "generated/sv2v_out.v:1450.23-1450.44" */
wire _112_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1450.23-1450.44" */
wire _113_;
/* src = "generated/sv2v_out.v:1451.21-1451.57" */
wire _114_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1451.21-1451.57" */
wire _115_;
/* src = "generated/sv2v_out.v:1453.36-1453.53" */
wire _116_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1453.36-1453.53" */
wire _117_;
/* src = "generated/sv2v_out.v:1450.49-1450.58" */
wire _118_;
/* src = "generated/sv2v_out.v:1451.33-1451.56" */
wire _119_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1451.33-1451.56" */
wire _120_;
wire _121_;
/* cellift = 32'd1 */
wire _122_;
wire _123_;
/* cellift = 32'd1 */
wire _124_;
wire _125_;
/* cellift = 32'd1 */
wire _126_;
/* src = "generated/sv2v_out.v:1442.13-1442.22" */
wire [31:0] byte_data;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1442.13-1442.22" */
wire [31:0] byte_data_t0;
/* src = "generated/sv2v_out.v:1434.13-1434.21" */
input data_ack;
wire data_ack;
/* cellift = 32'd1 */
input data_ack_t0;
wire data_ack_t0;
/* src = "generated/sv2v_out.v:1428.21-1428.30" */
output [31:0] data_addr;
wire [31:0] data_addr;
/* cellift = 32'd1 */
output [31:0] data_addr_t0;
wire [31:0] data_addr_t0;
/* src = "generated/sv2v_out.v:1431.20-1431.29" */
output [3:0] data_mask;
wire [3:0] data_mask;
/* cellift = 32'd1 */
output [3:0] data_mask_t0;
wire [3:0] data_mask_t0;
/* src = "generated/sv2v_out.v:1429.20-1429.32" */
input [31:0] data_rd_data;
wire [31:0] data_rd_data;
/* cellift = 32'd1 */
input [31:0] data_rd_data_t0;
wire [31:0] data_rd_data_t0;
/* src = "generated/sv2v_out.v:1433.14-1433.22" */
output data_req;
wire data_req;
/* cellift = 32'd1 */
output data_req_t0;
wire data_req_t0;
/* src = "generated/sv2v_out.v:1430.21-1430.33" */
output [31:0] data_wr_data;
wire [31:0] data_wr_data;
/* cellift = 32'd1 */
output [31:0] data_wr_data_t0;
wire [31:0] data_wr_data_t0;
/* src = "generated/sv2v_out.v:1432.14-1432.24" */
output data_wr_en;
wire data_wr_en;
/* cellift = 32'd1 */
output data_wr_en_t0;
wire data_wr_en_t0;
/* src = "generated/sv2v_out.v:1423.21-1423.27" */
input [180:0] decode;
wire [180:0] decode;
/* cellift = 32'd1 */
input [180:0] decode_t0;
wire [180:0] decode_t0;
/* src = "generated/sv2v_out.v:1441.13-1441.22" */
wire [31:0] half_data;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1441.13-1441.22" */
wire [31:0] half_data_t0;
/* src = "generated/sv2v_out.v:1426.20-1426.29" */
output [31:0] load_data;
wire [31:0] load_data;
/* cellift = 32'd1 */
output [31:0] load_data_t0;
wire [31:0] load_data_t0;
/* src = "generated/sv2v_out.v:1425.14-1425.21" */
output lsu_rdy;
wire lsu_rdy;
/* cellift = 32'd1 */
output lsu_rdy_t0;
wire lsu_rdy_t0;
/* src = "generated/sv2v_out.v:1424.13-1424.20" */
input lsu_vld;
wire lsu_vld;
/* cellift = 32'd1 */
input lsu_vld_t0;
wire lsu_vld_t0;
/* src = "generated/sv2v_out.v:1427.14-1427.23" */
output regwr_lsu;
wire regwr_lsu;
/* cellift = 32'd1 */
output regwr_lsu_t0;
wire regwr_lsu_t0;
/* src = "generated/sv2v_out.v:1440.13-1440.22" */
wire [31:0] word_data;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1440.13-1440.22" */
wire [31:0] word_data_t0;
assign _015_ = | decode_t0[130:129];
assign _017_ = | decode_t0[22:21];
assign _007_ = ~ decode_t0[130:129];
assign _014_ = ~ decode_t0[22:21];
assign _032_ = decode[130:129] & _007_;
assign _064_ = decode[22:21] & _014_;
assign _100_ = _032_ == { 1'h0, _007_[0] };
assign _101_ = _064_ == _014_;
assign _102_ = _064_ == { _014_[1], 1'h0 };
assign _103_ = _064_ == { 1'h0, _014_[0] };
assign _111_ = _100_ & _015_;
assign _122_ = _101_ & _017_;
assign _124_ = _102_ & _017_;
assign _126_ = _103_ & _017_;
assign _033_ = lsu_vld_t0 & decode[11];
assign _036_ = _113_ & _118_;
assign _039_ = lsu_vld_t0 & _119_;
assign _042_ = _115_ & _118_;
assign _045_ = decode_t0[12] & _116_;
assign _034_ = decode_t0[11] & lsu_vld;
assign _037_ = data_ack_t0 & _112_;
assign _040_ = _120_ & lsu_vld;
assign _043_ = data_ack_t0 & _114_;
assign _046_ = _117_ & decode[12];
assign _035_ = lsu_vld_t0 & decode_t0[11];
assign _038_ = _113_ & data_ack_t0;
assign _041_ = lsu_vld_t0 & _120_;
assign _044_ = _115_ & data_ack_t0;
assign _047_ = decode_t0[12] & _117_;
assign _077_ = _033_ | _034_;
assign _078_ = _036_ | _037_;
assign _079_ = _039_ | _040_;
assign _080_ = _042_ | _043_;
assign _081_ = _045_ | _046_;
assign _113_ = _077_ | _035_;
assign data_wr_en_t0 = _078_ | _038_;
assign _115_ = _079_ | _041_;
assign data_req_t0 = _080_ | _044_;
assign regwr_lsu_t0 = _081_ | _047_;
assign _016_ = | decode_t0[128:124];
assign _008_ = ~ decode_t0[128:124];
assign _048_ = decode[128:124] & _008_;
assign _018_ = ! _032_;
assign _019_ = ! _048_;
assign _109_ = _018_ & _015_;
assign _117_ = _019_ & _016_;
assign _004_ = ~ { _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_ };
assign _005_ = ~ { _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_ };
assign _006_ = ~ { _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_ };
assign _011_ = ~ { _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_ };
assign _012_ = ~ { _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_ };
assign _013_ = ~ { decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131] };
assign _068_ = { _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_ } | _004_;
assign _071_ = { _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_ } | _005_;
assign _074_ = { _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_ } | _006_;
assign _083_ = { _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_ } | _011_;
assign _086_ = { _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_ } | _012_;
assign _089_ = { decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131] } | _013_;
assign _069_ = { _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_ } | { _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_ };
assign _072_ = { _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_ } | { _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_, _125_ };
assign _075_ = { _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_ } | { _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_, _065_ };
assign _084_ = { _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_ } | { _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_, _110_ };
assign _087_ = { _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_ } | { _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_ };
assign _090_ = { decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131] } | { decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131], decode[131] };
assign _023_ = { data_rd_data_t0[15:0], data_rd_data_t0[31:16] } & _068_;
assign _026_ = data_rd_data_t0 & _071_;
assign _029_ = _107_ & _074_;
assign _052_ = word_data_t0 & _083_;
assign _055_ = _001_ & _086_;
assign _058_ = { word_data_t0[15], word_data_t0[15], word_data_t0[15], word_data_t0[15], word_data_t0[15], word_data_t0[15], word_data_t0[15], word_data_t0[15], word_data_t0[15], word_data_t0[15], word_data_t0[15], word_data_t0[15], word_data_t0[15], word_data_t0[15], word_data_t0[15], word_data_t0[15], word_data_t0[15:0] } & _089_;
assign _061_ = { word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7], word_data_t0[7:0] } & _089_;
assign _024_ = { data_rd_data_t0[23:0], data_rd_data_t0[31:24] } & _069_;
assign _027_ = { data_rd_data_t0[7:0], data_rd_data_t0[31:8] } & _072_;
assign _030_ = _105_ & _075_;
assign _053_ = half_data_t0 & _084_;
assign _056_ = byte_data_t0 & _087_;
assign _059_ = { 16'h0000, word_data_t0[15:0] } & _090_;
assign _062_ = { 24'h000000, word_data_t0[7:0] } & _090_;
assign _070_ = _023_ | _024_;
assign _073_ = _026_ | _027_;
assign _076_ = _029_ | _030_;
assign _085_ = _052_ | _053_;
assign _088_ = _055_ | _056_;
assign _091_ = _058_ | _059_;
assign _092_ = _061_ | _062_;
assign _093_ = { data_rd_data[15:0], data_rd_data[31:16] } ^ { data_rd_data[23:0], data_rd_data[31:24] };
assign _094_ = data_rd_data ^ { data_rd_data[7:0], data_rd_data[31:8] };
assign _095_ = _106_ ^ _104_;
assign _096_ = word_data ^ half_data;
assign _097_ = _000_ ^ byte_data;
assign _098_ = { word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15:0] } ^ { 16'h0000, word_data[15:0] };
assign _099_ = { word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7:0] } ^ { 24'h000000, word_data[7:0] };
assign _025_ = { _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_, _122_ } & _093_;
assign _028_ = { _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_, _126_ } & _094_;
assign _031_ = { _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_, _066_ } & _095_;
assign _054_ = { _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_, _111_ } & _096_;
assign _057_ = { _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_ } & _097_;
assign _060_ = { decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131] } & _098_;
assign _063_ = { decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131], decode_t0[131] } & _099_;
assign _105_ = _025_ | _070_;
assign _107_ = _028_ | _073_;
assign word_data_t0 = _031_ | _076_;
assign _001_ = _054_ | _085_;
assign load_data_t0 = _057_ | _088_;
assign half_data_t0 = _060_ | _091_;
assign byte_data_t0 = _063_ | _092_;
assign _002_ = ~ _123_;
assign _009_ = ~ decode[12];
assign _003_ = ~ _121_;
assign _010_ = ~ decode[11];
assign _020_ = _124_ & _003_;
assign _049_ = decode_t0[12] & _010_;
assign _021_ = _122_ & _002_;
assign _050_ = decode_t0[11] & _009_;
assign _022_ = _124_ & _122_;
assign _051_ = decode_t0[12] & decode_t0[11];
assign _067_ = _020_ | _021_;
assign _082_ = _049_ | _050_;
assign _066_ = _067_ | _022_;
assign _120_ = _082_ | _051_;
assign _065_ = _123_ | _121_;
assign _104_ = _121_ ? { data_rd_data[23:0], data_rd_data[31:24] } : { data_rd_data[15:0], data_rd_data[31:16] };
assign _106_ = _125_ ? { data_rd_data[7:0], data_rd_data[31:8] } : data_rd_data;
assign word_data = _065_ ? _104_ : _106_;
assign _108_ = ! /* src = "generated/sv2v_out.v:1475.7-1475.37" */ decode[130:129];
assign _110_ = decode[130:129] == /* src = "generated/sv2v_out.v:1477.12-1477.42" */ 2'h1;
assign _112_ = lsu_vld && /* src = "generated/sv2v_out.v:1450.23-1450.44" */ decode[11];
assign data_wr_en = _112_ && /* src = "generated/sv2v_out.v:1450.22-1450.58" */ _118_;
assign _114_ = lsu_vld && /* src = "generated/sv2v_out.v:1451.21-1451.57" */ _119_;
assign data_req = _114_ && /* src = "generated/sv2v_out.v:1451.20-1451.71" */ _118_;
assign regwr_lsu = decode[12] && /* src = "generated/sv2v_out.v:1453.21-1453.54" */ _116_;
assign _116_ = | /* src = "generated/sv2v_out.v:1453.36-1453.53" */ decode[128:124];
assign _118_ = ~ /* src = "generated/sv2v_out.v:1451.62-1451.71" */ data_ack;
assign _119_ = decode[12] | /* src = "generated/sv2v_out.v:1451.33-1451.56" */ decode[11];
assign _000_ = _110_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1477.12-1477.42|generated/sv2v_out.v:1477.8-1480.26" */ half_data : word_data;
assign load_data = _108_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1475.7-1475.37|generated/sv2v_out.v:1475.3-1480.26" */ byte_data : _000_;
assign half_data = decode[131] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1467.7-1467.15|generated/sv2v_out.v:1467.3-1470.56" */ { 16'h0000, word_data[15:0] } : { word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15], word_data[15:0] };
assign byte_data = decode[131] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:1463.7-1463.15|generated/sv2v_out.v:1463.3-1466.54" */ { 24'h000000, word_data[7:0] } : { word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7], word_data[7:0] };
assign _121_ = decode[22:21] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1456.3-1461.10" */ 2'h3;
assign _123_ = decode[22:21] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1456.3-1461.10" */ 2'h2;
assign _125_ = decode[22:21] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:1456.3-1461.10" */ 2'h1;
assign data_addr = { decode[52:23], 2'h0 };
assign data_addr_t0 = { decode_t0[52:23], 2'h0 };
assign data_mask = decode[10:7];
assign data_mask_t0 = decode_t0[10:7];
assign data_wr_data = decode[84:53];
assign data_wr_data_t0 = decode_t0[84:53];
assign lsu_rdy = data_ack;
assign lsu_rdy_t0 = data_ack_t0;
endmodule

module kronos_mem_top(clk_i, rst_ni, data_mem_req, data_mem_gnt, data_mem_addr, data_mem_wdata, data_mem_strb, data_mem_we, data_mem_rdata, instr_mem_req, instr_mem_gnt, instr_mem_addr, instr_mem_wdata, instr_mem_strb, instr_mem_we, instr_mem_rdata, software_interrupt, timer_interrupt, external_interrupt, timer_interrupt_t0, software_interrupt_t0
, external_interrupt_t0, data_mem_addr_t0, data_mem_gnt_t0, data_mem_rdata_t0, data_mem_req_t0, data_mem_strb_t0, data_mem_wdata_t0, data_mem_we_t0, instr_mem_addr_t0, instr_mem_gnt_t0, instr_mem_rdata_t0, instr_mem_req_t0, instr_mem_strb_t0, instr_mem_wdata_t0, instr_mem_we_t0);
/* src = "generated/sv2v_out.v:1720.8-1720.13" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:1749.7-1749.15" */
reg data_ack;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1749.7-1749.15" */
reg data_ack_t0;
/* src = "generated/sv2v_out.v:1743.14-1743.23" */
/* unused_bits = "20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] data_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1743.14-1743.23" */
/* unused_bits = "20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] data_addr_t0;
/* src = "generated/sv2v_out.v:1746.13-1746.22" */
wire [3:0] data_mask;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1746.13-1746.22" */
wire [3:0] data_mask_t0;
/* src = "generated/sv2v_out.v:1724.21-1724.34" */
output [19:0] data_mem_addr;
wire [19:0] data_mem_addr;
/* cellift = 32'd1 */
output [19:0] data_mem_addr_t0;
wire [19:0] data_mem_addr_t0;
/* src = "generated/sv2v_out.v:1723.13-1723.25" */
input data_mem_gnt;
wire data_mem_gnt;
/* cellift = 32'd1 */
input data_mem_gnt_t0;
wire data_mem_gnt_t0;
/* src = "generated/sv2v_out.v:1728.20-1728.34" */
input [31:0] data_mem_rdata;
wire [31:0] data_mem_rdata;
/* cellift = 32'd1 */
input [31:0] data_mem_rdata_t0;
wire [31:0] data_mem_rdata_t0;
/* src = "generated/sv2v_out.v:1722.14-1722.26" */
output data_mem_req;
wire data_mem_req;
/* cellift = 32'd1 */
output data_mem_req_t0;
wire data_mem_req_t0;
/* src = "generated/sv2v_out.v:1726.21-1726.34" */
output [31:0] data_mem_strb;
wire [31:0] data_mem_strb;
/* cellift = 32'd1 */
output [31:0] data_mem_strb_t0;
wire [31:0] data_mem_strb_t0;
/* src = "generated/sv2v_out.v:1725.21-1725.35" */
output [31:0] data_mem_wdata;
wire [31:0] data_mem_wdata;
/* cellift = 32'd1 */
output [31:0] data_mem_wdata_t0;
wire [31:0] data_mem_wdata_t0;
/* src = "generated/sv2v_out.v:1727.14-1727.25" */
output data_mem_we;
wire data_mem_we;
/* cellift = 32'd1 */
output data_mem_we_t0;
wire data_mem_we_t0;
/* src = "generated/sv2v_out.v:1738.13-1738.31" */
input external_interrupt;
wire external_interrupt;
/* cellift = 32'd1 */
input external_interrupt_t0;
wire external_interrupt_t0;
/* src = "generated/sv2v_out.v:1742.7-1742.16" */
reg instr_ack;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1742.7-1742.16" */
reg instr_ack_t0;
/* src = "generated/sv2v_out.v:1739.14-1739.24" */
/* unused_bits = "20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] instr_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:1739.14-1739.24" */
/* unused_bits = "20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] instr_addr_t0;
/* src = "generated/sv2v_out.v:1731.21-1731.35" */
output [19:0] instr_mem_addr;
wire [19:0] instr_mem_addr;
/* cellift = 32'd1 */
output [19:0] instr_mem_addr_t0;
wire [19:0] instr_mem_addr_t0;
/* src = "generated/sv2v_out.v:1730.13-1730.26" */
input instr_mem_gnt;
wire instr_mem_gnt;
/* cellift = 32'd1 */
input instr_mem_gnt_t0;
wire instr_mem_gnt_t0;
/* src = "generated/sv2v_out.v:1735.20-1735.35" */
input [31:0] instr_mem_rdata;
wire [31:0] instr_mem_rdata;
/* cellift = 32'd1 */
input [31:0] instr_mem_rdata_t0;
wire [31:0] instr_mem_rdata_t0;
/* src = "generated/sv2v_out.v:1729.14-1729.27" */
output instr_mem_req;
wire instr_mem_req;
/* cellift = 32'd1 */
output instr_mem_req_t0;
wire instr_mem_req_t0;
/* src = "generated/sv2v_out.v:1733.21-1733.35" */
output [31:0] instr_mem_strb;
wire [31:0] instr_mem_strb;
/* cellift = 32'd1 */
output [31:0] instr_mem_strb_t0;
wire [31:0] instr_mem_strb_t0;
/* src = "generated/sv2v_out.v:1732.21-1732.36" */
output [31:0] instr_mem_wdata;
wire [31:0] instr_mem_wdata;
/* cellift = 32'd1 */
output [31:0] instr_mem_wdata_t0;
wire [31:0] instr_mem_wdata_t0;
/* src = "generated/sv2v_out.v:1734.14-1734.26" */
output instr_mem_we;
wire instr_mem_we;
/* cellift = 32'd1 */
output instr_mem_we_t0;
wire instr_mem_we_t0;
/* src = "generated/sv2v_out.v:1721.8-1721.14" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:1736.13-1736.31" */
input software_interrupt;
wire software_interrupt;
/* cellift = 32'd1 */
input software_interrupt_t0;
wire software_interrupt_t0;
/* src = "generated/sv2v_out.v:1737.13-1737.28" */
input timer_interrupt;
wire timer_interrupt;
/* cellift = 32'd1 */
input timer_interrupt_t0;
wire timer_interrupt_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_mem_top */
/* PC_TAINT_INFO STATE_NAME instr_ack_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_ack_t0 <= 1'h0;
else instr_ack_t0 <= instr_mem_req_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME kronos_mem_top */
/* PC_TAINT_INFO STATE_NAME data_ack_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) data_ack_t0 <= 1'h0;
else data_ack_t0 <= data_mem_req_t0;
/* src = "generated/sv2v_out.v:1756.2-1764.6" */
/* PC_TAINT_INFO MODULE_NAME kronos_mem_top */
/* PC_TAINT_INFO STATE_NAME instr_ack */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_ack <= 1'h0;
else instr_ack <= instr_mem_req;
/* src = "generated/sv2v_out.v:1756.2-1764.6" */
/* PC_TAINT_INFO MODULE_NAME kronos_mem_top */
/* PC_TAINT_INFO STATE_NAME data_ack */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) data_ack <= 1'h0;
else data_ack <= data_mem_req;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:1787.4-1804.3" */
paramodsimplif_1b215dccbb32fdcc253c  i_kronos_core (
.clk(clk_i),
.data_ack(data_ack),
.data_ack_t0(data_ack_t0),
.data_addr(data_addr),
.data_addr_t0(data_addr_t0),
.data_mask(data_mask),
.data_mask_t0(data_mask_t0),
.data_rd_data(data_mem_rdata),
.data_rd_data_t0(data_mem_rdata_t0),
.data_req(data_mem_req),
.data_req_t0(data_mem_req_t0),
.data_wr_data(data_mem_wdata),
.data_wr_data_t0(data_mem_wdata_t0),
.data_wr_en(data_mem_we),
.data_wr_en_t0(data_mem_we_t0),
.external_interrupt(external_interrupt),
.external_interrupt_t0(external_interrupt_t0),
.instr_ack(instr_ack),
.instr_ack_t0(instr_ack_t0),
.instr_addr(instr_addr),
.instr_addr_t0(instr_addr_t0),
.instr_data(instr_mem_rdata),
.instr_data_t0(instr_mem_rdata_t0),
.instr_req(instr_mem_req),
.instr_req_t0(instr_mem_req_t0),
.rstz(rst_ni),
.software_interrupt(software_interrupt),
.software_interrupt_t0(software_interrupt_t0),
.timer_interrupt(timer_interrupt),
.timer_interrupt_t0(timer_interrupt_t0)
);
assign data_mem_addr = data_addr[19:0];
assign data_mem_addr_t0 = data_addr_t0[19:0];
assign data_mem_strb = { data_mask[3], data_mask[3], data_mask[3], data_mask[3], data_mask[3], data_mask[3], data_mask[3], data_mask[3:2], data_mask[2], data_mask[2], data_mask[2], data_mask[2], data_mask[2], data_mask[2], data_mask[2:1], data_mask[1], data_mask[1], data_mask[1], data_mask[1], data_mask[1], data_mask[1], data_mask[1:0], data_mask[0], data_mask[0], data_mask[0], data_mask[0], data_mask[0], data_mask[0], data_mask[0] };
assign data_mem_strb_t0 = { data_mask_t0[3], data_mask_t0[3], data_mask_t0[3], data_mask_t0[3], data_mask_t0[3], data_mask_t0[3], data_mask_t0[3], data_mask_t0[3:2], data_mask_t0[2], data_mask_t0[2], data_mask_t0[2], data_mask_t0[2], data_mask_t0[2], data_mask_t0[2], data_mask_t0[2:1], data_mask_t0[1], data_mask_t0[1], data_mask_t0[1], data_mask_t0[1], data_mask_t0[1], data_mask_t0[1], data_mask_t0[1:0], data_mask_t0[0], data_mask_t0[0], data_mask_t0[0], data_mask_t0[0], data_mask_t0[0], data_mask_t0[0], data_mask_t0[0] };
assign instr_mem_addr = instr_addr[19:0];
assign instr_mem_addr_t0 = instr_addr_t0[19:0];
assign instr_mem_strb = 32'd0;
assign instr_mem_strb_t0 = 32'd0;
assign instr_mem_wdata = 32'd0;
assign instr_mem_wdata_t0 = 32'd0;
assign instr_mem_we = 1'h0;
assign instr_mem_we_t0 = 1'h0;
endmodule