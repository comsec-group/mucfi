
`ifdef CRYPTO
`include "../common/formal/signal_defs/crypto_start_cond_reg.sv"
`endif

bit taint_start_cond_DIV_op1;
assign taint_start_cond_DIV_op1 = cpuregs_rs1_start_cond && DIV(instr_word);

bit taint_start_cond_DIV_op2;
assign taint_start_cond_DIV_op2 = cpuregs_rs2_start_cond && DIV(instr_word);

bit taint_start_cond_DIVU_op1;
assign taint_start_cond_DIVU_op1 = cpuregs_rs1_start_cond && DIVU(instr_word);

bit taint_start_cond_DIVU_op2;
assign taint_start_cond_DIVU_op2 = cpuregs_rs2_start_cond && DIV(instr_word);

bit taint_start_cond_MUL_op1;
assign taint_start_cond_MUL_op1 = cpuregs_rs1_start_cond && MUL(instr_word);

bit taint_start_cond_MUL_op2;
assign taint_start_cond_MUL_op2 = cpuregs_rs2_start_cond && MUL(instr_word);

bit taint_start_cond_MULH_op1;
assign taint_start_cond_MULH_op1 = cpuregs_rs1_start_cond && MULH(instr_word);

bit taint_start_cond_MULH_op2;
assign taint_start_cond_MULH_op2 = cpuregs_rs2_start_cond && MULH(instr_word);

bit taint_start_cond_MULHSU_op1;
assign taint_start_cond_MULHSU_op1 = cpuregs_rs1_start_cond && MULHSU(instr_word);

bit taint_start_cond_MULHSU_op2;
assign taint_start_cond_MULHSU_op2 = cpuregs_rs2_start_cond && MULHSU(instr_word);

bit taint_start_cond_MULHU_op1;
assign taint_start_cond_MULHU_op1 = cpuregs_rs1_start_cond && MULHU(instr_word);

bit taint_start_cond_MULHU_op2;
assign taint_start_cond_MULHU_op2 = cpuregs_rs2_start_cond && MULHU(instr_word);


bit taint_start_cond_REM_op1;
assign taint_start_cond_REM_op1 = cpuregs_rs1_start_cond && REM(instr_word);

bit taint_start_cond_REM_op2;
assign taint_start_cond_REM_op2 = cpuregs_rs2_start_cond && REM(instr_word);

bit taint_start_cond_REMU_op1;
assign taint_start_cond_REMU_op1 = cpuregs_rs1_start_cond && REMU(instr_word);

bit taint_start_cond_REMU_op2;
assign taint_start_cond_REMU_op2 = cpuregs_rs2_start_cond && REMU(instr_word);





// Generated by gen_checker_inst.py
bit taint_start_cond_CSRRS_op1;
assign taint_start_cond_CSRRS_op1 = cpuregs_rs1_start_cond && CSRRS(instr_word);

bit taint_start_cond_SRLI_op1;
assign taint_start_cond_SRLI_op1 = cpuregs_rs1_start_cond && SRLI(instr_word);

bit taint_start_cond_BEQ_op1;
assign taint_start_cond_BEQ_op1 = cpuregs_rs1_start_cond && BEQ(instr_word);

bit taint_start_cond_BEQ_op2;
assign taint_start_cond_BEQ_op2 = cpuregs_rs2_start_cond && BEQ(instr_word);

bit taint_start_cond_SLT_op1;
assign taint_start_cond_SLT_op1 = cpuregs_rs1_start_cond && SLT(instr_word);

bit taint_start_cond_SLT_op2;
assign taint_start_cond_SLT_op2 = cpuregs_rs2_start_cond && SLT(instr_word);

bit taint_start_cond_ADDI_op1;
assign taint_start_cond_ADDI_op1 = cpuregs_rs1_start_cond && ADDI(instr_word);

bit taint_start_cond_ORI_op1;
assign taint_start_cond_ORI_op1 = cpuregs_rs1_start_cond && ORI(instr_word);

bit taint_start_cond_SUB_op1;
assign taint_start_cond_SUB_op1 = cpuregs_rs1_start_cond && SUB(instr_word);

bit taint_start_cond_SUB_op2;
assign taint_start_cond_SUB_op2 = cpuregs_rs2_start_cond && SUB(instr_word);

bit taint_start_cond_AND_op1;
assign taint_start_cond_AND_op1 = cpuregs_rs1_start_cond && AND(instr_word);

bit taint_start_cond_AND_op2;
assign taint_start_cond_AND_op2 = cpuregs_rs2_start_cond && AND(instr_word);

bit taint_start_cond_ADD_op1;
assign taint_start_cond_ADD_op1 = cpuregs_rs1_start_cond && ADD(instr_word);

bit taint_start_cond_ADD_op2;
assign taint_start_cond_ADD_op2 = cpuregs_rs2_start_cond && ADD(instr_word);

bit taint_start_cond_CSRRC_op1;
assign taint_start_cond_CSRRC_op1 = cpuregs_rs1_start_cond && CSRRC(instr_word);

bit taint_start_cond_FENCE_op1;
assign taint_start_cond_FENCE_op1 = cpuregs_rs1_start_cond && FENCE(instr_word);

bit taint_start_cond_LH_op1;
assign taint_start_cond_LH_op1 = cpuregs_rs1_start_cond && LH(instr_word);

bit taint_start_cond_ANDI_op1;
assign taint_start_cond_ANDI_op1 = cpuregs_rs1_start_cond && ANDI(instr_word);

bit taint_start_cond_SLLI_op1;
assign taint_start_cond_SLLI_op1 = cpuregs_rs1_start_cond && SLLI(instr_word);

bit taint_start_cond_CSRRWI_op1;
assign taint_start_cond_CSRRWI_op1 = cpuregs_rs1_start_cond && CSRRWI(instr_word);

bit taint_start_cond_SRA_op1;
assign taint_start_cond_SRA_op1 = cpuregs_rs1_start_cond && SRA(instr_word);

bit taint_start_cond_SRA_op2;
assign taint_start_cond_SRA_op2 = cpuregs_rs2_start_cond && SRA(instr_word);

bit taint_start_cond_JALR_op1;
assign taint_start_cond_JALR_op1 = cpuregs_rs1_start_cond && JALR(instr_word);

bit taint_start_cond_OR_op1;
assign taint_start_cond_OR_op1 = cpuregs_rs1_start_cond && OR(instr_word);

bit taint_start_cond_OR_op2;
assign taint_start_cond_OR_op2 = cpuregs_rs2_start_cond && OR(instr_word);

bit taint_start_cond_FENCE_I_op1;
assign taint_start_cond_FENCE_I_op1 = cpuregs_rs1_start_cond && FENCE_I(instr_word);

bit taint_start_cond_CSRRSI_op1;
assign taint_start_cond_CSRRSI_op1 = cpuregs_rs1_start_cond && CSRRSI(instr_word);

bit taint_start_cond_SW_op1;
assign taint_start_cond_SW_op1 = cpuregs_rs1_start_cond && SW(instr_word);

bit taint_start_cond_SLL_op1;
assign taint_start_cond_SLL_op1 = cpuregs_rs1_start_cond && SLL(instr_word);

bit taint_start_cond_SLL_op2;
assign taint_start_cond_SLL_op2 = cpuregs_rs2_start_cond && SLL(instr_word);

bit taint_start_cond_CSRRW_op1;
assign taint_start_cond_CSRRW_op1 = cpuregs_rs1_start_cond && CSRRW(instr_word);

bit taint_start_cond_SH_op1;
assign taint_start_cond_SH_op1 = cpuregs_rs1_start_cond && SH(instr_word);

bit taint_start_cond_SLTI_op1;
assign taint_start_cond_SLTI_op1 = cpuregs_rs1_start_cond && SLTI(instr_word);

bit taint_start_cond_LBU_op1;
assign taint_start_cond_LBU_op1 = cpuregs_rs1_start_cond && LBU(instr_word);

bit taint_start_cond_XOR_op1;
assign taint_start_cond_XOR_op1 = cpuregs_rs1_start_cond && XOR(instr_word);

bit taint_start_cond_XOR_op2;
assign taint_start_cond_XOR_op2 = cpuregs_rs2_start_cond && XOR(instr_word);

bit taint_start_cond_EBREAK_op1;
assign taint_start_cond_EBREAK_op1 = cpuregs_rs1_start_cond && EBREAK(instr_word);

bit taint_start_cond_SRAI_op1;
assign taint_start_cond_SRAI_op1 = cpuregs_rs1_start_cond && SRAI(instr_word);

bit taint_start_cond_LB_op1;
assign taint_start_cond_LB_op1 = cpuregs_rs1_start_cond && LB(instr_word);

bit taint_start_cond_BLT_op1;
assign taint_start_cond_BLT_op1 = cpuregs_rs1_start_cond && BLT(instr_word);

bit taint_start_cond_BLT_op2;
assign taint_start_cond_BLT_op2 = cpuregs_rs2_start_cond && BLT(instr_word);

bit taint_start_cond_SLTIU_op1;
assign taint_start_cond_SLTIU_op1 = cpuregs_rs1_start_cond && SLTIU(instr_word);

bit taint_start_cond_LHU_op1;
assign taint_start_cond_LHU_op1 = cpuregs_rs1_start_cond && LHU(instr_word);

bit taint_start_cond_BGE_op1;
assign taint_start_cond_BGE_op1 = cpuregs_rs1_start_cond && BGE(instr_word);

bit taint_start_cond_BGE_op2;
assign taint_start_cond_BGE_op2 = cpuregs_rs2_start_cond && BGE(instr_word);

bit taint_start_cond_BNE_op1;
assign taint_start_cond_BNE_op1 = cpuregs_rs1_start_cond && BNE(instr_word);

bit taint_start_cond_BNE_op2;
assign taint_start_cond_BNE_op2 = cpuregs_rs2_start_cond && BNE(instr_word);

bit taint_start_cond_XORI_op1;
assign taint_start_cond_XORI_op1 = cpuregs_rs1_start_cond && XORI(instr_word);

bit taint_start_cond_SRL_op1;
assign taint_start_cond_SRL_op1 = cpuregs_rs1_start_cond && SRL(instr_word);

bit taint_start_cond_SRL_op2;
assign taint_start_cond_SRL_op2 = cpuregs_rs2_start_cond && SRL(instr_word);

bit taint_start_cond_SB_op1;
assign taint_start_cond_SB_op1 = cpuregs_rs1_start_cond && SB(instr_word);

bit taint_start_cond_BGEU_op1;
assign taint_start_cond_BGEU_op1 = cpuregs_rs1_start_cond && BGEU(instr_word);

bit taint_start_cond_BGEU_op2;
assign taint_start_cond_BGEU_op2 = cpuregs_rs2_start_cond && BGEU(instr_word);

bit taint_start_cond_LW_op1;
assign taint_start_cond_LW_op1 = cpuregs_rs1_start_cond && LW(instr_word);

bit taint_start_cond_CSRRCI_op1;
assign taint_start_cond_CSRRCI_op1 = cpuregs_rs1_start_cond && CSRRCI(instr_word);

bit taint_start_cond_BLTU_op1;
assign taint_start_cond_BLTU_op1 = cpuregs_rs1_start_cond && BLTU(instr_word);

bit taint_start_cond_BLTU_op2;
assign taint_start_cond_BLTU_op2 = cpuregs_rs2_start_cond && BLTU(instr_word);

bit taint_start_cond_ECALL_op1;
assign taint_start_cond_ECALL_op1 = cpuregs_rs1_start_cond && EBREAK(instr_word);

bit taint_start_cond_SLTU_op1;
assign taint_start_cond_SLTU_op1 = cpuregs_rs1_start_cond && SLTU(instr_word);

bit taint_start_cond_SLTU_op2;
assign taint_start_cond_SLTU_op2 = cpuregs_rs2_start_cond && SLTU(instr_word);

