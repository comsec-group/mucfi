module \$paramod$34601000fe8707ce2501f5ed778e152043201712\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _0_;
wire [6:0] _1_;
wire [6:0] _2_;
wire [6:0] _3_;
/* src = "generated/sv2v_out.v:14894.13-14894.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14898.28-14898.37" */
output [6:0] rd_data_o;
reg [6:0] rd_data_o;
/* cellift = 32'd1 */
output [6:0] rd_data_o_t0;
reg [6:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14899.14-14899.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14895.13-14895.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14896.27-14896.36" */
input [6:0] wr_data_i;
wire [6:0] wr_data_i;
/* cellift = 32'd1 */
input [6:0] wr_data_i_t0;
wire [6:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14897.13-14897.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _0_ = ~ wr_en_i;
assign _1_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _2_ = { _0_, _0_, _0_, _0_, _0_, _0_, _0_ } & rd_data_o_t0;
assign _3_ = _1_ | _2_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$34601000fe8707ce2501f5ed778e152043201712\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 7'h00;
else rd_data_o_t0 <= _3_;
/* src = "generated/sv2v_out.v:14901.2-14905.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$34601000fe8707ce2501f5ed778e152043201712\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 7'h00;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$410b37fbfbfa994790f1902c150d2be939cadb3b\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _0_;
wire [2:0] _1_;
wire [2:0] _2_;
wire [2:0] _3_;
/* src = "generated/sv2v_out.v:14894.13-14894.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14898.28-14898.37" */
output [2:0] rd_data_o;
reg [2:0] rd_data_o;
/* cellift = 32'd1 */
output [2:0] rd_data_o_t0;
reg [2:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14899.14-14899.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14895.13-14895.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14896.27-14896.36" */
input [2:0] wr_data_i;
wire [2:0] wr_data_i;
/* cellift = 32'd1 */
input [2:0] wr_data_i_t0;
wire [2:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14897.13-14897.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _0_ = ~ wr_en_i;
assign _1_ = { wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _2_ = { _0_, _0_, _0_ } & rd_data_o_t0;
assign _3_ = _1_ | _2_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$410b37fbfbfa994790f1902c150d2be939cadb3b\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 3'h0;
else rd_data_o_t0 <= _3_;
/* src = "generated/sv2v_out.v:14901.2-14905.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$410b37fbfbfa994790f1902c150d2be939cadb3b\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 3'h4;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_flop (clk_i, rst_ni, d_i, q_o, d_i_t0, q_o_t0);
/* src = "generated/sv2v_out.v:24678.8-24678.13" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:24680.22-24680.25" */
input [3:0] d_i;
wire [3:0] d_i;
/* cellift = 32'd1 */
input [3:0] d_i_t0;
wire [3:0] d_i_t0;
/* src = "generated/sv2v_out.v:24681.28-24681.31" */
output [3:0] q_o;
wire [3:0] q_o;
/* cellift = 32'd1 */
output [3:0] q_o_t0;
wire [3:0] q_o_t0;
/* src = "generated/sv2v_out.v:24679.8-24679.14" */
input rst_ni;
wire rst_ni;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:24699.6-24704.5" */
\$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_generic_flop  \gen_generic.u_impl_generic  (
.clk_i(clk_i),
.d_i(d_i),
.d_i_t0(d_i_t0),
.q_o(q_o),
.q_o_t0(q_o_t0),
.rst_ni(rst_ni)
);
endmodule

module \$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_generic_flop (clk_i, rst_ni, d_i, q_o, d_i_t0, q_o_t0);
/* src = "generated/sv2v_out.v:24938.8-24938.13" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:24940.22-24940.25" */
input [3:0] d_i;
wire [3:0] d_i;
/* cellift = 32'd1 */
input [3:0] d_i_t0;
wire [3:0] d_i_t0;
/* src = "generated/sv2v_out.v:24941.27-24941.30" */
output [3:0] q_o;
reg [3:0] q_o;
/* cellift = 32'd1 */
output [3:0] q_o_t0;
reg [3:0] q_o_t0;
/* src = "generated/sv2v_out.v:24939.8-24939.14" */
input rst_ni;
wire rst_ni;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_generic_flop  */
/* PC_TAINT_INFO STATE_NAME q_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) q_o_t0 <= 4'h0;
else q_o_t0 <= d_i_t0;
/* src = "generated/sv2v_out.v:24942.2-24946.15" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_generic_flop  */
/* PC_TAINT_INFO STATE_NAME q_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) q_o <= 4'ha;
else q_o <= d_i;
endmodule

module \$paramod$4f46e25470a27719ee9ca03cee1a0827eff766f7\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _0_;
wire [31:0] _1_;
wire [31:0] _2_;
wire [31:0] _3_;
/* src = "generated/sv2v_out.v:14894.13-14894.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14898.28-14898.37" */
output [31:0] rd_data_o;
reg [31:0] rd_data_o;
/* cellift = 32'd1 */
output [31:0] rd_data_o_t0;
reg [31:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14899.14-14899.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14895.13-14895.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14896.27-14896.36" */
input [31:0] wr_data_i;
wire [31:0] wr_data_i;
/* cellift = 32'd1 */
input [31:0] wr_data_i_t0;
wire [31:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14897.13-14897.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _0_ = ~ wr_en_i;
assign _1_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _2_ = { _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_ } & rd_data_o_t0;
assign _3_ = _1_ | _2_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$4f46e25470a27719ee9ca03cee1a0827eff766f7\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 32'd0;
else rd_data_o_t0 <= _3_;
/* src = "generated/sv2v_out.v:14901.2-14905.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$4f46e25470a27719ee9ca03cee1a0827eff766f7\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 32'd1;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$501c60d7519704ee720c78ef16ad88cf05835059\ibex_dummy_instr (clk_i, rst_ni, dummy_instr_en_i, dummy_instr_mask_i, dummy_instr_seed_en_i, dummy_instr_seed_i, fetch_valid_i, id_in_ready_i, insert_dummy_instr_o, dummy_instr_data_o, insert_dummy_instr_o_t0, id_in_ready_i_t0, fetch_valid_i_t0, dummy_instr_seed_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_mask_i_t0, dummy_instr_en_i_t0, dummy_instr_data_o_t0);
/* src = "generated/sv2v_out.v:15874.25-15874.57" */
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire [31:0] _06_;
wire [31:0] _07_;
wire _08_;
wire [31:0] _09_;
wire [2:0] _10_;
/* src = "generated/sv2v_out.v:15880.50-15880.84" */
wire _11_;
/* src = "generated/sv2v_out.v:15874.62-15874.96" */
wire _12_;
wire _13_;
wire _14_;
wire _15_;
/* src = "generated/sv2v_out.v:15817.13-15817.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:15833.13-15833.24" */
wire [4:0] dummy_cnt_d;
/* src = "generated/sv2v_out.v:15835.7-15835.19" */
wire dummy_cnt_en;
/* src = "generated/sv2v_out.v:15831.13-15831.27" */
wire [4:0] dummy_cnt_incr;
/* src = "generated/sv2v_out.v:15834.12-15834.23" */
reg [4:0] dummy_cnt_q;
/* src = "generated/sv2v_out.v:15832.13-15832.32" */
wire [4:0] dummy_cnt_threshold;
/* src = "generated/sv2v_out.v:15826.21-15826.39" */
output [31:0] dummy_instr_data_o;
wire [31:0] dummy_instr_data_o;
/* cellift = 32'd1 */
output [31:0] dummy_instr_data_o_t0;
wire [31:0] dummy_instr_data_o_t0;
/* src = "generated/sv2v_out.v:15819.13-15819.29" */
input dummy_instr_en_i;
wire dummy_instr_en_i;
/* cellift = 32'd1 */
input dummy_instr_en_i_t0;
wire dummy_instr_en_i_t0;
/* src = "generated/sv2v_out.v:15820.19-15820.37" */
input [2:0] dummy_instr_mask_i;
wire [2:0] dummy_instr_mask_i;
/* cellift = 32'd1 */
input [2:0] dummy_instr_mask_i_t0;
wire [2:0] dummy_instr_mask_i_t0;
/* src = "generated/sv2v_out.v:15843.14-15843.32" */
wire [31:0] dummy_instr_seed_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15843.14-15843.32" */
wire [31:0] dummy_instr_seed_d_t0;
/* src = "generated/sv2v_out.v:15821.13-15821.34" */
input dummy_instr_seed_en_i;
wire dummy_instr_seed_en_i;
/* cellift = 32'd1 */
input dummy_instr_seed_en_i_t0;
wire dummy_instr_seed_en_i_t0;
/* src = "generated/sv2v_out.v:15822.20-15822.38" */
input [31:0] dummy_instr_seed_i;
wire [31:0] dummy_instr_seed_i;
/* cellift = 32'd1 */
input [31:0] dummy_instr_seed_i_t0;
wire [31:0] dummy_instr_seed_i_t0;
/* src = "generated/sv2v_out.v:15842.13-15842.31" */
reg [31:0] dummy_instr_seed_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15842.13-15842.31" */
reg [31:0] dummy_instr_seed_q_t0;
/* src = "generated/sv2v_out.v:15840.12-15840.24" */
wire [2:0] dummy_opcode;
/* src = "generated/sv2v_out.v:15839.12-15839.21" */
wire [6:0] dummy_set;
/* src = "generated/sv2v_out.v:15823.13-15823.26" */
input fetch_valid_i;
wire fetch_valid_i;
/* cellift = 32'd1 */
input fetch_valid_i_t0;
wire fetch_valid_i_t0;
/* src = "generated/sv2v_out.v:15824.13-15824.26" */
input id_in_ready_i;
wire id_in_ready_i;
/* cellift = 32'd1 */
input id_in_ready_i_t0;
wire id_in_ready_i_t0;
/* src = "generated/sv2v_out.v:15825.14-15825.34" */
output insert_dummy_instr_o;
wire insert_dummy_instr_o;
/* cellift = 32'd1 */
output insert_dummy_instr_o_t0;
wire insert_dummy_instr_o_t0;
/* src = "generated/sv2v_out.v:15830.14-15830.23" */
wire [16:0] lfsr_data;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15830.14-15830.23" */
/* unused_bits = "0 1 2 3 4 15 16" */
wire [16:0] lfsr_data_t0;
/* src = "generated/sv2v_out.v:15836.7-15836.14" */
wire lfsr_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15836.7-15836.14" */
wire lfsr_en_t0;
/* src = "generated/sv2v_out.v:15818.13-15818.19" */
input rst_ni;
wire rst_ni;
assign dummy_cnt_incr = dummy_cnt_q + /* src = "generated/sv2v_out.v:15872.26-15872.58" */ 5'h01;
assign lfsr_en = insert_dummy_instr_o & /* src = "generated/sv2v_out.v:15844.19-15844.53" */ id_in_ready_i;
assign dummy_cnt_threshold = lfsr_data[4:0] & /* src = "generated/sv2v_out.v:15871.31-15871.93" */ { dummy_instr_mask_i, 2'h3 };
assign _00_ = dummy_instr_en_i & /* src = "generated/sv2v_out.v:15874.25-15874.57" */ id_in_ready_i;
assign dummy_cnt_en = _00_ & /* src = "generated/sv2v_out.v:15874.24-15874.97" */ _12_;
assign insert_dummy_instr_o = dummy_instr_en_i & /* src = "generated/sv2v_out.v:15880.30-15880.85" */ _11_;
assign _01_ = ~ dummy_instr_seed_en_i;
assign _06_ = { dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i } & dummy_instr_seed_d_t0;
assign _07_ = { _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_ } & dummy_instr_seed_q_t0;
assign _09_ = _06_ | _07_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$501c60d7519704ee720c78ef16ad88cf05835059\ibex_dummy_instr  */
/* PC_TAINT_INFO STATE_NAME dummy_instr_seed_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_instr_seed_q_t0 <= 32'd0;
else dummy_instr_seed_q_t0 <= _09_;
assign _03_ = insert_dummy_instr_o_t0 & id_in_ready_i;
assign insert_dummy_instr_o_t0 = dummy_instr_en_i_t0 & _11_;
assign _04_ = id_in_ready_i_t0 & insert_dummy_instr_o;
assign _05_ = insert_dummy_instr_o_t0 & id_in_ready_i_t0;
assign _08_ = _03_ | _04_;
assign lfsr_en_t0 = _08_ | _05_;
/* src = "generated/sv2v_out.v:15875.2-15879.31" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$501c60d7519704ee720c78ef16ad88cf05835059\ibex_dummy_instr  */
/* PC_TAINT_INFO STATE_NAME dummy_cnt_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_cnt_q <= 5'h00;
else if (dummy_cnt_en) dummy_cnt_q <= dummy_cnt_d;
/* src = "generated/sv2v_out.v:15846.2-15850.45" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$501c60d7519704ee720c78ef16ad88cf05835059\ibex_dummy_instr  */
/* PC_TAINT_INFO STATE_NAME dummy_instr_seed_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_instr_seed_q <= 32'd0;
else if (dummy_instr_seed_en_i) dummy_instr_seed_q <= dummy_instr_seed_d;
assign _02_ = | { _15_, _13_ };
assign _10_ = _14_ ? 3'h4 : 3'h0;
assign dummy_opcode = _13_ ? 3'h7 : _10_;
assign dummy_set = _02_ ? 7'h00 : 7'h01;
assign dummy_instr_seed_d_t0 = dummy_instr_seed_q_t0 | dummy_instr_seed_i_t0;
assign _11_ = dummy_cnt_q == /* src = "generated/sv2v_out.v:15880.50-15880.84" */ dummy_cnt_threshold;
assign _12_ = fetch_valid_i | /* src = "generated/sv2v_out.v:15874.62-15874.96" */ insert_dummy_instr_o;
assign _13_ = lfsr_data[16:15] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15882.3-15903.10" */ 2'h3;
assign _14_ = lfsr_data[16:15] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15882.3-15903.10" */ 2'h2;
assign _15_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15882.3-15903.10" */ lfsr_data[16:15];
assign dummy_cnt_d = insert_dummy_instr_o ? /* src = "generated/sv2v_out.v:15873.24-15873.73" */ 5'h00 : dummy_cnt_incr;
assign dummy_instr_seed_d = dummy_instr_seed_q ^ /* src = "generated/sv2v_out.v:15845.30-15845.69" */ dummy_instr_seed_i;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:15857.4-15865.3" */
\$paramod$5fd3ce2f8a67228d339c5f62898ff83b3c2a14f0\prim_lfsr  lfsr_i (
.clk_i(clk_i),
.entropy_i(8'h00),
.entropy_i_t0(8'h00),
.lfsr_en_i(lfsr_en),
.lfsr_en_i_t0(lfsr_en_t0),
.rst_ni(rst_ni),
.seed_en_i(dummy_instr_seed_en_i),
.seed_en_i_t0(dummy_instr_seed_en_i_t0),
.seed_i(dummy_instr_seed_d),
.seed_i_t0(dummy_instr_seed_d_t0),
.state_o(lfsr_data),
.state_o_t0(lfsr_data_t0)
);
assign dummy_instr_data_o = { dummy_set, lfsr_data[14:5], dummy_opcode, 12'h033 };
assign dummy_instr_data_o_t0 = { 7'h00, lfsr_data_t0[14:5], 15'h0000 };
endmodule

module \$paramod$5714e31d82f2b8816750797f158ebea69a089104\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _0_;
wire [5:0] _1_;
wire [5:0] _2_;
wire [5:0] _3_;
/* src = "generated/sv2v_out.v:14894.13-14894.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14898.28-14898.37" */
output [5:0] rd_data_o;
reg [5:0] rd_data_o;
/* cellift = 32'd1 */
output [5:0] rd_data_o_t0;
reg [5:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14899.14-14899.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14895.13-14895.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14896.27-14896.36" */
input [5:0] wr_data_i;
wire [5:0] wr_data_i;
/* cellift = 32'd1 */
input [5:0] wr_data_i_t0;
wire [5:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14897.13-14897.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _0_ = ~ wr_en_i;
assign _1_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _2_ = { _0_, _0_, _0_, _0_, _0_, _0_ } & rd_data_o_t0;
assign _3_ = _1_ | _2_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$5714e31d82f2b8816750797f158ebea69a089104\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 6'h00;
else rd_data_o_t0 <= _3_;
/* src = "generated/sv2v_out.v:14901.2-14905.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$5714e31d82f2b8816750797f158ebea69a089104\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 6'h10;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$5c0dc9f9e0551018f7d8916b4fcabdef94a17390\ibex_core (clk_i, rst_ni, hart_id_i, boot_addr_i, instr_req_o, instr_gnt_i, instr_rvalid_i, instr_addr_o, instr_rdata_i, instr_err_i, data_req_o, data_gnt_i, data_rvalid_i, data_we_o, data_be_o, data_addr_o, data_wdata_o, data_rdata_i, data_err_i, dummy_instr_id_o, dummy_instr_wb_o
, rf_raddr_a_o, rf_raddr_b_o, rf_waddr_wb_o, rf_we_wb_o, rf_wdata_wb_ecc_o, rf_rdata_a_ecc_i, rf_rdata_b_ecc_i, ic_tag_req_o, ic_tag_write_o, ic_tag_addr_o, ic_tag_wdata_o, ic_tag_rdata_i, ic_data_req_o, ic_data_write_o, ic_data_addr_o, ic_data_wdata_o, ic_data_rdata_i, ic_scr_key_valid_i, ic_scr_key_req_o, irq_software_i, irq_timer_i
, irq_external_i, irq_fast_i, irq_nm_i, irq_pending_o, debug_req_i, crash_dump_o, double_fault_seen_o, fetch_enable_i, alert_minor_o, alert_major_internal_o, alert_major_bus_o, core_busy_o, instr_rvalid_i_t0, instr_req_o_t0, instr_rdata_i_t0, instr_gnt_i_t0, instr_err_i_t0, instr_addr_o_t0, rf_raddr_b_o_t0, rf_raddr_a_o_t0, data_we_o_t0
, data_req_o_t0, debug_req_i_t0, data_rdata_i_t0, data_gnt_i_t0, data_be_o_t0, data_addr_o_t0, data_rvalid_i_t0, data_wdata_o_t0, irq_nm_i_t0, ic_tag_write_o_t0, ic_tag_wdata_o_t0, ic_tag_req_o_t0, ic_tag_rdata_i_t0, ic_tag_addr_o_t0, ic_scr_key_valid_i_t0, ic_scr_key_req_o_t0, ic_data_write_o_t0, ic_data_wdata_o_t0, ic_data_req_o_t0, ic_data_rdata_i_t0, ic_data_addr_o_t0
, dummy_instr_id_o_t0, boot_addr_i_t0, dummy_instr_wb_o_t0, rf_waddr_wb_o_t0, rf_we_wb_o_t0, double_fault_seen_o_t0, hart_id_i_t0, irq_external_i_t0, irq_fast_i_t0, irq_pending_o_t0, irq_software_i_t0, irq_timer_i_t0, alert_major_bus_o_t0, alert_major_internal_o_t0, alert_minor_o_t0, core_busy_o_t0, crash_dump_o_t0, data_err_i_t0, fetch_enable_i_t0, rf_rdata_a_ecc_i_t0, rf_rdata_b_ecc_i_t0
, rf_wdata_wb_ecc_o_t0);
/* src = "generated/sv2v_out.v:13437.30-13437.54" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13437.30-13437.54" */
wire _001_;
/* src = "generated/sv2v_out.v:13438.30-13438.54" */
wire _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13438.30-13438.54" */
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
/* src = "generated/sv2v_out.v:13146.41-13146.56" */
wire _080_;
/* src = "generated/sv2v_out.v:13437.58-13437.75" */
wire _081_;
/* src = "generated/sv2v_out.v:13438.58-13438.75" */
wire _082_;
/* src = "generated/sv2v_out.v:13397.46-13397.90" */
wire _083_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13397.46-13397.90" */
wire _084_;
/* src = "generated/sv2v_out.v:13398.48-13398.94" */
wire _085_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13398.48-13398.94" */
wire _086_;
/* src = "generated/sv2v_out.v:13439.47-13439.80" */
wire _087_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13439.47-13439.80" */
wire _088_;
/* src = "generated/sv2v_out.v:13463.35-13463.70" */
wire _089_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13463.35-13463.70" */
wire _090_;
/* src = "generated/sv2v_out.v:13464.30-13464.78" */
wire _091_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13464.30-13464.78" */
wire _092_;
/* src = "generated/sv2v_out.v:13058.30-13058.81" */
wire _093_;
/* src = "generated/sv2v_out.v:13058.30-13058.81" */
wire _094_;
/* src = "generated/sv2v_out.v:13437.30-13437.43" */
wire _095_;
/* src = "generated/sv2v_out.v:13438.30-13438.43" */
wire _096_;
/* src = "generated/sv2v_out.v:12874.14-12874.31" */
output alert_major_bus_o;
wire alert_major_bus_o;
/* cellift = 32'd1 */
output alert_major_bus_o_t0;
wire alert_major_bus_o_t0;
/* src = "generated/sv2v_out.v:12873.14-12873.36" */
output alert_major_internal_o;
wire alert_major_internal_o;
/* cellift = 32'd1 */
output alert_major_internal_o_t0;
wire alert_major_internal_o_t0;
/* src = "generated/sv2v_out.v:12872.14-12872.27" */
output alert_minor_o;
wire alert_minor_o;
/* cellift = 32'd1 */
output alert_minor_o_t0;
wire alert_minor_o_t0;
/* src = "generated/sv2v_out.v:12955.14-12955.33" */
wire [31:0] alu_adder_result_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12955.14-12955.33" */
wire [31:0] alu_adder_result_ex_t0;
/* src = "generated/sv2v_out.v:12951.14-12951.30" */
wire [31:0] alu_operand_a_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12951.14-12951.30" */
wire [31:0] alu_operand_a_ex_t0;
/* src = "generated/sv2v_out.v:12952.14-12952.30" */
wire [31:0] alu_operand_b_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12952.14-12952.30" */
wire [31:0] alu_operand_b_ex_t0;
/* src = "generated/sv2v_out.v:12950.13-12950.28" */
wire [6:0] alu_operator_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12950.13-12950.28" */
wire [6:0] alu_operator_ex_t0;
/* src = "generated/sv2v_out.v:12825.20-12825.31" */
input [31:0] boot_addr_i;
wire [31:0] boot_addr_i;
/* cellift = 32'd1 */
input [31:0] boot_addr_i_t0;
wire [31:0] boot_addr_i_t0;
/* src = "generated/sv2v_out.v:12928.7-12928.22" */
wire branch_decision;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12928.7-12928.22" */
wire branch_decision_t0;
/* src = "generated/sv2v_out.v:12927.14-12927.30" */
wire [31:0] branch_target_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12927.14-12927.30" */
wire [31:0] branch_target_ex_t0;
/* src = "generated/sv2v_out.v:12953.14-12953.26" */
wire [31:0] bt_a_operand;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12953.14-12953.26" */
wire [31:0] bt_a_operand_t0;
/* src = "generated/sv2v_out.v:12954.14-12954.26" */
wire [31:0] bt_b_operand;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12954.14-12954.26" */
wire [31:0] bt_b_operand_t0;
/* src = "generated/sv2v_out.v:12822.13-12822.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:12875.20-12875.31" */
output [3:0] core_busy_o;
wire [3:0] core_busy_o;
/* cellift = 32'd1 */
output [3:0] core_busy_o_t0;
wire [3:0] core_busy_o_t0;
/* src = "generated/sv2v_out.v:13456.14-13456.30" */
wire [31:0] crash_dump_mtval;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13456.14-13456.30" */
wire [31:0] crash_dump_mtval_t0;
/* src = "generated/sv2v_out.v:12869.22-12869.34" */
output [159:0] crash_dump_o;
wire [159:0] crash_dump_o;
/* cellift = 32'd1 */
output [159:0] crash_dump_o_t0;
wire [159:0] crash_dump_o_t0;
/* src = "generated/sv2v_out.v:12966.7-12966.17" */
wire csr_access;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12966.7-12966.17" */
wire csr_access_t0;
/* src = "generated/sv2v_out.v:12969.14-12969.22" */
wire [11:0] csr_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12969.14-12969.22" */
wire [11:0] csr_addr_t0;
/* src = "generated/sv2v_out.v:12998.14-12998.22" */
wire [31:0] csr_depc;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12998.14-12998.22" */
wire [31:0] csr_depc_t0;
/* src = "generated/sv2v_out.v:12997.14-12997.22" */
wire [31:0] csr_mepc;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12997.14-12997.22" */
wire [31:0] csr_mepc_t0;
/* src = "generated/sv2v_out.v:12996.7-12996.22" */
wire csr_mstatus_mie;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12996.7-12996.22" */
wire csr_mstatus_mie_t0;
/* src = "generated/sv2v_out.v:13013.7-13013.21" */
wire csr_mstatus_tw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13013.7-13013.21" */
wire csr_mstatus_tw_t0;
/* src = "generated/sv2v_out.v:13012.14-13012.23" */
wire [31:0] csr_mtval;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13012.14-13012.23" */
wire [31:0] csr_mtval_t0;
/* src = "generated/sv2v_out.v:13011.14-13011.23" */
wire [31:0] csr_mtvec;
/* src = "generated/sv2v_out.v:13010.7-13010.21" */
wire csr_mtvec_init;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13010.7-13010.21" */
wire csr_mtvec_init_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13011.14-13011.23" */
wire [31:0] csr_mtvec_t0;
/* src = "generated/sv2v_out.v:12967.13-12967.19" */
wire [1:0] csr_op;
/* src = "generated/sv2v_out.v:12968.7-12968.16" */
wire csr_op_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12968.7-12968.16" */
wire csr_op_en_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12967.13-12967.19" */
wire [1:0] csr_op_t0;
/* src = "generated/sv2v_out.v:12999.36-12999.48" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135" */
wire [135:0] csr_pmp_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12999.36-12999.48" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135" */
wire [135:0] csr_pmp_addr_t0;
/* src = "generated/sv2v_out.v:13000.35-13000.46" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23" */
wire [23:0] csr_pmp_cfg;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13000.35-13000.46" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23" */
wire [23:0] csr_pmp_cfg_t0;
/* src = "generated/sv2v_out.v:13001.13-13001.28" */
/* unused_bits = "0 1 2" */
wire [2:0] csr_pmp_mseccfg;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13001.13-13001.28" */
/* unused_bits = "0 1 2" */
wire [2:0] csr_pmp_mseccfg_t0;
/* src = "generated/sv2v_out.v:12970.14-12970.23" */
wire [31:0] csr_rdata;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12970.14-12970.23" */
wire [31:0] csr_rdata_t0;
/* src = "generated/sv2v_out.v:13008.7-13008.26" */
wire csr_restore_dret_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13008.7-13008.26" */
wire csr_restore_dret_id_t0;
/* src = "generated/sv2v_out.v:13007.7-13007.26" */
wire csr_restore_mret_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13007.7-13007.26" */
wire csr_restore_mret_id_t0;
/* src = "generated/sv2v_out.v:13009.7-13009.21" */
wire csr_save_cause;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13009.7-13009.21" */
wire csr_save_cause_t0;
/* src = "generated/sv2v_out.v:13005.7-13005.18" */
wire csr_save_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13005.7-13005.18" */
wire csr_save_id_t0;
/* src = "generated/sv2v_out.v:13004.7-13004.18" */
wire csr_save_if;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13004.7-13004.18" */
wire csr_save_if_t0;
/* src = "generated/sv2v_out.v:13006.7-13006.18" */
wire csr_save_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13006.7-13006.18" */
wire csr_save_wb_t0;
/* src = "generated/sv2v_out.v:12907.7-12907.21" */
wire csr_shadow_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12907.7-12907.21" */
wire csr_shadow_err_t0;
/* src = "generated/sv2v_out.v:12929.7-12929.16" */
wire ctrl_busy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12929.7-12929.16" */
wire ctrl_busy_t0;
/* src = "generated/sv2v_out.v:12837.21-12837.32" */
output [31:0] data_addr_o;
wire [31:0] data_addr_o;
/* cellift = 32'd1 */
output [31:0] data_addr_o_t0;
wire [31:0] data_addr_o_t0;
/* src = "generated/sv2v_out.v:12836.20-12836.29" */
output [3:0] data_be_o;
wire [3:0] data_be_o;
/* cellift = 32'd1 */
output [3:0] data_be_o_t0;
wire [3:0] data_be_o_t0;
/* src = "generated/sv2v_out.v:12840.13-12840.23" */
input data_err_i;
wire data_err_i;
/* cellift = 32'd1 */
input data_err_i_t0;
wire data_err_i_t0;
/* src = "generated/sv2v_out.v:12833.13-12833.23" */
input data_gnt_i;
wire data_gnt_i;
/* cellift = 32'd1 */
input data_gnt_i_t0;
wire data_gnt_i_t0;
/* src = "generated/sv2v_out.v:12898.7-12898.22" */
wire data_ind_timing;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12898.7-12898.22" */
wire data_ind_timing_t0;
/* src = "generated/sv2v_out.v:12839.34-12839.46" */
input [38:0] data_rdata_i;
wire [38:0] data_rdata_i;
/* cellift = 32'd1 */
input [38:0] data_rdata_i_t0;
wire [38:0] data_rdata_i_t0;
/* src = "generated/sv2v_out.v:12832.14-12832.24" */
output data_req_o;
wire data_req_o;
/* cellift = 32'd1 */
output data_req_o_t0;
wire data_req_o_t0;
/* src = "generated/sv2v_out.v:12834.13-12834.26" */
input data_rvalid_i;
wire data_rvalid_i;
/* cellift = 32'd1 */
input data_rvalid_i_t0;
wire data_rvalid_i_t0;
/* src = "generated/sv2v_out.v:12838.35-12838.47" */
output [38:0] data_wdata_o;
wire [38:0] data_wdata_o;
/* cellift = 32'd1 */
output [38:0] data_wdata_o_t0;
wire [38:0] data_wdata_o_t0;
/* src = "generated/sv2v_out.v:12835.14-12835.23" */
output data_we_o;
wire data_we_o;
/* cellift = 32'd1 */
output data_we_o_t0;
wire data_we_o_t0;
/* src = "generated/sv2v_out.v:13018.13-13018.24" */
wire [2:0] debug_cause;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13018.13-13018.24" */
wire [2:0] debug_cause_t0;
/* src = "generated/sv2v_out.v:13019.7-13019.21" */
wire debug_csr_save;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13019.7-13019.21" */
wire debug_csr_save_t0;
/* src = "generated/sv2v_out.v:13021.7-13021.20" */
wire debug_ebreakm;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13021.7-13021.20" */
wire debug_ebreakm_t0;
/* src = "generated/sv2v_out.v:13022.7-13022.20" */
wire debug_ebreaku;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13022.7-13022.20" */
wire debug_ebreaku_t0;
/* src = "generated/sv2v_out.v:13016.7-13016.17" */
wire debug_mode;
/* src = "generated/sv2v_out.v:13017.7-13017.26" */
wire debug_mode_entering;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13017.7-13017.26" */
wire debug_mode_entering_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13016.7-13016.17" */
wire debug_mode_t0;
/* src = "generated/sv2v_out.v:12868.13-12868.24" */
input debug_req_i;
wire debug_req_i;
/* cellift = 32'd1 */
input debug_req_i_t0;
wire debug_req_i_t0;
/* src = "generated/sv2v_out.v:13020.7-13020.24" */
wire debug_single_step;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13020.7-13020.24" */
wire debug_single_step_t0;
/* src = "generated/sv2v_out.v:12958.7-12958.16" */
wire div_en_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12958.7-12958.16" */
wire div_en_ex_t0;
/* src = "generated/sv2v_out.v:12960.7-12960.17" */
wire div_sel_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12960.7-12960.17" */
wire div_sel_ex_t0;
/* src = "generated/sv2v_out.v:12870.14-12870.33" */
output double_fault_seen_o;
wire double_fault_seen_o;
/* cellift = 32'd1 */
output double_fault_seen_o_t0;
wire double_fault_seen_o_t0;
/* src = "generated/sv2v_out.v:12899.7-12899.21" */
wire dummy_instr_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12899.7-12899.21" */
wire dummy_instr_en_t0;
/* src = "generated/sv2v_out.v:12841.14-12841.30" */
output dummy_instr_id_o;
wire dummy_instr_id_o;
/* cellift = 32'd1 */
output dummy_instr_id_o_t0;
wire dummy_instr_id_o_t0;
/* src = "generated/sv2v_out.v:12900.13-12900.29" */
wire [2:0] dummy_instr_mask;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12900.13-12900.29" */
wire [2:0] dummy_instr_mask_t0;
/* src = "generated/sv2v_out.v:12902.14-12902.30" */
wire [31:0] dummy_instr_seed;
/* src = "generated/sv2v_out.v:12901.7-12901.26" */
wire dummy_instr_seed_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12901.7-12901.26" */
wire dummy_instr_seed_en_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12902.14-12902.30" */
wire [31:0] dummy_instr_seed_t0;
/* src = "generated/sv2v_out.v:12842.14-12842.30" */
output dummy_instr_wb_o;
wire dummy_instr_wb_o;
/* cellift = 32'd1 */
output dummy_instr_wb_o_t0;
wire dummy_instr_wb_o_t0;
/* src = "generated/sv2v_out.v:12987.7-12987.12" */
wire en_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12987.7-12987.12" */
wire en_wb_t0;
/* src = "generated/sv2v_out.v:12981.7-12981.15" */
wire ex_valid;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12981.7-12981.15" */
wire ex_valid_t0;
/* src = "generated/sv2v_out.v:12915.13-12915.22" */
wire [6:0] exc_cause;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12915.13-12915.22" */
wire [6:0] exc_cause_t0;
/* src = "generated/sv2v_out.v:12914.13-12914.26" */
wire [1:0] exc_pc_mux_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12914.13-12914.26" */
wire [1:0] exc_pc_mux_id_t0;
/* src = "generated/sv2v_out.v:12923.7-12923.29" */
wire expecting_load_resp_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12923.7-12923.29" */
wire expecting_load_resp_id_t0;
/* src = "generated/sv2v_out.v:12924.7-12924.30" */
wire expecting_store_resp_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12924.7-12924.30" */
wire expecting_store_resp_id_t0;
/* src = "generated/sv2v_out.v:12871.19-12871.33" */
input [3:0] fetch_enable_i;
wire [3:0] fetch_enable_i;
/* cellift = 32'd1 */
input [3:0] fetch_enable_i_t0;
wire [3:0] fetch_enable_i_t0;
/* src = "generated/sv2v_out.v:13047.16-13047.29" */
wire [11:0] \g_core_busy_secure.busy_bits_buf ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13047.16-13047.29" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11" */
wire [11:0] \g_core_busy_secure.busy_bits_buf_t0 ;
/* src = "generated/sv2v_out.v:13590.15-13590.33" */
/* unused_bits = "0 1" */
wire [1:0] \g_no_pmp.unused_priv_lvl_ls ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13590.15-13590.33" */
/* unused_bits = "0 1" */
wire [1:0] \g_no_pmp.unused_priv_lvl_ls_t0 ;
/* src = "generated/sv2v_out.v:13419.15-13419.27" */
wire [1:0] \gen_regfile_ecc.rf_ecc_err_a ;
/* src = "generated/sv2v_out.v:13421.9-13421.24" */
wire \gen_regfile_ecc.rf_ecc_err_a_id ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13421.9-13421.24" */
wire \gen_regfile_ecc.rf_ecc_err_a_id_t0 ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13419.15-13419.27" */
/* unused_bits = "0 1" */
wire [1:0] \gen_regfile_ecc.rf_ecc_err_a_t0 ;
/* src = "generated/sv2v_out.v:13420.15-13420.27" */
wire [1:0] \gen_regfile_ecc.rf_ecc_err_b ;
/* src = "generated/sv2v_out.v:13422.9-13422.24" */
wire \gen_regfile_ecc.rf_ecc_err_b_id ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13422.9-13422.24" */
wire \gen_regfile_ecc.rf_ecc_err_b_id_t0 ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13420.15-13420.27" */
/* unused_bits = "0 1" */
wire [1:0] \gen_regfile_ecc.rf_ecc_err_b_t0 ;
/* src = "generated/sv2v_out.v:12824.20-12824.29" */
input [31:0] hart_id_i;
wire [31:0] hart_id_i;
/* cellift = 32'd1 */
input [31:0] hart_id_i_t0;
wire [31:0] hart_id_i_t0;
/* src = "generated/sv2v_out.v:12857.42-12857.56" */
output [7:0] ic_data_addr_o;
wire [7:0] ic_data_addr_o;
/* cellift = 32'd1 */
output [7:0] ic_data_addr_o_t0;
wire [7:0] ic_data_addr_o_t0;
/* src = "generated/sv2v_out.v:12859.58-12859.73" */
input [127:0] ic_data_rdata_i;
wire [127:0] ic_data_rdata_i;
/* cellift = 32'd1 */
input [127:0] ic_data_rdata_i_t0;
wire [127:0] ic_data_rdata_i_t0;
/* src = "generated/sv2v_out.v:12855.20-12855.33" */
output [1:0] ic_data_req_o;
wire [1:0] ic_data_req_o;
/* cellift = 32'd1 */
output [1:0] ic_data_req_o_t0;
wire [1:0] ic_data_req_o_t0;
/* src = "generated/sv2v_out.v:12858.34-12858.49" */
output [63:0] ic_data_wdata_o;
wire [63:0] ic_data_wdata_o;
/* cellift = 32'd1 */
output [63:0] ic_data_wdata_o_t0;
wire [63:0] ic_data_wdata_o_t0;
/* src = "generated/sv2v_out.v:12856.14-12856.29" */
output ic_data_write_o;
wire ic_data_write_o;
/* cellift = 32'd1 */
output ic_data_write_o_t0;
wire ic_data_write_o_t0;
/* src = "generated/sv2v_out.v:12861.14-12861.30" */
output ic_scr_key_req_o;
wire ic_scr_key_req_o;
/* cellift = 32'd1 */
output ic_scr_key_req_o_t0;
wire ic_scr_key_req_o_t0;
/* src = "generated/sv2v_out.v:12860.13-12860.31" */
input ic_scr_key_valid_i;
wire ic_scr_key_valid_i;
/* cellift = 32'd1 */
input ic_scr_key_valid_i_t0;
wire ic_scr_key_valid_i_t0;
/* src = "generated/sv2v_out.v:12852.42-12852.55" */
output [7:0] ic_tag_addr_o;
wire [7:0] ic_tag_addr_o;
/* cellift = 32'd1 */
output [7:0] ic_tag_addr_o_t0;
wire [7:0] ic_tag_addr_o_t0;
/* src = "generated/sv2v_out.v:12854.57-12854.71" */
input [43:0] ic_tag_rdata_i;
wire [43:0] ic_tag_rdata_i;
/* cellift = 32'd1 */
input [43:0] ic_tag_rdata_i_t0;
wire [43:0] ic_tag_rdata_i_t0;
/* src = "generated/sv2v_out.v:12850.20-12850.32" */
output [1:0] ic_tag_req_o;
wire [1:0] ic_tag_req_o;
/* cellift = 32'd1 */
output [1:0] ic_tag_req_o_t0;
wire [1:0] ic_tag_req_o_t0;
/* src = "generated/sv2v_out.v:12853.33-12853.47" */
output [21:0] ic_tag_wdata_o;
wire [21:0] ic_tag_wdata_o;
/* cellift = 32'd1 */
output [21:0] ic_tag_wdata_o_t0;
wire [21:0] ic_tag_wdata_o_t0;
/* src = "generated/sv2v_out.v:12851.14-12851.28" */
output ic_tag_write_o;
wire ic_tag_write_o;
/* cellift = 32'd1 */
output ic_tag_write_o_t0;
wire ic_tag_write_o_t0;
/* src = "generated/sv2v_out.v:12903.7-12903.20" */
wire icache_enable;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12903.7-12903.20" */
wire icache_enable_t0;
/* src = "generated/sv2v_out.v:12904.7-12904.19" */
wire icache_inval;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12904.7-12904.19" */
wire icache_inval_t0;
/* src = "generated/sv2v_out.v:12980.7-12980.18" */
wire id_in_ready;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12980.7-12980.18" */
wire id_in_ready_t0;
/* src = "generated/sv2v_out.v:12930.7-12930.14" */
wire if_busy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12930.7-12930.14" */
wire if_busy_t0;
/* src = "generated/sv2v_out.v:12891.7-12891.24" */
wire illegal_c_insn_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12891.7-12891.24" */
wire illegal_c_insn_id_t0;
/* src = "generated/sv2v_out.v:12972.7-12972.26" */
wire illegal_csr_insn_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12972.7-12972.26" */
wire illegal_csr_insn_id_t0;
/* src = "generated/sv2v_out.v:13039.7-13039.22" */
/* unused_bits = "0" */
wire illegal_insn_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13039.7-13039.22" */
/* unused_bits = "0" */
wire illegal_insn_id_t0;
/* src = "generated/sv2v_out.v:12895.14-12895.26" */
wire [67:0] imd_val_d_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12895.14-12895.26" */
wire [67:0] imd_val_d_ex_t0;
/* src = "generated/sv2v_out.v:12896.14-12896.26" */
wire [67:0] imd_val_q_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12896.14-12896.26" */
wire [67:0] imd_val_q_ex_t0;
/* src = "generated/sv2v_out.v:12897.13-12897.26" */
wire [1:0] imd_val_we_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12897.13-12897.26" */
wire [1:0] imd_val_we_ex_t0;
/* src = "generated/sv2v_out.v:12829.21-12829.33" */
output [31:0] instr_addr_o;
wire [31:0] instr_addr_o;
/* cellift = 32'd1 */
output [31:0] instr_addr_o_t0;
wire [31:0] instr_addr_o_t0;
/* src = "generated/sv2v_out.v:12888.7-12888.24" */
wire instr_bp_taken_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12888.7-12888.24" */
wire instr_bp_taken_id_t0;
/* src = "generated/sv2v_out.v:13025.7-13025.20" */
/* unused_bits = "0" */
wire instr_done_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13025.7-13025.20" */
/* unused_bits = "0" */
wire instr_done_wb_t0;
/* src = "generated/sv2v_out.v:12831.13-12831.24" */
input instr_err_i;
wire instr_err_i;
/* cellift = 32'd1 */
input instr_err_i_t0;
wire instr_err_i_t0;
/* src = "generated/sv2v_out.v:12986.7-12986.17" */
wire instr_exec;
/* src = "generated/sv2v_out.v:12889.7-12889.22" */
wire instr_fetch_err;
/* src = "generated/sv2v_out.v:12890.7-12890.28" */
wire instr_fetch_err_plus2;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12890.7-12890.28" */
wire instr_fetch_err_plus2_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12889.7-12889.22" */
wire instr_fetch_err_t0;
/* src = "generated/sv2v_out.v:12908.7-12908.27" */
wire instr_first_cycle_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12908.7-12908.27" */
wire instr_first_cycle_id_t0;
/* src = "generated/sv2v_out.v:12827.13-12827.24" */
input instr_gnt_i;
wire instr_gnt_i;
/* cellift = 32'd1 */
input instr_gnt_i_t0;
wire instr_gnt_i_t0;
/* src = "generated/sv2v_out.v:13024.7-13024.20" */
/* unused_bits = "0" */
wire instr_id_done;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13024.7-13024.20" */
/* unused_bits = "0" */
wire instr_id_done_t0;
/* src = "generated/sv2v_out.v:12916.7-12916.21" */
wire instr_intg_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12916.7-12916.21" */
wire instr_intg_err_t0;
/* src = "generated/sv2v_out.v:12886.7-12886.29" */
wire instr_is_compressed_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12886.7-12886.29" */
wire instr_is_compressed_id_t0;
/* src = "generated/sv2v_out.v:12882.7-12882.19" */
/* unused_bits = "0" */
wire instr_new_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12882.7-12882.19" */
/* unused_bits = "0" */
wire instr_new_id_t0;
/* src = "generated/sv2v_out.v:12887.7-12887.26" */
wire instr_perf_count_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12887.7-12887.26" */
wire instr_perf_count_id_t0;
/* src = "generated/sv2v_out.v:12884.14-12884.32" */
wire [31:0] instr_rdata_alu_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12884.14-12884.32" */
wire [31:0] instr_rdata_alu_id_t0;
/* src = "generated/sv2v_out.v:12885.14-12885.30" */
wire [15:0] instr_rdata_c_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12885.14-12885.30" */
wire [15:0] instr_rdata_c_id_t0;
/* src = "generated/sv2v_out.v:12830.34-12830.47" */
input [38:0] instr_rdata_i;
wire [38:0] instr_rdata_i;
/* cellift = 32'd1 */
input [38:0] instr_rdata_i_t0;
wire [38:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:12883.14-12883.28" */
wire [31:0] instr_rdata_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12883.14-12883.28" */
wire [31:0] instr_rdata_id_t0;
/* src = "generated/sv2v_out.v:12985.7-12985.22" */
wire instr_req_gated;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12985.7-12985.22" */
wire instr_req_gated_t0;
/* src = "generated/sv2v_out.v:12984.7-12984.20" */
wire instr_req_int;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12984.7-12984.20" */
wire instr_req_int_t0;
/* src = "generated/sv2v_out.v:12826.14-12826.25" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:12828.13-12828.27" */
input instr_rvalid_i;
wire instr_rvalid_i;
/* cellift = 32'd1 */
input instr_rvalid_i_t0;
wire instr_rvalid_i_t0;
/* src = "generated/sv2v_out.v:12988.13-12988.26" */
wire [1:0] instr_type_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12988.13-12988.26" */
wire [1:0] instr_type_wb_t0;
/* src = "generated/sv2v_out.v:12909.7-12909.24" */
wire instr_valid_clear;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12909.7-12909.24" */
wire instr_valid_clear_t0;
/* src = "generated/sv2v_out.v:12881.7-12881.21" */
wire instr_valid_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12881.7-12881.21" */
wire instr_valid_id_t0;
/* src = "generated/sv2v_out.v:12864.13-12864.27" */
input irq_external_i;
wire irq_external_i;
/* cellift = 32'd1 */
input irq_external_i_t0;
wire irq_external_i_t0;
/* src = "generated/sv2v_out.v:12865.20-12865.30" */
input [14:0] irq_fast_i;
wire [14:0] irq_fast_i;
/* cellift = 32'd1 */
input [14:0] irq_fast_i_t0;
wire [14:0] irq_fast_i_t0;
/* src = "generated/sv2v_out.v:12866.13-12866.21" */
input irq_nm_i;
wire irq_nm_i;
/* cellift = 32'd1 */
input irq_nm_i_t0;
wire irq_nm_i_t0;
/* src = "generated/sv2v_out.v:12867.14-12867.27" */
output irq_pending_o;
wire irq_pending_o;
/* cellift = 32'd1 */
output irq_pending_o_t0;
wire irq_pending_o_t0;
/* src = "generated/sv2v_out.v:12862.13-12862.27" */
input irq_software_i;
wire irq_software_i;
/* cellift = 32'd1 */
input irq_software_i_t0;
wire irq_software_i_t0;
/* src = "generated/sv2v_out.v:12863.13-12863.24" */
input irq_timer_i;
wire irq_timer_i;
/* cellift = 32'd1 */
input irq_timer_i_t0;
wire irq_timer_i_t0;
/* src = "generated/sv2v_out.v:12995.14-12995.18" */
wire [17:0] irqs;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12995.14-12995.18" */
wire [17:0] irqs_t0;
/* src = "generated/sv2v_out.v:12925.7-12925.24" */
wire lsu_addr_incr_req;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12925.7-12925.24" */
wire lsu_addr_incr_req_t0;
/* src = "generated/sv2v_out.v:12926.14-12926.27" */
wire [31:0] lsu_addr_last;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12926.14-12926.27" */
wire [31:0] lsu_addr_last_t0;
/* src = "generated/sv2v_out.v:12931.7-12931.15" */
wire lsu_busy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12931.7-12931.15" */
wire lsu_busy_t0;
/* src = "generated/sv2v_out.v:12917.7-12917.19" */
wire lsu_load_err;
/* src = "generated/sv2v_out.v:12918.7-12918.23" */
wire lsu_load_err_raw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12918.7-12918.23" */
wire lsu_load_err_raw_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12917.7-12917.19" */
wire lsu_load_err_t0;
/* src = "generated/sv2v_out.v:12921.7-12921.29" */
wire lsu_load_resp_intg_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12921.7-12921.29" */
wire lsu_load_resp_intg_err_t0;
/* src = "generated/sv2v_out.v:12977.7-12977.22" */
wire lsu_rdata_valid;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12977.7-12977.22" */
wire lsu_rdata_valid_t0;
/* src = "generated/sv2v_out.v:12976.7-12976.14" */
wire lsu_req;
/* src = "generated/sv2v_out.v:12979.7-12979.19" */
wire lsu_req_done;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12979.7-12979.19" */
wire lsu_req_done_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12976.7-12976.14" */
wire lsu_req_t0;
/* src = "generated/sv2v_out.v:12983.7-12983.19" */
wire lsu_resp_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12983.7-12983.19" */
wire lsu_resp_err_t0;
/* src = "generated/sv2v_out.v:12982.7-12982.21" */
wire lsu_resp_valid;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12982.7-12982.21" */
wire lsu_resp_valid_t0;
/* src = "generated/sv2v_out.v:12975.7-12975.19" */
wire lsu_sign_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12975.7-12975.19" */
wire lsu_sign_ext_t0;
/* src = "generated/sv2v_out.v:12919.7-12919.20" */
wire lsu_store_err;
/* src = "generated/sv2v_out.v:12920.7-12920.24" */
wire lsu_store_err_raw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12920.7-12920.24" */
wire lsu_store_err_raw_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12919.7-12919.20" */
wire lsu_store_err_t0;
/* src = "generated/sv2v_out.v:12922.7-12922.30" */
wire lsu_store_resp_intg_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12922.7-12922.30" */
wire lsu_store_resp_intg_err_t0;
/* src = "generated/sv2v_out.v:12974.13-12974.21" */
wire [1:0] lsu_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12974.13-12974.21" */
wire [1:0] lsu_type_t0;
/* src = "generated/sv2v_out.v:12978.14-12978.23" */
wire [31:0] lsu_wdata;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12978.14-12978.23" */
wire [31:0] lsu_wdata_t0;
/* src = "generated/sv2v_out.v:12973.7-12973.13" */
wire lsu_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12973.7-12973.13" */
wire lsu_we_t0;
/* src = "generated/sv2v_out.v:12957.7-12957.17" */
wire mult_en_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12957.7-12957.17" */
wire mult_en_ex_t0;
/* src = "generated/sv2v_out.v:12959.7-12959.18" */
wire mult_sel_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12959.7-12959.18" */
wire mult_sel_ex_t0;
/* src = "generated/sv2v_out.v:12963.14-12963.34" */
wire [31:0] multdiv_operand_a_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12963.14-12963.34" */
wire [31:0] multdiv_operand_a_ex_t0;
/* src = "generated/sv2v_out.v:12964.14-12964.34" */
wire [31:0] multdiv_operand_b_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12964.14-12964.34" */
wire [31:0] multdiv_operand_b_ex_t0;
/* src = "generated/sv2v_out.v:12961.13-12961.32" */
wire [1:0] multdiv_operator_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12961.13-12961.32" */
wire [1:0] multdiv_operator_ex_t0;
/* src = "generated/sv2v_out.v:12965.7-12965.23" */
wire multdiv_ready_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12965.7-12965.23" */
wire multdiv_ready_id_t0;
/* src = "generated/sv2v_out.v:12962.13-12962.35" */
wire [1:0] multdiv_signed_mode_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12962.13-12962.35" */
wire [1:0] multdiv_signed_mode_ex_t0;
/* src = "generated/sv2v_out.v:12994.7-12994.15" */
wire nmi_mode;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12994.7-12994.15" */
wire nmi_mode_t0;
/* src = "generated/sv2v_out.v:12912.14-12912.28" */
wire [31:0] nt_branch_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12912.14-12912.28" */
wire [31:0] nt_branch_addr_t0;
/* src = "generated/sv2v_out.v:12911.7-12911.27" */
wire nt_branch_mispredict;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12911.7-12911.27" */
wire nt_branch_mispredict_t0;
/* src = "generated/sv2v_out.v:12991.7-12991.26" */
wire outstanding_load_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12991.7-12991.26" */
wire outstanding_load_wb_t0;
/* src = "generated/sv2v_out.v:12992.7-12992.27" */
wire outstanding_store_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12992.7-12992.27" */
wire outstanding_store_wb_t0;
/* src = "generated/sv2v_out.v:12893.14-12893.19" */
wire [31:0] pc_id /* verilator public */;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12893.14-12893.19" */
wire [31:0] pc_id_t0 /* verilator public */;
/* src = "generated/sv2v_out.v:12892.14-12892.19" */
wire [31:0] pc_if;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12892.14-12892.19" */
wire [31:0] pc_if_t0;
/* src = "generated/sv2v_out.v:12906.7-12906.24" */
wire pc_mismatch_alert;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12906.7-12906.24" */
wire pc_mismatch_alert_t0;
/* src = "generated/sv2v_out.v:12913.13-12913.22" */
wire [2:0] pc_mux_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12913.13-12913.22" */
wire [2:0] pc_mux_id_t0;
/* src = "generated/sv2v_out.v:12910.7-12910.13" */
wire pc_set;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12910.7-12910.13" */
wire pc_set_t0;
/* src = "generated/sv2v_out.v:12894.14-12894.19" */
wire [31:0] pc_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12894.14-12894.19" */
wire [31:0] pc_wb_t0;
/* src = "generated/sv2v_out.v:13035.7-13035.18" */
wire perf_branch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13035.7-13035.18" */
wire perf_branch_t0;
/* src = "generated/sv2v_out.v:13033.7-13033.20" */
wire perf_div_wait;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13033.7-13033.20" */
wire perf_div_wait_t0;
/* src = "generated/sv2v_out.v:13031.7-13031.22" */
wire perf_dside_wait;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13031.7-13031.22" */
wire perf_dside_wait_t0;
/* src = "generated/sv2v_out.v:13027.7-13027.35" */
wire perf_instr_ret_compressed_wb;
/* src = "generated/sv2v_out.v:13029.7-13029.40" */
wire perf_instr_ret_compressed_wb_spec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13029.7-13029.40" */
wire perf_instr_ret_compressed_wb_spec_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13027.7-13027.35" */
wire perf_instr_ret_compressed_wb_t0;
/* src = "generated/sv2v_out.v:13026.7-13026.24" */
wire perf_instr_ret_wb;
/* src = "generated/sv2v_out.v:13028.7-13028.29" */
wire perf_instr_ret_wb_spec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13028.7-13028.29" */
wire perf_instr_ret_wb_spec_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13026.7-13026.24" */
wire perf_instr_ret_wb_t0;
/* src = "generated/sv2v_out.v:13030.7-13030.22" */
wire perf_iside_wait;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13030.7-13030.22" */
wire perf_iside_wait_t0;
/* src = "generated/sv2v_out.v:13034.7-13034.16" */
wire perf_jump;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13034.7-13034.16" */
wire perf_jump_t0;
/* src = "generated/sv2v_out.v:13037.7-13037.16" */
wire perf_load;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13037.7-13037.16" */
wire perf_load_t0;
/* src = "generated/sv2v_out.v:13032.7-13032.20" */
wire perf_mul_wait;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13032.7-13032.20" */
wire perf_mul_wait_t0;
/* src = "generated/sv2v_out.v:13038.7-13038.17" */
wire perf_store;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13038.7-13038.17" */
wire perf_store_t0;
/* src = "generated/sv2v_out.v:13036.7-13036.19" */
wire perf_tbranch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13036.7-13036.19" */
wire perf_tbranch_t0;
/* src = "generated/sv2v_out.v:13014.13-13014.25" */
wire [1:0] priv_mode_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13014.13-13014.25" */
wire [1:0] priv_mode_id_t0;
/* src = "generated/sv2v_out.v:12989.7-12989.15" */
wire ready_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12989.7-12989.15" */
wire ready_wb_t0;
/* src = "generated/sv2v_out.v:12956.14-12956.23" */
wire [31:0] result_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12956.14-12956.23" */
wire [31:0] result_ex_t0;
/* src = "generated/sv2v_out.v:12944.7-12944.22" */
wire rf_ecc_err_comb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12944.7-12944.22" */
wire rf_ecc_err_comb_t0;
/* src = "generated/sv2v_out.v:12843.20-12843.32" */
output [4:0] rf_raddr_a_o;
wire [4:0] rf_raddr_a_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_a_o_t0;
wire [4:0] rf_raddr_a_o_t0;
/* src = "generated/sv2v_out.v:12844.20-12844.32" */
output [4:0] rf_raddr_b_o;
wire [4:0] rf_raddr_b_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_b_o_t0;
wire [4:0] rf_raddr_b_o_t0;
/* src = "generated/sv2v_out.v:12948.7-12948.23" */
wire rf_rd_a_wb_match;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12948.7-12948.23" */
wire rf_rd_a_wb_match_t0;
/* src = "generated/sv2v_out.v:12949.7-12949.23" */
wire rf_rd_b_wb_match;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12949.7-12949.23" */
wire rf_rd_b_wb_match_t0;
/* src = "generated/sv2v_out.v:12848.38-12848.54" */
input [38:0] rf_rdata_a_ecc_i;
wire [38:0] rf_rdata_a_ecc_i;
/* cellift = 32'd1 */
input [38:0] rf_rdata_a_ecc_i_t0;
wire [38:0] rf_rdata_a_ecc_i_t0;
/* src = "generated/sv2v_out.v:12849.38-12849.54" */
input [38:0] rf_rdata_b_ecc_i;
wire [38:0] rf_rdata_b_ecc_i;
/* cellift = 32'd1 */
input [38:0] rf_rdata_b_ecc_i_t0;
wire [38:0] rf_rdata_b_ecc_i_t0;
/* src = "generated/sv2v_out.v:12936.7-12936.15" */
wire rf_ren_a;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12936.7-12936.15" */
wire rf_ren_a_t0;
/* src = "generated/sv2v_out.v:12937.7-12937.15" */
wire rf_ren_b;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12937.7-12937.15" */
wire rf_ren_b_t0;
/* src = "generated/sv2v_out.v:12945.13-12945.24" */
wire [4:0] rf_waddr_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12945.13-12945.24" */
wire [4:0] rf_waddr_id_t0;
/* src = "generated/sv2v_out.v:12845.20-12845.33" */
output [4:0] rf_waddr_wb_o;
wire [4:0] rf_waddr_wb_o;
/* cellift = 32'd1 */
output [4:0] rf_waddr_wb_o_t0;
wire [4:0] rf_waddr_wb_o_t0;
/* src = "generated/sv2v_out.v:12940.14-12940.29" */
wire [31:0] rf_wdata_fwd_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12940.14-12940.29" */
wire [31:0] rf_wdata_fwd_wb_t0;
/* src = "generated/sv2v_out.v:12946.14-12946.25" */
wire [31:0] rf_wdata_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12946.14-12946.25" */
wire [31:0] rf_wdata_id_t0;
/* src = "generated/sv2v_out.v:12941.14-12941.26" */
wire [31:0] rf_wdata_lsu;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12941.14-12941.26" */
wire [31:0] rf_wdata_lsu_t0;
/* src = "generated/sv2v_out.v:12939.14-12939.25" */
wire [31:0] rf_wdata_wb;
/* src = "generated/sv2v_out.v:12847.39-12847.56" */
output [38:0] rf_wdata_wb_ecc_o;
wire [38:0] rf_wdata_wb_ecc_o;
/* cellift = 32'd1 */
output [38:0] rf_wdata_wb_ecc_o_t0;
wire [38:0] rf_wdata_wb_ecc_o_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12939.14-12939.25" */
wire [31:0] rf_wdata_wb_t0;
/* src = "generated/sv2v_out.v:12947.7-12947.15" */
wire rf_we_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12947.7-12947.15" */
wire rf_we_id_t0;
/* src = "generated/sv2v_out.v:12943.7-12943.16" */
wire rf_we_lsu;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12943.7-12943.16" */
wire rf_we_lsu_t0;
/* src = "generated/sv2v_out.v:12846.14-12846.24" */
output rf_we_wb_o;
wire rf_we_wb_o;
/* cellift = 32'd1 */
output rf_we_wb_o_t0;
wire rf_we_wb_o_t0;
/* src = "generated/sv2v_out.v:12990.7-12990.18" */
wire rf_write_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12990.7-12990.18" */
wire rf_write_wb_t0;
/* src = "generated/sv2v_out.v:12823.13-12823.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:13023.7-13023.20" */
wire trigger_match;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13023.7-13023.20" */
wire trigger_match_t0;
assign perf_iside_wait = id_in_ready & /* src = "generated/sv2v_out.v:13146.27-13146.56" */ _080_;
assign instr_req_gated = instr_req_int & /* src = "generated/sv2v_out.v:13149.29-13149.84" */ instr_exec;
assign lsu_load_err = lsu_load_err_raw & /* src = "generated/sv2v_out.v:13397.26-13397.91" */ _083_;
assign lsu_store_err = lsu_store_err_raw & /* src = "generated/sv2v_out.v:13398.27-13398.95" */ _085_;
assign rf_we_lsu = lsu_rdata_valid & /* src = "generated/sv2v_out.v:13399.23-13399.87" */ _083_;
assign _000_ = _095_ & /* src = "generated/sv2v_out.v:13437.30-13437.54" */ rf_ren_a;
assign \gen_regfile_ecc.rf_ecc_err_a_id  = _000_ & /* src = "generated/sv2v_out.v:13437.29-13437.75" */ _081_;
assign _002_ = _096_ & /* src = "generated/sv2v_out.v:13438.30-13438.54" */ rf_ren_b;
assign \gen_regfile_ecc.rf_ecc_err_b_id  = _002_ & /* src = "generated/sv2v_out.v:13438.29-13438.75" */ _082_;
assign rf_ecc_err_comb = instr_valid_id & /* src = "generated/sv2v_out.v:13439.29-13439.81" */ _087_;
assign _020_ = id_in_ready_t0 & _080_;
assign instr_req_gated_t0 = instr_req_int_t0 & instr_exec;
assign _023_ = lsu_load_err_raw_t0 & _083_;
assign _026_ = lsu_store_err_raw_t0 & _085_;
assign _029_ = lsu_rdata_valid_t0 & _083_;
assign _032_ = _001_ & _081_;
assign _035_ = _003_ & _082_;
assign _038_ = instr_valid_id_t0 & _087_;
assign _021_ = instr_valid_id_t0 & id_in_ready;
assign _024_ = _084_ & lsu_load_err_raw;
assign _027_ = _086_ & lsu_store_err_raw;
assign _030_ = _084_ & lsu_rdata_valid;
assign _001_ = rf_ren_a_t0 & _095_;
assign _033_ = rf_rd_a_wb_match_t0 & _000_;
assign _003_ = rf_ren_b_t0 & _096_;
assign _036_ = rf_rd_b_wb_match_t0 & _002_;
assign _039_ = _088_ & instr_valid_id;
assign _022_ = id_in_ready_t0 & instr_valid_id_t0;
assign _025_ = lsu_load_err_raw_t0 & _084_;
assign _028_ = lsu_store_err_raw_t0 & _086_;
assign _031_ = lsu_rdata_valid_t0 & _084_;
assign _034_ = _001_ & rf_rd_a_wb_match_t0;
assign _037_ = _003_ & rf_rd_b_wb_match_t0;
assign _040_ = instr_valid_id_t0 & _088_;
assign _065_ = _020_ | _021_;
assign _066_ = _023_ | _024_;
assign _067_ = _026_ | _027_;
assign _068_ = _029_ | _030_;
assign _069_ = _032_ | _033_;
assign _070_ = _035_ | _036_;
assign _071_ = _038_ | _039_;
assign perf_iside_wait_t0 = _065_ | _022_;
assign lsu_load_err_t0 = _066_ | _025_;
assign lsu_store_err_t0 = _067_ | _028_;
assign rf_we_lsu_t0 = _068_ | _031_;
assign \gen_regfile_ecc.rf_ecc_err_a_id_t0  = _069_ | _034_;
assign \gen_regfile_ecc.rf_ecc_err_b_id_t0  = _070_ | _037_;
assign rf_ecc_err_comb_t0 = _071_ | _040_;
assign csr_addr_t0 = { csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access } & alu_operand_b_ex_t0[11:0];
assign _004_ = ~ lsu_load_err;
assign _005_ = ~ outstanding_store_wb;
assign _006_ = ~ outstanding_load_wb;
assign _007_ = ~ \gen_regfile_ecc.rf_ecc_err_a_id ;
assign _008_ = ~ rf_ecc_err_comb;
assign _009_ = ~ _089_;
assign _010_ = ~ lsu_load_resp_intg_err;
assign _011_ = ~ _091_;
assign _012_ = ~ lsu_store_err;
assign _013_ = ~ expecting_store_resp_id;
assign _014_ = ~ expecting_load_resp_id;
assign _015_ = ~ \gen_regfile_ecc.rf_ecc_err_b_id ;
assign _016_ = ~ pc_mismatch_alert;
assign _017_ = ~ csr_shadow_err;
assign _018_ = ~ lsu_store_resp_intg_err;
assign _019_ = ~ instr_intg_err;
assign _041_ = lsu_load_err_t0 & _012_;
assign _044_ = outstanding_store_wb_t0 & _013_;
assign _047_ = outstanding_load_wb_t0 & _014_;
assign _050_ = \gen_regfile_ecc.rf_ecc_err_a_id_t0  & _015_;
assign _053_ = rf_ecc_err_comb_t0 & _016_;
assign _056_ = _090_ & _017_;
assign _059_ = lsu_load_resp_intg_err_t0 & _018_;
assign _062_ = _092_ & _019_;
assign _042_ = lsu_store_err_t0 & _004_;
assign _045_ = expecting_store_resp_id_t0 & _005_;
assign _048_ = expecting_load_resp_id_t0 & _006_;
assign _051_ = \gen_regfile_ecc.rf_ecc_err_b_id_t0  & _007_;
assign _054_ = pc_mismatch_alert_t0 & _008_;
assign _057_ = csr_shadow_err_t0 & _009_;
assign _060_ = lsu_store_resp_intg_err_t0 & _010_;
assign _063_ = instr_intg_err_t0 & _011_;
assign _043_ = lsu_load_err_t0 & lsu_store_err_t0;
assign _046_ = outstanding_store_wb_t0 & expecting_store_resp_id_t0;
assign _049_ = outstanding_load_wb_t0 & expecting_load_resp_id_t0;
assign _052_ = \gen_regfile_ecc.rf_ecc_err_a_id_t0  & \gen_regfile_ecc.rf_ecc_err_b_id_t0 ;
assign _055_ = rf_ecc_err_comb_t0 & pc_mismatch_alert_t0;
assign _058_ = _090_ & csr_shadow_err_t0;
assign _061_ = lsu_load_resp_intg_err_t0 & lsu_store_resp_intg_err_t0;
assign _064_ = _092_ & instr_intg_err_t0;
assign _072_ = _041_ | _042_;
assign _073_ = _044_ | _045_;
assign _074_ = _047_ | _048_;
assign _075_ = _050_ | _051_;
assign _076_ = _053_ | _054_;
assign _077_ = _056_ | _057_;
assign _078_ = _059_ | _060_;
assign _079_ = _062_ | _063_;
assign lsu_resp_err_t0 = _072_ | _043_;
assign _086_ = _073_ | _046_;
assign _084_ = _074_ | _049_;
assign _088_ = _075_ | _052_;
assign _090_ = _076_ | _055_;
assign alert_major_internal_o_t0 = _077_ | _058_;
assign _092_ = _078_ | _061_;
assign alert_major_bus_o_t0 = _079_ | _064_;
assign instr_exec = fetch_enable_i == /* src = "generated/sv2v_out.v:13150.24-13150.61" */ 4'h5;
assign core_busy_o[1] = ! /* src = "generated/sv2v_out.v:13058.30-13058.81" */ _093_;
assign core_busy_o[3] = ! /* src = "generated/sv2v_out.v:13058.30-13058.81" */ _094_;
assign _080_ = ~ /* src = "generated/sv2v_out.v:13146.41-13146.56" */ instr_valid_id;
assign _081_ = ~ /* src = "generated/sv2v_out.v:13437.58-13437.75" */ rf_rd_a_wb_match;
assign _082_ = ~ /* src = "generated/sv2v_out.v:13438.58-13438.75" */ rf_rd_b_wb_match;
assign lsu_resp_err = lsu_load_err | /* src = "generated/sv2v_out.v:13322.24-13322.52" */ lsu_store_err;
assign _085_ = outstanding_store_wb | /* src = "generated/sv2v_out.v:13398.48-13398.94" */ expecting_store_resp_id;
assign _083_ = outstanding_load_wb | /* src = "generated/sv2v_out.v:13399.42-13399.86" */ expecting_load_resp_id;
assign _087_ = \gen_regfile_ecc.rf_ecc_err_a_id  | /* src = "generated/sv2v_out.v:13439.47-13439.80" */ \gen_regfile_ecc.rf_ecc_err_b_id ;
assign _089_ = rf_ecc_err_comb | /* src = "generated/sv2v_out.v:13463.35-13463.70" */ pc_mismatch_alert;
assign alert_major_internal_o = _089_ | /* src = "generated/sv2v_out.v:13463.34-13463.88" */ csr_shadow_err;
assign _091_ = lsu_load_resp_intg_err | /* src = "generated/sv2v_out.v:13464.30-13464.78" */ lsu_store_resp_intg_err;
assign alert_major_bus_o = _091_ | /* src = "generated/sv2v_out.v:13464.29-13464.96" */ instr_intg_err;
assign core_busy_o[0] = | /* src = "generated/sv2v_out.v:13055.30-13055.80" */ \g_core_busy_secure.busy_bits_buf [2:0];
assign core_busy_o[2] = | /* src = "generated/sv2v_out.v:13055.30-13055.80" */ \g_core_busy_secure.busy_bits_buf [8:6];
assign _093_ = | /* src = "generated/sv2v_out.v:13058.30-13058.81" */ \g_core_busy_secure.busy_bits_buf [5:3];
assign _094_ = | /* src = "generated/sv2v_out.v:13058.30-13058.81" */ \g_core_busy_secure.busy_bits_buf [11:9];
assign _095_ = | /* src = "generated/sv2v_out.v:13437.30-13437.43" */ \gen_regfile_ecc.rf_ecc_err_a ;
assign _096_ = | /* src = "generated/sv2v_out.v:13438.30-13438.43" */ \gen_regfile_ecc.rf_ecc_err_b ;
assign csr_addr = csr_access ? /* src = "generated/sv2v_out.v:13470.34-13470.88" */ alu_operand_b_ex[11:0] : 12'h000;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13486.4-13558.3" */
\$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers  cs_registers_i (
.boot_addr_i(boot_addr_i),
.boot_addr_i_t0(boot_addr_i_t0),
.branch_i(perf_branch),
.branch_i_t0(perf_branch_t0),
.branch_taken_i(perf_tbranch),
.branch_taken_i_t0(perf_tbranch_t0),
.clk_i(clk_i),
.csr_access_i(csr_access),
.csr_access_i_t0(csr_access_t0),
.csr_addr_i(csr_addr),
.csr_addr_i_t0(csr_addr_t0),
.csr_depc_o(csr_depc),
.csr_depc_o_t0(csr_depc_t0),
.csr_mcause_i(exc_cause),
.csr_mcause_i_t0(exc_cause_t0),
.csr_mepc_o(csr_mepc),
.csr_mepc_o_t0(csr_mepc_t0),
.csr_mstatus_mie_o(csr_mstatus_mie),
.csr_mstatus_mie_o_t0(csr_mstatus_mie_t0),
.csr_mstatus_tw_o(csr_mstatus_tw),
.csr_mstatus_tw_o_t0(csr_mstatus_tw_t0),
.csr_mtval_i(csr_mtval),
.csr_mtval_i_t0(csr_mtval_t0),
.csr_mtval_o(crash_dump_mtval),
.csr_mtval_o_t0(crash_dump_mtval_t0),
.csr_mtvec_init_i(csr_mtvec_init),
.csr_mtvec_init_i_t0(csr_mtvec_init_t0),
.csr_mtvec_o(csr_mtvec),
.csr_mtvec_o_t0(csr_mtvec_t0),
.csr_op_en_i(csr_op_en),
.csr_op_en_i_t0(csr_op_en_t0),
.csr_op_i(csr_op),
.csr_op_i_t0(csr_op_t0),
.csr_pmp_addr_o(csr_pmp_addr),
.csr_pmp_addr_o_t0(csr_pmp_addr_t0),
.csr_pmp_cfg_o(csr_pmp_cfg),
.csr_pmp_cfg_o_t0(csr_pmp_cfg_t0),
.csr_pmp_mseccfg_o(csr_pmp_mseccfg),
.csr_pmp_mseccfg_o_t0(csr_pmp_mseccfg_t0),
.csr_rdata_o(csr_rdata),
.csr_rdata_o_t0(csr_rdata_t0),
.csr_restore_dret_i(csr_restore_dret_id),
.csr_restore_dret_i_t0(csr_restore_dret_id_t0),
.csr_restore_mret_i(csr_restore_mret_id),
.csr_restore_mret_i_t0(csr_restore_mret_id_t0),
.csr_save_cause_i(csr_save_cause),
.csr_save_cause_i_t0(csr_save_cause_t0),
.csr_save_id_i(csr_save_id),
.csr_save_id_i_t0(csr_save_id_t0),
.csr_save_if_i(csr_save_if),
.csr_save_if_i_t0(csr_save_if_t0),
.csr_save_wb_i(csr_save_wb),
.csr_save_wb_i_t0(csr_save_wb_t0),
.csr_shadow_err_o(csr_shadow_err),
.csr_shadow_err_o_t0(csr_shadow_err_t0),
.csr_wdata_i(alu_operand_a_ex),
.csr_wdata_i_t0(alu_operand_a_ex_t0),
.data_ind_timing_o(data_ind_timing),
.data_ind_timing_o_t0(data_ind_timing_t0),
.debug_cause_i(debug_cause),
.debug_cause_i_t0(debug_cause_t0),
.debug_csr_save_i(debug_csr_save),
.debug_csr_save_i_t0(debug_csr_save_t0),
.debug_ebreakm_o(debug_ebreakm),
.debug_ebreakm_o_t0(debug_ebreakm_t0),
.debug_ebreaku_o(debug_ebreaku),
.debug_ebreaku_o_t0(debug_ebreaku_t0),
.debug_mode_entering_i(debug_mode_entering),
.debug_mode_entering_i_t0(debug_mode_entering_t0),
.debug_mode_i(debug_mode),
.debug_mode_i_t0(debug_mode_t0),
.debug_single_step_o(debug_single_step),
.debug_single_step_o_t0(debug_single_step_t0),
.div_wait_i(perf_div_wait),
.div_wait_i_t0(perf_div_wait_t0),
.double_fault_seen_o(double_fault_seen_o),
.double_fault_seen_o_t0(double_fault_seen_o_t0),
.dside_wait_i(perf_dside_wait),
.dside_wait_i_t0(perf_dside_wait_t0),
.dummy_instr_en_o(dummy_instr_en),
.dummy_instr_en_o_t0(dummy_instr_en_t0),
.dummy_instr_mask_o(dummy_instr_mask),
.dummy_instr_mask_o_t0(dummy_instr_mask_t0),
.dummy_instr_seed_en_o(dummy_instr_seed_en),
.dummy_instr_seed_en_o_t0(dummy_instr_seed_en_t0),
.dummy_instr_seed_o(dummy_instr_seed),
.dummy_instr_seed_o_t0(dummy_instr_seed_t0),
.hart_id_i(hart_id_i),
.hart_id_i_t0(hart_id_i_t0),
.ic_scr_key_valid_i(ic_scr_key_valid_i),
.ic_scr_key_valid_i_t0(ic_scr_key_valid_i_t0),
.icache_enable_o(icache_enable),
.icache_enable_o_t0(icache_enable_t0),
.illegal_csr_insn_o(illegal_csr_insn_id),
.illegal_csr_insn_o_t0(illegal_csr_insn_id_t0),
.instr_ret_compressed_i(perf_instr_ret_compressed_wb),
.instr_ret_compressed_i_t0(perf_instr_ret_compressed_wb_t0),
.instr_ret_compressed_spec_i(perf_instr_ret_compressed_wb_spec),
.instr_ret_compressed_spec_i_t0(perf_instr_ret_compressed_wb_spec_t0),
.instr_ret_i(perf_instr_ret_wb),
.instr_ret_i_t0(perf_instr_ret_wb_t0),
.instr_ret_spec_i(perf_instr_ret_wb_spec),
.instr_ret_spec_i_t0(perf_instr_ret_wb_spec_t0),
.irq_external_i(irq_external_i),
.irq_external_i_t0(irq_external_i_t0),
.irq_fast_i(irq_fast_i),
.irq_fast_i_t0(irq_fast_i_t0),
.irq_pending_o(irq_pending_o),
.irq_pending_o_t0(irq_pending_o_t0),
.irq_software_i(irq_software_i),
.irq_software_i_t0(irq_software_i_t0),
.irq_timer_i(irq_timer_i),
.irq_timer_i_t0(irq_timer_i_t0),
.irqs_o(irqs),
.irqs_o_t0(irqs_t0),
.iside_wait_i(perf_iside_wait),
.iside_wait_i_t0(perf_iside_wait_t0),
.jump_i(perf_jump),
.jump_i_t0(perf_jump_t0),
.mem_load_i(perf_load),
.mem_load_i_t0(perf_load_t0),
.mem_store_i(perf_store),
.mem_store_i_t0(perf_store_t0),
.mul_wait_i(perf_mul_wait),
.mul_wait_i_t0(perf_mul_wait_t0),
.nmi_mode_i(nmi_mode),
.nmi_mode_i_t0(nmi_mode_t0),
.pc_id_i(pc_id),
.pc_id_i_t0(pc_id_t0),
.pc_if_i(pc_if),
.pc_if_i_t0(pc_if_t0),
.pc_wb_i(pc_wb),
.pc_wb_i_t0(pc_wb_t0),
.priv_mode_id_o(priv_mode_id),
.priv_mode_id_o_t0(priv_mode_id_t0),
.priv_mode_lsu_o(\g_no_pmp.unused_priv_lvl_ls ),
.priv_mode_lsu_o_t0(\g_no_pmp.unused_priv_lvl_ls_t0 ),
.rst_ni(rst_ni),
.trigger_match_o(trigger_match),
.trigger_match_o_t0(trigger_match_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13292.4-13319.3" */
\$paramod$a308247794889ee6093207090edbf289adef8be1\ibex_ex_block  ex_block_i (
.alu_adder_result_ex_o(alu_adder_result_ex),
.alu_adder_result_ex_o_t0(alu_adder_result_ex_t0),
.alu_instr_first_cycle_i(instr_first_cycle_id),
.alu_instr_first_cycle_i_t0(instr_first_cycle_id_t0),
.alu_operand_a_i(alu_operand_a_ex),
.alu_operand_a_i_t0(alu_operand_a_ex_t0),
.alu_operand_b_i(alu_operand_b_ex),
.alu_operand_b_i_t0(alu_operand_b_ex_t0),
.alu_operator_i(alu_operator_ex),
.alu_operator_i_t0(alu_operator_ex_t0),
.branch_decision_o(branch_decision),
.branch_decision_o_t0(branch_decision_t0),
.branch_target_o(branch_target_ex),
.branch_target_o_t0(branch_target_ex_t0),
.bt_a_operand_i(bt_a_operand),
.bt_a_operand_i_t0(bt_a_operand_t0),
.bt_b_operand_i(bt_b_operand),
.bt_b_operand_i_t0(bt_b_operand_t0),
.clk_i(clk_i),
.data_ind_timing_i(data_ind_timing),
.data_ind_timing_i_t0(data_ind_timing_t0),
.div_en_i(div_en_ex),
.div_en_i_t0(div_en_ex_t0),
.div_sel_i(div_sel_ex),
.div_sel_i_t0(div_sel_ex_t0),
.ex_valid_o(ex_valid),
.ex_valid_o_t0(ex_valid_t0),
.imd_val_d_o(imd_val_d_ex),
.imd_val_d_o_t0(imd_val_d_ex_t0),
.imd_val_q_i(imd_val_q_ex),
.imd_val_q_i_t0(imd_val_q_ex_t0),
.imd_val_we_o(imd_val_we_ex),
.imd_val_we_o_t0(imd_val_we_ex_t0),
.mult_en_i(mult_en_ex),
.mult_en_i_t0(mult_en_ex_t0),
.mult_sel_i(mult_sel_ex),
.mult_sel_i_t0(mult_sel_ex_t0),
.multdiv_operand_a_i(multdiv_operand_a_ex),
.multdiv_operand_a_i_t0(multdiv_operand_a_ex_t0),
.multdiv_operand_b_i(multdiv_operand_b_ex),
.multdiv_operand_b_i_t0(multdiv_operand_b_ex_t0),
.multdiv_operator_i(multdiv_operator_ex),
.multdiv_operator_i_t0(multdiv_operator_ex_t0),
.multdiv_ready_id_i(multdiv_ready_id),
.multdiv_ready_id_i_t0(multdiv_ready_id_t0),
.multdiv_signed_mode_i(multdiv_signed_mode_ex),
.multdiv_signed_mode_i_t0(multdiv_signed_mode_ex_t0),
.result_ex_o(result_ex),
.result_ex_o_t0(result_ex_t0),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13048.36-13051.5" */
\$paramod\prim_buf\Width=32'00000000000000000000000000001100  \g_core_busy_secure.u_fetch_enable_buf  (
.in_i({ ctrl_busy, if_busy, lsu_busy, ctrl_busy, if_busy, lsu_busy, ctrl_busy, if_busy, lsu_busy, ctrl_busy, if_busy, lsu_busy }),
.in_i_t0({ ctrl_busy_t0, if_busy_t0, lsu_busy_t0, ctrl_busy_t0, if_busy_t0, lsu_busy_t0, ctrl_busy_t0, if_busy_t0, lsu_busy_t0, ctrl_busy_t0, if_busy_t0, lsu_busy_t0 }),
.out_o(\g_core_busy_secure.busy_bits_buf ),
.out_o_t0(\g_core_busy_secure.busy_bits_buf_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13427.30-13430.5" */
prim_secded_inv_39_32_dec \gen_regfile_ecc.regfile_ecc_dec_a  (
.data_i(rf_rdata_a_ecc_i),
.data_i_t0(rf_rdata_a_ecc_i_t0),
.err_o(\gen_regfile_ecc.rf_ecc_err_a ),
.err_o_t0(\gen_regfile_ecc.rf_ecc_err_a_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13431.30-13434.5" */
prim_secded_inv_39_32_dec \gen_regfile_ecc.regfile_ecc_dec_b  (
.data_i(rf_rdata_b_ecc_i),
.data_i_t0(rf_rdata_b_ecc_i_t0),
.err_o(\gen_regfile_ecc.rf_ecc_err_b ),
.err_o_t0(\gen_regfile_ecc.rf_ecc_err_b_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13423.30-13426.5" */
prim_secded_inv_39_32_enc \gen_regfile_ecc.regfile_ecc_enc  (
.data_i(rf_wdata_wb),
.data_i_t0(rf_wdata_wb_t0),
.data_o(rf_wdata_wb_ecc_o),
.data_o_t0(rf_wdata_wb_ecc_o_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13168.4-13286.3" */
\$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  id_stage_i (
.alu_operand_a_ex_o(alu_operand_a_ex),
.alu_operand_a_ex_o_t0(alu_operand_a_ex_t0),
.alu_operand_b_ex_o(alu_operand_b_ex),
.alu_operand_b_ex_o_t0(alu_operand_b_ex_t0),
.alu_operator_ex_o(alu_operator_ex),
.alu_operator_ex_o_t0(alu_operator_ex_t0),
.branch_decision_i(branch_decision),
.branch_decision_i_t0(branch_decision_t0),
.bt_a_operand_o(bt_a_operand),
.bt_a_operand_o_t0(bt_a_operand_t0),
.bt_b_operand_o(bt_b_operand),
.bt_b_operand_o_t0(bt_b_operand_t0),
.clk_i(clk_i),
.csr_access_o(csr_access),
.csr_access_o_t0(csr_access_t0),
.csr_mstatus_mie_i(csr_mstatus_mie),
.csr_mstatus_mie_i_t0(csr_mstatus_mie_t0),
.csr_mstatus_tw_i(csr_mstatus_tw),
.csr_mstatus_tw_i_t0(csr_mstatus_tw_t0),
.csr_mtval_o(csr_mtval),
.csr_mtval_o_t0(csr_mtval_t0),
.csr_op_en_o(csr_op_en),
.csr_op_en_o_t0(csr_op_en_t0),
.csr_op_o(csr_op),
.csr_op_o_t0(csr_op_t0),
.csr_rdata_i(csr_rdata),
.csr_rdata_i_t0(csr_rdata_t0),
.csr_restore_dret_id_o(csr_restore_dret_id),
.csr_restore_dret_id_o_t0(csr_restore_dret_id_t0),
.csr_restore_mret_id_o(csr_restore_mret_id),
.csr_restore_mret_id_o_t0(csr_restore_mret_id_t0),
.csr_save_cause_o(csr_save_cause),
.csr_save_cause_o_t0(csr_save_cause_t0),
.csr_save_id_o(csr_save_id),
.csr_save_id_o_t0(csr_save_id_t0),
.csr_save_if_o(csr_save_if),
.csr_save_if_o_t0(csr_save_if_t0),
.csr_save_wb_o(csr_save_wb),
.csr_save_wb_o_t0(csr_save_wb_t0),
.ctrl_busy_o(ctrl_busy),
.ctrl_busy_o_t0(ctrl_busy_t0),
.data_ind_timing_i(data_ind_timing),
.data_ind_timing_i_t0(data_ind_timing_t0),
.debug_cause_o(debug_cause),
.debug_cause_o_t0(debug_cause_t0),
.debug_csr_save_o(debug_csr_save),
.debug_csr_save_o_t0(debug_csr_save_t0),
.debug_ebreakm_i(debug_ebreakm),
.debug_ebreakm_i_t0(debug_ebreakm_t0),
.debug_ebreaku_i(debug_ebreaku),
.debug_ebreaku_i_t0(debug_ebreaku_t0),
.debug_mode_entering_o(debug_mode_entering),
.debug_mode_entering_o_t0(debug_mode_entering_t0),
.debug_mode_o(debug_mode),
.debug_mode_o_t0(debug_mode_t0),
.debug_req_i(debug_req_i),
.debug_req_i_t0(debug_req_i_t0),
.debug_single_step_i(debug_single_step),
.debug_single_step_i_t0(debug_single_step_t0),
.div_en_ex_o(div_en_ex),
.div_en_ex_o_t0(div_en_ex_t0),
.div_sel_ex_o(div_sel_ex),
.div_sel_ex_o_t0(div_sel_ex_t0),
.en_wb_o(en_wb),
.en_wb_o_t0(en_wb_t0),
.ex_valid_i(ex_valid),
.ex_valid_i_t0(ex_valid_t0),
.exc_cause_o(exc_cause),
.exc_cause_o_t0(exc_cause_t0),
.exc_pc_mux_o(exc_pc_mux_id),
.exc_pc_mux_o_t0(exc_pc_mux_id_t0),
.expecting_load_resp_o(expecting_load_resp_id),
.expecting_load_resp_o_t0(expecting_load_resp_id_t0),
.expecting_store_resp_o(expecting_store_resp_id),
.expecting_store_resp_o_t0(expecting_store_resp_id_t0),
.icache_inval_o(icache_inval),
.icache_inval_o_t0(icache_inval_t0),
.id_in_ready_o(id_in_ready),
.id_in_ready_o_t0(id_in_ready_t0),
.illegal_c_insn_i(illegal_c_insn_id),
.illegal_c_insn_i_t0(illegal_c_insn_id_t0),
.illegal_csr_insn_i(illegal_csr_insn_id),
.illegal_csr_insn_i_t0(illegal_csr_insn_id_t0),
.illegal_insn_o(illegal_insn_id),
.illegal_insn_o_t0(illegal_insn_id_t0),
.imd_val_d_ex_i(imd_val_d_ex),
.imd_val_d_ex_i_t0(imd_val_d_ex_t0),
.imd_val_q_ex_o(imd_val_q_ex),
.imd_val_q_ex_o_t0(imd_val_q_ex_t0),
.imd_val_we_ex_i(imd_val_we_ex),
.imd_val_we_ex_i_t0(imd_val_we_ex_t0),
.instr_bp_taken_i(instr_bp_taken_id),
.instr_bp_taken_i_t0(instr_bp_taken_id_t0),
.instr_exec_i(instr_exec),
.instr_exec_i_t0(1'h0),
.instr_fetch_err_i(instr_fetch_err),
.instr_fetch_err_i_t0(instr_fetch_err_t0),
.instr_fetch_err_plus2_i(instr_fetch_err_plus2),
.instr_fetch_err_plus2_i_t0(instr_fetch_err_plus2_t0),
.instr_first_cycle_id_o(instr_first_cycle_id),
.instr_first_cycle_id_o_t0(instr_first_cycle_id_t0),
.instr_id_done_o(instr_id_done),
.instr_id_done_o_t0(instr_id_done_t0),
.instr_is_compressed_i(instr_is_compressed_id),
.instr_is_compressed_i_t0(instr_is_compressed_id_t0),
.instr_perf_count_id_o(instr_perf_count_id),
.instr_perf_count_id_o_t0(instr_perf_count_id_t0),
.instr_rdata_alu_i(instr_rdata_alu_id),
.instr_rdata_alu_i_t0(instr_rdata_alu_id_t0),
.instr_rdata_c_i(instr_rdata_c_id),
.instr_rdata_c_i_t0(instr_rdata_c_id_t0),
.instr_rdata_i(instr_rdata_id),
.instr_rdata_i_t0(instr_rdata_id_t0),
.instr_req_o(instr_req_int),
.instr_req_o_t0(instr_req_int_t0),
.instr_type_wb_o(instr_type_wb),
.instr_type_wb_o_t0(instr_type_wb_t0),
.instr_valid_clear_o(instr_valid_clear),
.instr_valid_clear_o_t0(instr_valid_clear_t0),
.instr_valid_i(instr_valid_id),
.instr_valid_i_t0(instr_valid_id_t0),
.irq_nm_i(irq_nm_i),
.irq_nm_i_t0(irq_nm_i_t0),
.irq_pending_i(irq_pending_o),
.irq_pending_i_t0(irq_pending_o_t0),
.irqs_i(irqs),
.irqs_i_t0(irqs_t0),
.lsu_addr_incr_req_i(lsu_addr_incr_req),
.lsu_addr_incr_req_i_t0(lsu_addr_incr_req_t0),
.lsu_addr_last_i(lsu_addr_last),
.lsu_addr_last_i_t0(lsu_addr_last_t0),
.lsu_load_err_i(lsu_load_err),
.lsu_load_err_i_t0(lsu_load_err_t0),
.lsu_load_resp_intg_err_i(lsu_load_resp_intg_err),
.lsu_load_resp_intg_err_i_t0(lsu_load_resp_intg_err_t0),
.lsu_req_done_i(lsu_req_done),
.lsu_req_done_i_t0(lsu_req_done_t0),
.lsu_req_o(lsu_req),
.lsu_req_o_t0(lsu_req_t0),
.lsu_resp_valid_i(lsu_resp_valid),
.lsu_resp_valid_i_t0(lsu_resp_valid_t0),
.lsu_sign_ext_o(lsu_sign_ext),
.lsu_sign_ext_o_t0(lsu_sign_ext_t0),
.lsu_store_err_i(lsu_store_err),
.lsu_store_err_i_t0(lsu_store_err_t0),
.lsu_store_resp_intg_err_i(lsu_store_resp_intg_err),
.lsu_store_resp_intg_err_i_t0(lsu_store_resp_intg_err_t0),
.lsu_type_o(lsu_type),
.lsu_type_o_t0(lsu_type_t0),
.lsu_wdata_o(lsu_wdata),
.lsu_wdata_o_t0(lsu_wdata_t0),
.lsu_we_o(lsu_we),
.lsu_we_o_t0(lsu_we_t0),
.mult_en_ex_o(mult_en_ex),
.mult_en_ex_o_t0(mult_en_ex_t0),
.mult_sel_ex_o(mult_sel_ex),
.mult_sel_ex_o_t0(mult_sel_ex_t0),
.multdiv_operand_a_ex_o(multdiv_operand_a_ex),
.multdiv_operand_a_ex_o_t0(multdiv_operand_a_ex_t0),
.multdiv_operand_b_ex_o(multdiv_operand_b_ex),
.multdiv_operand_b_ex_o_t0(multdiv_operand_b_ex_t0),
.multdiv_operator_ex_o(multdiv_operator_ex),
.multdiv_operator_ex_o_t0(multdiv_operator_ex_t0),
.multdiv_ready_id_o(multdiv_ready_id),
.multdiv_ready_id_o_t0(multdiv_ready_id_t0),
.multdiv_signed_mode_ex_o(multdiv_signed_mode_ex),
.multdiv_signed_mode_ex_o_t0(multdiv_signed_mode_ex_t0),
.nmi_mode_o(nmi_mode),
.nmi_mode_o_t0(nmi_mode_t0),
.nt_branch_addr_o(nt_branch_addr),
.nt_branch_addr_o_t0(nt_branch_addr_t0),
.nt_branch_mispredict_o(nt_branch_mispredict),
.nt_branch_mispredict_o_t0(nt_branch_mispredict_t0),
.outstanding_load_wb_i(outstanding_load_wb),
.outstanding_load_wb_i_t0(outstanding_load_wb_t0),
.outstanding_store_wb_i(outstanding_store_wb),
.outstanding_store_wb_i_t0(outstanding_store_wb_t0),
.pc_id_i(pc_id),
.pc_id_i_t0(pc_id_t0),
.pc_mux_o(pc_mux_id),
.pc_mux_o_t0(pc_mux_id_t0),
.pc_set_o(pc_set),
.pc_set_o_t0(pc_set_t0),
.perf_branch_o(perf_branch),
.perf_branch_o_t0(perf_branch_t0),
.perf_div_wait_o(perf_div_wait),
.perf_div_wait_o_t0(perf_div_wait_t0),
.perf_dside_wait_o(perf_dside_wait),
.perf_dside_wait_o_t0(perf_dside_wait_t0),
.perf_jump_o(perf_jump),
.perf_jump_o_t0(perf_jump_t0),
.perf_mul_wait_o(perf_mul_wait),
.perf_mul_wait_o_t0(perf_mul_wait_t0),
.perf_tbranch_o(perf_tbranch),
.perf_tbranch_o_t0(perf_tbranch_t0),
.priv_mode_i(priv_mode_id),
.priv_mode_i_t0(priv_mode_id_t0),
.ready_wb_i(ready_wb),
.ready_wb_i_t0(ready_wb_t0),
.result_ex_i(result_ex),
.result_ex_i_t0(result_ex_t0),
.rf_raddr_a_o(rf_raddr_a_o),
.rf_raddr_a_o_t0(rf_raddr_a_o_t0),
.rf_raddr_b_o(rf_raddr_b_o),
.rf_raddr_b_o_t0(rf_raddr_b_o_t0),
.rf_rd_a_wb_match_o(rf_rd_a_wb_match),
.rf_rd_a_wb_match_o_t0(rf_rd_a_wb_match_t0),
.rf_rd_b_wb_match_o(rf_rd_b_wb_match),
.rf_rd_b_wb_match_o_t0(rf_rd_b_wb_match_t0),
.rf_rdata_a_i(rf_rdata_a_ecc_i[31:0]),
.rf_rdata_a_i_t0(rf_rdata_a_ecc_i_t0[31:0]),
.rf_rdata_b_i(rf_rdata_b_ecc_i[31:0]),
.rf_rdata_b_i_t0(rf_rdata_b_ecc_i_t0[31:0]),
.rf_ren_a_o(rf_ren_a),
.rf_ren_a_o_t0(rf_ren_a_t0),
.rf_ren_b_o(rf_ren_b),
.rf_ren_b_o_t0(rf_ren_b_t0),
.rf_waddr_id_o(rf_waddr_id),
.rf_waddr_id_o_t0(rf_waddr_id_t0),
.rf_waddr_wb_i(rf_waddr_wb_o),
.rf_waddr_wb_i_t0(rf_waddr_wb_o_t0),
.rf_wdata_fwd_wb_i(rf_wdata_fwd_wb),
.rf_wdata_fwd_wb_i_t0(rf_wdata_fwd_wb_t0),
.rf_wdata_id_o(rf_wdata_id),
.rf_wdata_id_o_t0(rf_wdata_id_t0),
.rf_we_id_o(rf_we_id),
.rf_we_id_o_t0(rf_we_id_t0),
.rf_write_wb_i(rf_write_wb),
.rf_write_wb_i_t0(rf_write_wb_t0),
.rst_ni(rst_ni),
.trigger_match_i(trigger_match),
.trigger_match_i_t0(trigger_match_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13084.4-13145.3" */
\$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  if_stage_i (
.boot_addr_i(boot_addr_i),
.boot_addr_i_t0(boot_addr_i_t0),
.branch_target_ex_i(branch_target_ex),
.branch_target_ex_i_t0(branch_target_ex_t0),
.clk_i(clk_i),
.csr_depc_i(csr_depc),
.csr_depc_i_t0(csr_depc_t0),
.csr_mepc_i(csr_mepc),
.csr_mepc_i_t0(csr_mepc_t0),
.csr_mtvec_i(csr_mtvec),
.csr_mtvec_i_t0(csr_mtvec_t0),
.csr_mtvec_init_o(csr_mtvec_init),
.csr_mtvec_init_o_t0(csr_mtvec_init_t0),
.dummy_instr_en_i(dummy_instr_en),
.dummy_instr_en_i_t0(dummy_instr_en_t0),
.dummy_instr_id_o(dummy_instr_id_o),
.dummy_instr_id_o_t0(dummy_instr_id_o_t0),
.dummy_instr_mask_i(dummy_instr_mask),
.dummy_instr_mask_i_t0(dummy_instr_mask_t0),
.dummy_instr_seed_en_i(dummy_instr_seed_en),
.dummy_instr_seed_en_i_t0(dummy_instr_seed_en_t0),
.dummy_instr_seed_i(dummy_instr_seed),
.dummy_instr_seed_i_t0(dummy_instr_seed_t0),
.exc_cause(exc_cause),
.exc_cause_t0(exc_cause_t0),
.exc_pc_mux_i(exc_pc_mux_id),
.exc_pc_mux_i_t0(exc_pc_mux_id_t0),
.ic_data_addr_o(ic_data_addr_o),
.ic_data_addr_o_t0(ic_data_addr_o_t0),
.ic_data_rdata_i(ic_data_rdata_i),
.ic_data_rdata_i_t0(ic_data_rdata_i_t0),
.ic_data_req_o(ic_data_req_o),
.ic_data_req_o_t0(ic_data_req_o_t0),
.ic_data_wdata_o(ic_data_wdata_o),
.ic_data_wdata_o_t0(ic_data_wdata_o_t0),
.ic_data_write_o(ic_data_write_o),
.ic_data_write_o_t0(ic_data_write_o_t0),
.ic_scr_key_req_o(ic_scr_key_req_o),
.ic_scr_key_req_o_t0(ic_scr_key_req_o_t0),
.ic_scr_key_valid_i(ic_scr_key_valid_i),
.ic_scr_key_valid_i_t0(ic_scr_key_valid_i_t0),
.ic_tag_addr_o(ic_tag_addr_o),
.ic_tag_addr_o_t0(ic_tag_addr_o_t0),
.ic_tag_rdata_i(ic_tag_rdata_i),
.ic_tag_rdata_i_t0(ic_tag_rdata_i_t0),
.ic_tag_req_o(ic_tag_req_o),
.ic_tag_req_o_t0(ic_tag_req_o_t0),
.ic_tag_wdata_o(ic_tag_wdata_o),
.ic_tag_wdata_o_t0(ic_tag_wdata_o_t0),
.ic_tag_write_o(ic_tag_write_o),
.ic_tag_write_o_t0(ic_tag_write_o_t0),
.icache_ecc_error_o(alert_minor_o),
.icache_ecc_error_o_t0(alert_minor_o_t0),
.icache_enable_i(icache_enable),
.icache_enable_i_t0(icache_enable_t0),
.icache_inval_i(icache_inval),
.icache_inval_i_t0(icache_inval_t0),
.id_in_ready_i(id_in_ready),
.id_in_ready_i_t0(id_in_ready_t0),
.if_busy_o(if_busy),
.if_busy_o_t0(if_busy_t0),
.illegal_c_insn_id_o(illegal_c_insn_id),
.illegal_c_insn_id_o_t0(illegal_c_insn_id_t0),
.instr_addr_o(instr_addr_o),
.instr_addr_o_t0(instr_addr_o_t0),
.instr_bp_taken_o(instr_bp_taken_id),
.instr_bp_taken_o_t0(instr_bp_taken_id_t0),
.instr_bus_err_i(instr_err_i),
.instr_bus_err_i_t0(instr_err_i_t0),
.instr_fetch_err_o(instr_fetch_err),
.instr_fetch_err_o_t0(instr_fetch_err_t0),
.instr_fetch_err_plus2_o(instr_fetch_err_plus2),
.instr_fetch_err_plus2_o_t0(instr_fetch_err_plus2_t0),
.instr_gnt_i(instr_gnt_i),
.instr_gnt_i_t0(instr_gnt_i_t0),
.instr_intg_err_o(instr_intg_err),
.instr_intg_err_o_t0(instr_intg_err_t0),
.instr_is_compressed_id_o(instr_is_compressed_id),
.instr_is_compressed_id_o_t0(instr_is_compressed_id_t0),
.instr_new_id_o(instr_new_id),
.instr_new_id_o_t0(instr_new_id_t0),
.instr_rdata_alu_id_o(instr_rdata_alu_id),
.instr_rdata_alu_id_o_t0(instr_rdata_alu_id_t0),
.instr_rdata_c_id_o(instr_rdata_c_id),
.instr_rdata_c_id_o_t0(instr_rdata_c_id_t0),
.instr_rdata_i(instr_rdata_i),
.instr_rdata_i_t0(instr_rdata_i_t0),
.instr_rdata_id_o(instr_rdata_id),
.instr_rdata_id_o_t0(instr_rdata_id_t0),
.instr_req_o(instr_req_o),
.instr_req_o_t0(instr_req_o_t0),
.instr_rvalid_i(instr_rvalid_i),
.instr_rvalid_i_t0(instr_rvalid_i_t0),
.instr_valid_clear_i(instr_valid_clear),
.instr_valid_clear_i_t0(instr_valid_clear_t0),
.instr_valid_id_o(instr_valid_id),
.instr_valid_id_o_t0(instr_valid_id_t0),
.nt_branch_addr_i(nt_branch_addr),
.nt_branch_addr_i_t0(nt_branch_addr_t0),
.nt_branch_mispredict_i(nt_branch_mispredict),
.nt_branch_mispredict_i_t0(nt_branch_mispredict_t0),
.pc_id_o(pc_id),
.pc_id_o_t0(pc_id_t0),
.pc_if_o(pc_if),
.pc_if_o_t0(pc_if_t0),
.pc_mismatch_alert_o(pc_mismatch_alert),
.pc_mismatch_alert_o_t0(pc_mismatch_alert_t0),
.pc_mux_i(pc_mux_id),
.pc_mux_i_t0(pc_mux_id_t0),
.pc_set_i(pc_set),
.pc_set_i_t0(pc_set_t0),
.pmp_err_if_i(1'h0),
.pmp_err_if_i_t0(1'h0),
.pmp_err_if_plus2_i(1'h0),
.pmp_err_if_plus2_i_t0(1'h0),
.req_i(instr_req_gated),
.req_i_t0(instr_req_gated_t0),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13326.4-13358.3" */
\$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  load_store_unit_i (
.adder_result_ex_i(alu_adder_result_ex),
.adder_result_ex_i_t0(alu_adder_result_ex_t0),
.addr_incr_req_o(lsu_addr_incr_req),
.addr_incr_req_o_t0(lsu_addr_incr_req_t0),
.addr_last_o(lsu_addr_last),
.addr_last_o_t0(lsu_addr_last_t0),
.busy_o(lsu_busy),
.busy_o_t0(lsu_busy_t0),
.clk_i(clk_i),
.data_addr_o(data_addr_o),
.data_addr_o_t0(data_addr_o_t0),
.data_be_o(data_be_o),
.data_be_o_t0(data_be_o_t0),
.data_bus_err_i(data_err_i),
.data_bus_err_i_t0(data_err_i_t0),
.data_gnt_i(data_gnt_i),
.data_gnt_i_t0(data_gnt_i_t0),
.data_pmp_err_i(1'h0),
.data_pmp_err_i_t0(1'h0),
.data_rdata_i(data_rdata_i),
.data_rdata_i_t0(data_rdata_i_t0),
.data_req_o(data_req_o),
.data_req_o_t0(data_req_o_t0),
.data_rvalid_i(data_rvalid_i),
.data_rvalid_i_t0(data_rvalid_i_t0),
.data_wdata_o(data_wdata_o),
.data_wdata_o_t0(data_wdata_o_t0),
.data_we_o(data_we_o),
.data_we_o_t0(data_we_o_t0),
.load_err_o(lsu_load_err_raw),
.load_err_o_t0(lsu_load_err_raw_t0),
.load_resp_intg_err_o(lsu_load_resp_intg_err),
.load_resp_intg_err_o_t0(lsu_load_resp_intg_err_t0),
.lsu_rdata_o(rf_wdata_lsu),
.lsu_rdata_o_t0(rf_wdata_lsu_t0),
.lsu_rdata_valid_o(lsu_rdata_valid),
.lsu_rdata_valid_o_t0(lsu_rdata_valid_t0),
.lsu_req_done_o(lsu_req_done),
.lsu_req_done_o_t0(lsu_req_done_t0),
.lsu_req_i(lsu_req),
.lsu_req_i_t0(lsu_req_t0),
.lsu_resp_valid_o(lsu_resp_valid),
.lsu_resp_valid_o_t0(lsu_resp_valid_t0),
.lsu_sign_ext_i(lsu_sign_ext),
.lsu_sign_ext_i_t0(lsu_sign_ext_t0),
.lsu_type_i(lsu_type),
.lsu_type_i_t0(lsu_type_t0),
.lsu_wdata_i(lsu_wdata),
.lsu_wdata_i_t0(lsu_wdata_t0),
.lsu_we_i(lsu_we),
.lsu_we_i_t0(lsu_we_t0),
.perf_load_o(perf_load),
.perf_load_o_t0(perf_load_t0),
.perf_store_o(perf_store),
.perf_store_o_t0(perf_store_t0),
.rst_ni(rst_ni),
.store_err_o(lsu_store_err_raw),
.store_err_o_t0(lsu_store_err_raw_t0),
.store_resp_intg_err_o(lsu_store_resp_intg_err),
.store_resp_intg_err_o_t0(lsu_store_resp_intg_err_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13363.4-13394.3" */
\$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'0\DummyInstructions=1'1  wb_stage_i (
.clk_i(clk_i),
.dummy_instr_id_i(dummy_instr_id_o),
.dummy_instr_id_i_t0(dummy_instr_id_o_t0),
.dummy_instr_wb_o(dummy_instr_wb_o),
.dummy_instr_wb_o_t0(dummy_instr_wb_o_t0),
.en_wb_i(en_wb),
.en_wb_i_t0(en_wb_t0),
.instr_done_wb_o(instr_done_wb),
.instr_done_wb_o_t0(instr_done_wb_t0),
.instr_is_compressed_id_i(instr_is_compressed_id),
.instr_is_compressed_id_i_t0(instr_is_compressed_id_t0),
.instr_perf_count_id_i(instr_perf_count_id),
.instr_perf_count_id_i_t0(instr_perf_count_id_t0),
.instr_type_wb_i(instr_type_wb),
.instr_type_wb_i_t0(instr_type_wb_t0),
.lsu_resp_err_i(lsu_resp_err),
.lsu_resp_err_i_t0(lsu_resp_err_t0),
.lsu_resp_valid_i(lsu_resp_valid),
.lsu_resp_valid_i_t0(lsu_resp_valid_t0),
.outstanding_load_wb_o(outstanding_load_wb),
.outstanding_load_wb_o_t0(outstanding_load_wb_t0),
.outstanding_store_wb_o(outstanding_store_wb),
.outstanding_store_wb_o_t0(outstanding_store_wb_t0),
.pc_id_i(pc_id),
.pc_id_i_t0(pc_id_t0),
.pc_wb_o(pc_wb),
.pc_wb_o_t0(pc_wb_t0),
.perf_instr_ret_compressed_wb_o(perf_instr_ret_compressed_wb),
.perf_instr_ret_compressed_wb_o_t0(perf_instr_ret_compressed_wb_t0),
.perf_instr_ret_compressed_wb_spec_o(perf_instr_ret_compressed_wb_spec),
.perf_instr_ret_compressed_wb_spec_o_t0(perf_instr_ret_compressed_wb_spec_t0),
.perf_instr_ret_wb_o(perf_instr_ret_wb),
.perf_instr_ret_wb_o_t0(perf_instr_ret_wb_t0),
.perf_instr_ret_wb_spec_o(perf_instr_ret_wb_spec),
.perf_instr_ret_wb_spec_o_t0(perf_instr_ret_wb_spec_t0),
.ready_wb_o(ready_wb),
.ready_wb_o_t0(ready_wb_t0),
.rf_waddr_id_i(rf_waddr_id),
.rf_waddr_id_i_t0(rf_waddr_id_t0),
.rf_waddr_wb_o(rf_waddr_wb_o),
.rf_waddr_wb_o_t0(rf_waddr_wb_o_t0),
.rf_wdata_fwd_wb_o(rf_wdata_fwd_wb),
.rf_wdata_fwd_wb_o_t0(rf_wdata_fwd_wb_t0),
.rf_wdata_id_i(rf_wdata_id),
.rf_wdata_id_i_t0(rf_wdata_id_t0),
.rf_wdata_lsu_i(rf_wdata_lsu),
.rf_wdata_lsu_i_t0(rf_wdata_lsu_t0),
.rf_wdata_wb_o(rf_wdata_wb),
.rf_wdata_wb_o_t0(rf_wdata_wb_t0),
.rf_we_id_i(rf_we_id),
.rf_we_id_i_t0(rf_we_id_t0),
.rf_we_lsu_i(rf_we_lsu),
.rf_we_lsu_i_t0(rf_we_lsu_t0),
.rf_we_wb_o(rf_we_wb_o),
.rf_we_wb_o_t0(rf_we_wb_o_t0),
.rf_write_wb_o(rf_write_wb),
.rf_write_wb_o_t0(rf_write_wb_t0),
.rst_ni(rst_ni)
);
assign core_busy_o_t0 = 4'h0;
assign crash_dump_o = { pc_id, pc_if, lsu_addr_last, csr_mepc, crash_dump_mtval };
assign crash_dump_o_t0 = { pc_id_t0, pc_if_t0, lsu_addr_last_t0, csr_mepc_t0, crash_dump_mtval_t0 };
endmodule

module \$paramod$5fd3ce2f8a67228d339c5f62898ff83b3c2a14f0\prim_lfsr (clk_i, rst_ni, seed_en_i, seed_i, lfsr_en_i, entropy_i, state_o, state_o_t0, seed_i_t0, seed_en_i_t0, lfsr_en_i_t0, entropy_i_t0);
wire _00_;
wire [31:0] _01_;
wire [31:0] _02_;
wire _03_;
wire [31:0] _04_;
wire [31:0] _05_;
wire [31:0] _06_;
wire [31:0] _07_;
wire [31:0] _08_;
/* src = "generated/sv2v_out.v:25506.41-25506.60" */
wire _09_;
/* src = "generated/sv2v_out.v:25488.22-25488.29" */
wire _10_;
/* src = "generated/sv2v_out.v:25506.83-25506.119" */
wire [31:0] _11_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25506.83-25506.119" */
wire [31:0] _12_;
/* src = "generated/sv2v_out.v:25506.41-25506.120" */
wire [31:0] _13_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25506.41-25506.120" */
wire [31:0] _14_;
/* src = "generated/sv2v_out.v:25487.30-25487.90" */
wire [31:0] _15_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25487.30-25487.90" */
wire [31:0] _16_;
/* src = "generated/sv2v_out.v:25454.8-25454.13" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:25459.26-25459.35" */
input [7:0] entropy_i;
wire [7:0] entropy_i;
/* cellift = 32'd1 */
input [7:0] entropy_i_t0;
wire [7:0] entropy_i_t0;
/* src = "generated/sv2v_out.v:25466.22-25466.28" */
wire [31:0] lfsr_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25466.22-25466.28" */
wire [31:0] lfsr_d_t0;
/* src = "generated/sv2v_out.v:25458.8-25458.17" */
input lfsr_en_i;
wire lfsr_en_i;
/* cellift = 32'd1 */
input lfsr_en_i_t0;
wire lfsr_en_i_t0;
/* src = "generated/sv2v_out.v:25467.21-25467.27" */
reg [31:0] lfsr_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25467.21-25467.27" */
reg [31:0] lfsr_q_t0;
/* src = "generated/sv2v_out.v:25465.7-25465.13" */
wire lockup;
/* src = "generated/sv2v_out.v:25468.22-25468.37" */
wire [31:0] next_lfsr_state;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25468.22-25468.37" */
wire [31:0] next_lfsr_state_t0;
/* src = "generated/sv2v_out.v:25455.8-25455.14" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:25456.8-25456.17" */
input seed_en_i;
wire seed_en_i;
/* cellift = 32'd1 */
input seed_en_i_t0;
wire seed_en_i_t0;
/* src = "generated/sv2v_out.v:25457.23-25457.29" */
input [31:0] seed_i;
wire [31:0] seed_i;
/* cellift = 32'd1 */
input [31:0] seed_i_t0;
wire [31:0] seed_i_t0;
/* src = "generated/sv2v_out.v:25460.33-25460.40" */
output [16:0] state_o;
wire [16:0] state_o;
/* cellift = 32'd1 */
output [16:0] state_o_t0;
wire [16:0] state_o_t0;
assign _00_ = ~ _03_;
assign _04_ = { _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_ } & lfsr_d_t0;
assign _05_ = { _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_ } & lfsr_q_t0;
assign _08_ = _04_ | _05_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$5fd3ce2f8a67228d339c5f62898ff83b3c2a14f0\prim_lfsr  */
/* PC_TAINT_INFO STATE_NAME lfsr_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) lfsr_q_t0 <= 32'd0;
else lfsr_q_t0 <= _08_;
/* src = "generated/sv2v_out.v:25585.2-25590.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$5fd3ce2f8a67228d339c5f62898ff83b3c2a14f0\prim_lfsr  */
/* PC_TAINT_INFO STATE_NAME lfsr_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) lfsr_q <= 32'd2891135988;
else if (_03_) lfsr_q <= lfsr_d;
assign _01_ = ~ { _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_ };
assign _02_ = ~ { seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i };
assign _14_ = _01_ & _12_;
assign _06_ = _02_ & _14_;
assign _12_ = { lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i } & next_lfsr_state_t0;
assign _07_ = { seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i } & seed_i_t0;
assign lfsr_d_t0 = _06_ | _07_;
assign _03_ = | { lfsr_en_i, seed_en_i, _09_ };
assign _16_ = { 24'h000000, entropy_i_t0 } | { lfsr_q_t0[0], 24'h000000, lfsr_q_t0[0], 1'h0, lfsr_q_t0[0], 1'h0, lfsr_q_t0[0], lfsr_q_t0[0], lfsr_q_t0[0] };
assign next_lfsr_state_t0 = _16_ | { 1'h0, lfsr_q_t0[31:1] };
assign _09_ = lfsr_en_i && /* src = "generated/sv2v_out.v:25506.41-25506.60" */ lockup;
assign lockup = ~ /* src = "generated/sv2v_out.v:25488.20-25488.30" */ _10_;
assign _10_ = | /* src = "generated/sv2v_out.v:25488.22-25488.29" */ lfsr_q;
assign _11_ = lfsr_en_i ? /* src = "generated/sv2v_out.v:25506.83-25506.119" */ next_lfsr_state : 32'hxxxxxxxx;
assign _13_ = _09_ ? /* src = "generated/sv2v_out.v:25506.41-25506.120" */ 32'd2891135988 : _11_;
assign lfsr_d = seed_en_i ? /* src = "generated/sv2v_out.v:25506.19-25506.121" */ seed_i : _13_;
assign _15_ = { 24'h000000, entropy_i } ^ /* src = "generated/sv2v_out.v:25487.30-25487.90" */ { lfsr_q[0], 24'h000000, lfsr_q[0], 1'h0, lfsr_q[0], 1'h0, lfsr_q[0], lfsr_q[0], lfsr_q[0] };
assign next_lfsr_state = _15_ ^ /* src = "generated/sv2v_out.v:25487.29-25487.107" */ { 1'h0, lfsr_q[31:1] };
assign state_o = { lfsr_q[21], lfsr_q[16], lfsr_q[5], lfsr_q[9], lfsr_q[12], lfsr_q[0], lfsr_q[19], lfsr_q[29], lfsr_q[4], lfsr_q[7], lfsr_q[1], lfsr_q[28], lfsr_q[10], lfsr_q[17], lfsr_q[22], lfsr_q[23], lfsr_q[13] };
assign state_o_t0 = { lfsr_q_t0[21], lfsr_q_t0[16], lfsr_q_t0[5], lfsr_q_t0[9], lfsr_q_t0[12], lfsr_q_t0[0], lfsr_q_t0[19], lfsr_q_t0[29], lfsr_q_t0[4], lfsr_q_t0[7], lfsr_q_t0[1], lfsr_q_t0[28], lfsr_q_t0[10], lfsr_q_t0[17], lfsr_q_t0[22], lfsr_q_t0[23], lfsr_q_t0[13] };
endmodule

module \$paramod$5ffe4cc9ba21eb548f33468a0c4a93d38de3dae5\ibex_decoder (clk_i, rst_ni, illegal_insn_o, ebrk_insn_o, mret_insn_o, dret_insn_o, ecall_insn_o, wfi_insn_o, jump_set_o, branch_taken_i, icache_inval_o, instr_first_cycle_i, instr_rdata_i, instr_rdata_alu_i, illegal_c_insn_i, imm_a_mux_sel_o, imm_b_mux_sel_o, bt_a_mux_sel_o, bt_b_mux_sel_o, imm_i_type_o, imm_s_type_o
, imm_b_type_o, imm_u_type_o, imm_j_type_o, zimm_rs1_type_o, rf_wdata_sel_o, rf_we_o, rf_raddr_a_o, rf_raddr_b_o, rf_waddr_o, rf_ren_a_o, rf_ren_b_o, alu_operator_o, alu_op_a_mux_sel_o, alu_op_b_mux_sel_o, alu_multicycle_o, mult_en_o, div_en_o, mult_sel_o, div_sel_o, multdiv_operator_o, multdiv_signed_mode_o
, csr_access_o, csr_op_o, data_req_o, data_we_o, data_type_o, data_sign_extension_o, jump_in_dec_o, branch_in_dec_o, instr_rdata_i_t0, zimm_rs1_type_o_t0, wfi_insn_o_t0, rf_we_o_t0, rf_wdata_sel_o_t0, rf_waddr_o_t0, rf_ren_b_o_t0, rf_ren_a_o_t0, rf_raddr_b_o_t0, rf_raddr_a_o_t0, multdiv_signed_mode_o_t0, multdiv_operator_o_t0, mult_sel_o_t0
, mult_en_o_t0, mret_insn_o_t0, jump_set_o_t0, jump_in_dec_o_t0, instr_rdata_alu_i_t0, instr_first_cycle_i_t0, imm_u_type_o_t0, imm_s_type_o_t0, imm_j_type_o_t0, imm_i_type_o_t0, imm_b_type_o_t0, imm_b_mux_sel_o_t0, imm_a_mux_sel_o_t0, illegal_insn_o_t0, illegal_c_insn_i_t0, icache_inval_o_t0, ecall_insn_o_t0, ebrk_insn_o_t0, dret_insn_o_t0, div_sel_o_t0, div_en_o_t0
, data_we_o_t0, data_type_o_t0, data_sign_extension_o_t0, data_req_o_t0, csr_op_o_t0, csr_access_o_t0, bt_b_mux_sel_o_t0, bt_a_mux_sel_o_t0, branch_taken_i_t0, branch_in_dec_o_t0, alu_operator_o_t0, alu_op_b_mux_sel_o_t0, alu_op_a_mux_sel_o_t0, alu_multicycle_o_t0);
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [6:0] _000_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [6:0] _001_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [6:0] _002_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _003_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [6:0] _004_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _005_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [6:0] _006_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _007_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _008_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _009_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _010_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _011_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _012_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _013_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _014_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _015_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _016_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _017_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _018_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _019_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _020_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire [1:0] _021_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire [1:0] _022_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire _023_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _024_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _025_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _026_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _027_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _028_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire _029_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [2:0] _030_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _031_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _032_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _033_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire _034_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire [1:0] _035_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire [1:0] _036_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _037_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _038_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _039_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [1:0] _040_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _041_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire [1:0] _042_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire _043_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _044_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _045_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _046_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _047_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [2:0] _048_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _049_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire _050_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire [1:0] _051_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire [1:0] _052_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _053_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _054_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [6:0] _055_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _056_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [2:0] _057_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [6:0] _058_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _059_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [2:0] _060_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [1:0] _061_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire _062_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _063_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [2:0] _064_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [6:0] _065_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [2:0] _066_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [1:0] _067_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _068_;
/* src = "generated/sv2v_out.v:15342.2-15793.5" */
wire [1:0] _069_;
/* src = "generated/sv2v_out.v:15090.2-15341.5" */
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire [1:0] _114_;
wire [6:0] _115_;
wire [6:0] _116_;
wire [6:0] _117_;
wire [6:0] _118_;
wire [6:0] _119_;
wire [6:0] _120_;
wire [6:0] _121_;
wire [6:0] _122_;
wire [6:0] _123_;
wire [6:0] _124_;
wire [6:0] _125_;
wire [6:0] _126_;
wire [6:0] _127_;
wire [6:0] _128_;
wire [6:0] _129_;
wire [6:0] _130_;
wire [6:0] _131_;
wire [6:0] _132_;
wire [6:0] _133_;
wire _134_;
wire _135_;
wire [1:0] _136_;
wire [1:0] _137_;
wire [1:0] _138_;
wire [1:0] _139_;
wire [6:0] _140_;
wire [6:0] _141_;
wire [6:0] _142_;
wire [6:0] _143_;
wire [2:0] _144_;
wire [2:0] _145_;
wire [2:0] _146_;
wire [2:0] _147_;
wire [2:0] _148_;
wire [1:0] _149_;
wire [1:0] _150_;
wire [1:0] _151_;
wire [1:0] _152_;
wire [1:0] _153_;
wire _154_;
wire [1:0] _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
/* src = "generated/sv2v_out.v:15087.9-15087.23" */
wire _170_;
/* src = "generated/sv2v_out.v:15087.29-15087.43" */
wire _171_;
/* src = "generated/sv2v_out.v:15087.50-15087.74" */
wire _172_;
/* src = "generated/sv2v_out.v:15185.34-15185.55" */
wire _173_;
/* src = "generated/sv2v_out.v:15237.9-15237.44" */
wire _174_;
/* src = "generated/sv2v_out.v:15302.9-15302.31" */
wire _175_;
/* src = "generated/sv2v_out.v:15547.16-15547.44" */
wire _176_;
/* src = "generated/sv2v_out.v:15549.16-15549.44" */
wire _177_;
/* src = "generated/sv2v_out.v:15777.9-15777.35" */
wire _178_;
/* src = "generated/sv2v_out.v:15087.7-15087.75" */
wire _179_;
/* src = "generated/sv2v_out.v:15087.8-15087.44" */
wire _180_;
/* src = "generated/sv2v_out.v:15311.10-15311.59" */
wire _181_;
/* src = "generated/sv2v_out.v:15133.9-15133.31" */
wire _182_;
/* src = "generated/sv2v_out.v:15311.11-15311.32" */
wire _183_;
/* src = "generated/sv2v_out.v:15311.38-15311.58" */
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire [9:0] _239_;
wire _240_;
wire _241_;
wire _242_;
wire [1:0] _243_;
wire _244_;
/* unused_bits = "1 2" */
wire [5:0] _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
/* src = "generated/sv2v_out.v:15185.34-15185.69" */
wire _255_;
/* src = "generated/sv2v_out.v:15013.13-15013.29" */
output alu_multicycle_o;
wire alu_multicycle_o;
/* cellift = 32'd1 */
output alu_multicycle_o_t0;
wire alu_multicycle_o_t0;
/* src = "generated/sv2v_out.v:15011.19-15011.37" */
output [1:0] alu_op_a_mux_sel_o;
wire [1:0] alu_op_a_mux_sel_o;
/* cellift = 32'd1 */
output [1:0] alu_op_a_mux_sel_o_t0;
wire [1:0] alu_op_a_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:15012.13-15012.31" */
output alu_op_b_mux_sel_o;
wire alu_op_b_mux_sel_o;
/* cellift = 32'd1 */
output alu_op_b_mux_sel_o_t0;
wire alu_op_b_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:15010.19-15010.33" */
output [6:0] alu_operator_o;
wire [6:0] alu_operator_o;
/* cellift = 32'd1 */
output [6:0] alu_operator_o_t0;
wire [6:0] alu_operator_o_t0;
/* src = "generated/sv2v_out.v:15027.13-15027.28" */
output branch_in_dec_o;
wire branch_in_dec_o;
/* cellift = 32'd1 */
output branch_in_dec_o_t0;
wire branch_in_dec_o_t0;
/* src = "generated/sv2v_out.v:14987.13-14987.27" */
input branch_taken_i;
wire branch_taken_i;
/* cellift = 32'd1 */
input branch_taken_i_t0;
wire branch_taken_i_t0;
/* src = "generated/sv2v_out.v:14995.19-14995.33" */
output [1:0] bt_a_mux_sel_o;
wire [1:0] bt_a_mux_sel_o;
/* cellift = 32'd1 */
output [1:0] bt_a_mux_sel_o_t0;
wire [1:0] bt_a_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:14996.19-14996.33" */
output [2:0] bt_b_mux_sel_o;
wire [2:0] bt_b_mux_sel_o;
/* cellift = 32'd1 */
output [2:0] bt_b_mux_sel_o_t0;
wire [2:0] bt_b_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:14978.13-14978.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:15020.13-15020.25" */
output csr_access_o;
wire csr_access_o;
/* cellift = 32'd1 */
output csr_access_o_t0;
wire csr_access_o_t0;
/* src = "generated/sv2v_out.v:15041.12-15041.18" */
wire [1:0] csr_op;
/* src = "generated/sv2v_out.v:15021.19-15021.27" */
output [1:0] csr_op_o;
wire [1:0] csr_op_o;
/* cellift = 32'd1 */
output [1:0] csr_op_o_t0;
wire [1:0] csr_op_o_t0;
/* src = "generated/sv2v_out.v:15022.13-15022.23" */
output data_req_o;
wire data_req_o;
/* cellift = 32'd1 */
output data_req_o_t0;
wire data_req_o_t0;
/* src = "generated/sv2v_out.v:15025.13-15025.34" */
output data_sign_extension_o;
wire data_sign_extension_o;
/* cellift = 32'd1 */
output data_sign_extension_o_t0;
wire data_sign_extension_o_t0;
/* src = "generated/sv2v_out.v:15024.19-15024.30" */
output [1:0] data_type_o;
wire [1:0] data_type_o;
/* cellift = 32'd1 */
output [1:0] data_type_o_t0;
wire [1:0] data_type_o_t0;
/* src = "generated/sv2v_out.v:15023.13-15023.22" */
output data_we_o;
wire data_we_o;
/* cellift = 32'd1 */
output data_we_o_t0;
wire data_we_o_t0;
/* src = "generated/sv2v_out.v:15015.14-15015.22" */
output div_en_o;
wire div_en_o;
/* cellift = 32'd1 */
output div_en_o_t0;
wire div_en_o_t0;
/* src = "generated/sv2v_out.v:15017.13-15017.22" */
output div_sel_o;
wire div_sel_o;
/* cellift = 32'd1 */
output div_sel_o_t0;
wire div_sel_o_t0;
/* src = "generated/sv2v_out.v:14983.13-14983.24" */
output dret_insn_o;
wire dret_insn_o;
/* cellift = 32'd1 */
output dret_insn_o_t0;
wire dret_insn_o_t0;
/* src = "generated/sv2v_out.v:14981.13-14981.24" */
output ebrk_insn_o;
wire ebrk_insn_o;
/* cellift = 32'd1 */
output ebrk_insn_o_t0;
wire ebrk_insn_o_t0;
/* src = "generated/sv2v_out.v:14984.13-14984.25" */
output ecall_insn_o;
wire ecall_insn_o;
/* cellift = 32'd1 */
output ecall_insn_o_t0;
wire ecall_insn_o_t0;
/* src = "generated/sv2v_out.v:14988.13-14988.27" */
output icache_inval_o;
wire icache_inval_o;
/* cellift = 32'd1 */
output icache_inval_o_t0;
wire icache_inval_o_t0;
/* src = "generated/sv2v_out.v:14992.13-14992.29" */
input illegal_c_insn_i;
wire illegal_c_insn_i;
/* cellift = 32'd1 */
input illegal_c_insn_i_t0;
wire illegal_c_insn_i_t0;
/* src = "generated/sv2v_out.v:14980.14-14980.28" */
output illegal_insn_o;
wire illegal_insn_o;
/* cellift = 32'd1 */
output illegal_insn_o_t0;
wire illegal_insn_o_t0;
/* src = "generated/sv2v_out.v:14993.13-14993.28" */
output imm_a_mux_sel_o;
wire imm_a_mux_sel_o;
/* cellift = 32'd1 */
output imm_a_mux_sel_o_t0;
wire imm_a_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:14994.19-14994.34" */
output [2:0] imm_b_mux_sel_o;
wire [2:0] imm_b_mux_sel_o;
/* cellift = 32'd1 */
output [2:0] imm_b_mux_sel_o_t0;
wire [2:0] imm_b_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:14999.21-14999.33" */
output [31:0] imm_b_type_o;
wire [31:0] imm_b_type_o;
/* cellift = 32'd1 */
output [31:0] imm_b_type_o_t0;
wire [31:0] imm_b_type_o_t0;
/* src = "generated/sv2v_out.v:14997.21-14997.33" */
output [31:0] imm_i_type_o;
wire [31:0] imm_i_type_o;
/* cellift = 32'd1 */
output [31:0] imm_i_type_o_t0;
wire [31:0] imm_i_type_o_t0;
/* src = "generated/sv2v_out.v:15001.21-15001.33" */
output [31:0] imm_j_type_o;
wire [31:0] imm_j_type_o;
/* cellift = 32'd1 */
output [31:0] imm_j_type_o_t0;
wire [31:0] imm_j_type_o_t0;
/* src = "generated/sv2v_out.v:14998.21-14998.33" */
output [31:0] imm_s_type_o;
wire [31:0] imm_s_type_o;
/* cellift = 32'd1 */
output [31:0] imm_s_type_o_t0;
wire [31:0] imm_s_type_o_t0;
/* src = "generated/sv2v_out.v:15000.21-15000.33" */
output [31:0] imm_u_type_o;
wire [31:0] imm_u_type_o;
/* cellift = 32'd1 */
output [31:0] imm_u_type_o_t0;
wire [31:0] imm_u_type_o_t0;
/* src = "generated/sv2v_out.v:14989.13-14989.32" */
input instr_first_cycle_i;
wire instr_first_cycle_i;
/* cellift = 32'd1 */
input instr_first_cycle_i_t0;
wire instr_first_cycle_i_t0;
/* src = "generated/sv2v_out.v:14991.20-14991.37" */
input [31:0] instr_rdata_alu_i;
wire [31:0] instr_rdata_alu_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_alu_i_t0;
wire [31:0] instr_rdata_alu_i_t0;
/* src = "generated/sv2v_out.v:14990.20-14990.33" */
input [31:0] instr_rdata_i;
wire [31:0] instr_rdata_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_i_t0;
wire [31:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:15026.13-15026.26" */
output jump_in_dec_o;
wire jump_in_dec_o;
/* cellift = 32'd1 */
output jump_in_dec_o_t0;
wire jump_in_dec_o_t0;
/* src = "generated/sv2v_out.v:14986.13-14986.23" */
output jump_set_o;
wire jump_set_o;
/* cellift = 32'd1 */
output jump_set_o_t0;
wire jump_set_o_t0;
/* src = "generated/sv2v_out.v:14982.13-14982.24" */
output mret_insn_o;
wire mret_insn_o;
/* cellift = 32'd1 */
output mret_insn_o_t0;
wire mret_insn_o_t0;
/* src = "generated/sv2v_out.v:15014.14-15014.23" */
output mult_en_o;
wire mult_en_o;
/* cellift = 32'd1 */
output mult_en_o_t0;
wire mult_en_o_t0;
/* src = "generated/sv2v_out.v:15016.13-15016.23" */
output mult_sel_o;
wire mult_sel_o;
/* cellift = 32'd1 */
output mult_sel_o_t0;
wire mult_sel_o_t0;
/* src = "generated/sv2v_out.v:15018.19-15018.37" */
output [1:0] multdiv_operator_o;
wire [1:0] multdiv_operator_o;
/* cellift = 32'd1 */
output [1:0] multdiv_operator_o_t0;
wire [1:0] multdiv_operator_o_t0;
/* src = "generated/sv2v_out.v:15019.19-15019.40" */
output [1:0] multdiv_signed_mode_o;
wire [1:0] multdiv_signed_mode_o;
/* cellift = 32'd1 */
output [1:0] multdiv_signed_mode_o_t0;
wire [1:0] multdiv_signed_mode_o_t0;
/* src = "generated/sv2v_out.v:15005.20-15005.32" */
output [4:0] rf_raddr_a_o;
wire [4:0] rf_raddr_a_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_a_o_t0;
wire [4:0] rf_raddr_a_o_t0;
/* src = "generated/sv2v_out.v:15006.20-15006.32" */
output [4:0] rf_raddr_b_o;
wire [4:0] rf_raddr_b_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_b_o_t0;
wire [4:0] rf_raddr_b_o_t0;
/* src = "generated/sv2v_out.v:15008.13-15008.23" */
output rf_ren_a_o;
wire rf_ren_a_o;
/* cellift = 32'd1 */
output rf_ren_a_o_t0;
wire rf_ren_a_o_t0;
/* src = "generated/sv2v_out.v:15009.13-15009.23" */
output rf_ren_b_o;
wire rf_ren_b_o;
/* cellift = 32'd1 */
output rf_ren_b_o_t0;
wire rf_ren_b_o_t0;
/* src = "generated/sv2v_out.v:15007.20-15007.30" */
output [4:0] rf_waddr_o;
wire [4:0] rf_waddr_o;
/* cellift = 32'd1 */
output [4:0] rf_waddr_o_t0;
wire [4:0] rf_waddr_o_t0;
/* src = "generated/sv2v_out.v:15003.13-15003.27" */
output rf_wdata_sel_o;
wire rf_wdata_sel_o;
/* cellift = 32'd1 */
output rf_wdata_sel_o_t0;
wire rf_wdata_sel_o_t0;
/* src = "generated/sv2v_out.v:15004.14-15004.21" */
output rf_we_o;
wire rf_we_o;
/* cellift = 32'd1 */
output rf_we_o_t0;
wire rf_we_o_t0;
/* src = "generated/sv2v_out.v:14979.13-14979.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14985.13-14985.23" */
output wfi_insn_o;
wire wfi_insn_o;
/* cellift = 32'd1 */
output wfi_insn_o_t0;
wire wfi_insn_o_t0;
/* src = "generated/sv2v_out.v:15002.21-15002.36" */
output [31:0] zimm_rs1_type_o;
wire [31:0] zimm_rs1_type_o;
/* cellift = 32'd1 */
output [31:0] zimm_rs1_type_o_t0;
wire [31:0] zimm_rs1_type_o_t0;
assign _071_ = ~ instr_rdata_i[14];
assign data_sign_extension_o_t0 = _246_ & instr_rdata_i_t0[14];
assign _083_ = | { _229_, _175_ };
assign _084_ = | { _217_, _216_ };
assign _085_ = | { _250_, _248_, _240_ };
assign _086_ = | { _228_, _227_, _226_, _225_, _224_ };
assign _087_ = | { _254_, _253_, _242_, _240_ };
assign _089_ = | { _251_, _250_, _248_, _246_, _242_, _240_ };
assign _090_ = | { _195_, _194_, _193_, _192_ };
assign _091_ = | { _191_, _190_, _189_, _188_ };
assign _092_ = | { _232_, _231_ };
assign _093_ = | { _234_, _233_ };
assign _094_ = | { _237_, _236_, _235_ };
assign _095_ = | { _204_, _195_, _194_, _193_, _192_, _191_, _190_, _189_, _188_ };
assign _096_ = | { _237_, _234_, _232_ };
assign _097_ = | { _219_, _217_ };
assign _098_ = | { _219_, _218_, _217_, _216_, _215_, _213_ };
assign _100_ = | { _239_, _238_, _237_, _236_, _235_, _234_, _233_, _232_, _231_ };
assign _101_ = | { _215_, _214_ };
assign _088_ = | { _252_, _251_ };
assign _099_ = | { _248_, _246_ };
assign _072_ = | { _186_, _178_ };
assign _073_ = | { _222_, _221_, _220_ };
assign _074_ = | { _247_, _222_ };
assign _075_ = | { _247_, _222_, _221_ };
assign _102_ = _196_ | _095_;
assign _103_ = _201_ | _200_;
assign _104_ = _186_ | _206_;
assign _105_ = _211_ | _210_;
assign _106_ = _186_ | _210_;
assign _107_ = _213_ | _205_;
assign _108_ = _215_ | _214_;
assign _109_ = _221_ | _220_;
assign _110_ = _093_ | _092_;
assign _111_ = _087_ | _223_;
assign _112_ = _230_ | _223_;
assign _113_ = _248_ | _246_;
assign _076_ = | { _199_, _198_, _197_, _102_ };
assign _077_ = | { _209_, _208_, _104_ };
assign _078_ = | { _209_, _208_, _206_ };
assign _079_ = | { _218_, _213_, _207_, _205_, _187_, _185_ };
assign _080_ = | { _207_, _205_, _187_ };
assign _081_ = | { _219_, _217_, _213_, _187_ };
assign _082_ = | { _112_, _254_, _253_, _252_, _242_, _240_ };
assign _114_ = _178_ ? 2'h0 : 2'h3;
assign _061_ = _186_ ? 2'h2 : _114_;
assign _115_ = _095_ ? 7'h00 : 7'h08;
assign _116_ = _198_ ? 7'h0a : 7'h04;
assign _117_ = _197_ ? 7'h09 : _116_;
assign _118_ = _102_ ? _115_ : _117_;
assign _119_ = _200_ ? 7'h03 : 7'h02;
assign _120_ = _203_ ? 7'h01 : 7'h2c;
assign _121_ = _202_ ? 7'h2b : _120_;
assign _122_ = _103_ ? _119_ : _121_;
assign _004_ = _076_ ? _118_ : _122_;
assign _123_ = _206_ ? _000_ : 7'h0a;
assign _124_ = _208_ ? 7'h04 : 7'h03;
assign _125_ = _104_ ? _123_ : _124_;
assign _126_ = _210_ ? 7'h02 : 7'h2c;
assign _127_ = _212_ ? 7'h2b : 7'h00;
assign _128_ = _105_ ? _126_ : _127_;
assign _065_ = _077_ ? _125_ : _128_;
assign _129_ = _209_ ? 7'h1a : 7'h1b;
assign _130_ = _208_ ? 7'h1c : _129_;
assign _131_ = _210_ ? 7'h19 : 7'h1e;
assign _132_ = _178_ ? 7'h1d : 7'h2c;
assign _133_ = _106_ ? _131_ : _132_;
assign _055_ = _078_ ? _130_ : _133_;
assign _134_ = _205_ ? 1'h0 : _062_;
assign _135_ = _214_ ? _038_ : 1'h1;
assign alu_op_b_mux_sel_o = _107_ ? _134_ : _135_;
assign _136_ = _187_ ? _061_ : 2'h0;
assign _137_ = _185_ ? _067_ : _136_;
assign _138_ = _101_ ? _040_ : 2'h3;
assign _139_ = _084_ ? 2'h2 : _138_;
assign alu_op_a_mux_sel_o = _079_ ? _137_ : _139_;
assign _140_ = _205_ ? _002_ : _065_;
assign _141_ = _187_ ? _006_ : _140_;
assign _142_ = _214_ ? _058_ : 7'h2c;
assign _143_ = _098_ ? 7'h00 : _142_;
assign alu_operator_o = _080_ ? _141_ : _143_;
assign _144_ = _097_ ? 3'h3 : _064_;
assign _145_ = _187_ ? _066_ : _144_;
assign _146_ = _214_ ? _057_ : _048_;
assign _147_ = _216_ ? _030_ : 3'h0;
assign _148_ = _108_ ? _146_ : _147_;
assign imm_b_mux_sel_o = _081_ ? _145_ : _148_;
assign _149_ = _220_ ? 2'h3 : 2'h2;
assign _150_ = _222_ ? 2'h1 : 2'h0;
assign _042_ = _109_ ? _149_ : _150_;
assign _151_ = _236_ ? 2'h1 : 2'h0;
assign _052_ = _096_ ? 2'h3 : _151_;
assign _152_ = _092_ ? 2'h3 : 2'h2;
assign _153_ = _094_ ? 2'h1 : 2'h0;
assign _051_ = _110_ ? _152_ : _153_;
assign _154_ = _229_ ? _070_ : 1'h0;
assign _068_ = _241_ ? _003_ : _154_;
assign _155_ = _247_ ? 2'h2 : 2'h0;
assign _022_ = _222_ ? 2'h1 : _155_;
assign _156_ = _074_ ? 1'h0 : 1'h1;
assign _063_ = _221_ ? _056_ : _156_;
assign _157_ = _223_ ? _020_ : 1'h1;
assign _158_ = _088_ ? _038_ : 1'h0;
assign _014_ = _111_ ? _157_ : _158_;
assign _159_ = _088_ ? _032_ : 1'h0;
assign _013_ = _230_ ? _027_ : _159_;
assign _160_ = _088_ ? 1'h1 : 1'h0;
assign _012_ = _230_ ? _031_ : _160_;
assign _161_ = _223_ ? _017_ : _016_;
assign _162_ = _242_ ? _068_ : 1'h0;
assign _163_ = _240_ ? _007_ : _162_;
assign _164_ = _112_ ? _161_ : _163_;
assign _165_ = _246_ ? _063_ : _059_;
assign _166_ = _251_ ? _028_ : 1'h1;
assign _167_ = _250_ ? _047_ : _166_;
assign _168_ = _113_ ? _165_ : _167_;
assign _011_ = _082_ ? _164_ : _168_;
assign _169_ = _089_ ? 1'h1 : 1'h0;
assign rf_ren_a_o = _223_ ? _037_ : _169_;
assign _170_ = csr_op == /* src = "generated/sv2v_out.v:15087.9-15087.23" */ 2'h2;
assign _171_ = csr_op == /* src = "generated/sv2v_out.v:15087.29-15087.43" */ 2'h3;
assign _172_ = ! /* src = "generated/sv2v_out.v:15087.50-15087.74" */ instr_rdata_i[19:15];
assign _174_ = { instr_rdata_i[26], instr_rdata_i[13:12] } == /* src = "generated/sv2v_out.v:15237.9-15237.44" */ 3'h5;
assign _176_ = ! /* src = "generated/sv2v_out.v:15547.16-15547.44" */ instr_rdata_alu_i[31:27];
assign _177_ = instr_rdata_alu_i[31:27] == /* src = "generated/sv2v_out.v:15549.16-15549.44" */ 5'h08;
assign _179_ = _180_ && /* src = "generated/sv2v_out.v:15087.7-15087.75" */ _172_;
assign _180_ = _170_ || /* src = "generated/sv2v_out.v:15087.8-15087.44" */ _171_;
assign _181_ = _183_ || /* src = "generated/sv2v_out.v:15311.10-15311.59" */ _184_;
assign _182_ = | /* src = "generated/sv2v_out.v:15133.9-15133.31" */ instr_rdata_i[14:12];
assign _183_ = | /* src = "generated/sv2v_out.v:15311.11-15311.32" */ instr_rdata_i[19:15];
assign _184_ = | /* src = "generated/sv2v_out.v:15311.38-15311.58" */ instr_rdata_i[11:7];
assign _069_ = instr_rdata_alu_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15785.10-15785.23|generated/sv2v_out.v:15785.6-15788.33" */ 2'h3 : 2'h0;
assign _067_ = _178_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15777.9-15777.35|generated/sv2v_out.v:15777.5-15789.8" */ 2'h0 : _069_;
assign _029_ = _178_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15777.9-15777.35|generated/sv2v_out.v:15777.5-15789.8" */ 1'h1 : 1'h0;
assign _006_ = _072_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15756.5-15775.12" */ 7'h00 : 7'h2c;
assign _066_ = _186_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15756.5-15775.12" */ 3'h5 : 3'h0;
assign _196_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 10'h105;
assign _197_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 10'h005;
assign _198_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 10'h001;
assign _199_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 10'h007;
assign _200_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 10'h006;
assign _201_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 10'h004;
assign _202_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 10'h002;
assign _203_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 10'h100;
assign _204_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] };
assign _043_ = _091_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 1'h1 : 1'h0;
assign _188_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 10'h00f;
assign _189_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 10'h00e;
assign _190_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 10'h00d;
assign _191_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 10'h00c;
assign _050_ = _090_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 1'h1 : 1'h0;
assign _192_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 10'h00b;
assign _193_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 10'h00a;
assign _194_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 10'h009;
assign _195_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15598.6-15753.13" */ 10'h008;
assign _023_ = instr_rdata_alu_i[26] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15558.9-15558.22|generated/sv2v_out.v:15558.5-15753.13" */ 1'h0 : _043_;
assign _034_ = instr_rdata_alu_i[26] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15558.9-15558.22|generated/sv2v_out.v:15558.5-15753.13" */ 1'h0 : _050_;
assign _002_ = instr_rdata_alu_i[26] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15558.9-15558.22|generated/sv2v_out.v:15558.5-15753.13" */ 7'h2c : _004_;
assign _001_ = _177_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15549.16-15549.44|generated/sv2v_out.v:15549.12-15550.30" */ 7'h08 : 7'h2c;
assign _000_ = _176_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15547.16-15547.44|generated/sv2v_out.v:15547.12-15550.30" */ 7'h09 : _001_;
assign _211_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15450.5-15553.12" */ 3'h3;
assign _212_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15450.5-15553.12" */ 3'h2;
assign _062_ = instr_rdata_alu_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15422.9-15422.23|generated/sv2v_out.v:15422.5-15425.8" */ 1'h0 : 1'h1;
assign _064_ = instr_rdata_alu_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15422.9-15422.23|generated/sv2v_out.v:15422.5-15425.8" */ 3'h0 : 3'h1;
assign _038_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15407.9-15407.28|generated/sv2v_out.v:15407.5-15416.8" */ 1'h0 : 1'h1;
assign _058_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15407.9-15407.28|generated/sv2v_out.v:15407.5-15416.8" */ _055_ : 7'h00;
assign _057_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15407.9-15407.28|generated/sv2v_out.v:15407.5-15416.8" */ 3'h0 : _060_;
assign _208_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15393.5-15402.12" */ 3'h7;
assign _209_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15393.5-15402.12" */ 3'h6;
assign _206_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15393.5-15402.12" */ 3'h5;
assign _210_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15393.5-15402.12" */ 3'h4;
assign _186_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15393.5-15402.12" */ 3'h1;
assign _178_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15393.5-15402.12" */ instr_rdata_alu_i[14:12];
assign _048_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15379.9-15379.48|generated/sv2v_out.v:15379.5-15390.8" */ 3'h0 : 3'h5;
assign _040_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15379.9-15379.48|generated/sv2v_out.v:15379.5-15390.8" */ 2'h0 : 2'h2;
assign _030_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15361.9-15361.48|generated/sv2v_out.v:15361.5-15372.8" */ 3'h4 : 3'h5;
assign _207_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15355.3-15792.10" */ 7'h13;
assign _218_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15355.3-15792.10" */ 7'h03;
assign _187_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15355.3-15792.10" */ 7'h0f;
assign _217_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15355.3-15792.10" */ 7'h17;
assign _219_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15355.3-15792.10" */ 7'h37;
assign _213_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15355.3-15792.10" */ 7'h23;
assign _214_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15355.3-15792.10" */ 7'h63;
assign _215_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15355.3-15792.10" */ 7'h67;
assign _216_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15355.3-15792.10" */ 7'h6f;
assign div_sel_o = _205_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15355.3-15792.10" */ _023_ : 1'h0;
assign mult_sel_o = _205_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15355.3-15792.10" */ _034_ : 1'h0;
assign _205_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15355.3-15792.10" */ 7'h33;
assign imm_a_mux_sel_o = _185_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15355.3-15792.10" */ _029_ : 1'h1;
assign _185_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15355.3-15792.10" */ 7'h73;
assign csr_access_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15332.7-15332.19|generated/sv2v_out.v:15332.3-15340.6" */ 1'h0 : rf_wdata_sel_o;
assign branch_in_dec_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15332.7-15332.19|generated/sv2v_out.v:15332.3-15340.6" */ 1'h0 : _008_;
assign jump_set_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15332.7-15332.19|generated/sv2v_out.v:15332.3-15340.6" */ 1'h0 : _013_;
assign jump_in_dec_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15332.7-15332.19|generated/sv2v_out.v:15332.3-15340.6" */ 1'h0 : _012_;
assign data_we_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15332.7-15332.19|generated/sv2v_out.v:15332.3-15340.6" */ 1'h0 : _010_;
assign data_req_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15332.7-15332.19|generated/sv2v_out.v:15332.3-15340.6" */ 1'h0 : _009_;
assign rf_we_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15332.7-15332.19|generated/sv2v_out.v:15332.3-15340.6" */ 1'h0 : _014_;
assign illegal_insn_o = illegal_c_insn_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15330.7-15330.23|generated/sv2v_out.v:15330.3-15331.24" */ 1'h1 : _011_;
assign _041_ = _073_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15320.6-15325.13" */ 1'h0 : 1'h1;
assign _220_ = instr_rdata_i[13:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15320.6-15325.13" */ 2'h3;
assign _053_ = instr_rdata_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15318.10-15318.20|generated/sv2v_out.v:15318.6-15319.25" */ 1'h0 : 1'h1;
assign _019_ = _181_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15311.10-15311.59|generated/sv2v_out.v:15311.6-15312.27" */ 1'h1 : _018_;
assign _046_ = _224_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15303.6-15310.13" */ 1'h1 : 1'h0;
assign _018_ = _086_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15303.6-15310.13" */ 1'h0 : 1'h1;
assign _224_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15303.6-15310.13" */ instr_rdata_i[31:20];
assign _054_ = _225_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15303.6-15310.13" */ 1'h1 : 1'h0;
assign _225_ = instr_rdata_i[31:20] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15303.6-15310.13" */ 12'h105;
assign _044_ = _226_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15303.6-15310.13" */ 1'h1 : 1'h0;
assign _226_ = instr_rdata_i[31:20] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15303.6-15310.13" */ 12'h7b2;
assign _049_ = _227_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15303.6-15310.13" */ 1'h1 : 1'h0;
assign _227_ = instr_rdata_i[31:20] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15303.6-15310.13" */ 12'h302;
assign _045_ = _228_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15303.6-15310.13" */ 1'h1 : 1'h0;
assign _228_ = instr_rdata_i[31:20] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15303.6-15310.13" */ 12'h001;
assign _017_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15302.9-15302.31|generated/sv2v_out.v:15302.5-15327.8" */ _019_ : _041_;
assign _039_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15302.9-15302.31|generated/sv2v_out.v:15302.5-15327.8" */ _054_ : 1'h0;
assign _026_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15302.9-15302.31|generated/sv2v_out.v:15302.5-15327.8" */ _046_ : 1'h0;
assign _024_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15302.9-15302.31|generated/sv2v_out.v:15302.5-15327.8" */ _044_ : 1'h0;
assign _033_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15302.9-15302.31|generated/sv2v_out.v:15302.5-15327.8" */ _049_ : 1'h0;
assign _025_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15302.9-15302.31|generated/sv2v_out.v:15302.5-15327.8" */ _045_ : 1'h0;
assign _037_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15302.9-15302.31|generated/sv2v_out.v:15302.5-15327.8" */ 1'h0 : _053_;
assign _020_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15302.9-15302.31|generated/sv2v_out.v:15302.5-15327.8" */ 1'h0 : 1'h1;
assign _021_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15302.9-15302.31|generated/sv2v_out.v:15302.5-15327.8" */ 2'h0 : _042_;
assign _016_ = _083_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15289.5-15300.12" */ 1'h0 : 1'h1;
assign _031_ = _229_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15289.5-15300.12" */ 1'h1 : 1'h0;
assign _027_ = _229_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15289.5-15300.12" */ _032_ : 1'h0;
assign _015_ = _100_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 1'h0 : 1'h1;
assign _238_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h008;
assign _239_[0] = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ { instr_rdata_i[31:25], instr_rdata_i[14:12] };
assign _239_[1] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h100;
assign _239_[2] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h002;
assign _239_[3] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h003;
assign _239_[4] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h004;
assign _239_[5] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h006;
assign _239_[6] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h007;
assign _239_[7] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h001;
assign _239_[8] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h005;
assign _239_[9] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h105;
assign _231_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h00f;
assign _232_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h00e;
assign _233_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h00d;
assign _234_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h00c;
assign _235_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h00b;
assign _236_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h00a;
assign _237_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15240.6-15286.13" */ 10'h009;
assign _007_ = _174_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15237.9-15237.44|generated/sv2v_out.v:15237.5-15286.13" */ 1'h1 : _015_;
assign _036_ = _174_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15237.9-15237.44|generated/sv2v_out.v:15237.5-15286.13" */ 2'h0 : _052_;
assign _035_ = _174_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15237.9-15237.44|generated/sv2v_out.v:15237.5-15286.13" */ 2'h0 : _051_;
assign _005_ = _244_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15205.8-15229.15" */ _255_ : 1'h1;
assign _244_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15205.8-15229.15" */ _243_;
assign _243_[1] = instr_rdata_i[31:27] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15205.8-15229.15" */ 5'h08;
assign _003_ = instr_rdata_i[26] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15202.11-15202.20|generated/sv2v_out.v:15202.7-15229.15" */ 1'h1 : _005_;
assign _173_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15194.9-15198.16" */ instr_rdata_i[26:25];
assign _070_ = _243_[0] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15184.7-15200.14" */ _255_ : 1'h1;
assign _243_[0] = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15184.7-15200.14" */ instr_rdata_i[31:27];
assign _056_ = instr_rdata_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15170.11-15170.20|generated/sv2v_out.v:15170.7-15171.28" */ 1'h1 : 1'h0;
assign _059_ = _075_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15153.5-15158.12" */ _056_ : 1'h1;
assign _221_ = instr_rdata_i[13:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15153.5-15158.12" */ 2'h2;
assign _222_ = instr_rdata_i[13:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15153.5-15158.12" */ 2'h1;
assign _247_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15153.5-15158.12" */ instr_rdata_i[13:12];
assign _047_ = _249_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15139.5-15142.12" */ 1'h0 : 1'h1;
assign _249_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15139.5-15142.12" */ { _245_[5:3], _241_, _229_, _175_ };
assign _175_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15139.5-15142.12" */ instr_rdata_i[14:12];
assign _229_ = instr_rdata_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15139.5-15142.12" */ 3'h1;
assign _245_[3] = instr_rdata_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15139.5-15142.12" */ 3'h4;
assign _241_ = instr_rdata_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15139.5-15142.12" */ 3'h5;
assign _245_[4] = instr_rdata_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15139.5-15142.12" */ 3'h6;
assign _245_[5] = instr_rdata_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15139.5-15142.12" */ 3'h7;
assign _028_ = _182_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15133.9-15133.31|generated/sv2v_out.v:15133.5-15134.26" */ 1'h1 : 1'h0;
assign _032_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15127.9-15127.28|generated/sv2v_out.v:15127.5-15132.19" */ 1'h1 : 1'h0;
assign _253_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ 7'h17;
assign _254_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ 7'h37;
assign _252_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ 7'h6f;
assign _008_ = _250_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ 1'h1 : 1'h0;
assign data_sign_extension_o = _246_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ _071_ : 1'h0;
assign data_type_o = _099_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ _022_ : 2'h0;
assign multdiv_signed_mode_o = _240_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ _036_ : 2'h0;
assign multdiv_operator_o = _240_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ _035_ : 2'h0;
assign rf_wdata_sel_o = _223_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ _020_ : 1'h0;
assign wfi_insn_o = _223_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ _039_ : 1'h0;
assign ecall_insn_o = _223_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ _026_ : 1'h0;
assign dret_insn_o = _223_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ _024_ : 1'h0;
assign mret_insn_o = _223_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ _033_ : 1'h0;
assign ebrk_insn_o = _223_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ _025_ : 1'h0;
assign rf_ren_b_o = _085_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ 1'h1 : 1'h0;
assign _240_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ 7'h33;
assign _242_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ 7'h13;
assign _246_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ 7'h03;
assign _248_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ 7'h23;
assign _250_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ 7'h63;
assign _251_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ 7'h67;
assign icache_inval_o = _230_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ _027_ : 1'h0;
assign _230_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ 7'h0f;
assign csr_op = _223_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ _021_ : 2'h0;
assign _223_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ 7'h73;
assign _010_ = _248_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ 1'h1 : 1'h0;
assign _009_ = _099_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15115.3-15329.10" */ 1'h1 : 1'h0;
assign csr_op_o = _179_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15087.7-15087.75|generated/sv2v_out.v:15087.3-15088.20" */ 2'h0 : csr_op;
assign _255_ = _173_ ? /* src = "generated/sv2v_out.v:15206.45-15206.80" */ 1'h0 : 1'h1;
assign _060_ = branch_taken_i ? /* src = "generated/sv2v_out.v:15414.25-15414.53" */ 3'h2 : 3'h5;
assign mult_en_o = illegal_insn_o ? /* src = "generated/sv2v_out.v:15794.22-15794.54" */ 1'h0 : mult_sel_o;
assign div_en_o = illegal_insn_o ? /* src = "generated/sv2v_out.v:15795.21-15795.52" */ 1'h0 : div_sel_o;
assign _245_[0] = _175_;
assign alu_multicycle_o = 1'h0;
assign alu_multicycle_o_t0 = 1'h0;
assign alu_op_a_mux_sel_o_t0 = 2'h0;
assign alu_op_b_mux_sel_o_t0 = 1'h0;
assign alu_operator_o_t0 = 7'h00;
assign branch_in_dec_o_t0 = 1'h0;
assign bt_a_mux_sel_o = 2'h2;
assign bt_a_mux_sel_o_t0 = 2'h0;
assign bt_b_mux_sel_o = 3'h0;
assign bt_b_mux_sel_o_t0 = 3'h0;
assign csr_access_o_t0 = 1'h0;
assign csr_op_o_t0 = 2'h0;
assign data_req_o_t0 = 1'h0;
assign data_type_o_t0 = 2'h0;
assign data_we_o_t0 = 1'h0;
assign div_en_o_t0 = 1'h0;
assign div_sel_o_t0 = 1'h0;
assign dret_insn_o_t0 = 1'h0;
assign ebrk_insn_o_t0 = 1'h0;
assign ecall_insn_o_t0 = 1'h0;
assign icache_inval_o_t0 = 1'h0;
assign illegal_insn_o_t0 = 1'h0;
assign imm_a_mux_sel_o_t0 = 1'h0;
assign imm_b_mux_sel_o_t0 = 3'h0;
assign imm_b_type_o = { instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[7], instr_rdata_i[30:25], instr_rdata_i[11:8], 1'h0 };
assign imm_b_type_o_t0 = { instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[7], instr_rdata_i_t0[30:25], instr_rdata_i_t0[11:8], 1'h0 };
assign imm_i_type_o = { instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31:20] };
assign imm_i_type_o_t0 = { instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31:20] };
assign imm_j_type_o = { instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[19:12], instr_rdata_i[20], instr_rdata_i[30:21], 1'h0 };
assign imm_j_type_o_t0 = { instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[19:12], instr_rdata_i_t0[20], instr_rdata_i_t0[30:21], 1'h0 };
assign imm_s_type_o = { instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31:25], instr_rdata_i[11:7] };
assign imm_s_type_o_t0 = { instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31:25], instr_rdata_i_t0[11:7] };
assign imm_u_type_o = { instr_rdata_i[31:12], 12'h000 };
assign imm_u_type_o_t0 = { instr_rdata_i_t0[31:12], 12'h000 };
assign jump_in_dec_o_t0 = 1'h0;
assign jump_set_o_t0 = 1'h0;
assign mret_insn_o_t0 = 1'h0;
assign mult_en_o_t0 = 1'h0;
assign mult_sel_o_t0 = 1'h0;
assign multdiv_operator_o_t0 = 2'h0;
assign multdiv_signed_mode_o_t0 = 2'h0;
assign rf_raddr_a_o = instr_rdata_i[19:15];
assign rf_raddr_a_o_t0 = instr_rdata_i_t0[19:15];
assign rf_raddr_b_o = instr_rdata_i[24:20];
assign rf_raddr_b_o_t0 = instr_rdata_i_t0[24:20];
assign rf_ren_a_o_t0 = 1'h0;
assign rf_ren_b_o_t0 = 1'h0;
assign rf_waddr_o = instr_rdata_i[11:7];
assign rf_waddr_o_t0 = instr_rdata_i_t0[11:7];
assign rf_wdata_sel_o_t0 = 1'h0;
assign rf_we_o_t0 = 1'h0;
assign wfi_insn_o_t0 = 1'h0;
assign zimm_rs1_type_o = { 27'h0000000, instr_rdata_i[19:15] };
assign zimm_rs1_type_o_t0 = { 27'h0000000, instr_rdata_i_t0[19:15] };
endmodule

module \$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _0_;
wire [31:0] _1_;
wire [31:0] _2_;
wire [31:0] _3_;
/* src = "generated/sv2v_out.v:14894.13-14894.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14898.28-14898.37" */
output [31:0] rd_data_o;
reg [31:0] rd_data_o;
/* cellift = 32'd1 */
output [31:0] rd_data_o_t0;
reg [31:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14899.14-14899.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14895.13-14895.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14896.27-14896.36" */
input [31:0] wr_data_i;
wire [31:0] wr_data_i;
/* cellift = 32'd1 */
input [31:0] wr_data_i_t0;
wire [31:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14897.13-14897.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _0_ = ~ wr_en_i;
assign _1_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _2_ = { _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_ } & rd_data_o_t0;
assign _3_ = _1_ | _2_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 32'd0;
else rd_data_o_t0 <= _3_;
/* src = "generated/sv2v_out.v:14901.2-14905.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 32'd0;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage (clk_i, rst_ni, boot_addr_i, req_i, instr_req_o, instr_addr_o, instr_gnt_i, instr_rvalid_i, instr_rdata_i, instr_bus_err_i, instr_intg_err_o, ic_tag_req_o, ic_tag_write_o, ic_tag_addr_o, ic_tag_wdata_o, ic_tag_rdata_i, ic_data_req_o, ic_data_write_o, ic_data_addr_o, ic_data_wdata_o, ic_data_rdata_i
, ic_scr_key_valid_i, ic_scr_key_req_o, instr_valid_id_o, instr_new_id_o, instr_rdata_id_o, instr_rdata_alu_id_o, instr_rdata_c_id_o, instr_is_compressed_id_o, instr_bp_taken_o, instr_fetch_err_o, instr_fetch_err_plus2_o, illegal_c_insn_id_o, dummy_instr_id_o, pc_if_o, pc_id_o, pmp_err_if_i, pmp_err_if_plus2_i, instr_valid_clear_i, pc_set_i, pc_mux_i, nt_branch_mispredict_i
, nt_branch_addr_i, exc_pc_mux_i, exc_cause, dummy_instr_en_i, dummy_instr_mask_i, dummy_instr_seed_en_i, dummy_instr_seed_i, icache_enable_i, icache_inval_i, icache_ecc_error_o, branch_target_ex_i, csr_mepc_i, csr_depc_i, csr_mtvec_i, csr_mtvec_init_o, id_in_ready_i, pc_mismatch_alert_o, if_busy_o, req_i_t0, instr_rvalid_i_t0, instr_req_o_t0
, instr_rdata_i_t0, instr_gnt_i_t0, instr_addr_o_t0, pmp_err_if_plus2_i_t0, pmp_err_if_i_t0, pc_set_i_t0, pc_mux_i_t0, pc_mismatch_alert_o_t0, pc_if_o_t0, pc_id_o_t0, nt_branch_mispredict_i_t0, nt_branch_addr_i_t0, instr_valid_id_o_t0, instr_valid_clear_i_t0, instr_rdata_id_o_t0, instr_rdata_c_id_o_t0, instr_rdata_alu_id_o_t0, instr_new_id_o_t0, instr_is_compressed_id_o_t0, instr_intg_err_o_t0, instr_fetch_err_plus2_o_t0
, instr_fetch_err_o_t0, instr_bus_err_i_t0, instr_bp_taken_o_t0, illegal_c_insn_id_o_t0, if_busy_o_t0, icache_inval_i_t0, icache_enable_i_t0, icache_ecc_error_o_t0, ic_tag_write_o_t0, ic_tag_wdata_o_t0, ic_tag_req_o_t0, ic_tag_rdata_i_t0, ic_tag_addr_o_t0, ic_scr_key_valid_i_t0, ic_scr_key_req_o_t0, ic_data_write_o_t0, ic_data_wdata_o_t0, ic_data_req_o_t0, ic_data_rdata_i_t0, ic_data_addr_o_t0, exc_pc_mux_i_t0
, exc_cause_t0, dummy_instr_id_o_t0, csr_mtvec_init_o_t0, csr_mtvec_i_t0, csr_mepc_i_t0, csr_depc_i_t0, branch_target_ex_i_t0, boot_addr_i_t0, id_in_ready_i_t0, dummy_instr_seed_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_mask_i_t0, dummy_instr_en_i_t0);
/* src = "generated/sv2v_out.v:18127.45-18127.84" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18127.45-18127.84" */
wire _001_;
/* src = "generated/sv2v_out.v:18127.44-18127.106" */
wire _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18127.44-18127.106" */
wire _003_;
/* src = "generated/sv2v_out.v:18133.12-18133.36" */
wire _004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18133.12-18133.36" */
wire _005_;
/* src = "generated/sv2v_out.v:18188.29-18188.73" */
wire _006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18188.29-18188.73" */
wire _007_;
/* src = "generated/sv2v_out.v:18188.78-18188.117" */
wire _008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18188.78-18188.117" */
wire _009_;
/* src = "generated/sv2v_out.v:18244.32-18244.81" */
wire _010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18244.32-18244.81" */
wire _011_;
/* src = "generated/sv2v_out.v:18244.31-18244.98" */
wire _012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18244.31-18244.98" */
wire _013_;
wire [31:0] _014_;
wire _015_;
wire [31:0] _016_;
wire [31:0] _017_;
wire [31:0] _018_;
wire [31:0] _019_;
wire [31:0] _020_;
wire [31:0] _021_;
wire [4:0] _022_;
wire [31:0] _023_;
wire [31:0] _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire [31:0] _037_;
wire [31:0] _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire [31:0] _077_;
wire [31:0] _078_;
wire [31:0] _079_;
wire [31:0] _080_;
wire [15:0] _081_;
wire [15:0] _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire [31:0] _091_;
wire [31:0] _092_;
wire [31:0] _093_;
wire [31:0] _094_;
wire [31:0] _095_;
wire [31:0] _096_;
wire [31:0] _097_;
wire [31:0] _098_;
wire [31:0] _099_;
wire [31:0] _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire [31:0] _119_;
wire [31:0] _120_;
wire [31:0] _121_;
wire [31:0] _122_;
wire [31:0] _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire [31:0] _137_;
wire [31:0] _138_;
wire [15:0] _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire [31:0] _152_;
wire [31:0] _153_;
wire [31:0] _154_;
wire [31:0] _155_;
/* cellift = 32'd1 */
wire [31:0] _156_;
wire [31:0] _157_;
/* cellift = 32'd1 */
wire [31:0] _158_;
wire [31:0] _159_;
/* cellift = 32'd1 */
wire [31:0] _160_;
wire [31:0] _161_;
wire [31:0] _162_;
/* cellift = 32'd1 */
wire [31:0] _163_;
/* src = "generated/sv2v_out.v:18012.29-18012.45" */
wire _164_;
/* src = "generated/sv2v_out.v:18255.53-18255.88" */
wire _165_;
/* src = "generated/sv2v_out.v:18127.64-18127.84" */
wire _166_;
/* src = "generated/sv2v_out.v:18188.97-18188.117" */
wire _167_;
/* src = "generated/sv2v_out.v:18244.85-18244.98" */
wire _168_;
/* src = "generated/sv2v_out.v:18129.31-18129.113" */
wire _169_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18129.31-18129.113" */
wire _170_;
/* src = "generated/sv2v_out.v:18244.33-18244.66" */
wire _171_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18244.33-18244.66" */
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
/* src = "generated/sv2v_out.v:17883.20-17883.31" */
input [31:0] boot_addr_i;
wire [31:0] boot_addr_i;
/* cellift = 32'd1 */
input [31:0] boot_addr_i_t0;
wire [31:0] boot_addr_i_t0;
/* src = "generated/sv2v_out.v:17933.20-17933.38" */
input [31:0] branch_target_ex_i;
wire [31:0] branch_target_ex_i;
/* cellift = 32'd1 */
input [31:0] branch_target_ex_i_t0;
wire [31:0] branch_target_ex_i_t0;
/* src = "generated/sv2v_out.v:17881.13-17881.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:17935.20-17935.30" */
input [31:0] csr_depc_i;
wire [31:0] csr_depc_i;
/* cellift = 32'd1 */
input [31:0] csr_depc_i_t0;
wire [31:0] csr_depc_i_t0;
/* src = "generated/sv2v_out.v:17934.20-17934.30" */
input [31:0] csr_mepc_i;
wire [31:0] csr_mepc_i;
/* cellift = 32'd1 */
input [31:0] csr_mepc_i_t0;
wire [31:0] csr_mepc_i_t0;
/* src = "generated/sv2v_out.v:17936.20-17936.31" */
input [31:0] csr_mtvec_i;
wire [31:0] csr_mtvec_i;
/* cellift = 32'd1 */
input [31:0] csr_mtvec_i_t0;
wire [31:0] csr_mtvec_i_t0;
/* src = "generated/sv2v_out.v:17937.14-17937.30" */
output csr_mtvec_init_o;
wire csr_mtvec_init_o;
/* cellift = 32'd1 */
output csr_mtvec_init_o_t0;
wire csr_mtvec_init_o_t0;
/* src = "generated/sv2v_out.v:17926.13-17926.29" */
input dummy_instr_en_i;
wire dummy_instr_en_i;
/* cellift = 32'd1 */
input dummy_instr_en_i_t0;
wire dummy_instr_en_i_t0;
/* src = "generated/sv2v_out.v:17914.13-17914.29" */
output dummy_instr_id_o;
reg dummy_instr_id_o;
/* cellift = 32'd1 */
output dummy_instr_id_o_t0;
reg dummy_instr_id_o_t0;
/* src = "generated/sv2v_out.v:17927.19-17927.37" */
input [2:0] dummy_instr_mask_i;
wire [2:0] dummy_instr_mask_i;
/* cellift = 32'd1 */
input [2:0] dummy_instr_mask_i_t0;
wire [2:0] dummy_instr_mask_i_t0;
/* src = "generated/sv2v_out.v:17928.13-17928.34" */
input dummy_instr_seed_en_i;
wire dummy_instr_seed_en_i;
/* cellift = 32'd1 */
input dummy_instr_seed_en_i_t0;
wire dummy_instr_seed_en_i_t0;
/* src = "generated/sv2v_out.v:17929.20-17929.38" */
input [31:0] dummy_instr_seed_i;
wire [31:0] dummy_instr_seed_i;
/* cellift = 32'd1 */
input [31:0] dummy_instr_seed_i_t0;
wire [31:0] dummy_instr_seed_i_t0;
/* src = "generated/sv2v_out.v:17925.19-17925.28" */
input [6:0] exc_cause;
wire [6:0] exc_cause;
/* cellift = 32'd1 */
input [6:0] exc_cause_t0;
wire [6:0] exc_cause_t0;
/* src = "generated/sv2v_out.v:17970.13-17970.19" */
wire [31:0] exc_pc;
/* src = "generated/sv2v_out.v:17924.19-17924.31" */
input [1:0] exc_pc_mux_i;
wire [1:0] exc_pc_mux_i;
/* cellift = 32'd1 */
input [1:0] exc_pc_mux_i_t0;
wire [1:0] exc_pc_mux_i_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17970.13-17970.19" */
wire [31:0] exc_pc_t0;
/* src = "generated/sv2v_out.v:17949.13-17949.25" */
/* unused_bits = "0" */
wire [31:0] fetch_addr_n;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17949.13-17949.25" */
/* unused_bits = "0" */
wire [31:0] fetch_addr_n_t0;
/* src = "generated/sv2v_out.v:17958.7-17958.16" */
wire fetch_err;
/* src = "generated/sv2v_out.v:17959.7-17959.22" */
wire fetch_err_plus2;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17959.7-17959.22" */
wire fetch_err_plus2_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17958.7-17958.16" */
wire fetch_err_t0;
/* src = "generated/sv2v_out.v:17956.14-17956.25" */
wire [31:0] fetch_rdata;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17956.14-17956.25" */
wire [31:0] fetch_rdata_t0;
/* src = "generated/sv2v_out.v:17955.7-17955.18" */
wire fetch_ready;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17955.7-17955.18" */
wire fetch_ready_t0;
/* src = "generated/sv2v_out.v:17954.7-17954.18" */
wire fetch_valid;
/* src = "generated/sv2v_out.v:17953.7-17953.22" */
wire fetch_valid_raw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17953.7-17953.22" */
wire fetch_valid_raw_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17954.7-17954.18" */
wire fetch_valid_t0;
/* src = "generated/sv2v_out.v:18015.15-18015.22" */
wire [1:0] \g_mem_ecc.ecc_err ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18015.15-18015.22" */
/* unused_bits = "0 1" */
wire [1:0] \g_mem_ecc.ecc_err_t0 ;
/* src = "generated/sv2v_out.v:18016.30-18016.45" */
wire [38:0] \g_mem_ecc.instr_rdata_buf ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18016.30-18016.45" */
wire [38:0] \g_mem_ecc.instr_rdata_buf_t0 ;
/* src = "generated/sv2v_out.v:18240.16-18240.36" */
wire [31:0] \g_secure_pc.prev_instr_addr_incr ;
/* src = "generated/sv2v_out.v:18241.16-18241.40" */
wire [31:0] \g_secure_pc.prev_instr_addr_incr_buf ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18241.16-18241.40" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] \g_secure_pc.prev_instr_addr_incr_buf_t0 ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18240.16-18240.36" */
wire [31:0] \g_secure_pc.prev_instr_addr_incr_t0 ;
/* src = "generated/sv2v_out.v:18243.9-18243.25" */
wire \g_secure_pc.prev_instr_seq_d ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18243.9-18243.25" */
wire \g_secure_pc.prev_instr_seq_d_t0 ;
/* src = "generated/sv2v_out.v:18242.8-18242.24" */
reg \g_secure_pc.prev_instr_seq_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18242.8-18242.24" */
reg \g_secure_pc.prev_instr_seq_q_t0 ;
/* src = "generated/sv2v_out.v:18142.16-18142.32" */
wire [31:0] \gen_dummy_instr.dummy_instr_data ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18142.16-18142.32" */
wire [31:0] \gen_dummy_instr.dummy_instr_data_t0 ;
/* src = "generated/sv2v_out.v:18141.9-18141.27" */
wire \gen_dummy_instr.insert_dummy_instr ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18141.9-18141.27" */
wire \gen_dummy_instr.insert_dummy_instr_t0 ;
/* src = "generated/sv2v_out.v:17899.42-17899.56" */
output [7:0] ic_data_addr_o;
wire [7:0] ic_data_addr_o;
/* cellift = 32'd1 */
output [7:0] ic_data_addr_o_t0;
wire [7:0] ic_data_addr_o_t0;
/* src = "generated/sv2v_out.v:17901.58-17901.73" */
input [127:0] ic_data_rdata_i;
wire [127:0] ic_data_rdata_i;
/* cellift = 32'd1 */
input [127:0] ic_data_rdata_i_t0;
wire [127:0] ic_data_rdata_i_t0;
/* src = "generated/sv2v_out.v:17897.20-17897.33" */
output [1:0] ic_data_req_o;
wire [1:0] ic_data_req_o;
/* cellift = 32'd1 */
output [1:0] ic_data_req_o_t0;
wire [1:0] ic_data_req_o_t0;
/* src = "generated/sv2v_out.v:17900.34-17900.49" */
output [63:0] ic_data_wdata_o;
wire [63:0] ic_data_wdata_o;
/* cellift = 32'd1 */
output [63:0] ic_data_wdata_o_t0;
wire [63:0] ic_data_wdata_o_t0;
/* src = "generated/sv2v_out.v:17898.14-17898.29" */
output ic_data_write_o;
wire ic_data_write_o;
/* cellift = 32'd1 */
output ic_data_write_o_t0;
wire ic_data_write_o_t0;
/* src = "generated/sv2v_out.v:17903.14-17903.30" */
output ic_scr_key_req_o;
wire ic_scr_key_req_o;
/* cellift = 32'd1 */
output ic_scr_key_req_o_t0;
wire ic_scr_key_req_o_t0;
/* src = "generated/sv2v_out.v:17902.13-17902.31" */
input ic_scr_key_valid_i;
wire ic_scr_key_valid_i;
/* cellift = 32'd1 */
input ic_scr_key_valid_i_t0;
wire ic_scr_key_valid_i_t0;
/* src = "generated/sv2v_out.v:17894.42-17894.55" */
output [7:0] ic_tag_addr_o;
wire [7:0] ic_tag_addr_o;
/* cellift = 32'd1 */
output [7:0] ic_tag_addr_o_t0;
wire [7:0] ic_tag_addr_o_t0;
/* src = "generated/sv2v_out.v:17896.57-17896.71" */
input [43:0] ic_tag_rdata_i;
wire [43:0] ic_tag_rdata_i;
/* cellift = 32'd1 */
input [43:0] ic_tag_rdata_i_t0;
wire [43:0] ic_tag_rdata_i_t0;
/* src = "generated/sv2v_out.v:17892.20-17892.32" */
output [1:0] ic_tag_req_o;
wire [1:0] ic_tag_req_o;
/* cellift = 32'd1 */
output [1:0] ic_tag_req_o_t0;
wire [1:0] ic_tag_req_o_t0;
/* src = "generated/sv2v_out.v:17895.33-17895.47" */
output [21:0] ic_tag_wdata_o;
wire [21:0] ic_tag_wdata_o;
/* cellift = 32'd1 */
output [21:0] ic_tag_wdata_o_t0;
wire [21:0] ic_tag_wdata_o_t0;
/* src = "generated/sv2v_out.v:17893.14-17893.28" */
output ic_tag_write_o;
wire ic_tag_write_o;
/* cellift = 32'd1 */
output ic_tag_write_o_t0;
wire ic_tag_write_o_t0;
/* src = "generated/sv2v_out.v:17932.14-17932.32" */
output icache_ecc_error_o;
wire icache_ecc_error_o;
/* cellift = 32'd1 */
output icache_ecc_error_o_t0;
wire icache_ecc_error_o_t0;
/* src = "generated/sv2v_out.v:17930.13-17930.28" */
input icache_enable_i;
wire icache_enable_i;
/* cellift = 32'd1 */
input icache_enable_i_t0;
wire icache_enable_i_t0;
/* src = "generated/sv2v_out.v:17931.13-17931.27" */
input icache_inval_i;
wire icache_inval_i;
/* cellift = 32'd1 */
input icache_inval_i_t0;
wire icache_inval_i_t0;
/* src = "generated/sv2v_out.v:17938.13-17938.26" */
input id_in_ready_i;
wire id_in_ready_i;
/* cellift = 32'd1 */
input id_in_ready_i_t0;
wire id_in_ready_i_t0;
/* src = "generated/sv2v_out.v:17940.14-17940.23" */
output if_busy_o;
wire if_busy_o;
/* cellift = 32'd1 */
output if_busy_o_t0;
wire if_busy_o_t0;
/* src = "generated/sv2v_out.v:17971.7-17971.24" */
wire if_id_pipe_reg_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17971.7-17971.24" */
wire if_id_pipe_reg_we_t0;
/* src = "generated/sv2v_out.v:17968.7-17968.19" */
wire if_instr_err;
/* src = "generated/sv2v_out.v:17969.7-17969.25" */
wire if_instr_err_plus2;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17969.7-17969.25" */
wire if_instr_err_plus2_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17968.7-17968.19" */
wire if_instr_err_t0;
/* src = "generated/sv2v_out.v:17967.7-17967.23" */
wire if_instr_pmp_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17967.7-17967.23" */
wire if_instr_pmp_err_t0;
/* src = "generated/sv2v_out.v:17961.7-17961.21" */
wire illegal_c_insn;
/* src = "generated/sv2v_out.v:17913.13-17913.32" */
output illegal_c_insn_id_o;
reg illegal_c_insn_id_o;
/* cellift = 32'd1 */
output illegal_c_insn_id_o_t0;
reg illegal_c_insn_id_o_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17961.7-17961.21" */
wire illegal_c_insn_t0;
/* src = "generated/sv2v_out.v:17975.7-17975.26" */
wire illegal_c_instr_out;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17975.7-17975.26" */
wire illegal_c_instr_out_t0;
/* src = "generated/sv2v_out.v:17886.21-17886.33" */
output [31:0] instr_addr_o;
wire [31:0] instr_addr_o;
/* cellift = 32'd1 */
output [31:0] instr_addr_o_t0;
wire [31:0] instr_addr_o_t0;
/* src = "generated/sv2v_out.v:17910.14-17910.30" */
output instr_bp_taken_o;
wire instr_bp_taken_o;
/* cellift = 32'd1 */
output instr_bp_taken_o_t0;
wire instr_bp_taken_o_t0;
/* src = "generated/sv2v_out.v:17890.13-17890.28" */
input instr_bus_err_i;
wire instr_bus_err_i;
/* cellift = 32'd1 */
input instr_bus_err_i_t0;
wire instr_bus_err_i_t0;
/* src = "generated/sv2v_out.v:17960.14-17960.32" */
wire [31:0] instr_decompressed;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17960.14-17960.32" */
wire [31:0] instr_decompressed_t0;
/* src = "generated/sv2v_out.v:17945.7-17945.16" */
wire instr_err;
/* src = "generated/sv2v_out.v:17976.7-17976.20" */
wire instr_err_out;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17976.7-17976.20" */
wire instr_err_out_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17945.7-17945.16" */
wire instr_err_t0;
/* src = "generated/sv2v_out.v:17911.13-17911.30" */
output instr_fetch_err_o;
reg instr_fetch_err_o;
/* cellift = 32'd1 */
output instr_fetch_err_o_t0;
reg instr_fetch_err_o_t0;
/* src = "generated/sv2v_out.v:17912.13-17912.36" */
output instr_fetch_err_plus2_o;
reg instr_fetch_err_plus2_o;
/* cellift = 32'd1 */
output instr_fetch_err_plus2_o_t0;
reg instr_fetch_err_plus2_o_t0;
/* src = "generated/sv2v_out.v:17887.13-17887.24" */
input instr_gnt_i;
wire instr_gnt_i;
/* cellift = 32'd1 */
input instr_gnt_i_t0;
wire instr_gnt_i_t0;
/* src = "generated/sv2v_out.v:17946.7-17946.21" */
wire instr_intg_err;
/* src = "generated/sv2v_out.v:17891.14-17891.30" */
output instr_intg_err_o;
wire instr_intg_err_o;
/* cellift = 32'd1 */
output instr_intg_err_o_t0;
wire instr_intg_err_o_t0;
/* src = "generated/sv2v_out.v:17962.7-17962.26" */
wire instr_is_compressed;
/* src = "generated/sv2v_out.v:17909.13-17909.37" */
output instr_is_compressed_id_o;
reg instr_is_compressed_id_o;
/* cellift = 32'd1 */
output instr_is_compressed_id_o_t0;
reg instr_is_compressed_id_o_t0;
/* src = "generated/sv2v_out.v:17974.7-17974.30" */
wire instr_is_compressed_out;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17974.7-17974.30" */
wire instr_is_compressed_out_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17962.7-17962.26" */
wire instr_is_compressed_t0;
/* src = "generated/sv2v_out.v:17905.14-17905.28" */
output instr_new_id_o;
reg instr_new_id_o;
/* cellift = 32'd1 */
output instr_new_id_o_t0;
reg instr_new_id_o_t0;
/* src = "generated/sv2v_out.v:17973.14-17973.23" */
wire [31:0] instr_out;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17973.14-17973.23" */
wire [31:0] instr_out_t0;
/* src = "generated/sv2v_out.v:17907.20-17907.40" */
output [31:0] instr_rdata_alu_id_o;
reg [31:0] instr_rdata_alu_id_o;
/* cellift = 32'd1 */
output [31:0] instr_rdata_alu_id_o_t0;
reg [31:0] instr_rdata_alu_id_o_t0;
/* src = "generated/sv2v_out.v:17908.20-17908.38" */
output [15:0] instr_rdata_c_id_o;
reg [15:0] instr_rdata_c_id_o;
/* cellift = 32'd1 */
output [15:0] instr_rdata_c_id_o_t0;
reg [15:0] instr_rdata_c_id_o_t0;
/* src = "generated/sv2v_out.v:17889.34-17889.47" */
input [38:0] instr_rdata_i;
wire [38:0] instr_rdata_i;
/* cellift = 32'd1 */
input [38:0] instr_rdata_i_t0;
wire [38:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:17906.20-17906.36" */
output [31:0] instr_rdata_id_o;
wire [31:0] instr_rdata_id_o;
/* cellift = 32'd1 */
output [31:0] instr_rdata_id_o_t0;
wire [31:0] instr_rdata_id_o_t0;
/* src = "generated/sv2v_out.v:17885.14-17885.25" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:17888.13-17888.27" */
input instr_rvalid_i;
wire instr_rvalid_i;
/* cellift = 32'd1 */
input instr_rvalid_i_t0;
wire instr_rvalid_i_t0;
/* src = "generated/sv2v_out.v:17919.13-17919.32" */
input instr_valid_clear_i;
wire instr_valid_clear_i;
/* cellift = 32'd1 */
input instr_valid_clear_i_t0;
wire instr_valid_clear_i_t0;
/* src = "generated/sv2v_out.v:17941.7-17941.23" */
wire instr_valid_id_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17941.7-17941.23" */
wire instr_valid_id_d_t0;
/* src = "generated/sv2v_out.v:17904.14-17904.30" */
output instr_valid_id_o;
reg instr_valid_id_o;
/* cellift = 32'd1 */
output instr_valid_id_o_t0;
reg instr_valid_id_o_t0;
/* src = "generated/sv2v_out.v:17979.12-17979.19" */
wire [4:0] irq_vec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17979.12-17979.19" */
wire [4:0] irq_vec_t0;
/* src = "generated/sv2v_out.v:17923.20-17923.36" */
input [31:0] nt_branch_addr_i;
wire [31:0] nt_branch_addr_i;
/* cellift = 32'd1 */
input [31:0] nt_branch_addr_i_t0;
wire [31:0] nt_branch_addr_i_t0;
/* src = "generated/sv2v_out.v:17922.13-17922.35" */
input nt_branch_mispredict_i;
wire nt_branch_mispredict_i;
/* cellift = 32'd1 */
input nt_branch_mispredict_i_t0;
wire nt_branch_mispredict_i_t0;
/* src = "generated/sv2v_out.v:17916.20-17916.27" */
output [31:0] pc_id_o;
reg [31:0] pc_id_o;
/* cellift = 32'd1 */
output [31:0] pc_id_o_t0;
reg [31:0] pc_id_o_t0;
/* src = "generated/sv2v_out.v:17915.21-17915.28" */
output [31:0] pc_if_o;
wire [31:0] pc_if_o;
/* cellift = 32'd1 */
output [31:0] pc_if_o_t0;
wire [31:0] pc_if_o_t0;
/* src = "generated/sv2v_out.v:17939.14-17939.33" */
output pc_mismatch_alert_o;
wire pc_mismatch_alert_o;
/* cellift = 32'd1 */
output pc_mismatch_alert_o_t0;
wire pc_mismatch_alert_o_t0;
/* src = "generated/sv2v_out.v:17921.19-17921.27" */
input [2:0] pc_mux_i;
wire [2:0] pc_mux_i;
/* cellift = 32'd1 */
input [2:0] pc_mux_i_t0;
wire [2:0] pc_mux_i_t0;
/* src = "generated/sv2v_out.v:17920.13-17920.21" */
input pc_set_i;
wire pc_set_i;
/* cellift = 32'd1 */
input pc_set_i_t0;
wire pc_set_i_t0;
/* src = "generated/sv2v_out.v:17917.13-17917.25" */
input pmp_err_if_i;
wire pmp_err_if_i;
/* cellift = 32'd1 */
input pmp_err_if_i_t0;
wire pmp_err_if_i_t0;
/* src = "generated/sv2v_out.v:17918.13-17918.31" */
input pmp_err_if_plus2_i;
wire pmp_err_if_plus2_i;
/* cellift = 32'd1 */
input pmp_err_if_plus2_i_t0;
wire pmp_err_if_plus2_i_t0;
/* src = "generated/sv2v_out.v:17952.14-17952.27" */
wire [31:0] prefetch_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17952.14-17952.27" */
wire [31:0] prefetch_addr_t0;
/* src = "generated/sv2v_out.v:17951.7-17951.22" */
wire prefetch_branch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17951.7-17951.22" */
wire prefetch_branch_t0;
/* src = "generated/sv2v_out.v:17884.13-17884.18" */
input req_i;
wire req_i;
/* cellift = 32'd1 */
input req_i_t0;
wire req_i_t0;
/* src = "generated/sv2v_out.v:17882.13-17882.19" */
input rst_ni;
wire rst_ni;
assign \g_secure_pc.prev_instr_addr_incr  = pc_id_o + /* src = "generated/sv2v_out.v:18250.34-18250.86" */ _038_;
assign csr_mtvec_init_o = _164_ & /* src = "generated/sv2v_out.v:18012.28-18012.57" */ pc_set_i;
assign instr_intg_err_o = instr_intg_err & /* src = "generated/sv2v_out.v:18032.28-18032.59" */ instr_rvalid_i;
assign fetch_valid = fetch_valid_raw & /* src = "generated/sv2v_out.v:18035.23-18035.64" */ _033_;
assign _000_ = pc_if_o[1] & /* src = "generated/sv2v_out.v:18129.33-18129.72" */ _166_;
assign _002_ = _000_ & /* src = "generated/sv2v_out.v:18129.32-18129.94" */ pmp_err_if_plus2_i;
assign if_instr_err_plus2 = _169_ & /* src = "generated/sv2v_out.v:18129.30-18129.130" */ _028_;
assign _004_ = fetch_valid & /* src = "generated/sv2v_out.v:18133.12-18133.36" */ _029_;
assign _006_ = if_id_pipe_reg_we & /* src = "generated/sv2v_out.v:18188.29-18188.73" */ _027_;
assign _008_ = instr_valid_id_o & /* src = "generated/sv2v_out.v:18188.78-18188.117" */ _167_;
assign if_id_pipe_reg_we = fetch_valid & /* src = "generated/sv2v_out.v:18189.26-18189.56" */ id_in_ready_i;
assign _010_ = _171_ & /* src = "generated/sv2v_out.v:18244.32-18244.81" */ _027_;
assign _012_ = _010_ & /* src = "generated/sv2v_out.v:18244.31-18244.98" */ _168_;
assign \g_secure_pc.prev_instr_seq_d  = _012_ & /* src = "generated/sv2v_out.v:18244.30-18244.120" */ _025_;
assign pc_mismatch_alert_o = \g_secure_pc.prev_instr_seq_q  & /* src = "generated/sv2v_out.v:18255.33-18255.89" */ _165_;
assign fetch_ready = id_in_ready_i & /* src = "generated/sv2v_out.v:18336.25-18336.59" */ _025_;
assign _014_ = ~ pc_id_o_t0;
assign _037_ = pc_id_o & _014_;
assign _153_ = _037_ + _038_;
assign _123_ = pc_id_o | pc_id_o_t0;
assign _154_ = _123_ + _038_;
assign _152_ = _153_ ^ _154_;
assign \g_secure_pc.prev_instr_addr_incr_t0  = _152_ | pc_id_o_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME \g_secure_pc.prev_instr_seq_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_secure_pc.prev_instr_seq_q_t0  <= 1'h0;
else \g_secure_pc.prev_instr_seq_q_t0  <= \g_secure_pc.prev_instr_seq_d_t0 ;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_valid_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_valid_id_o_t0 <= 1'h0;
else instr_valid_id_o_t0 <= instr_valid_id_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_new_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_new_id_o_t0 <= 1'h0;
else instr_new_id_o_t0 <= if_id_pipe_reg_we_t0;
assign _015_ = ~ if_id_pipe_reg_we;
assign _075_ = if_id_pipe_reg_we & \gen_dummy_instr.insert_dummy_instr_t0 ;
assign _077_ = { if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we } & pc_if_o_t0;
assign _079_ = { if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we } & instr_out_t0;
assign _081_ = { if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we } & fetch_rdata_t0[15:0];
assign _083_ = if_id_pipe_reg_we & instr_is_compressed_out_t0;
assign _085_ = if_id_pipe_reg_we & instr_err_out_t0;
assign _087_ = if_id_pipe_reg_we & if_instr_err_plus2_t0;
assign _089_ = if_id_pipe_reg_we & illegal_c_instr_out_t0;
assign _076_ = _015_ & dummy_instr_id_o_t0;
assign _078_ = { _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_ } & pc_id_o_t0;
assign _080_ = { _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_ } & instr_rdata_alu_id_o_t0;
assign _082_ = { _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_, _015_ } & instr_rdata_c_id_o_t0;
assign _084_ = _015_ & instr_is_compressed_id_o_t0;
assign _086_ = _015_ & instr_fetch_err_o_t0;
assign _088_ = _015_ & instr_fetch_err_plus2_o_t0;
assign _090_ = _015_ & illegal_c_insn_id_o_t0;
assign _136_ = _075_ | _076_;
assign _137_ = _077_ | _078_;
assign _138_ = _079_ | _080_;
assign _139_ = _081_ | _082_;
assign _140_ = _083_ | _084_;
assign _141_ = _085_ | _086_;
assign _142_ = _087_ | _088_;
assign _143_ = _089_ | _090_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME dummy_instr_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_instr_id_o_t0 <= 1'h0;
else dummy_instr_id_o_t0 <= _136_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME pc_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) pc_id_o_t0 <= 32'd0;
else pc_id_o_t0 <= _137_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_rdata_alu_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_rdata_alu_id_o_t0 <= 32'd0;
else instr_rdata_alu_id_o_t0 <= _138_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_rdata_c_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_rdata_c_id_o_t0 <= 16'h0000;
else instr_rdata_c_id_o_t0 <= _139_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_is_compressed_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_is_compressed_id_o_t0 <= 1'h0;
else instr_is_compressed_id_o_t0 <= _140_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_fetch_err_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_fetch_err_o_t0 <= 1'h0;
else instr_fetch_err_o_t0 <= _141_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_fetch_err_plus2_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_fetch_err_plus2_o_t0 <= 1'h0;
else instr_fetch_err_plus2_o_t0 <= _142_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME illegal_c_insn_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) illegal_c_insn_id_o_t0 <= 1'h0;
else illegal_c_insn_id_o_t0 <= _143_;
assign _039_ = fetch_valid_raw_t0 & _033_;
assign _042_ = pc_if_o_t0[1] & _166_;
assign _045_ = _001_ & pmp_err_if_plus2_i;
assign _048_ = _170_ & _028_;
assign _051_ = fetch_valid_t0 & _029_;
assign _054_ = if_id_pipe_reg_we_t0 & _027_;
assign _057_ = instr_valid_id_o_t0 & _167_;
assign _060_ = fetch_valid_t0 & id_in_ready_i;
assign _063_ = _172_ & _027_;
assign _066_ = _011_ & _168_;
assign _069_ = _013_ & _025_;
assign pc_mismatch_alert_o_t0 = \g_secure_pc.prev_instr_seq_q_t0  & _165_;
assign _072_ = id_in_ready_i_t0 & _025_;
assign csr_mtvec_init_o_t0 = pc_set_i_t0 & _164_;
assign instr_intg_err_o_t0 = instr_rvalid_i_t0 & instr_intg_err;
assign _040_ = nt_branch_mispredict_i_t0 & fetch_valid_raw;
assign _043_ = instr_is_compressed_t0 & pc_if_o[1];
assign _046_ = pmp_err_if_plus2_i_t0 & _000_;
assign _049_ = pmp_err_if_i_t0 & _169_;
assign _052_ = fetch_err_t0 & fetch_valid;
assign _055_ = pc_set_i_t0 & if_id_pipe_reg_we;
assign _058_ = instr_valid_clear_i_t0 & instr_valid_id_o;
assign _061_ = id_in_ready_i_t0 & fetch_valid;
assign _064_ = pc_set_i_t0 & _171_;
assign _067_ = if_instr_err_t0 & _010_;
assign _070_ = \gen_dummy_instr.insert_dummy_instr_t0  & _012_;
assign _073_ = \gen_dummy_instr.insert_dummy_instr_t0  & id_in_ready_i;
assign _041_ = fetch_valid_raw_t0 & nt_branch_mispredict_i_t0;
assign _044_ = pc_if_o_t0[1] & instr_is_compressed_t0;
assign _047_ = _001_ & pmp_err_if_plus2_i_t0;
assign _050_ = _170_ & pmp_err_if_i_t0;
assign _053_ = fetch_valid_t0 & fetch_err_t0;
assign _056_ = if_id_pipe_reg_we_t0 & pc_set_i_t0;
assign _059_ = instr_valid_id_o_t0 & instr_valid_clear_i_t0;
assign _062_ = fetch_valid_t0 & id_in_ready_i_t0;
assign _065_ = _172_ & pc_set_i_t0;
assign _068_ = _011_ & if_instr_err_t0;
assign _071_ = _013_ & \gen_dummy_instr.insert_dummy_instr_t0 ;
assign _074_ = id_in_ready_i_t0 & \gen_dummy_instr.insert_dummy_instr_t0 ;
assign _124_ = _039_ | _040_;
assign _125_ = _042_ | _043_;
assign _126_ = _045_ | _046_;
assign _127_ = _048_ | _049_;
assign _128_ = _051_ | _052_;
assign _129_ = _054_ | _055_;
assign _130_ = _057_ | _058_;
assign _131_ = _060_ | _061_;
assign _132_ = _063_ | _064_;
assign _133_ = _066_ | _067_;
assign _134_ = _069_ | _070_;
assign _135_ = _072_ | _073_;
assign fetch_valid_t0 = _124_ | _041_;
assign _001_ = _125_ | _044_;
assign _003_ = _126_ | _047_;
assign if_instr_err_plus2_t0 = _127_ | _050_;
assign _005_ = _128_ | _053_;
assign _007_ = _129_ | _056_;
assign _009_ = _130_ | _059_;
assign if_id_pipe_reg_we_t0 = _131_ | _062_;
assign _011_ = _132_ | _065_;
assign _013_ = _133_ | _068_;
assign \g_secure_pc.prev_instr_seq_d_t0  = _134_ | _071_;
assign fetch_ready_t0 = _135_ | _074_;
/* src = "generated/sv2v_out.v:18163.4-18167.45" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME dummy_instr_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_instr_id_o <= 1'h0;
else if (if_id_pipe_reg_we) dummy_instr_id_o <= \gen_dummy_instr.insert_dummy_instr ;
/* src = "generated/sv2v_out.v:18204.4-18224.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME pc_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) pc_id_o <= 32'd0;
else if (if_id_pipe_reg_we) pc_id_o <= pc_if_o;
/* src = "generated/sv2v_out.v:18204.4-18224.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_rdata_alu_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_rdata_alu_id_o <= 32'd0;
else if (if_id_pipe_reg_we) instr_rdata_alu_id_o <= instr_out;
/* src = "generated/sv2v_out.v:18204.4-18224.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_rdata_c_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_rdata_c_id_o <= 16'h0000;
else if (if_id_pipe_reg_we) instr_rdata_c_id_o <= fetch_rdata[15:0];
/* src = "generated/sv2v_out.v:18204.4-18224.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_is_compressed_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_is_compressed_id_o <= 1'h0;
else if (if_id_pipe_reg_we) instr_is_compressed_id_o <= instr_is_compressed_out;
/* src = "generated/sv2v_out.v:18204.4-18224.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_fetch_err_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_fetch_err_o <= 1'h0;
else if (if_id_pipe_reg_we) instr_fetch_err_o <= instr_err_out;
/* src = "generated/sv2v_out.v:18204.4-18224.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_fetch_err_plus2_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_fetch_err_plus2_o <= 1'h0;
else if (if_id_pipe_reg_we) instr_fetch_err_plus2_o <= if_instr_err_plus2;
/* src = "generated/sv2v_out.v:18204.4-18224.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME illegal_c_insn_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) illegal_c_insn_id_o <= 1'h0;
else if (if_id_pipe_reg_we) illegal_c_insn_id_o <= illegal_c_instr_out;
assign _016_ = ~ { _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_ };
assign _017_ = ~ { _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_ };
assign _018_ = ~ { _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_ };
assign _019_ = ~ { _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_ };
assign _020_ = ~ { _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_ };
assign _021_ = ~ { _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_ };
assign _022_ = ~ { exc_cause[6], exc_cause[6], exc_cause[6], exc_cause[6], exc_cause[6] };
assign _023_ = ~ { pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i };
assign _024_ = ~ { \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr  };
assign _025_ = ~ \gen_dummy_instr.insert_dummy_instr ;
assign _091_ = _016_ & csr_mepc_i_t0;
assign _093_ = _017_ & { boot_addr_i_t0[31:8], 8'h00 };
assign _095_ = _018_ & _158_;
assign _097_ = _019_ & _160_;
assign _099_ = _020_ & { csr_mtvec_i_t0[31:8], 8'h00 };
assign exc_pc_t0 = _021_ & _163_;
assign irq_vec_t0 = _022_ & exc_cause_t0[4:0];
assign _119_ = _023_ & nt_branch_addr_i_t0;
assign _121_ = _024_ & instr_decompressed_t0;
assign instr_is_compressed_out_t0 = _025_ & instr_is_compressed_t0;
assign illegal_c_instr_out_t0 = _025_ & illegal_c_insn_t0;
assign instr_err_out_t0 = _025_ & if_instr_err_t0;
assign _092_ = { _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_, _173_ } & csr_depc_i_t0;
assign _094_ = { _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_, _176_ } & branch_target_ex_i_t0;
assign _096_ = { _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_, _175_ } & exc_pc_t0;
assign _098_ = { _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_, _150_ } & _156_;
assign _100_ = { _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_, _179_ } & { csr_mtvec_i_t0[31:8], 1'h0, irq_vec_t0, 2'h0 };
assign _120_ = { pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i } & { fetch_addr_n_t0[31:1], 1'h0 };
assign _122_ = { \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr  } & \gen_dummy_instr.dummy_instr_data_t0 ;
assign _156_ = _091_ | _092_;
assign _158_ = _093_ | _094_;
assign _160_ = _095_ | _096_;
assign fetch_addr_n_t0 = _097_ | _098_;
assign _163_ = _099_ | _100_;
assign prefetch_addr_t0 = _119_ | _120_;
assign instr_out_t0 = _121_ | _122_;
assign _026_ = ~ instr_intg_err;
assign _027_ = ~ pc_set_i;
assign _028_ = ~ pmp_err_if_i;
assign _029_ = ~ fetch_err;
assign _030_ = ~ _002_;
assign _031_ = ~ _006_;
assign _032_ = ~ \g_secure_pc.prev_instr_seq_q ;
assign _033_ = ~ nt_branch_mispredict_i;
assign _034_ = ~ if_instr_pmp_err;
assign _035_ = ~ fetch_err_plus2;
assign _036_ = ~ _008_;
assign _101_ = pc_set_i_t0 & _033_;
assign _104_ = pmp_err_if_i_t0 & _030_;
assign _107_ = fetch_err_t0 & _034_;
assign _110_ = _003_ & _035_;
assign _113_ = _007_ & _036_;
assign _116_ = \g_secure_pc.prev_instr_seq_q_t0  & _015_;
assign instr_err_t0 = instr_bus_err_i_t0 & _026_;
assign _102_ = nt_branch_mispredict_i_t0 & _027_;
assign _105_ = _003_ & _028_;
assign _108_ = if_instr_pmp_err_t0 & _029_;
assign _111_ = fetch_err_plus2_t0 & _030_;
assign _114_ = _009_ & _031_;
assign _117_ = if_id_pipe_reg_we_t0 & _032_;
assign _103_ = pc_set_i_t0 & nt_branch_mispredict_i_t0;
assign _106_ = pmp_err_if_i_t0 & _003_;
assign _109_ = fetch_err_t0 & if_instr_pmp_err_t0;
assign _112_ = _003_ & fetch_err_plus2_t0;
assign _115_ = _007_ & _009_;
assign _118_ = \g_secure_pc.prev_instr_seq_q_t0  & if_id_pipe_reg_we_t0;
assign _144_ = _101_ | _102_;
assign _145_ = _104_ | _105_;
assign _146_ = _107_ | _108_;
assign _147_ = _110_ | _111_;
assign _148_ = _113_ | _114_;
assign _149_ = _116_ | _117_;
assign prefetch_branch_t0 = _144_ | _103_;
assign if_instr_pmp_err_t0 = _145_ | _106_;
assign if_instr_err_t0 = _146_ | _109_;
assign _170_ = _147_ | _112_;
assign instr_valid_id_d_t0 = _148_ | _115_;
assign _172_ = _149_ | _118_;
assign _150_ = _174_ | _173_;
assign _151_ = _178_ | _177_;
assign _155_ = _173_ ? csr_depc_i : csr_mepc_i;
assign _157_ = _176_ ? branch_target_ex_i : { boot_addr_i[31:8], 8'h80 };
assign _159_ = _175_ ? exc_pc : _157_;
assign fetch_addr_n = _150_ ? _155_ : _159_;
assign _161_ = _177_ ? 32'd437323784 : 32'd437323776;
assign _162_ = _179_ ? { csr_mtvec_i[31:8], 1'h0, irq_vec, 2'h0 } : { csr_mtvec_i[31:8], 8'h00 };
assign exc_pc = _151_ ? _161_ : _162_;
assign _164_ = ! /* src = "generated/sv2v_out.v:18012.29-18012.45" */ pc_mux_i;
assign _165_ = pc_if_o != /* src = "generated/sv2v_out.v:18255.53-18255.88" */ \g_secure_pc.prev_instr_addr_incr_buf ;
assign _166_ = ~ /* src = "generated/sv2v_out.v:18129.52-18129.72" */ instr_is_compressed;
assign _167_ = ~ /* src = "generated/sv2v_out.v:18188.97-18188.117" */ instr_valid_clear_i;
assign _168_ = ~ /* src = "generated/sv2v_out.v:18244.85-18244.98" */ if_instr_err;
assign instr_err = instr_intg_err | /* src = "generated/sv2v_out.v:18031.21-18031.53" */ instr_bus_err_i;
assign prefetch_branch = pc_set_i | /* src = "generated/sv2v_out.v:18033.27-18033.62" */ nt_branch_mispredict_i;
assign if_instr_pmp_err = pmp_err_if_i | /* src = "generated/sv2v_out.v:18127.28-18127.107" */ _002_;
assign if_instr_err = fetch_err | /* src = "generated/sv2v_out.v:18128.24-18128.59" */ if_instr_pmp_err;
assign _169_ = _002_ | /* src = "generated/sv2v_out.v:18129.31-18129.113" */ fetch_err_plus2;
assign instr_valid_id_d = _006_ | /* src = "generated/sv2v_out.v:18188.28-18188.118" */ _008_;
assign _171_ = \g_secure_pc.prev_instr_seq_q  | /* src = "generated/sv2v_out.v:18244.33-18244.66" */ if_id_pipe_reg_we;
/* src = "generated/sv2v_out.v:18245.4-18249.43" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME \g_secure_pc.prev_instr_seq_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_secure_pc.prev_instr_seq_q  <= 1'h0;
else \g_secure_pc.prev_instr_seq_q  <= \g_secure_pc.prev_instr_seq_d ;
/* src = "generated/sv2v_out.v:18190.2-18198.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_valid_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_valid_id_o <= 1'h0;
else instr_valid_id_o <= instr_valid_id_d;
/* src = "generated/sv2v_out.v:18190.2-18198.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_new_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_new_id_o <= 1'h0;
else instr_new_id_o <= if_id_pipe_reg_we;
assign _173_ = pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18002.3-18010.10" */ 3'h4;
assign _174_ = pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18002.3-18010.10" */ 3'h3;
assign _175_ = pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18002.3-18010.10" */ 3'h2;
assign _176_ = pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18002.3-18010.10" */ 3'h1;
assign _177_ = exc_pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17992.3-17998.10" */ 2'h3;
assign _178_ = exc_pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17992.3-17998.10" */ 2'h2;
assign _179_ = exc_pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17992.3-17998.10" */ 2'h1;
assign irq_vec = exc_cause[6] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17990.7-17990.19|generated/sv2v_out.v:17990.3-17991.43" */ 5'h1f : exc_cause[4:0];
assign instr_intg_err = | /* src = "generated/sv2v_out.v:18025.28-18025.36" */ \g_mem_ecc.ecc_err ;
assign prefetch_addr = pc_set_i ? /* src = "generated/sv2v_out.v:18034.26-18034.84" */ { fetch_addr_n[31:1], 1'h0 } : nt_branch_addr_i;
assign instr_out = \gen_dummy_instr.insert_dummy_instr  ? /* src = "generated/sv2v_out.v:18158.24-18158.82" */ \gen_dummy_instr.dummy_instr_data  : instr_decompressed;
assign instr_is_compressed_out = \gen_dummy_instr.insert_dummy_instr  ? /* src = "generated/sv2v_out.v:18159.38-18159.85" */ 1'h0 : instr_is_compressed;
assign illegal_c_instr_out = \gen_dummy_instr.insert_dummy_instr  ? /* src = "generated/sv2v_out.v:18160.34-18160.76" */ 1'h0 : illegal_c_insn;
assign instr_err_out = \gen_dummy_instr.insert_dummy_instr  ? /* src = "generated/sv2v_out.v:18161.28-18161.68" */ 1'h0 : if_instr_err;
assign _038_ = instr_is_compressed_id_o ? /* src = "generated/sv2v_out.v:18250.45-18250.85" */ 32'd2 : 32'd4;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18130.26-18138.3" */
ibex_compressed_decoder compressed_decoder_i (
.clk_i(clk_i),
.illegal_instr_o(illegal_c_insn),
.illegal_instr_o_t0(illegal_c_insn_t0),
.instr_i(fetch_rdata),
.instr_i_t0(fetch_rdata_t0),
.instr_o(instr_decompressed),
.instr_o_t0(instr_decompressed_t0),
.is_compressed_o(instr_is_compressed),
.is_compressed_o_t0(instr_is_compressed_t0),
.rst_ni(rst_ni),
.valid_i(_004_),
.valid_i_t0(_005_)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18021.30-18024.5" */
prim_secded_inv_39_32_dec \g_mem_ecc.u_instr_intg_dec  (
.data_i(\g_mem_ecc.instr_rdata_buf ),
.data_i_t0(\g_mem_ecc.instr_rdata_buf_t0 ),
.err_o(\g_mem_ecc.ecc_err ),
.err_o_t0(\g_mem_ecc.ecc_err_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18017.37-18020.5" */
\$paramod\prim_buf\Width=32'00000000000000000000000000100111  \g_mem_ecc.u_prim_buf_instr_rdata  (
.in_i(instr_rdata_i),
.in_i_t0(instr_rdata_i_t0),
.out_o(\g_mem_ecc.instr_rdata_buf ),
.out_o_t0(\g_mem_ecc.instr_rdata_buf_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18251.27-18254.5" */
\$paramod\prim_buf\Width=s32'00000000000000000000000000100000  \g_secure_pc.u_prev_instr_addr_incr_buf  (
.in_i(\g_secure_pc.prev_instr_addr_incr ),
.in_i_t0(\g_secure_pc.prev_instr_addr_incr_t0 ),
.out_o(\g_secure_pc.prev_instr_addr_incr_buf ),
.out_o_t0(\g_secure_pc.prev_instr_addr_incr_buf_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18146.6-18157.5" */
\$paramod$501c60d7519704ee720c78ef16ad88cf05835059\ibex_dummy_instr  \gen_dummy_instr.dummy_instr_i  (
.clk_i(clk_i),
.dummy_instr_data_o(\gen_dummy_instr.dummy_instr_data ),
.dummy_instr_data_o_t0(\gen_dummy_instr.dummy_instr_data_t0 ),
.dummy_instr_en_i(dummy_instr_en_i),
.dummy_instr_en_i_t0(dummy_instr_en_i_t0),
.dummy_instr_mask_i(dummy_instr_mask_i),
.dummy_instr_mask_i_t0(dummy_instr_mask_i_t0),
.dummy_instr_seed_en_i(dummy_instr_seed_en_i),
.dummy_instr_seed_en_i_t0(dummy_instr_seed_en_i_t0),
.dummy_instr_seed_i(dummy_instr_seed_i),
.dummy_instr_seed_i_t0(dummy_instr_seed_i_t0),
.fetch_valid_i(fetch_valid),
.fetch_valid_i_t0(fetch_valid_t0),
.id_in_ready_i(id_in_ready_i),
.id_in_ready_i_t0(id_in_ready_i_t0),
.insert_dummy_instr_o(\gen_dummy_instr.insert_dummy_instr ),
.insert_dummy_instr_o_t0(\gen_dummy_instr.insert_dummy_instr_t0 ),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18081.48-18100.5" */
\$paramod\ibex_prefetch_buffer\ResetAll=1'1  \gen_prefetch_buffer.prefetch_buffer_i  (
.addr_i(prefetch_addr),
.addr_i_t0(prefetch_addr_t0),
.addr_o(pc_if_o),
.addr_o_t0(pc_if_o_t0),
.branch_i(prefetch_branch),
.branch_i_t0(prefetch_branch_t0),
.busy_o(if_busy_o),
.busy_o_t0(if_busy_o_t0),
.clk_i(clk_i),
.err_o(fetch_err),
.err_o_t0(fetch_err_t0),
.err_plus2_o(fetch_err_plus2),
.err_plus2_o_t0(fetch_err_plus2_t0),
.instr_addr_o(instr_addr_o),
.instr_addr_o_t0(instr_addr_o_t0),
.instr_err_i(instr_err),
.instr_err_i_t0(instr_err_t0),
.instr_gnt_i(instr_gnt_i),
.instr_gnt_i_t0(instr_gnt_i_t0),
.instr_rdata_i(instr_rdata_i[31:0]),
.instr_rdata_i_t0(instr_rdata_i_t0[31:0]),
.instr_req_o(instr_req_o),
.instr_req_o_t0(instr_req_o_t0),
.instr_rvalid_i(instr_rvalid_i),
.instr_rvalid_i_t0(instr_rvalid_i_t0),
.rdata_o(fetch_rdata),
.rdata_o_t0(fetch_rdata_t0),
.ready_i(fetch_ready),
.ready_i_t0(fetch_ready_t0),
.req_i(req_i),
.req_i_t0(req_i_t0),
.rst_ni(rst_ni),
.valid_o(fetch_valid_raw),
.valid_o_t0(fetch_valid_raw_t0)
);
assign ic_data_addr_o = 8'h00;
assign ic_data_addr_o_t0 = 8'h00;
assign ic_data_req_o = 2'h0;
assign ic_data_req_o_t0 = 2'h0;
assign ic_data_wdata_o = 64'h0000000000000000;
assign ic_data_wdata_o_t0 = 64'h0000000000000000;
assign ic_data_write_o = 1'h0;
assign ic_data_write_o_t0 = 1'h0;
assign ic_scr_key_req_o = 1'h0;
assign ic_scr_key_req_o_t0 = 1'h0;
assign ic_tag_addr_o = 8'h00;
assign ic_tag_addr_o_t0 = 8'h00;
assign ic_tag_req_o = 2'h0;
assign ic_tag_req_o_t0 = 2'h0;
assign ic_tag_wdata_o = 22'h000000;
assign ic_tag_wdata_o_t0 = 22'h000000;
assign ic_tag_write_o = 1'h0;
assign ic_tag_write_o_t0 = 1'h0;
assign icache_ecc_error_o = 1'h0;
assign icache_ecc_error_o_t0 = 1'h0;
assign instr_bp_taken_o = 1'h0;
assign instr_bp_taken_o_t0 = 1'h0;
assign instr_rdata_id_o = instr_rdata_alu_id_o;
assign instr_rdata_id_o_t0 = instr_rdata_alu_id_o_t0;
endmodule

module \$paramod$916c47de983e2a42946808797a4a11650abb788f\prim_onehot_check (clk_i, rst_ni, oh_i, addr_i, en_i, err_o, addr_i_t0, en_i_t0, err_o_t0, oh_i_t0);
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _000_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _001_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _002_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _003_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _004_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _005_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _006_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _007_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _008_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _009_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _010_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _011_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _012_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _013_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _014_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _015_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _016_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _017_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _018_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _019_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _020_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _021_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _022_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _023_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _024_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _025_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _026_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _027_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _028_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _029_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _030_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _031_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _032_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _033_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _034_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _035_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _036_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _037_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _038_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _039_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _040_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _041_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _042_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _043_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _044_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _045_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _046_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _047_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _048_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _049_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _050_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _051_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _052_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _053_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _054_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _055_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _056_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _057_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _058_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _059_;
/* src = "generated/sv2v_out.v:26515.83-26515.130" */
wire _060_;
/* src = "generated/sv2v_out.v:26515.29-26515.77" */
wire _061_;
/* src = "generated/sv2v_out.v:26516.30-26516.56" */
wire _062_;
/* src = "generated/sv2v_out.v:26516.30-26516.56" */
wire _063_;
/* src = "generated/sv2v_out.v:26516.30-26516.56" */
wire _064_;
/* src = "generated/sv2v_out.v:26516.30-26516.56" */
wire _065_;
/* src = "generated/sv2v_out.v:26516.30-26516.56" */
wire _066_;
/* src = "generated/sv2v_out.v:26516.30-26516.56" */
wire _067_;
/* src = "generated/sv2v_out.v:26516.30-26516.56" */
wire _068_;
/* src = "generated/sv2v_out.v:26516.30-26516.56" */
wire _069_;
/* src = "generated/sv2v_out.v:26516.30-26516.56" */
wire _070_;
/* src = "generated/sv2v_out.v:26516.30-26516.56" */
wire _071_;
/* src = "generated/sv2v_out.v:26516.30-26516.56" */
wire _072_;
/* src = "generated/sv2v_out.v:26516.30-26516.56" */
wire _073_;
/* src = "generated/sv2v_out.v:26516.30-26516.56" */
wire _074_;
/* src = "generated/sv2v_out.v:26516.30-26516.56" */
wire _075_;
/* src = "generated/sv2v_out.v:26516.30-26516.56" */
wire _076_;
/* src = "generated/sv2v_out.v:26515.29-26515.61" */
wire _077_;
/* src = "generated/sv2v_out.v:26515.29-26515.61" */
wire _078_;
/* src = "generated/sv2v_out.v:26515.29-26515.61" */
wire _079_;
/* src = "generated/sv2v_out.v:26515.29-26515.61" */
wire _080_;
/* src = "generated/sv2v_out.v:26515.29-26515.61" */
wire _081_;
/* src = "generated/sv2v_out.v:26516.29-26516.73" */
wire _082_;
/* src = "generated/sv2v_out.v:26516.29-26516.73" */
wire _083_;
/* src = "generated/sv2v_out.v:26516.29-26516.73" */
wire _084_;
/* src = "generated/sv2v_out.v:26516.29-26516.73" */
wire _085_;
/* src = "generated/sv2v_out.v:26516.29-26516.73" */
wire _086_;
/* src = "generated/sv2v_out.v:26516.29-26516.73" */
wire _087_;
/* src = "generated/sv2v_out.v:26516.29-26516.73" */
wire _088_;
/* src = "generated/sv2v_out.v:26516.29-26516.73" */
wire _089_;
/* src = "generated/sv2v_out.v:26516.29-26516.73" */
wire _090_;
/* src = "generated/sv2v_out.v:26516.29-26516.73" */
wire _091_;
/* src = "generated/sv2v_out.v:26516.29-26516.73" */
wire _092_;
/* src = "generated/sv2v_out.v:26516.29-26516.73" */
wire _093_;
/* src = "generated/sv2v_out.v:26516.29-26516.73" */
wire _094_;
/* src = "generated/sv2v_out.v:26516.29-26516.73" */
wire _095_;
/* src = "generated/sv2v_out.v:26516.29-26516.73" */
wire _096_;
/* src = "generated/sv2v_out.v:26524.18-26524.39" */
wire _097_;
/* src = "generated/sv2v_out.v:26522.7-26522.15" */
wire addr_err;
/* src = "generated/sv2v_out.v:26485.31-26485.37" */
input [4:0] addr_i;
wire [4:0] addr_i;
/* cellift = 32'd1 */
input [4:0] addr_i_t0;
wire [4:0] addr_i_t0;
/* src = "generated/sv2v_out.v:26490.38-26490.46" */
wire [62:0] and_tree;
/* src = "generated/sv2v_out.v:26482.8-26482.13" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:26486.13-26486.17" */
input en_i;
wire en_i;
/* cellift = 32'd1 */
input en_i_t0;
wire en_i_t0;
/* src = "generated/sv2v_out.v:26521.7-26521.17" */
wire enable_err;
/* src = "generated/sv2v_out.v:26487.14-26487.19" */
output err_o;
wire err_o;
/* cellift = 32'd1 */
output err_o_t0;
wire err_o_t0;
/* src = "generated/sv2v_out.v:26491.38-26491.46" */
wire [62:0] err_tree;
/* src = "generated/sv2v_out.v:26523.7-26523.14" */
wire oh0_err;
/* src = "generated/sv2v_out.v:26484.33-26484.37" */
input [31:0] oh_i;
wire [31:0] oh_i;
/* cellift = 32'd1 */
input [31:0] oh_i_t0;
wire [31:0] oh_i_t0;
/* src = "generated/sv2v_out.v:26489.38-26489.45" */
wire [62:0] or_tree;
/* src = "generated/sv2v_out.v:26483.8-26483.14" */
input rst_ni;
wire rst_ni;
assign _000_ = addr_i[2] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ and_tree[14];
assign _001_ = _077_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ and_tree[15];
assign _002_ = addr_i[1] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ and_tree[16];
assign _003_ = _077_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ and_tree[17];
assign _004_ = addr_i[1] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ and_tree[18];
assign _005_ = _077_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ and_tree[19];
assign _006_ = addr_i[1] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ and_tree[20];
assign _007_ = _077_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ and_tree[21];
assign _008_ = addr_i[1] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ and_tree[22];
assign _009_ = _077_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ and_tree[23];
assign _010_ = addr_i[1] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ and_tree[24];
assign _011_ = _077_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ and_tree[25];
assign _012_ = addr_i[1] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ and_tree[26];
assign _013_ = _077_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ and_tree[27];
assign _014_ = addr_i[1] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ and_tree[28];
assign _015_ = _077_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ and_tree[29];
assign _016_ = addr_i[1] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ and_tree[30];
assign _017_ = _078_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ oh_i[0];
assign _018_ = addr_i[0] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ oh_i[1];
assign _019_ = _078_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ oh_i[2];
assign _020_ = addr_i[0] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ oh_i[3];
assign _021_ = _078_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ oh_i[4];
assign _022_ = addr_i[0] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ oh_i[5];
assign _023_ = _078_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ oh_i[6];
assign _024_ = addr_i[0] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ oh_i[7];
assign _025_ = _078_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ oh_i[8];
assign _026_ = addr_i[0] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ oh_i[9];
assign _027_ = _078_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ oh_i[10];
assign _028_ = addr_i[0] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ oh_i[11];
assign _029_ = _078_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ oh_i[12];
assign _030_ = addr_i[0] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ oh_i[13];
assign _031_ = _078_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ oh_i[14];
assign _032_ = addr_i[0] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ oh_i[15];
assign _033_ = _078_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ oh_i[16];
assign _034_ = addr_i[0] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ oh_i[17];
assign _035_ = _078_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ oh_i[18];
assign _036_ = addr_i[0] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ oh_i[19];
assign _037_ = _078_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ oh_i[20];
assign _038_ = addr_i[0] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ oh_i[21];
assign _039_ = _078_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ oh_i[22];
assign _040_ = addr_i[0] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ oh_i[23];
assign _041_ = _078_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ oh_i[24];
assign _042_ = addr_i[0] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ oh_i[25];
assign _043_ = _078_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ oh_i[26];
assign _044_ = addr_i[0] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ oh_i[27];
assign _045_ = _078_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ oh_i[28];
assign _046_ = addr_i[0] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ oh_i[29];
assign _047_ = _078_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ oh_i[30];
assign _048_ = addr_i[0] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ oh_i[31];
assign _049_ = _079_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ and_tree[1];
assign _050_ = addr_i[4] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ and_tree[2];
assign _051_ = _080_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ and_tree[3];
assign _052_ = addr_i[3] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ and_tree[4];
assign _053_ = _080_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ and_tree[5];
assign _054_ = addr_i[3] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ and_tree[6];
assign _055_ = _081_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ and_tree[7];
assign _056_ = addr_i[2] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ and_tree[8];
assign _057_ = _081_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ and_tree[9];
assign _058_ = addr_i[2] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ and_tree[10];
assign _059_ = _081_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ and_tree[11];
assign _060_ = addr_i[2] && /* src = "generated/sv2v_out.v:26515.83-26515.130" */ and_tree[12];
assign _061_ = _081_ && /* src = "generated/sv2v_out.v:26515.29-26515.77" */ and_tree[13];
assign _062_ = or_tree[13] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ or_tree[14];
assign _063_ = or_tree[15] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ or_tree[16];
assign _064_ = or_tree[17] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ or_tree[18];
assign _065_ = or_tree[19] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ or_tree[20];
assign _066_ = or_tree[21] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ or_tree[22];
assign _067_ = or_tree[23] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ or_tree[24];
assign _068_ = or_tree[25] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ or_tree[26];
assign _069_ = or_tree[27] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ or_tree[28];
assign _070_ = or_tree[29] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ or_tree[30];
assign err_tree[15] = oh_i[0] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ oh_i[1];
assign err_tree[16] = oh_i[2] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ oh_i[3];
assign err_tree[17] = oh_i[4] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ oh_i[5];
assign err_tree[18] = oh_i[6] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ oh_i[7];
assign err_tree[19] = oh_i[8] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ oh_i[9];
assign err_tree[20] = oh_i[10] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ oh_i[11];
assign err_tree[21] = oh_i[12] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ oh_i[13];
assign err_tree[22] = oh_i[14] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ oh_i[15];
assign err_tree[23] = oh_i[16] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ oh_i[17];
assign err_tree[24] = oh_i[18] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ oh_i[19];
assign err_tree[25] = oh_i[20] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ oh_i[21];
assign err_tree[26] = oh_i[22] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ oh_i[23];
assign err_tree[27] = oh_i[24] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ oh_i[25];
assign err_tree[28] = oh_i[26] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ oh_i[27];
assign err_tree[29] = oh_i[28] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ oh_i[29];
assign err_tree[30] = oh_i[30] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ oh_i[31];
assign _071_ = or_tree[1] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ or_tree[2];
assign _072_ = or_tree[3] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ or_tree[4];
assign _073_ = or_tree[5] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ or_tree[6];
assign _074_ = or_tree[7] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ or_tree[8];
assign _075_ = or_tree[9] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ or_tree[10];
assign _076_ = or_tree[11] && /* src = "generated/sv2v_out.v:26516.30-26516.56" */ or_tree[12];
assign _077_ = ! /* src = "generated/sv2v_out.v:26515.29-26515.61" */ addr_i[1];
assign _078_ = ! /* src = "generated/sv2v_out.v:26515.29-26515.61" */ addr_i[0];
assign _079_ = ! /* src = "generated/sv2v_out.v:26515.29-26515.61" */ addr_i[4];
assign _080_ = ! /* src = "generated/sv2v_out.v:26515.29-26515.61" */ addr_i[3];
assign _081_ = ! /* src = "generated/sv2v_out.v:26515.29-26515.61" */ addr_i[2];
assign or_tree[7] = or_tree[15] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ or_tree[16];
assign or_tree[8] = or_tree[17] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ or_tree[18];
assign or_tree[9] = or_tree[19] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ or_tree[20];
assign or_tree[10] = or_tree[21] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ or_tree[22];
assign or_tree[11] = or_tree[23] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ or_tree[24];
assign or_tree[12] = or_tree[25] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ or_tree[26];
assign or_tree[13] = or_tree[27] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ or_tree[28];
assign or_tree[14] = or_tree[29] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ or_tree[30];
assign or_tree[15] = oh_i[0] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ oh_i[1];
assign or_tree[16] = oh_i[2] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ oh_i[3];
assign or_tree[17] = oh_i[4] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ oh_i[5];
assign or_tree[18] = oh_i[6] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ oh_i[7];
assign or_tree[19] = oh_i[8] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ oh_i[9];
assign or_tree[20] = oh_i[10] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ oh_i[11];
assign or_tree[21] = oh_i[12] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ oh_i[13];
assign or_tree[22] = oh_i[14] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ oh_i[15];
assign or_tree[23] = oh_i[16] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ oh_i[17];
assign or_tree[24] = oh_i[18] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ oh_i[19];
assign or_tree[25] = oh_i[20] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ oh_i[21];
assign or_tree[26] = oh_i[22] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ oh_i[23];
assign or_tree[27] = oh_i[24] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ oh_i[25];
assign or_tree[28] = oh_i[26] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ oh_i[27];
assign or_tree[29] = oh_i[28] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ oh_i[29];
assign or_tree[30] = oh_i[30] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ oh_i[31];
assign or_tree[0] = or_tree[1] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ or_tree[2];
assign or_tree[1] = or_tree[3] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ or_tree[4];
assign or_tree[2] = or_tree[5] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ or_tree[6];
assign or_tree[3] = or_tree[7] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ or_tree[8];
assign or_tree[4] = or_tree[9] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ or_tree[10];
assign or_tree[5] = or_tree[11] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ or_tree[12];
assign or_tree[6] = or_tree[13] || /* src = "generated/sv2v_out.v:26514.27-26514.53" */ or_tree[14];
assign and_tree[6] = _061_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _000_;
assign and_tree[7] = _001_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _002_;
assign and_tree[8] = _003_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _004_;
assign and_tree[9] = _005_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _006_;
assign and_tree[10] = _007_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _008_;
assign and_tree[11] = _009_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _010_;
assign and_tree[12] = _011_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _012_;
assign and_tree[13] = _013_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _014_;
assign and_tree[14] = _015_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _016_;
assign and_tree[15] = _017_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _018_;
assign and_tree[16] = _019_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _020_;
assign and_tree[17] = _021_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _022_;
assign and_tree[18] = _023_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _024_;
assign and_tree[19] = _025_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _026_;
assign and_tree[20] = _027_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _028_;
assign and_tree[21] = _029_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _030_;
assign and_tree[22] = _031_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _032_;
assign and_tree[23] = _033_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _034_;
assign and_tree[24] = _035_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _036_;
assign and_tree[25] = _037_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _038_;
assign and_tree[26] = _039_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _040_;
assign and_tree[27] = _041_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _042_;
assign and_tree[28] = _043_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _044_;
assign and_tree[29] = _045_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _046_;
assign and_tree[30] = _047_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _048_;
assign and_tree[0] = _049_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _050_;
assign and_tree[1] = _051_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _052_;
assign and_tree[2] = _053_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _054_;
assign and_tree[3] = _055_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _056_;
assign and_tree[4] = _057_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _058_;
assign and_tree[5] = _059_ || /* src = "generated/sv2v_out.v:26515.28-26515.131" */ _060_;
assign _082_ = _062_ || /* src = "generated/sv2v_out.v:26516.29-26516.73" */ err_tree[13];
assign err_tree[6] = _082_ || /* src = "generated/sv2v_out.v:26516.28-26516.90" */ err_tree[14];
assign _083_ = _063_ || /* src = "generated/sv2v_out.v:26516.29-26516.73" */ err_tree[15];
assign err_tree[7] = _083_ || /* src = "generated/sv2v_out.v:26516.28-26516.90" */ err_tree[16];
assign _084_ = _064_ || /* src = "generated/sv2v_out.v:26516.29-26516.73" */ err_tree[17];
assign err_tree[8] = _084_ || /* src = "generated/sv2v_out.v:26516.28-26516.90" */ err_tree[18];
assign _085_ = _065_ || /* src = "generated/sv2v_out.v:26516.29-26516.73" */ err_tree[19];
assign err_tree[9] = _085_ || /* src = "generated/sv2v_out.v:26516.28-26516.90" */ err_tree[20];
assign _086_ = _066_ || /* src = "generated/sv2v_out.v:26516.29-26516.73" */ err_tree[21];
assign err_tree[10] = _086_ || /* src = "generated/sv2v_out.v:26516.28-26516.90" */ err_tree[22];
assign _087_ = _067_ || /* src = "generated/sv2v_out.v:26516.29-26516.73" */ err_tree[23];
assign err_tree[11] = _087_ || /* src = "generated/sv2v_out.v:26516.28-26516.90" */ err_tree[24];
assign _088_ = _068_ || /* src = "generated/sv2v_out.v:26516.29-26516.73" */ err_tree[25];
assign err_tree[12] = _088_ || /* src = "generated/sv2v_out.v:26516.28-26516.90" */ err_tree[26];
assign _089_ = _069_ || /* src = "generated/sv2v_out.v:26516.29-26516.73" */ err_tree[27];
assign err_tree[13] = _089_ || /* src = "generated/sv2v_out.v:26516.28-26516.90" */ err_tree[28];
assign _090_ = _070_ || /* src = "generated/sv2v_out.v:26516.29-26516.73" */ err_tree[29];
assign err_tree[14] = _090_ || /* src = "generated/sv2v_out.v:26516.28-26516.90" */ err_tree[30];
assign _091_ = _071_ || /* src = "generated/sv2v_out.v:26516.29-26516.73" */ err_tree[1];
assign oh0_err = _091_ || /* src = "generated/sv2v_out.v:26516.28-26516.90" */ err_tree[2];
assign _092_ = _072_ || /* src = "generated/sv2v_out.v:26516.29-26516.73" */ err_tree[3];
assign err_tree[1] = _092_ || /* src = "generated/sv2v_out.v:26516.28-26516.90" */ err_tree[4];
assign _093_ = _073_ || /* src = "generated/sv2v_out.v:26516.29-26516.73" */ err_tree[5];
assign err_tree[2] = _093_ || /* src = "generated/sv2v_out.v:26516.28-26516.90" */ err_tree[6];
assign _094_ = _074_ || /* src = "generated/sv2v_out.v:26516.29-26516.73" */ err_tree[7];
assign err_tree[3] = _094_ || /* src = "generated/sv2v_out.v:26516.28-26516.90" */ err_tree[8];
assign _095_ = _075_ || /* src = "generated/sv2v_out.v:26516.29-26516.73" */ err_tree[9];
assign err_tree[4] = _095_ || /* src = "generated/sv2v_out.v:26516.28-26516.90" */ err_tree[10];
assign _096_ = _076_ || /* src = "generated/sv2v_out.v:26516.29-26516.73" */ err_tree[11];
assign err_tree[5] = _096_ || /* src = "generated/sv2v_out.v:26516.28-26516.90" */ err_tree[12];
assign _097_ = oh0_err || /* src = "generated/sv2v_out.v:26524.18-26524.39" */ enable_err;
assign err_o = _097_ || /* src = "generated/sv2v_out.v:26524.17-26524.52" */ addr_err;
assign enable_err = or_tree[0] ^ /* src = "generated/sv2v_out.v:26529.25-26529.42" */ en_i;
assign addr_err = or_tree[0] ^ /* src = "generated/sv2v_out.v:26541.22-26541.46" */ and_tree[0];
assign and_tree[62:31] = oh_i;
assign err_o_t0 = 1'h0;
assign { err_tree[62:31], err_tree[0] } = { 32'h00000000, oh0_err };
assign or_tree[62:31] = oh_i;
endmodule

module \$paramod$9a435d8f6db004a67362aa9a56f32ea481a74dbe\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _0_;
wire [31:0] _1_;
wire [31:0] _2_;
wire [31:0] _3_;
/* src = "generated/sv2v_out.v:14894.13-14894.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14898.28-14898.37" */
output [31:0] rd_data_o;
reg [31:0] rd_data_o;
/* cellift = 32'd1 */
output [31:0] rd_data_o_t0;
reg [31:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14899.14-14899.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14895.13-14895.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14896.27-14896.36" */
input [31:0] wr_data_i;
wire [31:0] wr_data_i;
/* cellift = 32'd1 */
input [31:0] wr_data_i_t0;
wire [31:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14897.13-14897.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _0_ = ~ wr_en_i;
assign _1_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _2_ = { _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_ } & rd_data_o_t0;
assign _3_ = _1_ | _2_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$9a435d8f6db004a67362aa9a56f32ea481a74dbe\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 32'd0;
else rd_data_o_t0 <= _3_;
/* src = "generated/sv2v_out.v:14901.2-14905.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$9a435d8f6db004a67362aa9a56f32ea481a74dbe\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 32'd1073741827;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$a088b13b9337f1e1fba58a671f47d7c7701ffa49\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _0_;
wire [7:0] _1_;
wire [7:0] _2_;
wire [7:0] _3_;
/* src = "generated/sv2v_out.v:14894.13-14894.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14898.28-14898.37" */
output [7:0] rd_data_o;
reg [7:0] rd_data_o;
/* cellift = 32'd1 */
output [7:0] rd_data_o_t0;
reg [7:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14899.14-14899.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14895.13-14895.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14896.27-14896.36" */
input [7:0] wr_data_i;
wire [7:0] wr_data_i;
/* cellift = 32'd1 */
input [7:0] wr_data_i_t0;
wire [7:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14897.13-14897.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _0_ = ~ wr_en_i;
assign _1_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _2_ = { _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_ } & rd_data_o_t0;
assign _3_ = _1_ | _2_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a088b13b9337f1e1fba58a671f47d7c7701ffa49\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 8'h00;
else rd_data_o_t0 <= _3_;
/* src = "generated/sv2v_out.v:14901.2-14905.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a088b13b9337f1e1fba58a671f47d7c7701ffa49\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 8'h00;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$a308247794889ee6093207090edbf289adef8be1\ibex_ex_block (clk_i, rst_ni, alu_operator_i, alu_operand_a_i, alu_operand_b_i, alu_instr_first_cycle_i, bt_a_operand_i, bt_b_operand_i, multdiv_operator_i, mult_en_i, div_en_i, mult_sel_i, div_sel_i, multdiv_signed_mode_i, multdiv_operand_a_i, multdiv_operand_b_i, multdiv_ready_id_i, data_ind_timing_i, imd_val_we_o, imd_val_d_o, imd_val_q_i
, alu_adder_result_ex_o, result_ex_o, branch_target_o, branch_decision_o, ex_valid_o, ex_valid_o_t0, bt_b_operand_i_t0, bt_a_operand_i_t0, branch_target_o_t0, branch_decision_o_t0, alu_operand_b_i_t0, alu_instr_first_cycle_i_t0, div_en_i_t0, div_sel_i_t0, imd_val_d_o_t0, imd_val_q_i_t0, imd_val_we_o_t0, mult_en_i_t0, mult_sel_i_t0, multdiv_ready_id_i_t0, multdiv_operand_a_i_t0
, multdiv_operand_b_i_t0, alu_adder_result_ex_o_t0, alu_operator_i_t0, alu_operand_a_i_t0, result_ex_o_t0, multdiv_signed_mode_i_t0, multdiv_operator_i_t0, data_ind_timing_i_t0);
wire [33:0] _00_;
wire [1:0] _01_;
wire [31:0] _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire [33:0] _08_;
wire [33:0] _09_;
wire [33:0] _10_;
wire [33:0] _11_;
wire [1:0] _12_;
wire [1:0] _13_;
wire [31:0] _14_;
wire [31:0] _15_;
wire _16_;
/* src = "generated/sv2v_out.v:16080.53-16080.71" */
wire _17_;
/* src = "generated/sv2v_out.v:16080.55-16080.70" */
wire _18_;
/* src = "generated/sv2v_out.v:15960.21-15960.42" */
output [31:0] alu_adder_result_ex_o;
wire [31:0] alu_adder_result_ex_o;
/* cellift = 32'd1 */
output [31:0] alu_adder_result_ex_o_t0;
wire [31:0] alu_adder_result_ex_o_t0;
/* src = "generated/sv2v_out.v:15969.14-15969.34" */
wire [33:0] alu_adder_result_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15969.14-15969.34" */
wire [33:0] alu_adder_result_ext_t0;
/* src = "generated/sv2v_out.v:15975.14-15975.27" */
wire [63:0] alu_imd_val_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15975.14-15975.27" */
wire [63:0] alu_imd_val_d_t0;
/* src = "generated/sv2v_out.v:15976.13-15976.27" */
wire [1:0] alu_imd_val_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15976.13-15976.27" */
wire [1:0] alu_imd_val_we_t0;
/* src = "generated/sv2v_out.v:15944.13-15944.36" */
input alu_instr_first_cycle_i;
wire alu_instr_first_cycle_i;
/* cellift = 32'd1 */
input alu_instr_first_cycle_i_t0;
wire alu_instr_first_cycle_i_t0;
/* src = "generated/sv2v_out.v:15971.7-15971.26" */
wire alu_is_equal_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15971.7-15971.26" */
wire alu_is_equal_result_t0;
/* src = "generated/sv2v_out.v:15942.20-15942.35" */
input [31:0] alu_operand_a_i;
wire [31:0] alu_operand_a_i;
/* cellift = 32'd1 */
input [31:0] alu_operand_a_i_t0;
wire [31:0] alu_operand_a_i_t0;
/* src = "generated/sv2v_out.v:15943.20-15943.35" */
input [31:0] alu_operand_b_i;
wire [31:0] alu_operand_b_i;
/* cellift = 32'd1 */
input [31:0] alu_operand_b_i_t0;
wire [31:0] alu_operand_b_i_t0;
/* src = "generated/sv2v_out.v:15941.19-15941.33" */
input [6:0] alu_operator_i;
wire [6:0] alu_operator_i;
/* cellift = 32'd1 */
input [6:0] alu_operator_i_t0;
wire [6:0] alu_operator_i_t0;
/* src = "generated/sv2v_out.v:15965.14-15965.24" */
wire [31:0] alu_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15965.14-15965.24" */
wire [31:0] alu_result_t0;
/* src = "generated/sv2v_out.v:15963.14-15963.31" */
output branch_decision_o;
wire branch_decision_o;
/* cellift = 32'd1 */
output branch_decision_o_t0;
wire branch_decision_o_t0;
/* src = "generated/sv2v_out.v:15962.21-15962.36" */
output [31:0] branch_target_o;
wire [31:0] branch_target_o;
/* cellift = 32'd1 */
output [31:0] branch_target_o_t0;
wire [31:0] branch_target_o_t0;
/* src = "generated/sv2v_out.v:15945.20-15945.34" */
input [31:0] bt_a_operand_i;
wire [31:0] bt_a_operand_i;
/* cellift = 32'd1 */
input [31:0] bt_a_operand_i_t0;
wire [31:0] bt_a_operand_i_t0;
/* src = "generated/sv2v_out.v:15946.20-15946.34" */
input [31:0] bt_b_operand_i;
wire [31:0] bt_b_operand_i;
/* cellift = 32'd1 */
input [31:0] bt_b_operand_i_t0;
wire [31:0] bt_b_operand_i_t0;
/* src = "generated/sv2v_out.v:15939.13-15939.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:15956.13-15956.30" */
input data_ind_timing_i;
wire data_ind_timing_i;
/* cellift = 32'd1 */
input data_ind_timing_i_t0;
wire data_ind_timing_i_t0;
/* src = "generated/sv2v_out.v:15949.13-15949.21" */
input div_en_i;
wire div_en_i;
/* cellift = 32'd1 */
input div_en_i_t0;
wire div_en_i_t0;
/* src = "generated/sv2v_out.v:15951.13-15951.22" */
input div_sel_i;
wire div_sel_i;
/* cellift = 32'd1 */
input div_sel_i_t0;
wire div_sel_i_t0;
/* src = "generated/sv2v_out.v:15964.14-15964.24" */
output ex_valid_o;
wire ex_valid_o;
/* cellift = 32'd1 */
output ex_valid_o_t0;
wire ex_valid_o_t0;
/* src = "generated/sv2v_out.v:15958.21-15958.32" */
output [67:0] imd_val_d_o;
wire [67:0] imd_val_d_o;
/* cellift = 32'd1 */
output [67:0] imd_val_d_o_t0;
wire [67:0] imd_val_d_o_t0;
/* src = "generated/sv2v_out.v:15959.20-15959.31" */
input [67:0] imd_val_q_i;
wire [67:0] imd_val_q_i;
/* cellift = 32'd1 */
input [67:0] imd_val_q_i_t0;
wire [67:0] imd_val_q_i_t0;
/* src = "generated/sv2v_out.v:15957.20-15957.32" */
output [1:0] imd_val_we_o;
wire [1:0] imd_val_we_o;
/* cellift = 32'd1 */
output [1:0] imd_val_we_o_t0;
wire [1:0] imd_val_we_o_t0;
/* src = "generated/sv2v_out.v:15948.13-15948.22" */
input mult_en_i;
wire mult_en_i;
/* cellift = 32'd1 */
input mult_en_i_t0;
wire mult_en_i_t0;
/* src = "generated/sv2v_out.v:15950.13-15950.23" */
input mult_sel_i;
wire mult_sel_i;
/* cellift = 32'd1 */
input mult_sel_i_t0;
wire mult_sel_i_t0;
/* src = "generated/sv2v_out.v:15968.14-15968.35" */
wire [32:0] multdiv_alu_operand_a;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15968.14-15968.35" */
wire [32:0] multdiv_alu_operand_a_t0;
/* src = "generated/sv2v_out.v:15967.14-15967.35" */
wire [32:0] multdiv_alu_operand_b;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15967.14-15967.35" */
wire [32:0] multdiv_alu_operand_b_t0;
/* src = "generated/sv2v_out.v:15977.14-15977.31" */
wire [67:0] multdiv_imd_val_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15977.14-15977.31" */
wire [67:0] multdiv_imd_val_d_t0;
/* src = "generated/sv2v_out.v:15978.13-15978.31" */
wire [1:0] multdiv_imd_val_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15978.13-15978.31" */
wire [1:0] multdiv_imd_val_we_t0;
/* src = "generated/sv2v_out.v:15953.20-15953.39" */
input [31:0] multdiv_operand_a_i;
wire [31:0] multdiv_operand_a_i;
/* cellift = 32'd1 */
input [31:0] multdiv_operand_a_i_t0;
wire [31:0] multdiv_operand_a_i_t0;
/* src = "generated/sv2v_out.v:15954.20-15954.39" */
input [31:0] multdiv_operand_b_i;
wire [31:0] multdiv_operand_b_i;
/* cellift = 32'd1 */
input [31:0] multdiv_operand_b_i_t0;
wire [31:0] multdiv_operand_b_i_t0;
/* src = "generated/sv2v_out.v:15947.19-15947.37" */
input [1:0] multdiv_operator_i;
wire [1:0] multdiv_operator_i;
/* cellift = 32'd1 */
input [1:0] multdiv_operator_i_t0;
wire [1:0] multdiv_operator_i_t0;
/* src = "generated/sv2v_out.v:15955.13-15955.31" */
input multdiv_ready_id_i;
wire multdiv_ready_id_i;
/* cellift = 32'd1 */
input multdiv_ready_id_i_t0;
wire multdiv_ready_id_i_t0;
/* src = "generated/sv2v_out.v:15966.14-15966.28" */
wire [31:0] multdiv_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15966.14-15966.28" */
wire [31:0] multdiv_result_t0;
/* src = "generated/sv2v_out.v:15973.7-15973.18" */
wire multdiv_sel;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15973.7-15973.18" */
wire multdiv_sel_t0;
/* src = "generated/sv2v_out.v:15952.19-15952.40" */
input [1:0] multdiv_signed_mode_i;
wire [1:0] multdiv_signed_mode_i;
/* cellift = 32'd1 */
input [1:0] multdiv_signed_mode_i_t0;
wire [1:0] multdiv_signed_mode_i_t0;
/* src = "generated/sv2v_out.v:15972.7-15972.20" */
wire multdiv_valid;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15972.7-15972.20" */
wire multdiv_valid_t0;
/* src = "generated/sv2v_out.v:15961.21-15961.32" */
output [31:0] result_ex_o;
wire [31:0] result_ex_o;
/* cellift = 32'd1 */
output [31:0] result_ex_o_t0;
wire [31:0] result_ex_o_t0;
/* src = "generated/sv2v_out.v:15940.13-15940.19" */
input rst_ni;
wire rst_ni;
assign _00_ = ~ { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel };
assign _01_ = ~ { multdiv_sel, multdiv_sel };
assign _02_ = ~ { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel };
assign _08_ = _00_ & { 2'h0, alu_imd_val_d_t0[63:32] };
assign _10_ = _00_ & { 2'h0, alu_imd_val_d_t0[31:0] };
assign _12_ = _01_ & alu_imd_val_we_t0;
assign _14_ = _02_ & alu_result_t0;
assign _09_ = { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel } & multdiv_imd_val_d_t0[67:34];
assign _11_ = { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel } & multdiv_imd_val_d_t0[33:0];
assign _13_ = { multdiv_sel, multdiv_sel } & multdiv_imd_val_we_t0;
assign _15_ = { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel } & multdiv_result_t0;
assign ex_valid_o_t0 = multdiv_sel & multdiv_valid_t0;
assign imd_val_d_o_t0[67:34] = _08_ | _09_;
assign imd_val_d_o_t0[33:0] = _10_ | _11_;
assign imd_val_we_o_t0 = _12_ | _13_;
assign result_ex_o_t0 = _14_ | _15_;
assign _03_ = ~ mult_sel_i;
assign _04_ = ~ div_sel_i;
assign _05_ = mult_sel_i_t0 & _04_;
assign _06_ = div_sel_i_t0 & _03_;
assign _07_ = mult_sel_i_t0 & div_sel_i_t0;
assign _16_ = _05_ | _06_;
assign multdiv_sel_t0 = _16_ | _07_;
assign _17_ = ~ /* src = "generated/sv2v_out.v:16080.53-16080.71" */ _18_;
assign multdiv_sel = mult_sel_i | /* src = "generated/sv2v_out.v:15981.25-15981.47" */ div_sel_i;
assign _18_ = | /* src = "generated/sv2v_out.v:16080.55-16080.70" */ alu_imd_val_we;
assign imd_val_d_o[67:34] = multdiv_sel ? /* src = "generated/sv2v_out.v:15987.32-15987.104" */ multdiv_imd_val_d[67:34] : { 2'h0, alu_imd_val_d[63:32] };
assign imd_val_d_o[33:0] = multdiv_sel ? /* src = "generated/sv2v_out.v:15988.31-15988.101" */ multdiv_imd_val_d[33:0] : { 2'h0, alu_imd_val_d[31:0] };
assign imd_val_we_o = multdiv_sel ? /* src = "generated/sv2v_out.v:15989.25-15989.74" */ multdiv_imd_val_we : alu_imd_val_we;
assign result_ex_o = multdiv_sel ? /* src = "generated/sv2v_out.v:15991.24-15991.65" */ multdiv_result : alu_result;
assign ex_valid_o = multdiv_sel ? /* src = "generated/sv2v_out.v:16080.23-16080.71" */ multdiv_valid : _17_;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:16009.28-16025.3" */
\$paramod\ibex_alu\RV32B=s32'00000000000000000000000000000000  alu_i (
.adder_result_ext_o(alu_adder_result_ext),
.adder_result_ext_o_t0(alu_adder_result_ext_t0),
.adder_result_o(alu_adder_result_ex_o),
.adder_result_o_t0(alu_adder_result_ex_o_t0),
.comparison_result_o(branch_decision_o),
.comparison_result_o_t0(branch_decision_o_t0),
.imd_val_d_o(alu_imd_val_d),
.imd_val_d_o_t0(alu_imd_val_d_t0),
.imd_val_q_i({ imd_val_q_i[65:34], imd_val_q_i[31:0] }),
.imd_val_q_i_t0({ imd_val_q_i_t0[65:34], imd_val_q_i_t0[31:0] }),
.imd_val_we_o(alu_imd_val_we),
.imd_val_we_o_t0(alu_imd_val_we_t0),
.instr_first_cycle_i(alu_instr_first_cycle_i),
.instr_first_cycle_i_t0(alu_instr_first_cycle_i_t0),
.is_equal_result_o(alu_is_equal_result),
.is_equal_result_o_t0(alu_is_equal_result_t0),
.multdiv_operand_a_i(multdiv_alu_operand_a),
.multdiv_operand_a_i_t0(multdiv_alu_operand_a_t0),
.multdiv_operand_b_i(multdiv_alu_operand_b),
.multdiv_operand_b_i_t0(multdiv_alu_operand_b_t0),
.multdiv_sel_i(multdiv_sel),
.multdiv_sel_i_t0(multdiv_sel_t0),
.operand_a_i(alu_operand_a_i),
.operand_a_i_t0(alu_operand_a_i_t0),
.operand_b_i(alu_operand_b_i),
.operand_b_i_t0(alu_operand_b_i_t0),
.operator_i(alu_operator_i),
.operator_i_t0(alu_operator_i_t0),
.result_o(alu_result),
.result_o_t0(alu_result_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:16028.22-16051.5" */
ibex_multdiv_slow \gen_multdiv_slow.multdiv_i  (
.alu_adder_ext_i(alu_adder_result_ext),
.alu_adder_ext_i_t0(alu_adder_result_ext_t0),
.alu_adder_i(alu_adder_result_ex_o),
.alu_adder_i_t0(alu_adder_result_ex_o_t0),
.alu_operand_a_o(multdiv_alu_operand_a),
.alu_operand_a_o_t0(multdiv_alu_operand_a_t0),
.alu_operand_b_o(multdiv_alu_operand_b),
.alu_operand_b_o_t0(multdiv_alu_operand_b_t0),
.clk_i(clk_i),
.data_ind_timing_i(data_ind_timing_i),
.data_ind_timing_i_t0(data_ind_timing_i_t0),
.div_en_i(div_en_i),
.div_en_i_t0(div_en_i_t0),
.div_sel_i(div_sel_i),
.div_sel_i_t0(div_sel_i_t0),
.equal_to_zero_i(alu_is_equal_result),
.equal_to_zero_i_t0(alu_is_equal_result_t0),
.imd_val_d_o(multdiv_imd_val_d),
.imd_val_d_o_t0(multdiv_imd_val_d_t0),
.imd_val_q_i(imd_val_q_i),
.imd_val_q_i_t0(imd_val_q_i_t0),
.imd_val_we_o(multdiv_imd_val_we),
.imd_val_we_o_t0(multdiv_imd_val_we_t0),
.mult_en_i(mult_en_i),
.mult_en_i_t0(mult_en_i_t0),
.mult_sel_i(mult_sel_i),
.mult_sel_i_t0(mult_sel_i_t0),
.multdiv_ready_id_i(multdiv_ready_id_i),
.multdiv_ready_id_i_t0(multdiv_ready_id_i_t0),
.multdiv_result_o(multdiv_result),
.multdiv_result_o_t0(multdiv_result_t0),
.op_a_i(multdiv_operand_a_i),
.op_a_i_t0(multdiv_operand_a_i_t0),
.op_b_i(multdiv_operand_b_i),
.op_b_i_t0(multdiv_operand_b_i_t0),
.operator_i(multdiv_operator_i),
.operator_i_t0(multdiv_operator_i_t0),
.rst_ni(rst_ni),
.signed_mode_i(multdiv_signed_mode_i),
.signed_mode_i_t0(multdiv_signed_mode_i_t0),
.valid_o(multdiv_valid),
.valid_o_t0(multdiv_valid_t0)
);
assign branch_target_o = alu_adder_result_ex_o;
assign branch_target_o_t0 = alu_adder_result_ex_o_t0;
endmodule

module \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff (clk_i, rst_ni, test_en_i, dummy_instr_id_i, dummy_instr_wb_i, raddr_a_i, rdata_a_o, raddr_b_i, rdata_b_o, waddr_a_i, wdata_a_i, we_a_i, err_o, test_en_i_t0, err_o_t0, dummy_instr_id_i_t0, dummy_instr_wb_i_t0, raddr_a_i_t0, raddr_b_i_t0, rdata_a_o_t0, rdata_b_o_t0
, waddr_a_i_t0, wdata_a_i_t0, we_a_i_t0);
wire _0000_;
wire _0001_;
wire _0002_;
wire _0003_;
wire _0004_;
wire _0005_;
wire _0006_;
wire _0007_;
wire _0008_;
wire _0009_;
wire _0010_;
wire _0011_;
wire _0012_;
wire _0013_;
wire _0014_;
wire _0015_;
wire _0016_;
wire _0017_;
wire _0018_;
wire _0019_;
wire _0020_;
wire _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire _0026_;
wire _0027_;
wire _0028_;
wire _0029_;
wire _0030_;
wire _0031_;
wire [38:0] _0032_;
wire [38:0] _0033_;
wire [38:0] _0034_;
wire [38:0] _0035_;
wire [38:0] _0036_;
wire [38:0] _0037_;
wire [38:0] _0038_;
wire [38:0] _0039_;
wire [38:0] _0040_;
wire [38:0] _0041_;
wire [38:0] _0042_;
wire [38:0] _0043_;
wire [38:0] _0044_;
wire [38:0] _0045_;
wire [38:0] _0046_;
wire [38:0] _0047_;
wire [38:0] _0048_;
wire [38:0] _0049_;
wire [38:0] _0050_;
wire [38:0] _0051_;
wire [38:0] _0052_;
wire [38:0] _0053_;
wire [38:0] _0054_;
wire [38:0] _0055_;
wire [38:0] _0056_;
wire [38:0] _0057_;
wire [38:0] _0058_;
wire [38:0] _0059_;
wire [38:0] _0060_;
wire [38:0] _0061_;
wire [38:0] _0062_;
wire [38:0] _0063_;
wire [38:0] _0064_;
wire [38:0] _0065_;
wire [38:0] _0066_;
wire [38:0] _0067_;
wire [38:0] _0068_;
wire [38:0] _0069_;
wire [38:0] _0070_;
wire [38:0] _0071_;
wire [38:0] _0072_;
wire [38:0] _0073_;
wire [38:0] _0074_;
wire [38:0] _0075_;
wire [38:0] _0076_;
wire [38:0] _0077_;
wire [38:0] _0078_;
wire [38:0] _0079_;
wire [38:0] _0080_;
wire [38:0] _0081_;
wire [38:0] _0082_;
wire [38:0] _0083_;
wire [38:0] _0084_;
wire [38:0] _0085_;
wire [38:0] _0086_;
wire [38:0] _0087_;
wire [38:0] _0088_;
wire [38:0] _0089_;
wire [38:0] _0090_;
wire [38:0] _0091_;
wire [38:0] _0092_;
wire [38:0] _0093_;
wire _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire [38:0] _0108_;
wire [38:0] _0109_;
wire [38:0] _0110_;
wire [38:0] _0111_;
wire [38:0] _0112_;
wire [38:0] _0113_;
wire [38:0] _0114_;
wire [38:0] _0115_;
wire [38:0] _0116_;
wire [38:0] _0117_;
wire [38:0] _0118_;
wire [38:0] _0119_;
wire [38:0] _0120_;
wire [38:0] _0121_;
wire [38:0] _0122_;
wire [38:0] _0123_;
wire [38:0] _0124_;
wire [38:0] _0125_;
wire [38:0] _0126_;
wire [38:0] _0127_;
wire [38:0] _0128_;
wire [38:0] _0129_;
wire [38:0] _0130_;
wire [38:0] _0131_;
wire [38:0] _0132_;
wire [38:0] _0133_;
wire [38:0] _0134_;
wire [38:0] _0135_;
wire [38:0] _0136_;
wire [38:0] _0137_;
wire [38:0] _0138_;
wire [38:0] _0139_;
wire [38:0] _0140_;
wire [38:0] _0141_;
wire [38:0] _0142_;
wire [38:0] _0143_;
wire [38:0] _0144_;
wire [38:0] _0145_;
wire [38:0] _0146_;
wire [38:0] _0147_;
wire [38:0] _0148_;
wire [38:0] _0149_;
wire [38:0] _0150_;
wire [38:0] _0151_;
wire [38:0] _0152_;
wire [38:0] _0153_;
wire [38:0] _0154_;
wire [38:0] _0155_;
wire [38:0] _0156_;
wire [38:0] _0157_;
wire [38:0] _0158_;
wire [38:0] _0159_;
wire [38:0] _0160_;
wire [38:0] _0161_;
wire [38:0] _0162_;
wire [38:0] _0163_;
wire [38:0] _0164_;
wire [38:0] _0165_;
wire [38:0] _0166_;
wire [38:0] _0167_;
wire [38:0] _0168_;
wire [38:0] _0169_;
wire [38:0] _0170_;
wire [38:0] _0171_;
wire [38:0] _0172_;
wire [38:0] _0173_;
wire [38:0] _0174_;
wire [38:0] _0175_;
wire [38:0] _0176_;
wire [38:0] _0177_;
wire [38:0] _0178_;
wire [38:0] _0179_;
wire [38:0] _0180_;
wire [38:0] _0181_;
wire [38:0] _0182_;
wire [38:0] _0183_;
wire [38:0] _0184_;
wire [38:0] _0185_;
wire [38:0] _0186_;
wire [38:0] _0187_;
wire [38:0] _0188_;
wire [38:0] _0189_;
wire [38:0] _0190_;
wire [38:0] _0191_;
wire [38:0] _0192_;
wire [38:0] _0193_;
wire [38:0] _0194_;
wire [38:0] _0195_;
wire [38:0] _0196_;
wire [38:0] _0197_;
wire [38:0] _0198_;
wire [38:0] _0199_;
wire [38:0] _0200_;
wire [38:0] _0201_;
wire [38:0] _0202_;
wire [38:0] _0203_;
wire [38:0] _0204_;
wire [38:0] _0205_;
wire [38:0] _0206_;
wire [38:0] _0207_;
wire [38:0] _0208_;
wire [38:0] _0209_;
wire [38:0] _0210_;
wire [38:0] _0211_;
wire [38:0] _0212_;
wire [38:0] _0213_;
wire [38:0] _0214_;
wire [38:0] _0215_;
wire [38:0] _0216_;
wire [38:0] _0217_;
wire [38:0] _0218_;
wire [38:0] _0219_;
wire [38:0] _0220_;
wire [38:0] _0221_;
wire [38:0] _0222_;
wire [38:0] _0223_;
wire [38:0] _0224_;
wire [38:0] _0225_;
wire [38:0] _0226_;
wire [38:0] _0227_;
wire [38:0] _0228_;
wire [38:0] _0229_;
wire [38:0] _0230_;
wire [38:0] _0231_;
wire [38:0] _0232_;
wire [38:0] _0233_;
wire [38:0] _0234_;
wire [38:0] _0235_;
wire [38:0] _0236_;
wire [38:0] _0237_;
wire [38:0] _0238_;
wire [38:0] _0239_;
wire [38:0] _0240_;
wire [38:0] _0241_;
wire [38:0] _0242_;
wire [38:0] _0243_;
wire [38:0] _0244_;
wire [38:0] _0245_;
wire [38:0] _0246_;
wire [38:0] _0247_;
wire [38:0] _0248_;
wire [38:0] _0249_;
wire [38:0] _0250_;
wire [38:0] _0251_;
wire [38:0] _0252_;
wire [38:0] _0253_;
wire [38:0] _0254_;
wire [38:0] _0255_;
wire [38:0] _0256_;
wire [38:0] _0257_;
wire [38:0] _0258_;
wire [38:0] _0259_;
wire [38:0] _0260_;
wire [38:0] _0261_;
wire [38:0] _0262_;
wire [38:0] _0263_;
wire [38:0] _0264_;
wire [38:0] _0265_;
wire [38:0] _0266_;
wire [38:0] _0267_;
wire [38:0] _0268_;
wire [38:0] _0269_;
wire [38:0] _0270_;
wire [38:0] _0271_;
wire [38:0] _0272_;
wire [38:0] _0273_;
wire [38:0] _0274_;
wire [38:0] _0275_;
wire [38:0] _0276_;
wire [38:0] _0277_;
wire [38:0] _0278_;
wire [38:0] _0279_;
wire [38:0] _0280_;
wire [38:0] _0281_;
wire [38:0] _0282_;
wire [38:0] _0283_;
wire [38:0] _0284_;
wire [38:0] _0285_;
wire [38:0] _0286_;
wire [38:0] _0287_;
wire [38:0] _0288_;
wire [38:0] _0289_;
wire [38:0] _0290_;
wire [38:0] _0291_;
wire [38:0] _0292_;
wire [38:0] _0293_;
wire [38:0] _0294_;
wire [38:0] _0295_;
wire [38:0] _0296_;
wire [38:0] _0297_;
wire [38:0] _0298_;
wire [38:0] _0299_;
wire [38:0] _0300_;
wire [38:0] _0301_;
wire [38:0] _0302_;
wire [38:0] _0303_;
wire [38:0] _0304_;
wire [38:0] _0305_;
wire [38:0] _0306_;
wire [38:0] _0307_;
wire [38:0] _0308_;
wire [38:0] _0309_;
wire [38:0] _0310_;
wire [38:0] _0311_;
wire [38:0] _0312_;
wire [38:0] _0313_;
wire [38:0] _0314_;
wire [38:0] _0315_;
wire [38:0] _0316_;
wire [38:0] _0317_;
wire [38:0] _0318_;
wire [38:0] _0319_;
wire [38:0] _0320_;
wire [38:0] _0321_;
wire [38:0] _0322_;
wire [38:0] _0323_;
wire [38:0] _0324_;
wire [38:0] _0325_;
wire [38:0] _0326_;
wire [38:0] _0327_;
wire _0328_;
wire _0329_;
wire _0330_;
wire _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire _0335_;
wire _0336_;
wire _0337_;
wire _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire [38:0] _0344_;
/* cellift = 32'd1 */
wire [38:0] _0345_;
wire [38:0] _0346_;
/* cellift = 32'd1 */
wire [38:0] _0347_;
wire [38:0] _0348_;
/* cellift = 32'd1 */
wire [38:0] _0349_;
wire [38:0] _0350_;
/* cellift = 32'd1 */
wire [38:0] _0351_;
wire [38:0] _0352_;
/* cellift = 32'd1 */
wire [38:0] _0353_;
wire [38:0] _0354_;
/* cellift = 32'd1 */
wire [38:0] _0355_;
wire [38:0] _0356_;
/* cellift = 32'd1 */
wire [38:0] _0357_;
wire [38:0] _0358_;
/* cellift = 32'd1 */
wire [38:0] _0359_;
wire [38:0] _0360_;
/* cellift = 32'd1 */
wire [38:0] _0361_;
wire [38:0] _0362_;
/* cellift = 32'd1 */
wire [38:0] _0363_;
wire [38:0] _0364_;
/* cellift = 32'd1 */
wire [38:0] _0365_;
wire [38:0] _0366_;
/* cellift = 32'd1 */
wire [38:0] _0367_;
wire [38:0] _0368_;
/* cellift = 32'd1 */
wire [38:0] _0369_;
wire [38:0] _0370_;
/* cellift = 32'd1 */
wire [38:0] _0371_;
wire [38:0] _0372_;
/* cellift = 32'd1 */
wire [38:0] _0373_;
wire [38:0] _0374_;
/* cellift = 32'd1 */
wire [38:0] _0375_;
wire [38:0] _0376_;
/* cellift = 32'd1 */
wire [38:0] _0377_;
wire [38:0] _0378_;
/* cellift = 32'd1 */
wire [38:0] _0379_;
wire [38:0] _0380_;
/* cellift = 32'd1 */
wire [38:0] _0381_;
wire [38:0] _0382_;
/* cellift = 32'd1 */
wire [38:0] _0383_;
wire [38:0] _0384_;
/* cellift = 32'd1 */
wire [38:0] _0385_;
wire [38:0] _0386_;
/* cellift = 32'd1 */
wire [38:0] _0387_;
wire [38:0] _0388_;
/* cellift = 32'd1 */
wire [38:0] _0389_;
wire [38:0] _0390_;
/* cellift = 32'd1 */
wire [38:0] _0391_;
wire [38:0] _0392_;
/* cellift = 32'd1 */
wire [38:0] _0393_;
wire [38:0] _0394_;
/* cellift = 32'd1 */
wire [38:0] _0395_;
wire [38:0] _0396_;
/* cellift = 32'd1 */
wire [38:0] _0397_;
wire [38:0] _0398_;
/* cellift = 32'd1 */
wire [38:0] _0399_;
wire [38:0] _0400_;
/* cellift = 32'd1 */
wire [38:0] _0401_;
wire [38:0] _0402_;
/* cellift = 32'd1 */
wire [38:0] _0403_;
wire [38:0] _0404_;
/* cellift = 32'd1 */
wire [38:0] _0405_;
wire [38:0] _0406_;
/* cellift = 32'd1 */
wire [38:0] _0407_;
wire [38:0] _0408_;
/* cellift = 32'd1 */
wire [38:0] _0409_;
wire [38:0] _0410_;
/* cellift = 32'd1 */
wire [38:0] _0411_;
wire [38:0] _0412_;
/* cellift = 32'd1 */
wire [38:0] _0413_;
wire [38:0] _0414_;
/* cellift = 32'd1 */
wire [38:0] _0415_;
wire [38:0] _0416_;
/* cellift = 32'd1 */
wire [38:0] _0417_;
wire [38:0] _0418_;
/* cellift = 32'd1 */
wire [38:0] _0419_;
wire [38:0] _0420_;
/* cellift = 32'd1 */
wire [38:0] _0421_;
wire [38:0] _0422_;
/* cellift = 32'd1 */
wire [38:0] _0423_;
wire [38:0] _0424_;
/* cellift = 32'd1 */
wire [38:0] _0425_;
wire [38:0] _0426_;
/* cellift = 32'd1 */
wire [38:0] _0427_;
wire [38:0] _0428_;
/* cellift = 32'd1 */
wire [38:0] _0429_;
wire [38:0] _0430_;
/* cellift = 32'd1 */
wire [38:0] _0431_;
wire [38:0] _0432_;
/* cellift = 32'd1 */
wire [38:0] _0433_;
wire [38:0] _0434_;
/* cellift = 32'd1 */
wire [38:0] _0435_;
wire [38:0] _0436_;
/* cellift = 32'd1 */
wire [38:0] _0437_;
wire [38:0] _0438_;
/* cellift = 32'd1 */
wire [38:0] _0439_;
wire [38:0] _0440_;
/* cellift = 32'd1 */
wire [38:0] _0441_;
wire [38:0] _0442_;
/* cellift = 32'd1 */
wire [38:0] _0443_;
wire [38:0] _0444_;
/* cellift = 32'd1 */
wire [38:0] _0445_;
wire [38:0] _0446_;
/* cellift = 32'd1 */
wire [38:0] _0447_;
wire [38:0] _0448_;
/* cellift = 32'd1 */
wire [38:0] _0449_;
wire [38:0] _0450_;
/* cellift = 32'd1 */
wire [38:0] _0451_;
wire [38:0] _0452_;
/* cellift = 32'd1 */
wire [38:0] _0453_;
wire [38:0] _0454_;
/* cellift = 32'd1 */
wire [38:0] _0455_;
wire [38:0] _0456_;
/* cellift = 32'd1 */
wire [38:0] _0457_;
wire [38:0] _0458_;
/* cellift = 32'd1 */
wire [38:0] _0459_;
wire [38:0] _0460_;
/* cellift = 32'd1 */
wire [38:0] _0461_;
wire [38:0] _0462_;
/* cellift = 32'd1 */
wire [38:0] _0463_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0464_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0465_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0466_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0467_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0468_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0469_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0470_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0471_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0472_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0473_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0474_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0475_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0476_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0477_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0478_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0479_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0480_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0481_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0482_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0483_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0484_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0485_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0486_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0487_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0488_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0489_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0490_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0491_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0492_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0493_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0494_;
/* src = "generated/sv2v_out.v:20105.20-20105.47" */
wire _0495_;
wire _0496_;
wire _0497_;
wire _0498_;
wire _0499_;
wire _0500_;
wire _0501_;
wire _0502_;
wire _0503_;
wire _0504_;
wire _0505_;
wire _0506_;
wire _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0517_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
wire _0525_;
wire _0526_;
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire _0534_;
wire _0535_;
wire _0536_;
wire _0537_;
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0542_;
wire _0543_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
/* src = "generated/sv2v_out.v:20080.13-20080.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:20083.13-20083.29" */
input dummy_instr_id_i;
wire dummy_instr_id_i;
/* cellift = 32'd1 */
input dummy_instr_id_i_t0;
wire dummy_instr_id_i_t0;
/* src = "generated/sv2v_out.v:20084.13-20084.29" */
input dummy_instr_wb_i;
wire dummy_instr_wb_i;
/* cellift = 32'd1 */
input dummy_instr_wb_i_t0;
wire dummy_instr_wb_i_t0;
/* src = "generated/sv2v_out.v:20092.14-20092.19" */
output err_o;
wire err_o;
/* cellift = 32'd1 */
output err_o_t0;
wire err_o_t0;
/* src = "generated/sv2v_out.v:20147.26-20147.33" */
reg [38:0] \g_dummy_r0.rf_r0_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20147.26-20147.33" */
reg [38:0] \g_dummy_r0.rf_r0_q_t0 ;
/* src = "generated/sv2v_out.v:20146.9-20146.20" */
wire \g_dummy_r0.we_r0_dummy ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[10].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[10].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[11].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[11].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[12].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[12].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[13].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[13].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[14].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[14].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[15].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[15].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[16].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[16].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[17].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[17].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[18].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[18].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[19].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[19].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[1].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[1].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[20].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[20].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[21].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[21].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[22].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[22].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[23].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[23].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[24].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[24].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[25].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[25].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[26].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[26].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[27].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[27].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[28].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[28].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[29].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[29].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[2].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[2].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[30].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[30].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[31].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[31].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[3].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[3].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[4].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[4].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[5].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[5].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[6].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[6].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[7].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[7].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[8].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[8].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[9].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20137.26-20137.34" */
reg [38:0] \g_rf_flops[9].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20110.27-20110.39" */
wire [31:0] \gen_wren_check.we_a_dec_buf ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20110.27-20110.39" */
wire [31:0] \gen_wren_check.we_a_dec_buf_t0 ;
/* src = "generated/sv2v_out.v:20085.19-20085.28" */
input [4:0] raddr_a_i;
wire [4:0] raddr_a_i;
/* cellift = 32'd1 */
input [4:0] raddr_a_i_t0;
wire [4:0] raddr_a_i_t0;
/* src = "generated/sv2v_out.v:20087.19-20087.28" */
input [4:0] raddr_b_i;
wire [4:0] raddr_b_i;
/* cellift = 32'd1 */
input [4:0] raddr_b_i_t0;
wire [4:0] raddr_b_i_t0;
/* src = "generated/sv2v_out.v:20086.32-20086.41" */
output [38:0] rdata_a_o;
wire [38:0] rdata_a_o;
/* cellift = 32'd1 */
output [38:0] rdata_a_o_t0;
wire [38:0] rdata_a_o_t0;
/* src = "generated/sv2v_out.v:20088.32-20088.41" */
output [38:0] rdata_b_o;
wire [38:0] rdata_b_o;
/* cellift = 32'd1 */
output [38:0] rdata_b_o_t0;
wire [38:0] rdata_b_o_t0;
/* src = "generated/sv2v_out.v:20095.25-20095.31" */
wire [38:0] \rf_reg[0] ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20095.25-20095.31" */
wire [38:0] \rf_reg[0]_t0 ;
/* src = "generated/sv2v_out.v:20081.13-20081.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:20082.13-20082.22" */
input test_en_i;
wire test_en_i;
/* cellift = 32'd1 */
input test_en_i_t0;
wire test_en_i_t0;
/* src = "generated/sv2v_out.v:20089.19-20089.28" */
input [4:0] waddr_a_i;
wire [4:0] waddr_a_i;
/* cellift = 32'd1 */
input [4:0] waddr_a_i_t0;
wire [4:0] waddr_a_i_t0;
/* src = "generated/sv2v_out.v:20090.31-20090.40" */
input [38:0] wdata_a_i;
wire [38:0] wdata_a_i;
/* cellift = 32'd1 */
input [38:0] wdata_a_i_t0;
wire [38:0] wdata_a_i_t0;
/* src = "generated/sv2v_out.v:20096.24-20096.32" */
wire [31:0] we_a_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20096.24-20096.32" */
wire [31:0] we_a_dec_t0;
/* src = "generated/sv2v_out.v:20091.13-20091.19" */
input we_a_i;
wire we_a_i;
/* cellift = 32'd1 */
input we_a_i_t0;
wire we_a_i_t0;
assign \g_dummy_r0.we_r0_dummy  = we_a_i & /* src = "generated/sv2v_out.v:20148.25-20148.50" */ dummy_instr_wb_i;
assign _0000_ = ~ we_a_dec[31];
assign _0001_ = ~ we_a_dec[30];
assign _0002_ = ~ we_a_dec[29];
assign _0003_ = ~ we_a_dec[28];
assign _0004_ = ~ we_a_dec[27];
assign _0005_ = ~ we_a_dec[26];
assign _0006_ = ~ we_a_dec[25];
assign _0007_ = ~ we_a_dec[24];
assign _0008_ = ~ we_a_dec[23];
assign _0009_ = ~ we_a_dec[22];
assign _0010_ = ~ we_a_dec[21];
assign _0011_ = ~ we_a_dec[20];
assign _0012_ = ~ we_a_dec[19];
assign _0013_ = ~ we_a_dec[18];
assign _0014_ = ~ we_a_dec[17];
assign _0015_ = ~ we_a_dec[16];
assign _0016_ = ~ we_a_dec[15];
assign _0017_ = ~ we_a_dec[14];
assign _0018_ = ~ we_a_dec[13];
assign _0019_ = ~ we_a_dec[12];
assign _0020_ = ~ we_a_dec[11];
assign _0021_ = ~ we_a_dec[10];
assign _0022_ = ~ we_a_dec[9];
assign _0023_ = ~ we_a_dec[8];
assign _0024_ = ~ we_a_dec[7];
assign _0025_ = ~ we_a_dec[6];
assign _0026_ = ~ we_a_dec[5];
assign _0027_ = ~ we_a_dec[4];
assign _0028_ = ~ we_a_dec[3];
assign _0029_ = ~ we_a_dec[2];
assign _0030_ = ~ we_a_dec[1];
assign _0031_ = ~ \g_dummy_r0.we_r0_dummy ;
assign _0108_ = { we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31] } & wdata_a_i_t0;
assign _0110_ = { we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30] } & wdata_a_i_t0;
assign _0112_ = { we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29] } & wdata_a_i_t0;
assign _0114_ = { we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28] } & wdata_a_i_t0;
assign _0116_ = { we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27] } & wdata_a_i_t0;
assign _0118_ = { we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26] } & wdata_a_i_t0;
assign _0120_ = { we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25] } & wdata_a_i_t0;
assign _0122_ = { we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24] } & wdata_a_i_t0;
assign _0124_ = { we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23] } & wdata_a_i_t0;
assign _0126_ = { we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22] } & wdata_a_i_t0;
assign _0128_ = { we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21] } & wdata_a_i_t0;
assign _0130_ = { we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20] } & wdata_a_i_t0;
assign _0132_ = { we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19] } & wdata_a_i_t0;
assign _0134_ = { we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18] } & wdata_a_i_t0;
assign _0136_ = { we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17] } & wdata_a_i_t0;
assign _0138_ = { we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16] } & wdata_a_i_t0;
assign _0140_ = { we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15] } & wdata_a_i_t0;
assign _0142_ = { we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14] } & wdata_a_i_t0;
assign _0144_ = { we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13] } & wdata_a_i_t0;
assign _0146_ = { we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12] } & wdata_a_i_t0;
assign _0148_ = { we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11] } & wdata_a_i_t0;
assign _0150_ = { we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10] } & wdata_a_i_t0;
assign _0152_ = { we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9] } & wdata_a_i_t0;
assign _0154_ = { we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8] } & wdata_a_i_t0;
assign _0156_ = { we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7] } & wdata_a_i_t0;
assign _0158_ = { we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6] } & wdata_a_i_t0;
assign _0160_ = { we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5] } & wdata_a_i_t0;
assign _0162_ = { we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4] } & wdata_a_i_t0;
assign _0164_ = { we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3] } & wdata_a_i_t0;
assign _0166_ = { we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2] } & wdata_a_i_t0;
assign _0168_ = { we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1] } & wdata_a_i_t0;
assign _0170_ = { \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy  } & wdata_a_i_t0;
assign _0109_ = { _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_ } & \g_rf_flops[31].rf_reg_q_t0 ;
assign _0111_ = { _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_ } & \g_rf_flops[30].rf_reg_q_t0 ;
assign _0113_ = { _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_ } & \g_rf_flops[29].rf_reg_q_t0 ;
assign _0115_ = { _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_ } & \g_rf_flops[28].rf_reg_q_t0 ;
assign _0117_ = { _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_ } & \g_rf_flops[27].rf_reg_q_t0 ;
assign _0119_ = { _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_ } & \g_rf_flops[26].rf_reg_q_t0 ;
assign _0121_ = { _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_ } & \g_rf_flops[25].rf_reg_q_t0 ;
assign _0123_ = { _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_ } & \g_rf_flops[24].rf_reg_q_t0 ;
assign _0125_ = { _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_ } & \g_rf_flops[23].rf_reg_q_t0 ;
assign _0127_ = { _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_ } & \g_rf_flops[22].rf_reg_q_t0 ;
assign _0129_ = { _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_ } & \g_rf_flops[21].rf_reg_q_t0 ;
assign _0131_ = { _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_ } & \g_rf_flops[20].rf_reg_q_t0 ;
assign _0133_ = { _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_ } & \g_rf_flops[19].rf_reg_q_t0 ;
assign _0135_ = { _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_ } & \g_rf_flops[18].rf_reg_q_t0 ;
assign _0137_ = { _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_ } & \g_rf_flops[17].rf_reg_q_t0 ;
assign _0139_ = { _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_ } & \g_rf_flops[16].rf_reg_q_t0 ;
assign _0141_ = { _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_ } & \g_rf_flops[15].rf_reg_q_t0 ;
assign _0143_ = { _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_ } & \g_rf_flops[14].rf_reg_q_t0 ;
assign _0145_ = { _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_ } & \g_rf_flops[13].rf_reg_q_t0 ;
assign _0147_ = { _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_ } & \g_rf_flops[12].rf_reg_q_t0 ;
assign _0149_ = { _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_ } & \g_rf_flops[11].rf_reg_q_t0 ;
assign _0151_ = { _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_ } & \g_rf_flops[10].rf_reg_q_t0 ;
assign _0153_ = { _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_ } & \g_rf_flops[9].rf_reg_q_t0 ;
assign _0155_ = { _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_ } & \g_rf_flops[8].rf_reg_q_t0 ;
assign _0157_ = { _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_ } & \g_rf_flops[7].rf_reg_q_t0 ;
assign _0159_ = { _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_ } & \g_rf_flops[6].rf_reg_q_t0 ;
assign _0161_ = { _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_ } & \g_rf_flops[5].rf_reg_q_t0 ;
assign _0163_ = { _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_ } & \g_rf_flops[4].rf_reg_q_t0 ;
assign _0165_ = { _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_ } & \g_rf_flops[3].rf_reg_q_t0 ;
assign _0167_ = { _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_ } & \g_rf_flops[2].rf_reg_q_t0 ;
assign _0169_ = { _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_ } & \g_rf_flops[1].rf_reg_q_t0 ;
assign _0171_ = { _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_ } & \g_dummy_r0.rf_r0_q_t0 ;
assign _0296_ = _0108_ | _0109_;
assign _0297_ = _0110_ | _0111_;
assign _0298_ = _0112_ | _0113_;
assign _0299_ = _0114_ | _0115_;
assign _0300_ = _0116_ | _0117_;
assign _0301_ = _0118_ | _0119_;
assign _0302_ = _0120_ | _0121_;
assign _0303_ = _0122_ | _0123_;
assign _0304_ = _0124_ | _0125_;
assign _0305_ = _0126_ | _0127_;
assign _0306_ = _0128_ | _0129_;
assign _0307_ = _0130_ | _0131_;
assign _0308_ = _0132_ | _0133_;
assign _0309_ = _0134_ | _0135_;
assign _0310_ = _0136_ | _0137_;
assign _0311_ = _0138_ | _0139_;
assign _0312_ = _0140_ | _0141_;
assign _0313_ = _0142_ | _0143_;
assign _0314_ = _0144_ | _0145_;
assign _0315_ = _0146_ | _0147_;
assign _0316_ = _0148_ | _0149_;
assign _0317_ = _0150_ | _0151_;
assign _0318_ = _0152_ | _0153_;
assign _0319_ = _0154_ | _0155_;
assign _0320_ = _0156_ | _0157_;
assign _0321_ = _0158_ | _0159_;
assign _0322_ = _0160_ | _0161_;
assign _0323_ = _0162_ | _0163_;
assign _0324_ = _0164_ | _0165_;
assign _0325_ = _0166_ | _0167_;
assign _0326_ = _0168_ | _0169_;
assign _0327_ = _0170_ | _0171_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[31].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[31].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[31].rf_reg_q_t0  <= _0296_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[30].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[30].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[30].rf_reg_q_t0  <= _0297_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[29].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[29].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[29].rf_reg_q_t0  <= _0298_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[28].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[28].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[28].rf_reg_q_t0  <= _0299_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[27].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[27].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[27].rf_reg_q_t0  <= _0300_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[26].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[26].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[26].rf_reg_q_t0  <= _0301_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[25].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[25].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[25].rf_reg_q_t0  <= _0302_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[24].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[24].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[24].rf_reg_q_t0  <= _0303_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[23].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[23].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[23].rf_reg_q_t0  <= _0304_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[22].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[22].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[22].rf_reg_q_t0  <= _0305_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[21].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[21].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[21].rf_reg_q_t0  <= _0306_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[20].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[20].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[20].rf_reg_q_t0  <= _0307_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[19].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[19].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[19].rf_reg_q_t0  <= _0308_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[18].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[18].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[18].rf_reg_q_t0  <= _0309_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[17].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[17].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[17].rf_reg_q_t0  <= _0310_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[16].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[16].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[16].rf_reg_q_t0  <= _0311_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[15].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[15].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[15].rf_reg_q_t0  <= _0312_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[14].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[14].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[14].rf_reg_q_t0  <= _0313_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[13].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[13].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[13].rf_reg_q_t0  <= _0314_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[12].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[12].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[12].rf_reg_q_t0  <= _0315_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[11].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[11].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[11].rf_reg_q_t0  <= _0316_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[10].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[10].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[10].rf_reg_q_t0  <= _0317_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[9].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[9].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[9].rf_reg_q_t0  <= _0318_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[8].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[8].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[8].rf_reg_q_t0  <= _0319_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[7].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[7].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[7].rf_reg_q_t0  <= _0320_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[6].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[6].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[6].rf_reg_q_t0  <= _0321_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[5].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[5].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[5].rf_reg_q_t0  <= _0322_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[4].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[4].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[4].rf_reg_q_t0  <= _0323_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[3].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[3].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[3].rf_reg_q_t0  <= _0324_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[2].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[2].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[2].rf_reg_q_t0  <= _0325_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[1].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[1].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[1].rf_reg_q_t0  <= _0326_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_dummy_r0.rf_r0_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_dummy_r0.rf_r0_q_t0  <= 39'h0000000000;
else \g_dummy_r0.rf_r0_q_t0  <= _0327_;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[31].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[31].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[31]) \g_rf_flops[31].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[30].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[30].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[30]) \g_rf_flops[30].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[29].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[29].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[29]) \g_rf_flops[29].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[28].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[28].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[28]) \g_rf_flops[28].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[27].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[27].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[27]) \g_rf_flops[27].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[26].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[26].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[26]) \g_rf_flops[26].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[25].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[25].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[25]) \g_rf_flops[25].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[24].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[24].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[24]) \g_rf_flops[24].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[23].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[23].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[23]) \g_rf_flops[23].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[22].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[22].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[22]) \g_rf_flops[22].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[21].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[21].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[21]) \g_rf_flops[21].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[20].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[20].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[20]) \g_rf_flops[20].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[19].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[19].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[19]) \g_rf_flops[19].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[18].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[18].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[18]) \g_rf_flops[18].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[17].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[17].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[17]) \g_rf_flops[17].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[16].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[16].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[16]) \g_rf_flops[16].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[15].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[15].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[15]) \g_rf_flops[15].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[14].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[14].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[14]) \g_rf_flops[14].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[13].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[13].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[13]) \g_rf_flops[13].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[12].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[12].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[12]) \g_rf_flops[12].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[11].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[11].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[11]) \g_rf_flops[11].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[10].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[10].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[10]) \g_rf_flops[10].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[9].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[9].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[9]) \g_rf_flops[9].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[8].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[8].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[8]) \g_rf_flops[8].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[7].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[7].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[7]) \g_rf_flops[7].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[6].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[6].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[6]) \g_rf_flops[6].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[5].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[5].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[5]) \g_rf_flops[5].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[4].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[4].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[4]) \g_rf_flops[4].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[3].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[3].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[3]) \g_rf_flops[3].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[2].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[2].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[2]) \g_rf_flops[2].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20138.4-20142.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[1].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[1].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[1]) \g_rf_flops[1].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20149.4-20153.27" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_dummy_r0.rf_r0_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_dummy_r0.rf_r0_q  <= 39'h2a00000000;
else if (\g_dummy_r0.we_r0_dummy ) \g_dummy_r0.rf_r0_q  <= wdata_a_i;
assign _0032_ = ~ { _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_ };
assign _0033_ = ~ { _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_ };
assign _0034_ = ~ { _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_ };
assign _0035_ = ~ { _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_ };
assign _0036_ = ~ { _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_ };
assign _0037_ = ~ { _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_ };
assign _0038_ = ~ { _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_ };
assign _0039_ = ~ { _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_ };
assign _0040_ = ~ { _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_ };
assign _0041_ = ~ { _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_ };
assign _0042_ = ~ { _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_ };
assign _0043_ = ~ { _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_ };
assign _0044_ = ~ { _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_ };
assign _0045_ = ~ { _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_ };
assign _0046_ = ~ { _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_ };
assign _0047_ = ~ { _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_ };
assign _0048_ = ~ { _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_ };
assign _0049_ = ~ { _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_ };
assign _0050_ = ~ { _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_ };
assign _0051_ = ~ { _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_ };
assign _0052_ = ~ { _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_ };
assign _0053_ = ~ { _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_ };
assign _0054_ = ~ { _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_ };
assign _0055_ = ~ { _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_ };
assign _0056_ = ~ { _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_ };
assign _0057_ = ~ { _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_ };
assign _0058_ = ~ { _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_ };
assign _0059_ = ~ { _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_ };
assign _0060_ = ~ { _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_ };
assign _0061_ = ~ { _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_ };
assign _0062_ = ~ { _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_ };
assign _0063_ = ~ { _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_ };
assign _0064_ = ~ { _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_ };
assign _0065_ = ~ { _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_ };
assign _0066_ = ~ { _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_ };
assign _0067_ = ~ { _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_ };
assign _0068_ = ~ { _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_ };
assign _0069_ = ~ { _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_ };
assign _0070_ = ~ { _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_ };
assign _0071_ = ~ { _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_ };
assign _0072_ = ~ { _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_ };
assign _0073_ = ~ { _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_ };
assign _0074_ = ~ { _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_ };
assign _0075_ = ~ { _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_ };
assign _0076_ = ~ { _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_ };
assign _0077_ = ~ { _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_ };
assign _0078_ = ~ { _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_ };
assign _0079_ = ~ { _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_ };
assign _0080_ = ~ { _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_ };
assign _0081_ = ~ { _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_ };
assign _0082_ = ~ { _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_ };
assign _0083_ = ~ { _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_ };
assign _0084_ = ~ { _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_ };
assign _0085_ = ~ { _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_ };
assign _0086_ = ~ { _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_ };
assign _0087_ = ~ { _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_ };
assign _0088_ = ~ { _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_ };
assign _0089_ = ~ { _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_ };
assign _0090_ = ~ { _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_ };
assign _0091_ = ~ { _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_ };
assign _0092_ = ~ { _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_ };
assign _0093_ = ~ { _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_ };
assign _0172_ = _0032_ & \g_rf_flops[30].rf_reg_q_t0 ;
assign _0174_ = _0033_ & \g_rf_flops[28].rf_reg_q_t0 ;
assign _0176_ = _0034_ & _0347_;
assign _0178_ = _0035_ & \g_rf_flops[26].rf_reg_q_t0 ;
assign _0180_ = _0036_ & \g_rf_flops[24].rf_reg_q_t0 ;
assign _0182_ = _0037_ & _0353_;
assign _0184_ = _0038_ & _0355_;
assign _0186_ = _0039_ & \g_rf_flops[22].rf_reg_q_t0 ;
assign _0188_ = _0040_ & \g_rf_flops[20].rf_reg_q_t0 ;
assign _0190_ = _0041_ & _0361_;
assign _0192_ = _0042_ & \g_rf_flops[18].rf_reg_q_t0 ;
assign _0194_ = _0043_ & \g_rf_flops[16].rf_reg_q_t0 ;
assign _0196_ = _0044_ & _0367_;
assign _0198_ = _0045_ & _0369_;
assign _0200_ = _0046_ & _0371_;
assign _0202_ = _0047_ & \g_rf_flops[14].rf_reg_q_t0 ;
assign _0204_ = _0048_ & \g_rf_flops[12].rf_reg_q_t0 ;
assign _0206_ = _0049_ & _0377_;
assign _0208_ = _0050_ & \g_rf_flops[10].rf_reg_q_t0 ;
assign _0210_ = _0051_ & \g_rf_flops[8].rf_reg_q_t0 ;
assign _0212_ = _0052_ & _0383_;
assign _0214_ = _0053_ & _0385_;
assign _0216_ = _0054_ & \g_rf_flops[6].rf_reg_q_t0 ;
assign _0218_ = _0055_ & \g_rf_flops[4].rf_reg_q_t0 ;
assign _0220_ = _0056_ & _0391_;
assign _0222_ = _0057_ & \g_rf_flops[2].rf_reg_q_t0 ;
assign _0224_ = _0058_ & \rf_reg[0]_t0 ;
assign _0226_ = _0059_ & _0397_;
assign _0228_ = _0060_ & _0399_;
assign _0230_ = _0061_ & _0401_;
assign _0232_ = _0062_ & _0403_;
assign _0234_ = _0063_ & \g_rf_flops[30].rf_reg_q_t0 ;
assign _0236_ = _0064_ & \g_rf_flops[28].rf_reg_q_t0 ;
assign _0238_ = _0065_ & _0407_;
assign _0240_ = _0066_ & \g_rf_flops[26].rf_reg_q_t0 ;
assign _0242_ = _0067_ & \g_rf_flops[24].rf_reg_q_t0 ;
assign _0244_ = _0068_ & _0413_;
assign _0246_ = _0069_ & _0415_;
assign _0248_ = _0070_ & \g_rf_flops[22].rf_reg_q_t0 ;
assign _0250_ = _0071_ & \g_rf_flops[20].rf_reg_q_t0 ;
assign _0252_ = _0072_ & _0421_;
assign _0254_ = _0073_ & \g_rf_flops[18].rf_reg_q_t0 ;
assign _0256_ = _0074_ & \g_rf_flops[16].rf_reg_q_t0 ;
assign _0258_ = _0075_ & _0427_;
assign _0260_ = _0076_ & _0429_;
assign _0262_ = _0077_ & _0431_;
assign _0264_ = _0078_ & \g_rf_flops[14].rf_reg_q_t0 ;
assign _0266_ = _0079_ & \g_rf_flops[12].rf_reg_q_t0 ;
assign _0268_ = _0080_ & _0437_;
assign _0270_ = _0081_ & \g_rf_flops[10].rf_reg_q_t0 ;
assign _0272_ = _0082_ & \g_rf_flops[8].rf_reg_q_t0 ;
assign _0274_ = _0083_ & _0443_;
assign _0276_ = _0084_ & _0445_;
assign _0278_ = _0085_ & \g_rf_flops[6].rf_reg_q_t0 ;
assign _0280_ = _0086_ & \g_rf_flops[4].rf_reg_q_t0 ;
assign _0282_ = _0087_ & _0451_;
assign _0284_ = _0088_ & \g_rf_flops[2].rf_reg_q_t0 ;
assign _0286_ = _0089_ & \rf_reg[0]_t0 ;
assign _0288_ = _0090_ & _0457_;
assign _0290_ = _0091_ & _0459_;
assign _0292_ = _0092_ & _0461_;
assign _0294_ = _0093_ & _0463_;
assign _0173_ = { _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_ } & \g_rf_flops[31].rf_reg_q_t0 ;
assign _0175_ = { _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_ } & \g_rf_flops[29].rf_reg_q_t0 ;
assign _0177_ = { _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_, _0328_ } & _0345_;
assign _0179_ = { _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_ } & \g_rf_flops[27].rf_reg_q_t0 ;
assign _0181_ = { _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_ } & \g_rf_flops[25].rf_reg_q_t0 ;
assign _0183_ = { _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_, _0329_ } & _0351_;
assign _0185_ = { _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_ } & _0349_;
assign _0187_ = { _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_ } & \g_rf_flops[23].rf_reg_q_t0 ;
assign _0189_ = { _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_ } & \g_rf_flops[21].rf_reg_q_t0 ;
assign _0191_ = { _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_, _0330_ } & _0359_;
assign _0193_ = { _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_ } & \g_rf_flops[19].rf_reg_q_t0 ;
assign _0195_ = { _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_ } & \g_rf_flops[17].rf_reg_q_t0 ;
assign _0197_ = { _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_, _0331_ } & _0365_;
assign _0199_ = { _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_ } & _0363_;
assign _0201_ = { _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_ } & _0357_;
assign _0203_ = { _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_ } & \g_rf_flops[15].rf_reg_q_t0 ;
assign _0205_ = { _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_ } & \g_rf_flops[13].rf_reg_q_t0 ;
assign _0207_ = { _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_, _0332_ } & _0375_;
assign _0209_ = { _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_ } & \g_rf_flops[11].rf_reg_q_t0 ;
assign _0211_ = { _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_ } & \g_rf_flops[9].rf_reg_q_t0 ;
assign _0213_ = { _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_, _0333_ } & _0381_;
assign _0215_ = { _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_ } & _0379_;
assign _0217_ = { _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_ } & \g_rf_flops[7].rf_reg_q_t0 ;
assign _0219_ = { _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_ } & \g_rf_flops[5].rf_reg_q_t0 ;
assign _0221_ = { _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_, _0334_ } & _0389_;
assign _0223_ = { _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_ } & \g_rf_flops[3].rf_reg_q_t0 ;
assign _0225_ = { _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_ } & \g_rf_flops[1].rf_reg_q_t0 ;
assign _0227_ = { _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_, _0335_ } & _0395_;
assign _0229_ = { _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_ } & _0393_;
assign _0231_ = { _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_ } & _0387_;
assign _0233_ = { _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_ } & _0373_;
assign _0235_ = { _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_ } & \g_rf_flops[31].rf_reg_q_t0 ;
assign _0237_ = { _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_ } & \g_rf_flops[29].rf_reg_q_t0 ;
assign _0239_ = { _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_, _0336_ } & _0405_;
assign _0241_ = { _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_ } & \g_rf_flops[27].rf_reg_q_t0 ;
assign _0243_ = { _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_ } & \g_rf_flops[25].rf_reg_q_t0 ;
assign _0245_ = { _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_, _0337_ } & _0411_;
assign _0247_ = { _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_ } & _0409_;
assign _0249_ = { _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_ } & \g_rf_flops[23].rf_reg_q_t0 ;
assign _0251_ = { _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_ } & \g_rf_flops[21].rf_reg_q_t0 ;
assign _0253_ = { _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_, _0338_ } & _0419_;
assign _0255_ = { _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_ } & \g_rf_flops[19].rf_reg_q_t0 ;
assign _0257_ = { _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_ } & \g_rf_flops[17].rf_reg_q_t0 ;
assign _0259_ = { _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_, _0339_ } & _0425_;
assign _0261_ = { _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_ } & _0423_;
assign _0263_ = { _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_ } & _0417_;
assign _0265_ = { _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_ } & \g_rf_flops[15].rf_reg_q_t0 ;
assign _0267_ = { _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_ } & \g_rf_flops[13].rf_reg_q_t0 ;
assign _0269_ = { _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_, _0340_ } & _0435_;
assign _0271_ = { _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_ } & \g_rf_flops[11].rf_reg_q_t0 ;
assign _0273_ = { _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_ } & \g_rf_flops[9].rf_reg_q_t0 ;
assign _0275_ = { _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_, _0341_ } & _0441_;
assign _0277_ = { _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_ } & _0439_;
assign _0279_ = { _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_ } & \g_rf_flops[7].rf_reg_q_t0 ;
assign _0281_ = { _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_ } & \g_rf_flops[5].rf_reg_q_t0 ;
assign _0283_ = { _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_ } & _0449_;
assign _0285_ = { _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_ } & \g_rf_flops[3].rf_reg_q_t0 ;
assign _0287_ = { _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_ } & \g_rf_flops[1].rf_reg_q_t0 ;
assign _0289_ = { _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_ } & _0455_;
assign _0291_ = { _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_ } & _0453_;
assign _0293_ = { _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_ } & _0447_;
assign _0295_ = { _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_ } & _0433_;
assign we_a_dec_t0[0] = _0464_ & we_a_i_t0;
assign we_a_dec_t0[1] = _0465_ & we_a_i_t0;
assign we_a_dec_t0[2] = _0466_ & we_a_i_t0;
assign we_a_dec_t0[3] = _0467_ & we_a_i_t0;
assign we_a_dec_t0[4] = _0468_ & we_a_i_t0;
assign we_a_dec_t0[5] = _0469_ & we_a_i_t0;
assign we_a_dec_t0[6] = _0470_ & we_a_i_t0;
assign we_a_dec_t0[7] = _0471_ & we_a_i_t0;
assign we_a_dec_t0[8] = _0472_ & we_a_i_t0;
assign we_a_dec_t0[9] = _0473_ & we_a_i_t0;
assign we_a_dec_t0[10] = _0474_ & we_a_i_t0;
assign we_a_dec_t0[11] = _0475_ & we_a_i_t0;
assign we_a_dec_t0[12] = _0476_ & we_a_i_t0;
assign we_a_dec_t0[13] = _0477_ & we_a_i_t0;
assign we_a_dec_t0[14] = _0478_ & we_a_i_t0;
assign we_a_dec_t0[15] = _0479_ & we_a_i_t0;
assign we_a_dec_t0[16] = _0480_ & we_a_i_t0;
assign we_a_dec_t0[17] = _0481_ & we_a_i_t0;
assign we_a_dec_t0[18] = _0482_ & we_a_i_t0;
assign we_a_dec_t0[19] = _0483_ & we_a_i_t0;
assign we_a_dec_t0[20] = _0484_ & we_a_i_t0;
assign we_a_dec_t0[21] = _0485_ & we_a_i_t0;
assign we_a_dec_t0[22] = _0486_ & we_a_i_t0;
assign we_a_dec_t0[23] = _0487_ & we_a_i_t0;
assign we_a_dec_t0[24] = _0488_ & we_a_i_t0;
assign we_a_dec_t0[25] = _0489_ & we_a_i_t0;
assign we_a_dec_t0[26] = _0490_ & we_a_i_t0;
assign we_a_dec_t0[27] = _0491_ & we_a_i_t0;
assign we_a_dec_t0[28] = _0492_ & we_a_i_t0;
assign we_a_dec_t0[29] = _0493_ & we_a_i_t0;
assign we_a_dec_t0[30] = _0494_ & we_a_i_t0;
assign we_a_dec_t0[31] = _0495_ & we_a_i_t0;
assign \rf_reg[0]_t0  = { dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i } & \g_dummy_r0.rf_r0_q_t0 ;
assign _0345_ = _0172_ | _0173_;
assign _0347_ = _0174_ | _0175_;
assign _0349_ = _0176_ | _0177_;
assign _0351_ = _0178_ | _0179_;
assign _0353_ = _0180_ | _0181_;
assign _0355_ = _0182_ | _0183_;
assign _0357_ = _0184_ | _0185_;
assign _0359_ = _0186_ | _0187_;
assign _0361_ = _0188_ | _0189_;
assign _0363_ = _0190_ | _0191_;
assign _0365_ = _0192_ | _0193_;
assign _0367_ = _0194_ | _0195_;
assign _0369_ = _0196_ | _0197_;
assign _0371_ = _0198_ | _0199_;
assign _0373_ = _0200_ | _0201_;
assign _0375_ = _0202_ | _0203_;
assign _0377_ = _0204_ | _0205_;
assign _0379_ = _0206_ | _0207_;
assign _0381_ = _0208_ | _0209_;
assign _0383_ = _0210_ | _0211_;
assign _0385_ = _0212_ | _0213_;
assign _0387_ = _0214_ | _0215_;
assign _0389_ = _0216_ | _0217_;
assign _0391_ = _0218_ | _0219_;
assign _0393_ = _0220_ | _0221_;
assign _0395_ = _0222_ | _0223_;
assign _0397_ = _0224_ | _0225_;
assign _0399_ = _0226_ | _0227_;
assign _0401_ = _0228_ | _0229_;
assign _0403_ = _0230_ | _0231_;
assign rdata_b_o_t0 = _0232_ | _0233_;
assign _0405_ = _0234_ | _0235_;
assign _0407_ = _0236_ | _0237_;
assign _0409_ = _0238_ | _0239_;
assign _0411_ = _0240_ | _0241_;
assign _0413_ = _0242_ | _0243_;
assign _0415_ = _0244_ | _0245_;
assign _0417_ = _0246_ | _0247_;
assign _0419_ = _0248_ | _0249_;
assign _0421_ = _0250_ | _0251_;
assign _0423_ = _0252_ | _0253_;
assign _0425_ = _0254_ | _0255_;
assign _0427_ = _0256_ | _0257_;
assign _0429_ = _0258_ | _0259_;
assign _0431_ = _0260_ | _0261_;
assign _0433_ = _0262_ | _0263_;
assign _0435_ = _0264_ | _0265_;
assign _0437_ = _0266_ | _0267_;
assign _0439_ = _0268_ | _0269_;
assign _0441_ = _0270_ | _0271_;
assign _0443_ = _0272_ | _0273_;
assign _0445_ = _0274_ | _0275_;
assign _0447_ = _0276_ | _0277_;
assign _0449_ = _0278_ | _0279_;
assign _0451_ = _0280_ | _0281_;
assign _0453_ = _0282_ | _0283_;
assign _0455_ = _0284_ | _0285_;
assign _0457_ = _0286_ | _0287_;
assign _0459_ = _0288_ | _0289_;
assign _0461_ = _0290_ | _0291_;
assign _0463_ = _0292_ | _0293_;
assign rdata_a_o_t0 = _0294_ | _0295_;
assign _0328_ = _0497_ | _0496_;
assign _0329_ = _0501_ | _0500_;
assign _0330_ = _0505_ | _0504_;
assign _0331_ = _0509_ | _0508_;
assign _0332_ = _0513_ | _0512_;
assign _0333_ = _0517_ | _0516_;
assign _0334_ = _0521_ | _0520_;
assign _0335_ = _0525_ | _0524_;
assign _0336_ = _0528_ | _0527_;
assign _0337_ = _0532_ | _0531_;
assign _0338_ = _0536_ | _0535_;
assign _0339_ = _0540_ | _0539_;
assign _0340_ = _0544_ | _0543_;
assign _0341_ = _0548_ | _0547_;
assign _0342_ = _0552_ | _0551_;
assign _0343_ = _0556_ | _0555_;
assign _0094_ = | { _0328_, _0499_, _0498_ };
assign _0095_ = | { _0330_, _0507_, _0506_ };
assign _0096_ = | { _0328_, _0329_, _0503_, _0502_, _0499_, _0498_ };
assign _0097_ = | { _0332_, _0515_, _0514_ };
assign _0098_ = | { _0334_, _0523_, _0522_ };
assign _0099_ = | { _0332_, _0333_, _0519_, _0518_, _0515_, _0514_ };
assign _0100_ = | { _0328_, _0329_, _0330_, _0331_, _0510_, _0511_, _0507_, _0506_, _0503_, _0502_, _0499_, _0498_ };
assign _0101_ = | { _0336_, _0529_, _0530_ };
assign _0102_ = | { _0338_, _0538_, _0537_ };
assign _0103_ = | { _0336_, _0337_, _0534_, _0533_, _0529_, _0530_ };
assign _0104_ = | { _0340_, _0546_, _0545_ };
assign _0105_ = | { _0342_, _0554_, _0553_ };
assign _0106_ = | { _0340_, _0341_, _0550_, _0549_, _0546_, _0545_ };
assign _0107_ = | { _0336_, _0337_, _0338_, _0339_, _0542_, _0541_, _0538_, _0537_, _0534_, _0533_, _0529_, _0530_ };
assign _0344_ = _0496_ ? \g_rf_flops[31].rf_reg_q  : \g_rf_flops[30].rf_reg_q ;
assign _0346_ = _0498_ ? \g_rf_flops[29].rf_reg_q  : \g_rf_flops[28].rf_reg_q ;
assign _0348_ = _0328_ ? _0344_ : _0346_;
assign _0350_ = _0500_ ? \g_rf_flops[27].rf_reg_q  : \g_rf_flops[26].rf_reg_q ;
assign _0352_ = _0502_ ? \g_rf_flops[25].rf_reg_q  : \g_rf_flops[24].rf_reg_q ;
assign _0354_ = _0329_ ? _0350_ : _0352_;
assign _0356_ = _0094_ ? _0348_ : _0354_;
assign _0358_ = _0504_ ? \g_rf_flops[23].rf_reg_q  : \g_rf_flops[22].rf_reg_q ;
assign _0360_ = _0506_ ? \g_rf_flops[21].rf_reg_q  : \g_rf_flops[20].rf_reg_q ;
assign _0362_ = _0330_ ? _0358_ : _0360_;
assign _0364_ = _0508_ ? \g_rf_flops[19].rf_reg_q  : \g_rf_flops[18].rf_reg_q ;
assign _0366_ = _0510_ ? \g_rf_flops[17].rf_reg_q  : \g_rf_flops[16].rf_reg_q ;
assign _0368_ = _0331_ ? _0364_ : _0366_;
assign _0370_ = _0095_ ? _0362_ : _0368_;
assign _0372_ = _0096_ ? _0356_ : _0370_;
assign _0374_ = _0512_ ? \g_rf_flops[15].rf_reg_q  : \g_rf_flops[14].rf_reg_q ;
assign _0376_ = _0514_ ? \g_rf_flops[13].rf_reg_q  : \g_rf_flops[12].rf_reg_q ;
assign _0378_ = _0332_ ? _0374_ : _0376_;
assign _0380_ = _0516_ ? \g_rf_flops[11].rf_reg_q  : \g_rf_flops[10].rf_reg_q ;
assign _0382_ = _0518_ ? \g_rf_flops[9].rf_reg_q  : \g_rf_flops[8].rf_reg_q ;
assign _0384_ = _0333_ ? _0380_ : _0382_;
assign _0386_ = _0097_ ? _0378_ : _0384_;
assign _0388_ = _0520_ ? \g_rf_flops[7].rf_reg_q  : \g_rf_flops[6].rf_reg_q ;
assign _0390_ = _0522_ ? \g_rf_flops[5].rf_reg_q  : \g_rf_flops[4].rf_reg_q ;
assign _0392_ = _0334_ ? _0388_ : _0390_;
assign _0394_ = _0524_ ? \g_rf_flops[3].rf_reg_q  : \g_rf_flops[2].rf_reg_q ;
assign _0396_ = _0526_ ? \g_rf_flops[1].rf_reg_q  : \rf_reg[0] ;
assign _0398_ = _0335_ ? _0394_ : _0396_;
assign _0400_ = _0098_ ? _0392_ : _0398_;
assign _0402_ = _0099_ ? _0386_ : _0400_;
assign rdata_b_o = _0100_ ? _0372_ : _0402_;
assign _0404_ = _0527_ ? \g_rf_flops[31].rf_reg_q  : \g_rf_flops[30].rf_reg_q ;
assign _0406_ = _0529_ ? \g_rf_flops[29].rf_reg_q  : \g_rf_flops[28].rf_reg_q ;
assign _0408_ = _0336_ ? _0404_ : _0406_;
assign _0410_ = _0531_ ? \g_rf_flops[27].rf_reg_q  : \g_rf_flops[26].rf_reg_q ;
assign _0412_ = _0533_ ? \g_rf_flops[25].rf_reg_q  : \g_rf_flops[24].rf_reg_q ;
assign _0414_ = _0337_ ? _0410_ : _0412_;
assign _0416_ = _0101_ ? _0408_ : _0414_;
assign _0418_ = _0535_ ? \g_rf_flops[23].rf_reg_q  : \g_rf_flops[22].rf_reg_q ;
assign _0420_ = _0537_ ? \g_rf_flops[21].rf_reg_q  : \g_rf_flops[20].rf_reg_q ;
assign _0422_ = _0338_ ? _0418_ : _0420_;
assign _0424_ = _0539_ ? \g_rf_flops[19].rf_reg_q  : \g_rf_flops[18].rf_reg_q ;
assign _0426_ = _0541_ ? \g_rf_flops[17].rf_reg_q  : \g_rf_flops[16].rf_reg_q ;
assign _0428_ = _0339_ ? _0424_ : _0426_;
assign _0430_ = _0102_ ? _0422_ : _0428_;
assign _0432_ = _0103_ ? _0416_ : _0430_;
assign _0434_ = _0543_ ? \g_rf_flops[15].rf_reg_q  : \g_rf_flops[14].rf_reg_q ;
assign _0436_ = _0545_ ? \g_rf_flops[13].rf_reg_q  : \g_rf_flops[12].rf_reg_q ;
assign _0438_ = _0340_ ? _0434_ : _0436_;
assign _0440_ = _0547_ ? \g_rf_flops[11].rf_reg_q  : \g_rf_flops[10].rf_reg_q ;
assign _0442_ = _0549_ ? \g_rf_flops[9].rf_reg_q  : \g_rf_flops[8].rf_reg_q ;
assign _0444_ = _0341_ ? _0440_ : _0442_;
assign _0446_ = _0104_ ? _0438_ : _0444_;
assign _0448_ = _0551_ ? \g_rf_flops[7].rf_reg_q  : \g_rf_flops[6].rf_reg_q ;
assign _0450_ = _0553_ ? \g_rf_flops[5].rf_reg_q  : \g_rf_flops[4].rf_reg_q ;
assign _0452_ = _0342_ ? _0448_ : _0450_;
assign _0454_ = _0555_ ? \g_rf_flops[3].rf_reg_q  : \g_rf_flops[2].rf_reg_q ;
assign _0456_ = _0557_ ? \g_rf_flops[1].rf_reg_q  : \rf_reg[0] ;
assign _0458_ = _0343_ ? _0454_ : _0456_;
assign _0460_ = _0105_ ? _0452_ : _0458_;
assign _0462_ = _0106_ ? _0446_ : _0460_;
assign rdata_a_o = _0107_ ? _0432_ : _0462_;
assign _0464_ = ! /* src = "generated/sv2v_out.v:20105.20-20105.47" */ waddr_a_i;
assign _0465_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h01;
assign _0466_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h02;
assign _0467_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h03;
assign _0468_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h04;
assign _0469_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h05;
assign _0470_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h06;
assign _0471_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h07;
assign _0472_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h08;
assign _0473_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h09;
assign _0474_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h0a;
assign _0475_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h0b;
assign _0476_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h0c;
assign _0477_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h0d;
assign _0478_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h0e;
assign _0479_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h0f;
assign _0480_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h10;
assign _0481_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h11;
assign _0482_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h12;
assign _0483_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h13;
assign _0484_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h14;
assign _0485_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h15;
assign _0486_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h16;
assign _0487_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h17;
assign _0488_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h18;
assign _0489_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h19;
assign _0490_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h1a;
assign _0491_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h1b;
assign _0492_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h1c;
assign _0493_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h1d;
assign _0494_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h1e;
assign _0495_ = waddr_a_i == /* src = "generated/sv2v_out.v:20105.20-20105.47" */ 5'h1f;
assign _0496_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1f;
assign _0497_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1e;
assign _0498_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1d;
assign _0499_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1c;
assign _0500_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1b;
assign _0501_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1a;
assign _0502_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h19;
assign _0503_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h18;
assign _0504_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h17;
assign _0505_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h16;
assign _0506_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h15;
assign _0507_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h14;
assign _0508_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h13;
assign _0509_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h12;
assign _0510_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h11;
assign _0511_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h10;
assign _0512_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0f;
assign _0513_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0e;
assign _0514_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0d;
assign _0515_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0c;
assign _0516_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0b;
assign _0517_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0a;
assign _0518_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h09;
assign _0519_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h08;
assign _0520_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h07;
assign _0521_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h06;
assign _0522_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h05;
assign _0523_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h04;
assign _0524_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h03;
assign _0525_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h02;
assign _0526_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h01;
assign _0527_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1f;
assign _0528_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1e;
assign _0529_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1d;
assign _0530_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1c;
assign _0531_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1b;
assign _0532_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1a;
assign _0533_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h19;
assign _0534_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h18;
assign _0535_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h17;
assign _0536_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h16;
assign _0537_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h15;
assign _0538_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h14;
assign _0539_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h13;
assign _0540_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h12;
assign _0541_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h11;
assign _0542_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h10;
assign _0543_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0f;
assign _0544_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0e;
assign _0545_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0d;
assign _0546_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0c;
assign _0547_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0b;
assign _0548_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0a;
assign _0549_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h09;
assign _0550_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h08;
assign _0551_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h07;
assign _0552_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h06;
assign _0553_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h05;
assign _0554_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h04;
assign _0555_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h03;
assign _0556_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h02;
assign _0557_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h01;
assign we_a_dec[0] = _0464_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[1] = _0465_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[2] = _0466_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[3] = _0467_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[4] = _0468_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[5] = _0469_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[6] = _0470_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[7] = _0471_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[8] = _0472_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[9] = _0473_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[10] = _0474_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[11] = _0475_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[12] = _0476_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[13] = _0477_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[14] = _0478_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[15] = _0479_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[16] = _0480_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[17] = _0481_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[18] = _0482_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[19] = _0483_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[20] = _0484_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[21] = _0485_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[22] = _0486_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[23] = _0487_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[24] = _0488_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[25] = _0489_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[26] = _0490_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[27] = _0491_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[28] = _0492_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[29] = _0493_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[30] = _0494_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign we_a_dec[31] = _0495_ ? /* src = "generated/sv2v_out.v:20105.20-20105.63" */ we_a_i : 1'h0;
assign \rf_reg[0]  = dummy_instr_id_i ? /* src = "generated/sv2v_out.v:20154.24-20154.64" */ \g_dummy_r0.rf_r0_q  : 39'h2a00000000;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20111.34-20114.5" */
\$paramod\prim_buf\Width=32'00000000000000000000000000100000  \gen_wren_check.u_prim_buf  (
.in_i(we_a_dec),
.in_i_t0(we_a_dec_t0),
.out_o(\gen_wren_check.we_a_dec_buf ),
.out_o_t0(\gen_wren_check.we_a_dec_buf_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20119.6-20126.5" */
\$paramod$916c47de983e2a42946808797a4a11650abb788f\prim_onehot_check  \gen_wren_check.u_prim_onehot_check  (
.addr_i(waddr_a_i),
.addr_i_t0(waddr_a_i_t0),
.clk_i(clk_i),
.en_i(we_a_i),
.en_i_t0(we_a_i_t0),
.err_o(err_o),
.err_o_t0(err_o_t0),
.oh_i(\gen_wren_check.we_a_dec_buf ),
.oh_i_t0(\gen_wren_check.we_a_dec_buf_t0 ),
.rst_ni(rst_ni)
);
endmodule

module \$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers (clk_i, rst_ni, hart_id_i, priv_mode_id_o, priv_mode_lsu_o, csr_mstatus_tw_o, csr_mtvec_o, csr_mtvec_init_i, boot_addr_i, csr_access_i, csr_addr_i, csr_wdata_i, csr_op_i, csr_op_en_i, csr_rdata_o, irq_software_i, irq_timer_i, irq_external_i, irq_fast_i, nmi_mode_i, irq_pending_o
, irqs_o, csr_mstatus_mie_o, csr_mepc_o, csr_mtval_o, csr_pmp_cfg_o, csr_pmp_addr_o, csr_pmp_mseccfg_o, debug_mode_i, debug_mode_entering_i, debug_cause_i, debug_csr_save_i, csr_depc_o, debug_single_step_o, debug_ebreakm_o, debug_ebreaku_o, trigger_match_o, pc_if_i, pc_id_i, pc_wb_i, data_ind_timing_o, dummy_instr_en_o
, dummy_instr_mask_o, dummy_instr_seed_en_o, dummy_instr_seed_o, icache_enable_o, csr_shadow_err_o, ic_scr_key_valid_i, csr_save_if_i, csr_save_id_i, csr_save_wb_i, csr_restore_mret_i, csr_restore_dret_i, csr_save_cause_i, csr_mcause_i, csr_mtval_i, illegal_csr_insn_o, double_fault_seen_o, instr_ret_i, instr_ret_compressed_i, instr_ret_spec_i, instr_ret_compressed_spec_i, iside_wait_i
, jump_i, branch_i, branch_taken_i, mem_load_i, mem_store_i, dside_wait_i, mul_wait_i, div_wait_i, csr_mtval_o_t0, branch_i_t0, branch_taken_i_t0, pc_id_i_t0, ic_scr_key_valid_i_t0, boot_addr_i_t0, csr_access_i_t0, csr_addr_i_t0, csr_depc_o_t0, csr_mcause_i_t0, csr_mepc_o_t0, csr_mstatus_mie_o_t0, csr_mstatus_tw_o_t0
, csr_mtval_i_t0, csr_mtvec_init_i_t0, csr_mtvec_o_t0, csr_op_en_i_t0, csr_op_i_t0, csr_pmp_addr_o_t0, csr_pmp_cfg_o_t0, csr_pmp_mseccfg_o_t0, csr_rdata_o_t0, csr_restore_dret_i_t0, csr_restore_mret_i_t0, csr_save_cause_i_t0, csr_save_id_i_t0, csr_save_if_i_t0, csr_save_wb_i_t0, csr_shadow_err_o_t0, csr_wdata_i_t0, data_ind_timing_o_t0, debug_cause_i_t0, debug_csr_save_i_t0, debug_ebreakm_o_t0
, debug_ebreaku_o_t0, debug_mode_entering_i_t0, debug_mode_i_t0, debug_single_step_o_t0, div_wait_i_t0, double_fault_seen_o_t0, dside_wait_i_t0, dummy_instr_en_o_t0, dummy_instr_mask_o_t0, dummy_instr_seed_en_o_t0, dummy_instr_seed_o_t0, hart_id_i_t0, icache_enable_o_t0, illegal_csr_insn_o_t0, instr_ret_compressed_i_t0, instr_ret_compressed_spec_i_t0, instr_ret_i_t0, instr_ret_spec_i_t0, irq_external_i_t0, irq_fast_i_t0, irq_pending_o_t0
, irq_software_i_t0, irq_timer_i_t0, irqs_o_t0, iside_wait_i_t0, jump_i_t0, mem_load_i_t0, mem_store_i_t0, mul_wait_i_t0, nmi_mode_i_t0, pc_if_i_t0, pc_wb_i_t0, priv_mode_id_o_t0, priv_mode_lsu_o_t0, trigger_match_o_t0);
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [7:0] _0000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [7:0] _0001_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0002_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0003_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0004_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0005_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0006_;
/* src = "generated/sv2v_out.v:13982.2-14112.5" */
wire _0007_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0008_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0009_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [5:0] _0010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [5:0] _0011_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0012_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0013_;
/* src = "generated/sv2v_out.v:13982.2-14112.5" */
wire [63:0] _0014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13982.2-14112.5" */
wire [63:0] _0015_;
/* src = "generated/sv2v_out.v:13982.2-14112.5" */
wire [31:0] _0016_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [7:0] _0017_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [7:0] _0018_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0019_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0021_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0022_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0023_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0024_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0025_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0026_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0027_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0028_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0029_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0030_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [6:0] _0031_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [6:0] _0032_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0033_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0034_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0035_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0036_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0037_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0038_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0039_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0040_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0041_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0042_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0043_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0044_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [5:0] _0045_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [5:0] _0046_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0047_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0048_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0049_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0050_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0051_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0052_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [1:0] _0053_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [1:0] _0054_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0055_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [6:0] _0056_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [6:0] _0057_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0058_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0059_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0060_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [1:0] _0061_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [1:0] _0062_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0063_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0064_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [1:0] _0065_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [1:0] _0066_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0067_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0068_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0069_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0070_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [6:0] _0071_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [6:0] _0072_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0073_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0074_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [31:0] _0075_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0076_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0077_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0078_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [1:0] _0079_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [1:0] _0080_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0081_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0082_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0083_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0084_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [3:0] _0085_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [3:0] _0086_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0087_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0088_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [1:0] _0089_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [1:0] _0090_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0091_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [1:0] _0092_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [1:0] _0093_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0094_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0095_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [3:0] _0096_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [3:0] _0097_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0098_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0099_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [2:0] _0100_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [2:0] _0101_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0102_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire _0103_;
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [2:0] _0104_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14117.2-14256.5" */
wire [2:0] _0105_;
/* src = "generated/sv2v_out.v:14268.26-14268.52" */
wire [31:0] _0106_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14268.26-14268.52" */
wire [31:0] _0107_;
/* src = "generated/sv2v_out.v:14273.23-14273.43" */
wire _0108_;
/* src = "generated/sv2v_out.v:14645.18-14645.57" */
wire _0109_;
/* src = "generated/sv2v_out.v:14657.18-14657.57" */
wire _0110_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14657.18-14657.57" */
wire _0111_;
/* src = "generated/sv2v_out.v:14664.27-14664.63" */
wire _0112_;
wire _0113_;
wire _0114_;
wire [2:0] _0115_;
wire [2:0] _0116_;
wire _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire [2:0] _0132_;
wire [2:0] _0133_;
wire [2:0] _0134_;
wire [2:0] _0135_;
wire [2:0] _0136_;
wire [2:0] _0137_;
wire [2:0] _0138_;
wire [2:0] _0139_;
wire [2:0] _0140_;
wire [2:0] _0141_;
wire [2:0] _0142_;
wire [2:0] _0143_;
wire [2:0] _0144_;
wire [2:0] _0145_;
wire [2:0] _0146_;
wire [2:0] _0147_;
wire [2:0] _0148_;
wire [2:0] _0149_;
wire [2:0] _0150_;
wire [2:0] _0151_;
wire [2:0] _0152_;
wire [2:0] _0153_;
wire [2:0] _0154_;
wire [2:0] _0155_;
wire [2:0] _0156_;
wire [2:0] _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire [2:0] _0172_;
wire [2:0] _0173_;
wire [2:0] _0174_;
wire [2:0] _0175_;
wire [8:0] _0176_;
wire [8:0] _0177_;
wire [8:0] _0178_;
wire [8:0] _0179_;
wire [8:0] _0180_;
wire [8:0] _0181_;
wire [8:0] _0182_;
wire [8:0] _0183_;
wire [8:0] _0184_;
wire [8:0] _0185_;
wire [8:0] _0186_;
wire [8:0] _0187_;
wire [8:0] _0188_;
wire [8:0] _0189_;
wire [63:0] _0190_;
wire [63:0] _0191_;
wire [31:0] _0192_;
wire [31:0] _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire [31:0] _0199_;
wire _0200_;
wire [2:0] _0201_;
wire [2:0] _0202_;
wire [2:0] _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire [1:0] _0209_;
wire [6:0] _0210_;
wire [31:0] _0211_;
wire [31:0] _0212_;
wire [2:0] _0213_;
wire [1:0] _0214_;
wire [6:0] _0215_;
wire [3:0] _0216_;
wire [31:0] _0217_;
wire [31:0] _0218_;
wire [31:0] _0219_;
wire [31:0] _0220_;
wire [1:0] _0221_;
wire [6:0] _0222_;
wire [6:0] _0223_;
wire [6:0] _0224_;
wire [31:0] _0225_;
wire [31:0] _0226_;
wire [6:0] _0227_;
wire [1:0] _0228_;
wire [3:0] _0229_;
wire [1:0] _0230_;
wire [11:0] _0231_;
wire [1:0] _0232_;
wire [1:0] _0233_;
wire [1:0] _0234_;
wire [7:0] _0235_;
wire _0236_;
wire [7:0] _0237_;
wire [31:0] _0238_;
wire [5:0] _0239_;
wire [31:0] _0240_;
wire [1:0] _0241_;
wire [63:0] _0242_;
wire _0243_;
wire _0244_;
wire [31:0] _0245_;
wire _0246_;
wire _0247_;
wire _0248_;
wire [31:0] _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire _0271_;
wire _0272_;
wire _0273_;
wire [31:0] _0274_;
wire [31:0] _0275_;
wire [31:0] _0276_;
wire [17:0] _0277_;
wire [17:0] _0278_;
wire [17:0] _0279_;
wire _0280_;
wire _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire _0285_;
wire [1:0] _0286_;
wire [1:0] _0287_;
wire [1:0] _0288_;
wire [1:0] _0289_;
wire [2:0] _0290_;
wire [2:0] _0291_;
wire [2:0] _0292_;
wire [2:0] _0293_;
wire _0294_;
wire _0295_;
wire _0296_;
wire _0297_;
wire _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire [2:0] _0324_;
wire [2:0] _0325_;
wire [2:0] _0326_;
wire [2:0] _0327_;
wire [2:0] _0328_;
wire [2:0] _0329_;
wire [2:0] _0330_;
wire [2:0] _0331_;
wire [2:0] _0332_;
wire [2:0] _0333_;
wire [2:0] _0334_;
wire [2:0] _0335_;
wire [2:0] _0336_;
wire [2:0] _0337_;
wire [2:0] _0338_;
wire [2:0] _0339_;
wire [2:0] _0340_;
wire [2:0] _0341_;
wire [2:0] _0342_;
wire [2:0] _0343_;
wire [2:0] _0344_;
wire [2:0] _0345_;
wire [2:0] _0346_;
wire [2:0] _0347_;
wire [2:0] _0348_;
wire [2:0] _0349_;
wire [2:0] _0350_;
wire [2:0] _0351_;
wire [2:0] _0352_;
wire [2:0] _0353_;
wire [2:0] _0354_;
wire [2:0] _0355_;
wire [2:0] _0356_;
wire [2:0] _0357_;
wire [2:0] _0358_;
wire [2:0] _0359_;
wire [2:0] _0360_;
wire [2:0] _0361_;
wire [2:0] _0362_;
wire [2:0] _0363_;
wire [2:0] _0364_;
wire [2:0] _0365_;
wire [2:0] _0366_;
wire [2:0] _0367_;
wire [2:0] _0368_;
wire [2:0] _0369_;
wire [2:0] _0370_;
wire [2:0] _0371_;
wire [2:0] _0372_;
wire [2:0] _0373_;
wire [2:0] _0374_;
wire [2:0] _0375_;
wire [2:0] _0376_;
wire [2:0] _0377_;
wire [2:0] _0378_;
wire [2:0] _0379_;
wire [2:0] _0380_;
wire [2:0] _0381_;
wire [2:0] _0382_;
wire [2:0] _0383_;
wire [2:0] _0384_;
wire [2:0] _0385_;
wire [2:0] _0386_;
wire [2:0] _0387_;
wire [2:0] _0388_;
wire [2:0] _0389_;
wire [2:0] _0390_;
wire [2:0] _0391_;
wire [2:0] _0392_;
wire [2:0] _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire _0398_;
wire _0399_;
wire _0400_;
wire _0401_;
wire _0402_;
wire _0403_;
wire _0404_;
wire _0405_;
wire _0406_;
wire _0407_;
wire _0408_;
wire _0409_;
wire _0410_;
wire _0411_;
wire _0412_;
wire _0413_;
wire _0414_;
wire _0415_;
wire _0416_;
wire _0417_;
wire _0418_;
wire _0419_;
wire _0420_;
wire _0421_;
wire _0422_;
wire _0423_;
wire _0424_;
wire _0425_;
wire _0426_;
wire _0427_;
wire _0428_;
wire _0429_;
wire _0430_;
wire _0431_;
wire _0432_;
wire _0433_;
wire _0434_;
wire _0435_;
wire _0436_;
wire _0437_;
wire _0438_;
wire _0439_;
wire _0440_;
wire _0441_;
wire [2:0] _0442_;
wire [2:0] _0443_;
wire [2:0] _0444_;
wire [2:0] _0445_;
wire [2:0] _0446_;
wire [2:0] _0447_;
wire [2:0] _0448_;
wire [2:0] _0449_;
wire [2:0] _0450_;
wire [2:0] _0451_;
wire [2:0] _0452_;
wire [2:0] _0453_;
wire [2:0] _0454_;
wire [2:0] _0455_;
wire [2:0] _0456_;
wire [2:0] _0457_;
wire [2:0] _0458_;
wire [2:0] _0459_;
wire [2:0] _0460_;
wire [2:0] _0461_;
wire _0462_;
wire _0463_;
wire _0464_;
wire _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire _0469_;
wire _0470_;
wire _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire _0477_;
wire _0478_;
wire _0479_;
wire _0480_;
wire _0481_;
wire _0482_;
wire _0483_;
wire _0484_;
wire _0485_;
wire [8:0] _0486_;
wire [8:0] _0487_;
wire [8:0] _0488_;
wire [8:0] _0489_;
wire [8:0] _0490_;
wire [8:0] _0491_;
wire [8:0] _0492_;
wire [8:0] _0493_;
wire [8:0] _0494_;
wire [8:0] _0495_;
wire [8:0] _0496_;
wire [8:0] _0497_;
wire [8:0] _0498_;
wire [8:0] _0499_;
wire [8:0] _0500_;
wire [8:0] _0501_;
wire [8:0] _0502_;
wire [8:0] _0503_;
wire [8:0] _0504_;
wire [8:0] _0505_;
wire [8:0] _0506_;
wire [8:0] _0507_;
wire [8:0] _0508_;
wire [8:0] _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0517_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
wire _0525_;
wire _0526_;
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire _0534_;
wire _0535_;
wire [63:0] _0536_;
wire [63:0] _0537_;
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0542_;
wire _0543_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire _0560_;
wire _0561_;
wire _0562_;
wire _0563_;
wire [31:0] _0564_;
wire [31:0] _0565_;
wire [31:0] _0566_;
wire [31:0] _0567_;
wire _0568_;
wire _0569_;
wire _0570_;
wire _0571_;
wire _0572_;
wire _0573_;
wire _0574_;
wire _0575_;
wire _0576_;
wire _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire _0596_;
wire _0597_;
wire _0598_;
wire _0599_;
wire _0600_;
wire _0601_;
wire _0602_;
wire _0603_;
wire _0604_;
wire _0605_;
wire _0606_;
wire _0607_;
wire _0608_;
wire _0609_;
wire _0610_;
wire _0611_;
wire _0612_;
wire _0613_;
wire _0614_;
wire _0615_;
wire _0616_;
wire _0617_;
wire [2:0] _0618_;
wire [2:0] _0619_;
wire [2:0] _0620_;
wire [2:0] _0621_;
wire [2:0] _0622_;
wire [2:0] _0623_;
wire [2:0] _0624_;
wire [2:0] _0625_;
wire [2:0] _0626_;
wire [2:0] _0627_;
wire [2:0] _0628_;
wire [2:0] _0629_;
wire [2:0] _0630_;
wire [2:0] _0631_;
wire [2:0] _0632_;
wire [2:0] _0633_;
wire [2:0] _0634_;
wire [2:0] _0635_;
wire [2:0] _0636_;
wire [2:0] _0637_;
wire _0638_;
wire _0639_;
wire _0640_;
wire [31:0] _0641_;
wire _0642_;
wire _0643_;
wire _0644_;
wire _0645_;
wire _0646_;
wire _0647_;
wire _0648_;
wire _0649_;
wire _0650_;
wire _0651_;
wire _0652_;
wire [31:0] _0653_;
wire [31:0] _0654_;
wire [2:0] _0655_;
wire [2:0] _0656_;
wire [2:0] _0657_;
wire [2:0] _0658_;
wire [2:0] _0659_;
wire [2:0] _0660_;
wire _0661_;
wire _0662_;
wire _0663_;
wire _0664_;
wire _0665_;
wire _0666_;
wire _0667_;
wire _0668_;
wire _0669_;
wire _0670_;
wire _0671_;
wire _0672_;
wire [1:0] _0673_;
wire [1:0] _0674_;
wire [6:0] _0675_;
wire [6:0] _0676_;
wire [31:0] _0677_;
wire [31:0] _0678_;
wire _0679_;
wire _0680_;
wire [1:0] _0681_;
wire [1:0] _0682_;
wire _0683_;
wire _0684_;
wire [31:0] _0685_;
wire [31:0] _0686_;
wire [31:0] _0687_;
wire [31:0] _0688_;
wire [2:0] _0689_;
wire [2:0] _0690_;
wire [1:0] _0691_;
wire [1:0] _0692_;
wire [1:0] _0693_;
wire [1:0] _0694_;
wire [31:0] _0695_;
wire [31:0] _0696_;
wire [6:0] _0697_;
wire [6:0] _0698_;
wire [31:0] _0699_;
wire [31:0] _0700_;
wire [3:0] _0701_;
wire [3:0] _0702_;
wire [31:0] _0703_;
wire [31:0] _0704_;
wire [31:0] _0705_;
wire [31:0] _0706_;
wire [31:0] _0707_;
wire [31:0] _0708_;
wire _0709_;
wire _0710_;
wire _0711_;
wire _0712_;
wire [31:0] _0713_;
wire [31:0] _0714_;
wire [2:0] _0715_;
wire [2:0] _0716_;
wire [1:0] _0717_;
wire [1:0] _0718_;
wire [31:0] _0719_;
wire [31:0] _0720_;
wire [6:0] _0721_;
wire [6:0] _0722_;
wire [6:0] _0723_;
wire [6:0] _0724_;
wire [6:0] _0725_;
wire [6:0] _0726_;
wire [31:0] _0727_;
wire [31:0] _0728_;
wire [31:0] _0729_;
wire [31:0] _0730_;
wire [31:0] _0731_;
wire [31:0] _0732_;
wire [6:0] _0733_;
wire [6:0] _0734_;
wire [1:0] _0735_;
wire [1:0] _0736_;
wire [1:0] _0737_;
wire [1:0] _0738_;
wire [1:0] _0739_;
wire [1:0] _0740_;
wire _0741_;
wire _0742_;
wire [1:0] _0743_;
wire [1:0] _0744_;
wire [1:0] _0745_;
wire [1:0] _0746_;
wire _0747_;
wire _0748_;
wire [1:0] _0749_;
wire [1:0] _0750_;
wire [7:0] _0751_;
wire [7:0] _0752_;
wire [7:0] _0753_;
wire [7:0] _0754_;
wire [31:0] _0755_;
wire [31:0] _0756_;
wire _0757_;
wire _0758_;
wire [5:0] _0759_;
wire [5:0] _0760_;
wire [31:0] _0761_;
wire [31:0] _0762_;
wire [1:0] _0763_;
wire [1:0] _0764_;
wire [63:0] _0765_;
wire [63:0] _0766_;
wire _0767_;
wire _0768_;
wire _0769_;
wire _0770_;
wire _0771_;
wire _0772_;
wire _0773_;
wire _0774_;
wire _0775_;
wire _0776_;
wire _0777_;
wire _0778_;
wire _0779_;
wire [31:0] _0780_;
wire [17:0] _0781_;
wire _0782_;
wire _0783_;
wire [1:0] _0784_;
wire [1:0] _0785_;
wire _0786_;
wire [31:0] _0787_;
wire _0788_;
wire _0789_;
wire _0790_;
wire [2:0] _0791_;
/* cellift = 32'd1 */
wire [2:0] _0792_;
wire [2:0] _0793_;
wire [2:0] _0794_;
/* cellift = 32'd1 */
wire [2:0] _0795_;
wire [2:0] _0796_;
/* cellift = 32'd1 */
wire [2:0] _0797_;
wire _0798_;
/* cellift = 32'd1 */
wire _0799_;
wire _0800_;
/* cellift = 32'd1 */
wire _0801_;
wire _0802_;
/* cellift = 32'd1 */
wire _0803_;
wire _0804_;
/* cellift = 32'd1 */
wire _0805_;
wire _0806_;
/* cellift = 32'd1 */
wire _0807_;
wire _0808_;
/* cellift = 32'd1 */
wire _0809_;
wire _0810_;
/* cellift = 32'd1 */
wire _0811_;
wire _0812_;
/* cellift = 32'd1 */
wire _0813_;
wire _0814_;
/* cellift = 32'd1 */
wire _0815_;
wire _0816_;
/* cellift = 32'd1 */
wire _0817_;
wire _0818_;
/* cellift = 32'd1 */
wire _0819_;
wire _0820_;
/* cellift = 32'd1 */
wire _0821_;
wire _0822_;
/* cellift = 32'd1 */
wire _0823_;
wire _0824_;
/* cellift = 32'd1 */
wire _0825_;
wire _0826_;
/* cellift = 32'd1 */
wire _0827_;
wire _0828_;
/* cellift = 32'd1 */
wire _0829_;
wire [2:0] _0830_;
/* cellift = 32'd1 */
wire [2:0] _0831_;
wire [2:0] _0832_;
/* cellift = 32'd1 */
wire [2:0] _0833_;
wire [2:0] _0834_;
/* cellift = 32'd1 */
wire [2:0] _0835_;
wire [2:0] _0836_;
/* cellift = 32'd1 */
wire [2:0] _0837_;
wire [2:0] _0838_;
/* cellift = 32'd1 */
wire [2:0] _0839_;
wire [2:0] _0840_;
/* cellift = 32'd1 */
wire [2:0] _0841_;
wire [2:0] _0842_;
/* cellift = 32'd1 */
wire [2:0] _0843_;
wire [2:0] _0844_;
/* cellift = 32'd1 */
wire [2:0] _0845_;
wire [2:0] _0846_;
/* cellift = 32'd1 */
wire [2:0] _0847_;
wire [2:0] _0848_;
/* cellift = 32'd1 */
wire [2:0] _0849_;
wire [2:0] _0850_;
/* cellift = 32'd1 */
wire [2:0] _0851_;
wire [2:0] _0852_;
/* cellift = 32'd1 */
wire [2:0] _0853_;
wire [2:0] _0854_;
wire [2:0] _0855_;
/* cellift = 32'd1 */
wire [2:0] _0856_;
wire [2:0] _0857_;
/* cellift = 32'd1 */
wire [2:0] _0858_;
wire [2:0] _0859_;
/* cellift = 32'd1 */
wire [2:0] _0860_;
wire [2:0] _0861_;
/* cellift = 32'd1 */
wire [2:0] _0862_;
wire [2:0] _0863_;
/* cellift = 32'd1 */
wire [2:0] _0864_;
wire [2:0] _0865_;
/* cellift = 32'd1 */
wire [2:0] _0866_;
wire [2:0] _0867_;
/* cellift = 32'd1 */
wire [2:0] _0868_;
wire [2:0] _0869_;
/* cellift = 32'd1 */
wire [2:0] _0870_;
wire [2:0] _0871_;
/* cellift = 32'd1 */
wire [2:0] _0872_;
wire [2:0] _0873_;
/* cellift = 32'd1 */
wire [2:0] _0874_;
wire [2:0] _0875_;
/* cellift = 32'd1 */
wire [2:0] _0876_;
wire [2:0] _0877_;
/* cellift = 32'd1 */
wire [2:0] _0878_;
wire [2:0] _0879_;
/* cellift = 32'd1 */
wire [2:0] _0880_;
wire [2:0] _0881_;
/* cellift = 32'd1 */
wire [2:0] _0882_;
wire [2:0] _0883_;
/* cellift = 32'd1 */
wire [2:0] _0884_;
wire [2:0] _0885_;
/* cellift = 32'd1 */
wire [2:0] _0886_;
wire [2:0] _0887_;
/* cellift = 32'd1 */
wire [2:0] _0888_;
wire [2:0] _0889_;
/* cellift = 32'd1 */
wire [2:0] _0890_;
wire [2:0] _0891_;
/* cellift = 32'd1 */
wire [2:0] _0892_;
wire [2:0] _0893_;
/* cellift = 32'd1 */
wire [2:0] _0894_;
wire [2:0] _0895_;
/* cellift = 32'd1 */
wire [2:0] _0896_;
wire [2:0] _0897_;
/* cellift = 32'd1 */
wire [2:0] _0898_;
wire [2:0] _0899_;
/* cellift = 32'd1 */
wire [2:0] _0900_;
wire [2:0] _0901_;
/* cellift = 32'd1 */
wire [2:0] _0902_;
wire [2:0] _0903_;
/* cellift = 32'd1 */
wire [2:0] _0904_;
wire [2:0] _0905_;
/* cellift = 32'd1 */
wire [2:0] _0906_;
wire [2:0] _0907_;
/* cellift = 32'd1 */
wire [2:0] _0908_;
wire [2:0] _0909_;
/* cellift = 32'd1 */
wire [2:0] _0910_;
wire [2:0] _0911_;
/* cellift = 32'd1 */
wire [2:0] _0912_;
wire [2:0] _0913_;
/* cellift = 32'd1 */
wire [2:0] _0914_;
wire [2:0] _0915_;
/* cellift = 32'd1 */
wire [2:0] _0916_;
wire _0917_;
/* cellift = 32'd1 */
wire _0918_;
wire _0919_;
/* cellift = 32'd1 */
wire _0920_;
wire _0921_;
/* cellift = 32'd1 */
wire _0922_;
wire _0923_;
/* cellift = 32'd1 */
wire _0924_;
wire _0925_;
/* cellift = 32'd1 */
wire _0926_;
wire _0927_;
/* cellift = 32'd1 */
wire _0928_;
wire _0929_;
/* cellift = 32'd1 */
wire _0930_;
wire _0931_;
/* cellift = 32'd1 */
wire _0932_;
wire _0933_;
/* cellift = 32'd1 */
wire _0934_;
wire _0935_;
/* cellift = 32'd1 */
wire _0936_;
wire _0937_;
/* cellift = 32'd1 */
wire _0938_;
wire _0939_;
/* cellift = 32'd1 */
wire _0940_;
wire _0941_;
/* cellift = 32'd1 */
wire _0942_;
wire _0943_;
/* cellift = 32'd1 */
wire _0944_;
wire _0945_;
/* cellift = 32'd1 */
wire _0946_;
wire _0947_;
/* cellift = 32'd1 */
wire _0948_;
wire _0949_;
/* cellift = 32'd1 */
wire _0950_;
wire _0951_;
/* cellift = 32'd1 */
wire _0952_;
wire _0953_;
/* cellift = 32'd1 */
wire _0954_;
wire _0955_;
/* cellift = 32'd1 */
wire _0956_;
wire _0957_;
/* cellift = 32'd1 */
wire _0958_;
wire _0959_;
/* cellift = 32'd1 */
wire _0960_;
wire _0961_;
/* cellift = 32'd1 */
wire _0962_;
wire _0963_;
/* cellift = 32'd1 */
wire _0964_;
wire _0965_;
/* cellift = 32'd1 */
wire _0966_;
wire _0967_;
/* cellift = 32'd1 */
wire _0968_;
wire _0969_;
/* cellift = 32'd1 */
wire _0970_;
wire _0971_;
/* cellift = 32'd1 */
wire _0972_;
wire _0973_;
/* cellift = 32'd1 */
wire _0974_;
wire [2:0] _0975_;
/* cellift = 32'd1 */
wire [2:0] _0976_;
wire [2:0] _0977_;
/* cellift = 32'd1 */
wire [2:0] _0978_;
wire [2:0] _0979_;
/* cellift = 32'd1 */
wire [2:0] _0980_;
wire [2:0] _0981_;
/* cellift = 32'd1 */
wire [2:0] _0982_;
wire [2:0] _0983_;
/* cellift = 32'd1 */
wire [2:0] _0984_;
wire [2:0] _0985_;
/* cellift = 32'd1 */
wire [2:0] _0986_;
wire [2:0] _0987_;
/* cellift = 32'd1 */
wire [2:0] _0988_;
wire [2:0] _0989_;
/* cellift = 32'd1 */
wire [2:0] _0990_;
wire [2:0] _0991_;
/* cellift = 32'd1 */
wire [2:0] _0992_;
wire [2:0] _0993_;
/* cellift = 32'd1 */
wire [2:0] _0994_;
wire [2:0] _0995_;
/* cellift = 32'd1 */
wire [2:0] _0996_;
wire [2:0] _0997_;
/* cellift = 32'd1 */
wire [2:0] _0998_;
wire _0999_;
/* cellift = 32'd1 */
wire _1000_;
wire _1001_;
/* cellift = 32'd1 */
wire _1002_;
wire _1003_;
/* cellift = 32'd1 */
wire _1004_;
wire _1005_;
/* cellift = 32'd1 */
wire _1006_;
wire _1007_;
/* cellift = 32'd1 */
wire _1008_;
wire _1009_;
/* cellift = 32'd1 */
wire _1010_;
wire _1011_;
/* cellift = 32'd1 */
wire _1012_;
wire _1013_;
/* cellift = 32'd1 */
wire _1014_;
wire _1015_;
/* cellift = 32'd1 */
wire _1016_;
wire _1017_;
/* cellift = 32'd1 */
wire _1018_;
wire _1019_;
/* cellift = 32'd1 */
wire _1020_;
wire _1021_;
/* cellift = 32'd1 */
wire _1022_;
wire _1023_;
/* cellift = 32'd1 */
wire _1024_;
wire _1025_;
/* cellift = 32'd1 */
wire _1026_;
wire [8:0] _1027_;
/* cellift = 32'd1 */
wire [8:0] _1028_;
wire [8:0] _1029_;
/* cellift = 32'd1 */
wire [8:0] _1030_;
wire [8:0] _1031_;
/* cellift = 32'd1 */
wire [8:0] _1032_;
wire [8:0] _1033_;
/* cellift = 32'd1 */
wire [8:0] _1034_;
wire [8:0] _1035_;
/* cellift = 32'd1 */
wire [8:0] _1036_;
wire [8:0] _1037_;
/* cellift = 32'd1 */
wire [8:0] _1038_;
wire [8:0] _1039_;
/* cellift = 32'd1 */
wire [8:0] _1040_;
wire [8:0] _1041_;
/* cellift = 32'd1 */
wire [8:0] _1042_;
wire [8:0] _1043_;
/* cellift = 32'd1 */
wire [8:0] _1044_;
wire [8:0] _1045_;
/* cellift = 32'd1 */
wire [8:0] _1046_;
wire [8:0] _1047_;
/* cellift = 32'd1 */
wire [8:0] _1048_;
wire [8:0] _1049_;
/* cellift = 32'd1 */
wire [8:0] _1050_;
wire [8:0] _1051_;
/* cellift = 32'd1 */
wire [8:0] _1052_;
wire [8:0] _1053_;
/* cellift = 32'd1 */
wire [8:0] _1054_;
wire [8:0] _1055_;
/* cellift = 32'd1 */
wire [8:0] _1056_;
wire _1057_;
/* cellift = 32'd1 */
wire _1058_;
wire _1059_;
/* cellift = 32'd1 */
wire _1060_;
wire _1061_;
/* cellift = 32'd1 */
wire _1062_;
wire _1063_;
/* cellift = 32'd1 */
wire _1064_;
wire _1065_;
/* cellift = 32'd1 */
wire _1066_;
wire _1067_;
/* cellift = 32'd1 */
wire _1068_;
wire _1069_;
/* cellift = 32'd1 */
wire _1070_;
wire _1071_;
/* cellift = 32'd1 */
wire _1072_;
wire _1073_;
/* cellift = 32'd1 */
wire _1074_;
wire _1075_;
/* cellift = 32'd1 */
wire _1076_;
wire _1077_;
/* cellift = 32'd1 */
wire _1078_;
wire _1079_;
/* cellift = 32'd1 */
wire _1080_;
wire _1081_;
/* cellift = 32'd1 */
wire _1082_;
wire _1083_;
/* cellift = 32'd1 */
wire _1084_;
wire _1085_;
/* cellift = 32'd1 */
wire _1086_;
wire [63:0] _1087_;
/* cellift = 32'd1 */
wire [63:0] _1088_;
wire _1089_;
/* cellift = 32'd1 */
wire _1090_;
wire _1091_;
/* cellift = 32'd1 */
wire _1092_;
wire _1093_;
/* cellift = 32'd1 */
wire _1094_;
wire _1095_;
/* cellift = 32'd1 */
wire _1096_;
wire _1097_;
/* cellift = 32'd1 */
wire _1098_;
wire _1099_;
/* cellift = 32'd1 */
wire _1100_;
wire _1101_;
/* cellift = 32'd1 */
wire _1102_;
wire _1103_;
/* cellift = 32'd1 */
wire _1104_;
wire _1105_;
/* cellift = 32'd1 */
wire _1106_;
wire _1107_;
/* cellift = 32'd1 */
wire _1108_;
wire _1109_;
/* cellift = 32'd1 */
wire _1110_;
wire _1111_;
/* cellift = 32'd1 */
wire _1112_;
wire _1113_;
/* cellift = 32'd1 */
wire _1114_;
wire _1115_;
/* cellift = 32'd1 */
wire _1116_;
wire _1117_;
/* cellift = 32'd1 */
wire _1118_;
wire [31:0] _1119_;
/* cellift = 32'd1 */
wire [31:0] _1120_;
wire _1121_;
/* cellift = 32'd1 */
wire _1122_;
wire _1123_;
/* cellift = 32'd1 */
wire _1124_;
wire _1125_;
/* cellift = 32'd1 */
wire _1126_;
wire _1127_;
/* cellift = 32'd1 */
wire _1128_;
wire _1129_;
/* cellift = 32'd1 */
wire _1130_;
wire _1131_;
/* cellift = 32'd1 */
wire _1132_;
wire _1133_;
/* cellift = 32'd1 */
wire _1134_;
wire _1135_;
/* cellift = 32'd1 */
wire _1136_;
wire _1137_;
/* cellift = 32'd1 */
wire _1138_;
wire _1139_;
/* cellift = 32'd1 */
wire _1140_;
wire _1141_;
/* cellift = 32'd1 */
wire _1142_;
wire _1143_;
/* cellift = 32'd1 */
wire _1144_;
wire _1145_;
/* cellift = 32'd1 */
wire _1146_;
wire _1147_;
/* cellift = 32'd1 */
wire _1148_;
wire _1149_;
/* cellift = 32'd1 */
wire _1150_;
wire _1151_;
/* cellift = 32'd1 */
wire _1152_;
wire _1153_;
/* cellift = 32'd1 */
wire _1154_;
wire _1155_;
/* cellift = 32'd1 */
wire _1156_;
wire _1157_;
/* cellift = 32'd1 */
wire _1158_;
wire _1159_;
/* cellift = 32'd1 */
wire _1160_;
wire _1161_;
/* cellift = 32'd1 */
wire _1162_;
wire _1163_;
/* cellift = 32'd1 */
wire _1164_;
wire _1165_;
/* cellift = 32'd1 */
wire _1166_;
wire _1167_;
/* cellift = 32'd1 */
wire _1168_;
wire _1169_;
/* cellift = 32'd1 */
wire _1170_;
wire _1171_;
/* cellift = 32'd1 */
wire _1172_;
wire _1173_;
/* cellift = 32'd1 */
wire _1174_;
wire _1175_;
/* cellift = 32'd1 */
wire _1176_;
wire [2:0] _1177_;
/* cellift = 32'd1 */
wire [2:0] _1178_;
wire [2:0] _1179_;
/* cellift = 32'd1 */
wire [2:0] _1180_;
wire [2:0] _1181_;
/* cellift = 32'd1 */
wire [2:0] _1182_;
wire [2:0] _1183_;
/* cellift = 32'd1 */
wire [2:0] _1184_;
wire [2:0] _1185_;
/* cellift = 32'd1 */
wire [2:0] _1186_;
wire [2:0] _1187_;
/* cellift = 32'd1 */
wire [2:0] _1188_;
wire [2:0] _1189_;
/* cellift = 32'd1 */
wire [2:0] _1190_;
wire [2:0] _1191_;
/* cellift = 32'd1 */
wire [2:0] _1192_;
wire [2:0] _1193_;
/* cellift = 32'd1 */
wire [2:0] _1194_;
wire [2:0] _1195_;
/* cellift = 32'd1 */
wire [2:0] _1196_;
/* src = "generated/sv2v_out.v:13958.30-13958.54" */
wire _1197_;
/* src = "generated/sv2v_out.v:14110.409-14110.428" */
wire _1198_;
/* src = "generated/sv2v_out.v:14110.388-14110.407" */
wire _1199_;
/* src = "generated/sv2v_out.v:14110.367-14110.386" */
wire _1200_;
/* src = "generated/sv2v_out.v:14110.346-14110.365" */
wire _1201_;
/* src = "generated/sv2v_out.v:14110.325-14110.344" */
wire _1202_;
/* src = "generated/sv2v_out.v:14110.304-14110.323" */
wire _1203_;
/* src = "generated/sv2v_out.v:14110.283-14110.302" */
wire _1204_;
/* src = "generated/sv2v_out.v:14110.262-14110.281" */
wire _1205_;
/* src = "generated/sv2v_out.v:14110.241-14110.260" */
wire _1206_;
/* src = "generated/sv2v_out.v:14110.220-14110.239" */
wire _1207_;
/* src = "generated/sv2v_out.v:14110.199-14110.218" */
wire _1208_;
/* src = "generated/sv2v_out.v:14110.178-14110.197" */
wire _1209_;
/* src = "generated/sv2v_out.v:14110.157-14110.176" */
wire _1210_;
/* src = "generated/sv2v_out.v:14110.136-14110.155" */
wire _1211_;
/* src = "generated/sv2v_out.v:14110.115-14110.134" */
wire _1212_;
/* src = "generated/sv2v_out.v:14110.94-14110.113" */
wire _1213_;
/* src = "generated/sv2v_out.v:14110.73-14110.92" */
wire _1214_;
/* src = "generated/sv2v_out.v:14110.52-14110.71" */
wire _1215_;
/* src = "generated/sv2v_out.v:14110.31-14110.50" */
wire _1216_;
/* src = "generated/sv2v_out.v:14110.10-14110.29" */
wire _1217_;
/* src = "generated/sv2v_out.v:14127.46-14127.75" */
wire _1218_;
/* src = "generated/sv2v_out.v:14127.15-14127.44" */
wire _1219_;
/* src = "generated/sv2v_out.v:14272.56-14272.72" */
wire _1220_;
/* src = "generated/sv2v_out.v:14272.38-14272.54" */
wire _1221_;
/* src = "generated/sv2v_out.v:14272.20-14272.36" */
wire _1222_;
/* src = "generated/sv2v_out.v:14824.50-14824.69" */
wire _1223_;
/* src = "generated/sv2v_out.v:14154.10-14154.66" */
wire _1224_;
/* src = "generated/sv2v_out.v:14166.10-14166.60" */
wire _1225_;
/* src = "generated/sv2v_out.v:14221.12-14221.38" */
wire _1226_;
/* src = "generated/sv2v_out.v:14154.11-14154.35" */
wire _1227_;
/* src = "generated/sv2v_out.v:14154.41-14154.65" */
wire _1228_;
/* src = "generated/sv2v_out.v:14166.11-14166.32" */
wire _1229_;
/* src = "generated/sv2v_out.v:14166.38-14166.59" */
wire _1230_;
/* src = "generated/sv2v_out.v:14236.9-14236.33" */
wire _1231_;
/* src = "generated/sv2v_out.v:0.0-0.0" */
wire [31:0] _1232_;
/* src = "generated/sv2v_out.v:14273.47-14273.66" */
wire _1233_;
/* src = "generated/sv2v_out.v:14657.40-14657.57" */
wire _1234_;
/* src = "generated/sv2v_out.v:14868.50-14868.89" */
wire _1235_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14868.50-14868.89" */
wire _1236_;
/* src = "generated/sv2v_out.v:0.0-0.0" */
wire [31:0] _1237_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:0.0-0.0" */
wire [31:0] _1238_;
/* src = "generated/sv2v_out.v:13959.48-13959.79" */
wire _1239_;
/* src = "generated/sv2v_out.v:13959.47-13959.99" */
wire _1240_;
/* src = "generated/sv2v_out.v:13959.46-13959.118" */
wire _1241_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13959.46-13959.118" */
wire _1242_;
/* src = "generated/sv2v_out.v:14014.30-14014.55" */
wire _1243_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14014.30-14014.55" */
wire _1244_;
/* src = "generated/sv2v_out.v:14267.26-14267.51" */
wire [31:0] _1245_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14267.26-14267.51" */
wire [31:0] _1246_;
/* src = "generated/sv2v_out.v:14868.52-14868.88" */
wire _1247_;
/* src = "generated/sv2v_out.v:14881.31-14881.54" */
wire _1248_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14881.31-14881.54" */
wire _1249_;
wire _1250_;
wire [2:0] _1251_;
/* cellift = 32'd1 */
wire [2:0] _1252_;
wire [2:0] _1253_;
/* cellift = 32'd1 */
wire [2:0] _1254_;
wire _1255_;
/* cellift = 32'd1 */
wire _1256_;
wire _1257_;
/* cellift = 32'd1 */
wire _1258_;
wire _1259_;
/* cellift = 32'd1 */
wire _1260_;
wire _1261_;
/* cellift = 32'd1 */
wire _1262_;
wire [31:0] _1263_;
/* cellift = 32'd1 */
wire [31:0] _1264_;
wire [31:0] _1265_;
/* cellift = 32'd1 */
wire [31:0] _1266_;
wire _1267_;
wire _1268_;
wire _1269_;
/* cellift = 32'd1 */
wire _1270_;
wire _1271_;
/* cellift = 32'd1 */
wire _1272_;
wire _1273_;
wire _1274_;
wire [6:0] _1275_;
/* cellift = 32'd1 */
wire [6:0] _1276_;
wire [6:0] _1277_;
/* cellift = 32'd1 */
wire [6:0] _1278_;
wire _1279_;
wire _1280_;
wire [31:0] _1281_;
/* cellift = 32'd1 */
wire [31:0] _1282_;
wire [31:0] _1283_;
/* cellift = 32'd1 */
wire [31:0] _1284_;
wire _1285_;
wire _1286_;
wire [1:0] _1287_;
/* cellift = 32'd1 */
wire [1:0] _1288_;
wire [1:0] _1289_;
/* cellift = 32'd1 */
wire [1:0] _1290_;
wire _1291_;
wire _1292_;
wire [30:0] _1293_;
wire _1294_;
wire [30:0] _1295_;
wire _1296_;
wire _1297_;
wire _1298_;
wire _1299_;
wire _1300_;
wire _1301_;
wire _1302_;
wire _1303_;
wire _1304_;
wire _1305_;
wire _1306_;
wire _1307_;
wire _1308_;
wire [28:0] _1309_;
wire _1310_;
wire _1311_;
wire _1312_;
wire _1313_;
wire _1314_;
wire _1315_;
wire _1316_;
wire _1317_;
wire _1318_;
wire _1319_;
wire _1320_;
wire _1321_;
wire _1322_;
wire _1323_;
wire _1324_;
wire _1325_;
wire _1326_;
wire _1327_;
wire _1328_;
wire _1329_;
wire _1330_;
wire _1331_;
wire _1332_;
wire _1333_;
wire _1334_;
wire _1335_;
wire _1336_;
wire _1337_;
wire _1338_;
wire _1339_;
wire _1340_;
wire _1341_;
wire _1342_;
wire _1343_;
wire _1344_;
wire _1345_;
wire _1346_;
wire _1347_;
wire [1:0] _1348_;
wire _1349_;
wire _1350_;
wire _1351_;
wire _1352_;
/* src = "generated/sv2v_out.v:14014.58-14014.116" */
wire [25:0] _1353_;
/* src = "generated/sv2v_out.v:13778.20-13778.31" */
input [31:0] boot_addr_i;
wire [31:0] boot_addr_i;
/* cellift = 32'd1 */
input [31:0] boot_addr_i_t0;
wire [31:0] boot_addr_i_t0;
/* src = "generated/sv2v_out.v:13834.13-13834.21" */
input branch_i;
wire branch_i;
/* cellift = 32'd1 */
input branch_i_t0;
wire branch_i_t0;
/* src = "generated/sv2v_out.v:13835.13-13835.27" */
input branch_taken_i;
wire branch_taken_i;
/* cellift = 32'd1 */
input branch_taken_i_t0;
wire branch_taken_i_t0;
/* src = "generated/sv2v_out.v:13770.13-13770.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:13933.12-13933.29" */
wire [7:0] cpuctrlsts_part_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13933.12-13933.29" */
wire [7:0] cpuctrlsts_part_d_t0;
/* src = "generated/sv2v_out.v:13937.7-13937.26" */
wire cpuctrlsts_part_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13937.7-13937.26" */
wire cpuctrlsts_part_err_t0;
/* src = "generated/sv2v_out.v:13932.13-13932.30" */
wire [7:0] cpuctrlsts_part_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13932.13-13932.30" */
wire [7:0] cpuctrlsts_part_q_t0;
/* src = "generated/sv2v_out.v:13936.6-13936.24" */
wire cpuctrlsts_part_we;
/* src = "generated/sv2v_out.v:13779.13-13779.25" */
input csr_access_i;
wire csr_access_i;
/* cellift = 32'd1 */
input csr_access_i_t0;
wire csr_access_i_t0;
/* src = "generated/sv2v_out.v:13780.20-13780.30" */
input [11:0] csr_addr_i;
wire [11:0] csr_addr_i;
/* cellift = 32'd1 */
input [11:0] csr_addr_i_t0;
wire [11:0] csr_addr_i_t0;
/* src = "generated/sv2v_out.v:13802.21-13802.31" */
output [31:0] csr_depc_o;
wire [31:0] csr_depc_o;
/* cellift = 32'd1 */
output [31:0] csr_depc_o_t0;
wire [31:0] csr_depc_o_t0;
/* src = "generated/sv2v_out.v:13824.19-13824.31" */
input [6:0] csr_mcause_i;
wire [6:0] csr_mcause_i;
/* cellift = 32'd1 */
input [6:0] csr_mcause_i_t0;
wire [6:0] csr_mcause_i_t0;
/* src = "generated/sv2v_out.v:13793.21-13793.31" */
output [31:0] csr_mepc_o;
wire [31:0] csr_mepc_o;
/* cellift = 32'd1 */
output [31:0] csr_mepc_o_t0;
wire [31:0] csr_mepc_o_t0;
/* src = "generated/sv2v_out.v:13792.14-13792.31" */
output csr_mstatus_mie_o;
wire csr_mstatus_mie_o;
/* cellift = 32'd1 */
output csr_mstatus_mie_o_t0;
wire csr_mstatus_mie_o_t0;
/* src = "generated/sv2v_out.v:13775.14-13775.30" */
output csr_mstatus_tw_o;
wire csr_mstatus_tw_o;
/* cellift = 32'd1 */
output csr_mstatus_tw_o_t0;
wire csr_mstatus_tw_o_t0;
/* src = "generated/sv2v_out.v:13825.20-13825.31" */
input [31:0] csr_mtval_i;
wire [31:0] csr_mtval_i;
/* cellift = 32'd1 */
input [31:0] csr_mtval_i_t0;
wire [31:0] csr_mtval_i_t0;
/* src = "generated/sv2v_out.v:13794.21-13794.32" */
output [31:0] csr_mtval_o;
wire [31:0] csr_mtval_o;
/* cellift = 32'd1 */
output [31:0] csr_mtval_o_t0;
wire [31:0] csr_mtval_o_t0;
/* src = "generated/sv2v_out.v:13777.13-13777.29" */
input csr_mtvec_init_i;
wire csr_mtvec_init_i;
/* cellift = 32'd1 */
input csr_mtvec_init_i_t0;
wire csr_mtvec_init_i_t0;
/* src = "generated/sv2v_out.v:13776.21-13776.32" */
output [31:0] csr_mtvec_o;
wire [31:0] csr_mtvec_o;
/* cellift = 32'd1 */
output [31:0] csr_mtvec_o_t0;
wire [31:0] csr_mtvec_o_t0;
/* src = "generated/sv2v_out.v:13783.8-13783.19" */
input csr_op_en_i;
wire csr_op_en_i;
/* cellift = 32'd1 */
input csr_op_en_i_t0;
wire csr_op_en_i_t0;
/* src = "generated/sv2v_out.v:13782.19-13782.27" */
input [1:0] csr_op_i;
wire [1:0] csr_op_i;
/* cellift = 32'd1 */
input [1:0] csr_op_i_t0;
wire [1:0] csr_op_i_t0;
/* src = "generated/sv2v_out.v:13796.43-13796.57" */
output [135:0] csr_pmp_addr_o;
wire [135:0] csr_pmp_addr_o;
/* cellift = 32'd1 */
output [135:0] csr_pmp_addr_o_t0;
wire [135:0] csr_pmp_addr_o_t0;
/* src = "generated/sv2v_out.v:13795.42-13795.55" */
output [23:0] csr_pmp_cfg_o;
wire [23:0] csr_pmp_cfg_o;
/* cellift = 32'd1 */
output [23:0] csr_pmp_cfg_o_t0;
wire [23:0] csr_pmp_cfg_o_t0;
/* src = "generated/sv2v_out.v:13797.20-13797.37" */
output [2:0] csr_pmp_mseccfg_o;
wire [2:0] csr_pmp_mseccfg_o;
/* cellift = 32'd1 */
output [2:0] csr_pmp_mseccfg_o_t0;
wire [2:0] csr_pmp_mseccfg_o_t0;
/* src = "generated/sv2v_out.v:13784.21-13784.32" */
output [31:0] csr_rdata_o;
wire [31:0] csr_rdata_o;
/* cellift = 32'd1 */
output [31:0] csr_rdata_o_t0;
wire [31:0] csr_rdata_o_t0;
/* src = "generated/sv2v_out.v:13822.13-13822.31" */
input csr_restore_dret_i;
wire csr_restore_dret_i;
/* cellift = 32'd1 */
input csr_restore_dret_i_t0;
wire csr_restore_dret_i_t0;
/* src = "generated/sv2v_out.v:13821.13-13821.31" */
input csr_restore_mret_i;
wire csr_restore_mret_i;
/* cellift = 32'd1 */
input csr_restore_mret_i_t0;
wire csr_restore_mret_i_t0;
/* src = "generated/sv2v_out.v:13823.13-13823.29" */
input csr_save_cause_i;
wire csr_save_cause_i;
/* cellift = 32'd1 */
input csr_save_cause_i_t0;
wire csr_save_cause_i_t0;
/* src = "generated/sv2v_out.v:13819.13-13819.26" */
input csr_save_id_i;
wire csr_save_id_i;
/* cellift = 32'd1 */
input csr_save_id_i_t0;
wire csr_save_id_i_t0;
/* src = "generated/sv2v_out.v:13818.13-13818.26" */
input csr_save_if_i;
wire csr_save_if_i;
/* cellift = 32'd1 */
input csr_save_if_i_t0;
wire csr_save_if_i_t0;
/* src = "generated/sv2v_out.v:13820.13-13820.26" */
input csr_save_wb_i;
wire csr_save_wb_i;
/* cellift = 32'd1 */
input csr_save_wb_i_t0;
wire csr_save_wb_i_t0;
/* src = "generated/sv2v_out.v:13816.14-13816.30" */
output csr_shadow_err_o;
wire csr_shadow_err_o;
/* cellift = 32'd1 */
output csr_shadow_err_o_t0;
wire csr_shadow_err_o_t0;
/* src = "generated/sv2v_out.v:13781.20-13781.31" */
input [31:0] csr_wdata_i;
wire [31:0] csr_wdata_i;
/* cellift = 32'd1 */
input [31:0] csr_wdata_i_t0;
wire [31:0] csr_wdata_i_t0;
/* src = "generated/sv2v_out.v:13942.7-13942.17" */
wire csr_we_int;
/* src = "generated/sv2v_out.v:13943.7-13943.13" */
wire csr_wr;
/* src = "generated/sv2v_out.v:13810.14-13810.31" */
output data_ind_timing_o;
wire data_ind_timing_o;
/* cellift = 32'd1 */
output data_ind_timing_o_t0;
wire data_ind_timing_o_t0;
/* src = "generated/sv2v_out.v:13944.6-13944.13" */
wire dbg_csr;
/* src = "generated/sv2v_out.v:13892.13-13892.19" */
wire [31:0] dcsr_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13892.13-13892.19" */
wire [31:0] dcsr_d_t0;
/* src = "generated/sv2v_out.v:13893.6-13893.13" */
wire dcsr_en;
/* src = "generated/sv2v_out.v:13891.14-13891.20" */
wire [31:0] dcsr_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13891.14-13891.20" */
wire [31:0] dcsr_q_t0;
/* src = "generated/sv2v_out.v:13800.19-13800.32" */
input [2:0] debug_cause_i;
wire [2:0] debug_cause_i;
/* cellift = 32'd1 */
input [2:0] debug_cause_i_t0;
wire [2:0] debug_cause_i_t0;
/* src = "generated/sv2v_out.v:13801.13-13801.29" */
input debug_csr_save_i;
wire debug_csr_save_i;
/* cellift = 32'd1 */
input debug_csr_save_i_t0;
wire debug_csr_save_i_t0;
/* src = "generated/sv2v_out.v:13804.14-13804.29" */
output debug_ebreakm_o;
wire debug_ebreakm_o;
/* cellift = 32'd1 */
output debug_ebreakm_o_t0;
wire debug_ebreakm_o_t0;
/* src = "generated/sv2v_out.v:13805.14-13805.29" */
output debug_ebreaku_o;
wire debug_ebreaku_o;
/* cellift = 32'd1 */
output debug_ebreaku_o_t0;
wire debug_ebreaku_o_t0;
/* src = "generated/sv2v_out.v:13799.13-13799.34" */
input debug_mode_entering_i;
wire debug_mode_entering_i;
/* cellift = 32'd1 */
input debug_mode_entering_i_t0;
wire debug_mode_entering_i_t0;
/* src = "generated/sv2v_out.v:13798.13-13798.25" */
input debug_mode_i;
wire debug_mode_i;
/* cellift = 32'd1 */
input debug_mode_i_t0;
wire debug_mode_i_t0;
/* src = "generated/sv2v_out.v:13803.14-13803.33" */
output debug_single_step_o;
wire debug_single_step_o;
/* cellift = 32'd1 */
output debug_single_step_o_t0;
wire debug_single_step_o_t0;
/* src = "generated/sv2v_out.v:13895.13-13895.19" */
wire [31:0] depc_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13895.13-13895.19" */
wire [31:0] depc_d_t0;
/* src = "generated/sv2v_out.v:13896.6-13896.13" */
wire depc_en;
/* src = "generated/sv2v_out.v:13840.13-13840.23" */
input div_wait_i;
wire div_wait_i;
/* cellift = 32'd1 */
input div_wait_i_t0;
wire div_wait_i_t0;
/* src = "generated/sv2v_out.v:13827.13-13827.32" */
output double_fault_seen_o;
wire double_fault_seen_o;
/* cellift = 32'd1 */
output double_fault_seen_o_t0;
wire double_fault_seen_o_t0;
/* src = "generated/sv2v_out.v:13899.6-13899.18" */
wire dscratch0_en;
/* src = "generated/sv2v_out.v:13897.14-13897.25" */
wire [31:0] dscratch0_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13897.14-13897.25" */
wire [31:0] dscratch0_q_t0;
/* src = "generated/sv2v_out.v:13900.6-13900.18" */
wire dscratch1_en;
/* src = "generated/sv2v_out.v:13898.14-13898.25" */
wire [31:0] dscratch1_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13898.14-13898.25" */
wire [31:0] dscratch1_q_t0;
/* src = "generated/sv2v_out.v:13838.13-13838.25" */
input dside_wait_i;
wire dside_wait_i;
/* cellift = 32'd1 */
input dside_wait_i_t0;
wire dside_wait_i_t0;
/* src = "generated/sv2v_out.v:13811.14-13811.30" */
output dummy_instr_en_o;
wire dummy_instr_en_o;
/* cellift = 32'd1 */
output dummy_instr_en_o_t0;
wire dummy_instr_en_o_t0;
/* src = "generated/sv2v_out.v:13812.20-13812.38" */
output [2:0] dummy_instr_mask_o;
wire [2:0] dummy_instr_mask_o;
/* cellift = 32'd1 */
output [2:0] dummy_instr_mask_o_t0;
wire [2:0] dummy_instr_mask_o_t0;
/* src = "generated/sv2v_out.v:13813.14-13813.35" */
output dummy_instr_seed_en_o;
wire dummy_instr_seed_en_o;
/* cellift = 32'd1 */
output dummy_instr_seed_en_o_t0;
wire dummy_instr_seed_en_o_t0;
/* src = "generated/sv2v_out.v:13814.21-13814.39" */
output [31:0] dummy_instr_seed_o;
wire [31:0] dummy_instr_seed_o;
/* cellift = 32'd1 */
output [31:0] dummy_instr_seed_o_t0;
wire [31:0] dummy_instr_seed_o_t0;
/* src = "generated/sv2v_out.v:13772.20-13772.29" */
input [31:0] hart_id_i;
wire [31:0] hart_id_i;
/* cellift = 32'd1 */
input [31:0] hart_id_i_t0;
wire [31:0] hart_id_i_t0;
/* src = "generated/sv2v_out.v:13817.13-13817.31" */
input ic_scr_key_valid_i;
wire ic_scr_key_valid_i;
/* cellift = 32'd1 */
input ic_scr_key_valid_i_t0;
wire ic_scr_key_valid_i_t0;
/* src = "generated/sv2v_out.v:13815.14-13815.29" */
output icache_enable_o;
wire icache_enable_o;
/* cellift = 32'd1 */
output icache_enable_o_t0;
wire icache_enable_o_t0;
/* src = "generated/sv2v_out.v:13945.6-13945.17" */
wire illegal_csr;
/* src = "generated/sv2v_out.v:13947.7-13947.22" */
wire illegal_csr_dbg;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13947.7-13947.22" */
wire illegal_csr_dbg_t0;
/* src = "generated/sv2v_out.v:13826.14-13826.32" */
output illegal_csr_insn_o;
wire illegal_csr_insn_o;
/* cellift = 32'd1 */
output illegal_csr_insn_o_t0;
wire illegal_csr_insn_o_t0;
/* src = "generated/sv2v_out.v:13946.7-13946.23" */
wire illegal_csr_priv;
/* src = "generated/sv2v_out.v:13948.7-13948.24" */
wire illegal_csr_write;
/* src = "generated/sv2v_out.v:13829.13-13829.35" */
input instr_ret_compressed_i;
wire instr_ret_compressed_i;
/* cellift = 32'd1 */
input instr_ret_compressed_i_t0;
wire instr_ret_compressed_i_t0;
/* src = "generated/sv2v_out.v:13831.13-13831.40" */
input instr_ret_compressed_spec_i;
wire instr_ret_compressed_spec_i;
/* cellift = 32'd1 */
input instr_ret_compressed_spec_i_t0;
wire instr_ret_compressed_spec_i_t0;
/* src = "generated/sv2v_out.v:13828.13-13828.24" */
input instr_ret_i;
wire instr_ret_i;
/* cellift = 32'd1 */
input instr_ret_i_t0;
wire instr_ret_i_t0;
/* src = "generated/sv2v_out.v:13830.13-13830.29" */
input instr_ret_spec_i;
wire instr_ret_spec_i;
/* cellift = 32'd1 */
input instr_ret_spec_i_t0;
wire instr_ret_spec_i_t0;
/* src = "generated/sv2v_out.v:13787.13-13787.27" */
input irq_external_i;
wire irq_external_i;
/* cellift = 32'd1 */
input irq_external_i_t0;
wire irq_external_i_t0;
/* src = "generated/sv2v_out.v:13788.20-13788.30" */
input [14:0] irq_fast_i;
wire [14:0] irq_fast_i;
/* cellift = 32'd1 */
input [14:0] irq_fast_i_t0;
wire [14:0] irq_fast_i_t0;
/* src = "generated/sv2v_out.v:13790.14-13790.27" */
output irq_pending_o;
wire irq_pending_o;
/* cellift = 32'd1 */
output irq_pending_o_t0;
wire irq_pending_o_t0;
/* src = "generated/sv2v_out.v:13785.13-13785.27" */
input irq_software_i;
wire irq_software_i;
/* cellift = 32'd1 */
input irq_software_i_t0;
wire irq_software_i_t0;
/* src = "generated/sv2v_out.v:13786.13-13786.24" */
input irq_timer_i;
wire irq_timer_i;
/* cellift = 32'd1 */
input irq_timer_i_t0;
wire irq_timer_i_t0;
/* src = "generated/sv2v_out.v:13791.21-13791.27" */
output [17:0] irqs_o;
wire [17:0] irqs_o;
/* cellift = 32'd1 */
output [17:0] irqs_o_t0;
wire [17:0] irqs_o_t0;
/* src = "generated/sv2v_out.v:13832.13-13832.25" */
input iside_wait_i;
wire iside_wait_i;
/* cellift = 32'd1 */
input iside_wait_i_t0;
wire iside_wait_i_t0;
/* src = "generated/sv2v_out.v:13833.13-13833.19" */
input jump_i;
wire jump_i;
/* cellift = 32'd1 */
input jump_i_t0;
wire jump_i_t0;
/* src = "generated/sv2v_out.v:13881.12-13881.20" */
wire [6:0] mcause_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13881.12-13881.20" */
wire [6:0] mcause_d_t0;
/* src = "generated/sv2v_out.v:13882.6-13882.15" */
wire mcause_en;
/* src = "generated/sv2v_out.v:13880.13-13880.21" */
wire [6:0] mcause_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13880.13-13880.21" */
wire [6:0] mcause_q_t0;
/* src = "generated/sv2v_out.v:13914.14-13914.27" */
wire [31:0] mcountinhibit;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13914.14-13914.27" */
wire [31:0] mcountinhibit_t0;
/* src = "generated/sv2v_out.v:13917.6-13917.22" */
wire mcountinhibit_we;
/* src = "generated/sv2v_out.v:13836.13-13836.23" */
input mem_load_i;
wire mem_load_i;
/* cellift = 32'd1 */
input mem_load_i_t0;
wire mem_load_i_t0;
/* src = "generated/sv2v_out.v:13837.13-13837.24" */
input mem_store_i;
wire mem_store_i;
/* cellift = 32'd1 */
input mem_store_i_t0;
wire mem_store_i_t0;
/* src = "generated/sv2v_out.v:13878.13-13878.19" */
wire [31:0] mepc_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13878.13-13878.19" */
wire [31:0] mepc_d_t0;
/* src = "generated/sv2v_out.v:13879.6-13879.13" */
wire mepc_en;
/* src = "generated/sv2v_out.v:13918.14-13918.25" */
wire [63:0] \mhpmcounter[0] ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13918.14-13918.25" */
wire [63:0] \mhpmcounter[0]_t0 ;
/* src = "generated/sv2v_out.v:13918.14-13918.25" */
wire [63:0] \mhpmcounter[2] ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13918.14-13918.25" */
wire [63:0] \mhpmcounter[2]_t0 ;
/* src = "generated/sv2v_out.v:13919.13-13919.27" */
/* unused_bits = "1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] mhpmcounter_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13919.13-13919.27" */
/* unused_bits = "1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] mhpmcounter_we_t0;
/* src = "generated/sv2v_out.v:13920.13-13920.28" */
/* unused_bits = "1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] mhpmcounterh_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13920.13-13920.28" */
/* unused_bits = "1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] mhpmcounterh_we_t0;
/* src = "generated/sv2v_out.v:13874.6-13874.12" */
wire mie_en;
/* src = "generated/sv2v_out.v:13872.14-13872.19" */
wire [17:0] mie_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13872.14-13872.19" */
wire [17:0] mie_q_t0;
/* src = "generated/sv2v_out.v:13927.14-13927.27" */
wire [63:0] minstret_next;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13927.14-13927.27" */
wire [63:0] minstret_next_t0;
/* src = "generated/sv2v_out.v:13928.14-13928.26" */
wire [63:0] minstret_raw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13928.14-13928.26" */
wire [63:0] minstret_raw_t0;
/* src = "generated/sv2v_out.v:13876.6-13876.17" */
wire mscratch_en;
/* src = "generated/sv2v_out.v:13875.14-13875.24" */
wire [31:0] mscratch_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13875.14-13875.24" */
wire [31:0] mscratch_q_t0;
/* src = "generated/sv2v_out.v:13906.13-13906.27" */
wire [6:0] mstack_cause_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13906.13-13906.27" */
wire [6:0] mstack_cause_q_t0;
/* src = "generated/sv2v_out.v:13903.6-13903.15" */
wire mstack_en;
/* src = "generated/sv2v_out.v:13904.14-13904.26" */
wire [31:0] mstack_epc_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13904.14-13904.26" */
wire [31:0] mstack_epc_q_t0;
/* src = "generated/sv2v_out.v:13901.13-13901.21" */
wire [2:0] mstack_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13901.13-13901.21" */
wire [2:0] mstack_q_t0;
/* src = "generated/sv2v_out.v:13869.12-13869.21" */
wire [5:0] mstatus_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13869.12-13869.21" */
wire [5:0] mstatus_d_t0;
/* src = "generated/sv2v_out.v:13871.6-13871.16" */
wire mstatus_en;
/* src = "generated/sv2v_out.v:13870.7-13870.18" */
wire mstatus_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13870.7-13870.18" */
wire mstatus_err_t0;
/* src = "generated/sv2v_out.v:13868.13-13868.22" */
wire [5:0] mstatus_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13868.13-13868.22" */
wire [5:0] mstatus_q_t0;
/* src = "generated/sv2v_out.v:13884.13-13884.20" */
wire [31:0] mtval_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13884.13-13884.20" */
wire [31:0] mtval_d_t0;
/* src = "generated/sv2v_out.v:13885.6-13885.14" */
wire mtval_en;
/* src = "generated/sv2v_out.v:13887.13-13887.20" */
wire [31:0] mtvec_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13887.13-13887.20" */
wire [31:0] mtvec_d_t0;
/* src = "generated/sv2v_out.v:13889.6-13889.14" */
wire mtvec_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13889.6-13889.14" */
wire mtvec_en_t0;
/* src = "generated/sv2v_out.v:13888.7-13888.16" */
wire mtvec_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13888.7-13888.16" */
wire mtvec_err_t0;
/* src = "generated/sv2v_out.v:13839.13-13839.23" */
input mul_wait_i;
wire mul_wait_i;
/* cellift = 32'd1 */
input mul_wait_i_t0;
wire mul_wait_i_t0;
/* src = "generated/sv2v_out.v:13789.13-13789.23" */
input nmi_mode_i;
wire nmi_mode_i;
/* cellift = 32'd1 */
input nmi_mode_i_t0;
wire nmi_mode_i_t0;
/* src = "generated/sv2v_out.v:13808.20-13808.27" */
input [31:0] pc_id_i;
wire [31:0] pc_id_i;
/* cellift = 32'd1 */
input [31:0] pc_id_i_t0;
wire [31:0] pc_id_i_t0;
/* src = "generated/sv2v_out.v:13807.20-13807.27" */
input [31:0] pc_if_i;
wire [31:0] pc_if_i;
/* cellift = 32'd1 */
input [31:0] pc_if_i_t0;
wire [31:0] pc_if_i_t0;
/* src = "generated/sv2v_out.v:13809.20-13809.27" */
input [31:0] pc_wb_i;
wire [31:0] pc_wb_i;
/* cellift = 32'd1 */
input [31:0] pc_wb_i_t0;
wire [31:0] pc_wb_i_t0;
/* src = "generated/sv2v_out.v:13867.12-13867.22" */
wire [1:0] priv_lvl_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13867.12-13867.22" */
wire [1:0] priv_lvl_d_t0;
/* src = "generated/sv2v_out.v:13773.20-13773.34" */
output [1:0] priv_mode_id_o;
reg [1:0] priv_mode_id_o;
/* cellift = 32'd1 */
output [1:0] priv_mode_id_o_t0;
reg [1:0] priv_mode_id_o_t0;
/* src = "generated/sv2v_out.v:13774.20-13774.35" */
output [1:0] priv_mode_lsu_o;
wire [1:0] priv_mode_lsu_o;
/* cellift = 32'd1 */
output [1:0] priv_mode_lsu_o_t0;
wire [1:0] priv_mode_lsu_o_t0;
/* src = "generated/sv2v_out.v:13771.13-13771.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:13806.14-13806.29" */
output trigger_match_o;
wire trigger_match_o;
/* cellift = 32'd1 */
output trigger_match_o_t0;
wire trigger_match_o_t0;
assign illegal_csr_dbg = dbg_csr & /* src = "generated/sv2v_out.v:13956.27-13956.50" */ _0208_;
assign illegal_csr_insn_o = csr_access_i & /* src = "generated/sv2v_out.v:13959.30-13959.119" */ _1241_;
assign _0106_ = _0245_ & /* src = "generated/sv2v_out.v:14268.26-14268.52" */ csr_rdata_o;
assign _0108_ = csr_wr & /* src = "generated/sv2v_out.v:14273.23-14273.43" */ csr_op_en_i;
assign csr_we_int = _0108_ & /* src = "generated/sv2v_out.v:14273.22-14273.66" */ _1233_;
assign irqs_o = { irq_software_i, irq_timer_i, irq_external_i, irq_fast_i } & /* src = "generated/sv2v_out.v:14284.18-14284.29" */ mie_q;
assign _0110_ = instr_ret_i & /* src = "generated/sv2v_out.v:14657.18-14657.57" */ _1234_;
assign _0112_ = instr_ret_spec_i & /* src = "generated/sv2v_out.v:14664.27-14664.63" */ _1234_;
assign icache_enable_o = cpuctrlsts_part_q[0] & /* src = "generated/sv2v_out.v:14868.27-14868.89" */ _1235_;
assign _0113_ = ~ _0265_;
assign _0114_ = ~ mcountinhibit_we;
assign _0286_ = { _0265_, _0265_ } & priv_lvl_d_t0;
assign _0288_ = { mcountinhibit_we, mcountinhibit_we } & { dummy_instr_seed_o_t0[2], dummy_instr_seed_o_t0[0] };
assign _0287_ = { _0113_, _0113_ } & priv_mode_id_o_t0;
assign _0289_ = { _0114_, _0114_ } & { mcountinhibit_t0[2], mcountinhibit_t0[0] };
assign _0784_ = _0286_ | _0287_;
assign _0785_ = _0288_ | _0289_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers  */
/* PC_TAINT_INFO STATE_NAME priv_mode_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) priv_mode_id_o_t0 <= 2'h0;
else priv_mode_id_o_t0 <= _0784_;
reg [1:0] _1372_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers  */
/* PC_TAINT_INFO STATE_NAME _1372_ */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) _1372_ <= 2'h0;
else _1372_ <= _0785_;
assign { mcountinhibit_t0[2], mcountinhibit_t0[0] } = _1372_;
assign _0271_ = csr_access_i_t0 & _1241_;
assign _0274_ = csr_wdata_i_t0 & csr_rdata_o;
assign _0277_ = { irq_software_i_t0, irq_timer_i_t0, irq_external_i_t0, irq_fast_i_t0 } & mie_q;
assign _0280_ = instr_ret_i_t0 & _1234_;
assign _0283_ = cpuctrlsts_part_q_t0[0] & _1235_;
assign illegal_csr_dbg_t0 = debug_mode_i_t0 & dbg_csr;
assign _0272_ = _1242_ & csr_access_i;
assign _0278_ = mie_q_t0 & { irq_software_i, irq_timer_i, irq_external_i, irq_fast_i };
assign _0281_ = mcountinhibit_t0[2] & instr_ret_i;
assign _0284_ = _1236_ & cpuctrlsts_part_q[0];
assign _0273_ = csr_access_i_t0 & _1242_;
assign _0276_ = csr_wdata_i_t0 & csr_rdata_o_t0;
assign _0279_ = { irq_software_i_t0, irq_timer_i_t0, irq_external_i_t0, irq_fast_i_t0 } & mie_q_t0;
assign _0282_ = instr_ret_i_t0 & mcountinhibit_t0[2];
assign _0285_ = cpuctrlsts_part_q_t0[0] & _1236_;
assign _0779_ = _0271_ | _0272_;
assign _0780_ = _0274_ | _0275_;
assign _0781_ = _0277_ | _0278_;
assign _0782_ = _0280_ | _0281_;
assign _0783_ = _0283_ | _0284_;
assign illegal_csr_insn_o_t0 = _0779_ | _0273_;
assign _0107_ = _0780_ | _0276_;
assign irqs_o_t0 = _0781_ | _0279_;
assign _0111_ = _0782_ | _0282_;
assign icache_enable_o_t0 = _0783_ | _0285_;
/* src = "generated/sv2v_out.v:14257.2-14261.29" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers  */
/* PC_TAINT_INFO STATE_NAME priv_mode_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) priv_mode_id_o <= 2'h3;
else if (_0265_) priv_mode_id_o <= priv_lvl_d;
reg [1:0] _1399_;
/* src = "generated/sv2v_out.v:14719.2-14723.39" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers  */
/* PC_TAINT_INFO STATE_NAME _1399_ */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) _1399_ <= 2'h0;
else if (mcountinhibit_we) _1399_ <= { dummy_instr_seed_o[2], dummy_instr_seed_o[0] };
assign { mcountinhibit[2], mcountinhibit[0] } = _1399_;
assign _0116_ = ~ { _0254_, _0254_, _0254_ };
assign _0119_ = ~ _1299_;
assign _0123_ = ~ _0255_;
assign _0127_ = ~ _1306_;
assign _0128_ = ~ _1292_;
assign _0130_ = ~ _0253_;
assign _0131_ = ~ _0256_;
assign _0133_ = ~ { _0768_, _0768_, _0768_ };
assign _0134_ = ~ { _1298_, _1298_, _1298_ };
assign _0135_ = ~ { _1301_, _1301_, _1301_ };
assign _0137_ = ~ { _0772_, _0772_, _0772_ };
assign _0139_ = ~ { _1303_, _1303_, _1303_ };
assign _0141_ = ~ { _0770_, _0770_, _0770_ };
assign _0144_ = ~ { _0257_, _0257_, _0257_ };
assign _0145_ = ~ { _1294_, _1294_, _1294_ };
assign _0146_ = ~ { _1299_, _1299_, _1299_ };
assign _0147_ = ~ { _0769_, _0769_, _0769_ };
assign _0148_ = ~ { _0258_, _0258_, _0258_ };
assign _0140_ = ~ { _1305_, _1305_, _1305_ };
assign _0142_ = ~ { _1306_, _1306_, _1306_ };
assign _0143_ = ~ { _0773_, _0773_, _0773_ };
assign _0149_ = ~ { _0259_, _0259_, _0259_ };
assign _0150_ = ~ { _1310_, _1310_, _1310_ };
assign _0151_ = ~ { _0774_, _0774_, _0774_ };
assign _0136_ = ~ { _1300_, _1300_, _1300_ };
assign _0152_ = ~ { _1291_, _1291_, _1291_ };
assign _0153_ = ~ { _0775_, _0775_, _0775_ };
assign _0154_ = ~ { _0260_, _0260_, _0260_ };
assign _0155_ = ~ { _1346_, _1346_, _1346_ };
assign _0156_ = ~ { _0771_, _0771_, _0771_ };
assign _0115_ = ~ { _0253_, _0253_, _0253_ };
assign _0157_ = ~ { _0261_, _0261_, _0261_ };
assign _0166_ = ~ _0776_;
assign _0168_ = ~ _0777_;
assign _0169_ = ~ _0262_;
assign _0170_ = ~ _0263_;
assign _0172_ = ~ { _1304_, _1304_, _1304_ };
assign _0173_ = ~ { _1302_, _1302_, _1302_ };
assign _0174_ = ~ { _0778_, _0778_, _0778_ };
assign _0175_ = ~ { _0264_, _0264_, _0264_ };
assign _0176_ = ~ { _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_ };
assign _0177_ = ~ { _1310_, _1310_, _1310_, _1310_, _1310_, _1310_, _1310_, _1310_, _1310_ };
assign _0178_ = ~ { _0774_, _0774_, _0774_, _0774_, _0774_, _0774_, _0774_, _0774_, _0774_ };
assign _0179_ = ~ { _1300_, _1300_, _1300_, _1300_, _1300_, _1300_, _1300_, _1300_, _1300_ };
assign _0180_ = ~ { _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_ };
assign _0181_ = ~ { _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_ };
assign _0182_ = ~ { _0260_, _0260_, _0260_, _0260_, _0260_, _0260_, _0260_, _0260_, _0260_ };
assign _0183_ = ~ { _1305_, _1305_, _1305_, _1305_, _1305_, _1305_, _1305_, _1305_, _1305_ };
assign _0184_ = ~ { _0770_, _0770_, _0770_, _0770_, _0770_, _0770_, _0770_, _0770_, _0770_ };
assign _0185_ = ~ { _1306_, _1306_, _1306_, _1306_, _1306_, _1306_, _1306_, _1306_, _1306_ };
assign _0186_ = ~ { _1346_, _1346_, _1346_, _1346_, _1346_, _1346_, _1346_, _1346_, _1346_ };
assign _0187_ = ~ { _0771_, _0771_, _0771_, _0771_, _0771_, _0771_, _0771_, _0771_, _0771_ };
assign _0188_ = ~ { _0253_, _0253_, _0253_, _0253_, _0253_, _0253_, _0253_, _0253_, _0253_ };
assign _0189_ = ~ { _0261_, _0261_, _0261_, _0261_, _0261_, _0261_, _0261_, _0261_, _0261_ };
assign _0162_ = ~ _0775_;
assign _0125_ = ~ _1305_;
assign _0190_ = ~ { _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_ };
assign _0191_ = ~ { _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_ };
assign _0158_ = ~ _1294_;
assign _0159_ = ~ _1310_;
assign _0160_ = ~ _0774_;
assign _0161_ = ~ _1300_;
assign _0163_ = ~ _0260_;
assign _0129_ = ~ _0771_;
assign _0171_ = ~ _0261_;
assign _0192_ = ~ { _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_ };
assign _0193_ = ~ { _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_ };
assign _0121_ = ~ _1301_;
assign _0122_ = ~ _0769_;
assign _0194_ = ~ _0258_;
assign _0164_ = ~ _1304_;
assign _0165_ = ~ _1302_;
assign _0195_ = ~ _0778_;
assign _0196_ = ~ _0264_;
assign _0197_ = ~ _0259_;
assign _0118_ = ~ _0768_;
assign _0124_ = ~ _1303_;
assign _0126_ = ~ _0770_;
assign _0132_ = ~ { _1297_, _1297_, _1297_ };
assign _0138_ = ~ { _0255_, _0255_, _0255_ };
assign _0199_ = ~ { nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i };
assign _0200_ = ~ _1231_;
assign _0201_ = ~ { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
assign _0202_ = ~ { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
assign _0207_ = ~ _1226_;
assign _0206_ = ~ cpuctrlsts_part_q[6];
assign _0210_ = ~ { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i };
assign _0211_ = ~ { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i };
assign _0209_ = ~ { debug_mode_i, debug_mode_i };
assign _0212_ = ~ { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
assign _0213_ = ~ { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
assign _0214_ = ~ { debug_csr_save_i, debug_csr_save_i };
assign _0215_ = ~ { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
assign _0216_ = ~ { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
assign _0217_ = ~ { csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i };
assign _0218_ = ~ { csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i };
assign _0219_ = ~ { csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i };
assign _0204_ = ~ csr_restore_mret_i;
assign _0205_ = ~ csr_restore_dret_i;
assign _0198_ = ~ csr_save_cause_i;
assign _0203_ = ~ { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
assign _0221_ = ~ { csr_save_cause_i, csr_save_cause_i };
assign _0220_ = ~ { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
assign _0222_ = ~ { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
assign _0223_ = ~ { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
assign _0224_ = ~ { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
assign _0225_ = ~ { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
assign _0226_ = ~ { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
assign _0227_ = ~ { nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i };
assign _0228_ = ~ { csr_restore_dret_i, csr_restore_dret_i };
assign _0208_ = ~ debug_mode_i;
assign _0229_ = ~ { _1291_, _1291_, _1291_, _1291_ };
assign _0230_ = ~ { _1292_, _1292_ };
assign _0231_ = ~ { _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_ };
assign _0232_ = ~ { _1291_, _1291_ };
assign _0120_ = ~ _1291_;
assign _0233_ = ~ { _1225_, _1225_ };
assign _0234_ = ~ { _1224_, _1224_ };
assign _0117_ = ~ _1297_;
assign _0235_ = ~ { _1297_, _1297_, _1297_, _1297_, _1297_, _1297_, _1297_, _1297_ };
assign _0237_ = ~ { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int };
assign _0238_ = ~ { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int };
assign _0236_ = ~ csr_we_int;
assign _0239_ = ~ { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int };
assign _0240_ = ~ { csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i };
assign _0241_ = ~ { mstatus_q[1], mstatus_q[1] };
assign _0242_ = ~ { _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_ };
assign _0290_ = _0115_ & _0795_;
assign _0292_ = _0116_ & _0797_;
assign _0294_ = _0117_ & _0015_[35];
assign _0296_ = _0118_ & _0801_;
assign _0298_ = _0119_ & dscratch0_q_t0[3];
assign _0300_ = _0120_ & irq_software_i_t0;
assign _0302_ = _0121_ & _0807_;
assign _0304_ = _0122_ & _0809_;
assign _0306_ = _0123_ & _0811_;
assign _0308_ = _0124_ & mcause_q_t0[3];
assign _0310_ = _0125_ & csr_mtvec_o_t0[3];
assign _0312_ = _0126_ & _0817_;
assign _0314_ = _0127_ & mie_q_t0[17];
assign _0316_ = _0128_ & _0823_;
assign _0318_ = _0129_ & _0825_;
assign _0320_ = _0130_ & _0827_;
assign _0322_ = _0131_ & _0829_;
assign _0324_ = _0132_ & _0015_[34:32];
assign _0326_ = _0133_ & _0833_;
assign _0328_ = _0134_ & dscratch1_q_t0[2:0];
assign _0330_ = _0135_ & dcsr_q_t0[2:0];
assign _0332_ = _0136_ & _0839_;
assign _0334_ = _0137_ & _0841_;
assign _0336_ = _0138_ & _0843_;
assign _0338_ = _0139_ & mcause_q_t0[2:0];
assign _0340_ = _0140_ & csr_mtvec_o_t0[2:0];
assign _0342_ = _0141_ & _0849_;
assign _0344_ = _0143_ & _0856_;
assign _0346_ = _0115_ & _0858_;
assign _0348_ = _0144_ & _0860_;
assign _0350_ = _0145_ & _0862_;
assign _0352_ = _0146_ & dscratch0_q_t0[10:8];
assign _0354_ = _0135_ & dcsr_q_t0[10:8];
assign _0356_ = _0147_ & _0868_;
assign _0358_ = _0148_ & _0870_;
assign _0360_ = _0140_ & csr_mtvec_o_t0[10:8];
assign _0362_ = _0141_ & _0876_;
assign _0364_ = _0143_ & _0882_;
assign _0366_ = _0115_ & _0884_;
assign _0368_ = _0149_ & _0886_;
assign _0370_ = _0145_ & _0015_[20:18];
assign _0890_ = _0150_ & dscratch1_q_t0[20:18];
assign _0372_ = _0151_ & _0890_;
assign _0374_ = _0136_ & csr_depc_o_t0[20:18];
assign _0376_ = _0152_ & irq_fast_i_t0[4:2];
assign _0378_ = _0153_ & _0896_;
assign _0380_ = _0154_ & _0898_;
assign _0382_ = _0140_ & csr_mtvec_o_t0[20:18];
assign _0384_ = _0141_ & _0904_;
assign _0386_ = _0142_ & mie_q_t0[4:2];
assign _0912_ = _0155_ & _0910_;
assign _0388_ = _0156_ & _0912_;
assign _0390_ = _0115_ & _0914_;
assign _0392_ = _0157_ & _0916_;
assign _0394_ = _0158_ & _0015_[12];
assign _0920_ = _0159_ & dscratch1_q_t0[12];
assign _0396_ = _0160_ & _0920_;
assign _0398_ = _0161_ & csr_depc_o_t0[12];
assign _0400_ = _0120_ & csr_mtval_o_t0[12];
assign _0402_ = _0162_ & _0926_;
assign _0404_ = _0163_ & _0928_;
assign _0932_ = _0164_ & csr_mepc_o_t0[12];
assign _0406_ = _0165_ & mscratch_q_t0[12];
assign _0408_ = _0166_ & _0934_;
assign _0938_ = _0167_ & mstatus_q_t0[3];
assign _0410_ = _0168_ & _0940_;
assign _0412_ = _0169_ & _0942_;
assign _0414_ = _0170_ & _0944_;
assign _0416_ = _0158_ & _0015_[17];
assign _0948_ = _0159_ & dscratch1_q_t0[17];
assign _0418_ = _0160_ & _0948_;
assign _0420_ = _0161_ & csr_depc_o_t0[17];
assign _0422_ = _0120_ & irq_fast_i_t0[1];
assign _0424_ = _0162_ & _0954_;
assign _0426_ = _0163_ & _0956_;
assign _0428_ = _0125_ & csr_mtvec_o_t0[17];
assign _0430_ = _0126_ & _0962_;
assign _0432_ = _0127_ & mie_q_t0[1];
assign _0434_ = _0128_ & _0968_;
assign _0436_ = _0129_ & _0970_;
assign _0438_ = _0130_ & _0972_;
assign _0440_ = _0171_ & _0974_;
assign _0442_ = _0145_ & _0976_;
assign _0444_ = _0146_ & dscratch0_q_t0[15:13];
assign _0446_ = _0135_ & dcsr_q_t0[15:13];
assign _0448_ = _0147_ & _0982_;
assign _0450_ = _0148_ & _0984_;
assign _0988_ = _0172_ & csr_mepc_o_t0[15:13];
assign _0452_ = _0139_ & _0988_;
assign _0454_ = _0173_ & mscratch_q_t0[15:13];
assign _0456_ = _0174_ & _0994_;
assign _0458_ = _0175_ & _0996_;
assign _0460_ = _0149_ & _0998_;
assign _0462_ = _0158_ & _0015_[16];
assign _1002_ = _0159_ & dscratch1_q_t0[16];
assign _0464_ = _0160_ & _1002_;
assign _0466_ = _0161_ & csr_depc_o_t0[16];
assign _0468_ = _0120_ & irq_fast_i_t0[0];
assign _0470_ = _0162_ & _1008_;
assign _0472_ = _0163_ & _1010_;
assign _0474_ = _0125_ & csr_mtvec_o_t0[16];
assign _0476_ = _0126_ & _1016_;
assign _0478_ = _0127_ & mie_q_t0[0];
assign _0480_ = _0129_ & _1022_;
assign _0482_ = _0130_ & _1024_;
assign _0484_ = _0171_ & _1026_;
assign _0486_ = _0176_ & _0015_[30:22];
assign _1030_ = _0177_ & dscratch1_q_t0[30:22];
assign _0488_ = _0178_ & _1030_;
assign _0490_ = _0179_ & csr_depc_o_t0[30:22];
assign _0492_ = _0180_ & irq_fast_i_t0[14:6];
assign _0494_ = _0181_ & _1036_;
assign _0496_ = _0182_ & _1038_;
assign _0498_ = _0183_ & csr_mtvec_o_t0[30:22];
assign _0500_ = _0184_ & _1044_;
assign _0502_ = _0185_ & mie_q_t0[14:6];
assign _1052_ = _0186_ & _1050_;
assign _0504_ = _0187_ & _1052_;
assign _0506_ = _0188_ & _1054_;
assign _0508_ = _0189_ & _1056_;
assign _0510_ = _0158_ & _0015_[11];
assign _1060_ = _0159_ & dscratch1_q_t0[11];
assign _0512_ = _0160_ & _1060_;
assign _0514_ = _0161_ & csr_depc_o_t0[11];
assign _0516_ = _0120_ & irq_external_i_t0;
assign _0518_ = _0162_ & _1066_;
assign _0520_ = _0163_ & _1068_;
assign _0522_ = _0125_ & csr_mtvec_o_t0[11];
assign _0524_ = _0126_ & _1074_;
assign _0526_ = _0127_ & mie_q_t0[15];
assign _0528_ = _0128_ & _1080_;
assign _0530_ = _0129_ & _1082_;
assign _0532_ = _0130_ & _1084_;
assign _0534_ = _0171_ & _1086_;
assign _0536_ = _0190_ & \mhpmcounter[0]_t0 ;
assign _0015_ = _0191_ & _1088_;
assign _0538_ = _0158_ & _0015_[21];
assign _1092_ = _0159_ & dscratch1_q_t0[21];
assign _0540_ = _0160_ & _1092_;
assign _0542_ = _0161_ & csr_depc_o_t0[21];
assign _0544_ = _0120_ & irq_fast_i_t0[5];
assign _0546_ = _0162_ & _1098_;
assign _0548_ = _0163_ & _1100_;
assign _0550_ = _0125_ & csr_mtvec_o_t0[21];
assign _0552_ = _0126_ & _1106_;
assign _0554_ = _0127_ & mie_q_t0[5];
assign _0556_ = _0128_ & _1112_;
assign _0558_ = _0129_ & _1114_;
assign _0560_ = _0130_ & _1116_;
assign _0562_ = _0171_ & _1118_;
assign _0564_ = _0192_ & _1246_;
assign _0566_ = _0193_ & _1120_;
assign _0568_ = _0158_ & _1122_;
assign _0570_ = _0119_ & dscratch0_q_t0[31];
assign _0572_ = _0121_ & dcsr_q_t0[31];
assign _0574_ = _0122_ & _1128_;
assign _0576_ = _0194_ & _1130_;
assign _0578_ = _0164_ & csr_mepc_o_t0[31];
assign _0580_ = _0124_ & _1134_;
assign _0582_ = _0165_ & mscratch_q_t0[31];
assign _0584_ = _0195_ & _1140_;
assign _0586_ = _0196_ & _1142_;
assign _0588_ = _0197_ & _1144_;
assign _0590_ = _0117_ & _0015_[39];
assign _0592_ = _0118_ & _1148_;
assign _0594_ = _0119_ & dscratch0_q_t0[7];
assign _0596_ = _0120_ & irq_timer_i_t0;
assign _0598_ = _0121_ & _1154_;
assign _0600_ = _0122_ & _1156_;
assign _0602_ = _0123_ & _1158_;
assign _0604_ = _0125_ & csr_mtvec_o_t0[7];
assign _0606_ = _0126_ & _1164_;
assign _0608_ = _0127_ & mie_q_t0[16];
assign _0610_ = _0128_ & _1170_;
assign _0612_ = _0129_ & _1172_;
assign _0614_ = _0130_ & _1174_;
assign _0616_ = _0131_ & _1176_;
assign _0618_ = _0132_ & _0015_[38:36];
assign _0620_ = _0133_ & _1180_;
assign _0622_ = _0146_ & dscratch0_q_t0[6:4];
assign _0624_ = _0135_ & dcsr_q_t0[6:4];
assign _0626_ = _0147_ & _1186_;
assign _0628_ = _0138_ & _1188_;
assign _0630_ = _0139_ & { 2'h0, mcause_q_t0[4] };
assign _0632_ = _0140_ & csr_mtvec_o_t0[6:4];
assign _0634_ = _0141_ & _1194_;
assign _0636_ = _0142_ & hart_id_i_t0[6:4];
assign _0651_ = _0198_ & _0001_[7];
assign _0653_ = _0199_ & { dummy_instr_seed_o_t0[31:1], 1'h0 };
assign _0103_ = _0200_ & _0011_[1];
assign _0655_ = _0201_ & _0011_[4:2];
assign _0657_ = _0202_ & _1252_;
assign _0659_ = _0203_ & _1254_;
assign _0661_ = _0204_ & _0011_[1];
assign _0663_ = _0205_ & _1256_;
assign _0665_ = _0198_ & _1258_;
assign _0667_ = _0204_ & _0011_[5];
assign _0669_ = _0205_ & _1260_;
assign _0671_ = _0198_ & _1262_;
assign _0099_ = _0206_ & _0001_[7];
assign _0673_ = _0209_ & _0090_;
assign _0675_ = _0210_ & csr_mcause_i_t0;
assign _0677_ = _0211_ & _0030_;
assign _0679_ = _0207_ & _0099_;
assign _0681_ = _0209_ & priv_mode_id_o_t0;
assign _0683_ = _0208_ & mstatus_q_t0[5];
assign _0685_ = _0211_ & csr_mtval_i_t0;
assign _0687_ = _0212_ & { dummy_instr_seed_o_t0[31:1], 1'h0 };
assign _0689_ = _0213_ & _0004_[8:6];
assign _0691_ = _0214_ & _0004_[1:0];
assign _0693_ = _0214_ & _0080_;
assign _0695_ = _0212_ & _0064_;
assign _0697_ = _0215_ & _0057_;
assign _0699_ = _0212_ & _0059_;
assign _0701_ = _0216_ & _0097_;
assign _0703_ = _0217_ & pc_id_i_t0;
assign _0705_ = _0218_ & _1264_;
assign _0707_ = _0219_ & _1266_;
assign _1270_ = _0204_ & _0001_[6];
assign _0709_ = _0205_ & _1270_;
assign _0711_ = _0198_ & _1272_;
assign _0713_ = _0220_ & { dummy_instr_seed_o_t0[31:1], 1'h0 };
assign _0715_ = _0203_ & _0004_[8:6];
assign _0717_ = _0221_ & _0004_[1:0];
assign _0719_ = _0220_ & dummy_instr_seed_o_t0;
assign _0721_ = _0222_ & { 2'h0, dummy_instr_seed_o_t0[4:0] };
assign _0723_ = _0223_ & _1276_;
assign _0725_ = _0224_ & _1278_;
assign _0727_ = _0225_ & { dummy_instr_seed_o_t0[31:1], 1'h0 };
assign _0729_ = _0226_ & _1282_;
assign _0731_ = _0220_ & _1284_;
assign _0733_ = _0227_ & { 2'h0, dummy_instr_seed_o_t0[4:0] };
assign _0735_ = _0228_ & _1288_;
assign priv_lvl_d_t0 = _0221_ & _1290_;
assign _0021_[31:28] = _0229_ & dcsr_q_t0[31:28];
assign _0737_ = _0230_ & mstatus_q_t0[5:4];
assign _0739_ = _0230_ & mstatus_q_t0[3:2];
assign _0741_ = _0120_ & dcsr_q_t0[15];
assign _0021_[14] = _0120_ & dcsr_q_t0[14];
assign _0021_[27:16] = _0231_ & dcsr_q_t0[27:16];
assign _0743_ = _0230_ & mstatus_q_t0[1:0];
assign _0745_ = _0232_ & dcsr_q_t0[1:0];
assign _0021_[5] = _0120_ & dcsr_q_t0[5];
assign _0021_[4] = _0120_ & dcsr_q_t0[4];
assign _0021_[3] = _0120_ & dcsr_q_t0[3];
assign _0747_ = _0120_ & dcsr_q_t0[2];
assign _0749_ = _0232_ & dcsr_q_t0[13:12];
assign _0021_[11] = _0120_ & dcsr_q_t0[11];
assign _0054_ = _0233_ & dummy_instr_seed_o_t0[1:0];
assign _0021_[9] = _0120_ & dcsr_q_t0[9];
assign _0062_ = _0234_ & dummy_instr_seed_o_t0[12:11];
assign _0751_ = _0235_ & cpuctrlsts_part_q_t0;
assign _0021_[10] = _0120_ & dcsr_q_t0[10];
assign _0052_ = _0165_ & csr_mtvec_init_i_t0;
assign _0753_ = _0237_ & cpuctrlsts_part_q_t0;
assign _0755_ = _0238_ & dcsr_q_t0;
assign _0757_ = _0236_ & csr_mtvec_init_i_t0;
assign _0759_ = _0239_ & mstatus_q_t0;
assign _0761_ = _0240_ & { dummy_instr_seed_o_t0[31:8], 8'h00 };
assign _0763_ = _0241_ & priv_mode_id_o_t0;
assign _0765_ = _0242_ & minstret_raw_t0;
assign _0795_ = { _0767_, _0767_, _0767_ } & _0792_;
assign _0291_ = { _0253_, _0253_, _0253_ } & _1196_;
assign _0293_ = { _0254_, _0254_, _0254_ } & _1190_;
assign _0295_ = _1297_ & cpuctrlsts_part_q_t0[3];
assign _0801_ = _1296_ & _0015_[3];
assign _0297_ = _0768_ & _0799_;
assign _0299_ = _1299_ & dscratch1_q_t0[3];
assign _0301_ = _1291_ & dcsr_q_t0[3];
assign _0303_ = _1301_ & csr_depc_o_t0[3];
assign _0305_ = _0769_ & _0805_;
assign _0307_ = _0255_ & _0803_;
assign _0309_ = _1303_ & csr_mtval_o_t0[3];
assign _0311_ = _1305_ & csr_mepc_o_t0[3];
assign _0313_ = _0770_ & _0815_;
assign _0315_ = _1306_ & mscratch_q_t0[3];
assign _0823_ = _1311_ & hart_id_i_t0[3];
assign _0317_ = _1292_ & mstatus_q_t0[5];
assign _0319_ = _0771_ & _0821_;
assign _0321_ = _0253_ & _0819_;
assign _0323_ = _0256_ & _0813_;
assign _0325_ = { _1297_, _1297_, _1297_ } & cpuctrlsts_part_q_t0[2:0];
assign _0833_ = { _1296_, _1296_, _1296_ } & _0015_[2:0];
assign _0327_ = { _0768_, _0768_, _0768_ } & _0831_;
assign _0329_ = { _1298_, _1298_, _1298_ } & { mcountinhibit_t0[2], 1'h0, mcountinhibit_t0[0] };
assign _0331_ = { _1301_, _1301_, _1301_ } & csr_depc_o_t0[2:0];
assign _0333_ = { _1300_, _1300_, _1300_ } & dscratch0_q_t0[2:0];
assign _0335_ = { _0772_, _0772_, _0772_ } & _0837_;
assign _0337_ = { _0255_, _0255_, _0255_ } & _0835_;
assign _0339_ = { _1303_, _1303_, _1303_ } & csr_mtval_o_t0[2:0];
assign _0341_ = { _1305_, _1305_, _1305_ } & csr_mepc_o_t0[2:0];
assign _0343_ = { _0770_, _0770_, _0770_ } & _0847_;
assign _0853_ = { _1306_, _1306_, _1306_ } & mscratch_q_t0[2:0];
assign _0856_ = { _1311_, _1311_, _1311_ } & hart_id_i_t0[2:0];
assign _0345_ = { _0773_, _0773_, _0773_ } & _0853_;
assign _0347_ = { _0253_, _0253_, _0253_ } & _0851_;
assign _0349_ = { _0257_, _0257_, _0257_ } & _0845_;
assign _0862_ = { _1296_, _1296_, _1296_ } & _0015_[10:8];
assign _0351_ = { _1294_, _1294_, _1294_ } & _0015_[42:40];
assign _0353_ = { _1299_, _1299_, _1299_ } & dscratch1_q_t0[10:8];
assign _0355_ = { _1301_, _1301_, _1301_ } & csr_depc_o_t0[10:8];
assign _0357_ = { _0769_, _0769_, _0769_ } & _0866_;
assign _0359_ = { _0258_, _0258_, _0258_ } & _0864_;
assign _0874_ = { _1303_, _1303_, _1303_ } & csr_mtval_o_t0[10:8];
assign _0361_ = { _1305_, _1305_, _1305_ } & csr_mepc_o_t0[10:8];
assign _0363_ = { _0770_, _0770_, _0770_ } & _0874_;
assign _0880_ = { _1306_, _1306_, _1306_ } & mscratch_q_t0[10:8];
assign _0882_ = { _1311_, _1311_, _1311_ } & hart_id_i_t0[10:8];
assign _0365_ = { _0773_, _0773_, _0773_ } & _0880_;
assign _0367_ = { _0253_, _0253_, _0253_ } & _0878_;
assign _0369_ = { _0259_, _0259_, _0259_ } & _0872_;
assign _0371_ = { _1294_, _1294_, _1294_ } & _0015_[52:50];
assign _0373_ = { _0774_, _0774_, _0774_ } & _0888_;
assign _0375_ = { _1300_, _1300_, _1300_ } & dscratch0_q_t0[20:18];
assign _0377_ = { _1291_, _1291_, _1291_ } & dcsr_q_t0[20:18];
assign _0379_ = { _0775_, _0775_, _0775_ } & _0894_;
assign _0381_ = { _0260_, _0260_, _0260_ } & _0892_;
assign _0902_ = { _1303_, _1303_, _1303_ } & csr_mtval_o_t0[20:18];
assign _0383_ = { _1305_, _1305_, _1305_ } & csr_mepc_o_t0[20:18];
assign _0385_ = { _0770_, _0770_, _0770_ } & _0902_;
assign _0387_ = { _1306_, _1306_, _1306_ } & mscratch_q_t0[20:18];
assign _0910_ = { _1311_, _1311_, _1311_ } & hart_id_i_t0[20:18];
assign _0389_ = { _0771_, _0771_, _0771_ } & _0908_;
assign _0391_ = { _0253_, _0253_, _0253_ } & _0906_;
assign _0393_ = { _0261_, _0261_, _0261_ } & _0900_;
assign _0395_ = _1294_ & _0015_[44];
assign _0397_ = _0774_ & _0918_;
assign _0399_ = _1300_ & dscratch0_q_t0[12];
assign _0401_ = _1291_ & dcsr_q_t0[12];
assign _0403_ = _0775_ & _0924_;
assign _0405_ = _0260_ & _0922_;
assign _0407_ = _1302_ & csr_mtvec_o_t0[12];
assign _0409_ = _0776_ & _0932_;
assign _0940_ = _1311_ & hart_id_i_t0[12];
assign _0411_ = _0777_ & _0938_;
assign _0413_ = _0262_ & _0936_;
assign _0415_ = _0263_ & _0930_;
assign _0417_ = _1294_ & _0015_[49];
assign _0419_ = _0774_ & _0946_;
assign _0421_ = _1300_ & dscratch0_q_t0[17];
assign _0423_ = _1291_ & dcsr_q_t0[17];
assign _0425_ = _0775_ & _0952_;
assign _0427_ = _0260_ & _0950_;
assign _0960_ = _1303_ & csr_mtval_o_t0[17];
assign _0429_ = _1305_ & csr_mepc_o_t0[17];
assign _0431_ = _0770_ & _0960_;
assign _0433_ = _1306_ & mscratch_q_t0[17];
assign _0968_ = _1311_ & hart_id_i_t0[17];
assign _0435_ = _1292_ & mstatus_q_t0[1];
assign _0437_ = _0771_ & _0966_;
assign _0439_ = _0253_ & _0964_;
assign _0441_ = _0261_ & _0958_;
assign _0976_ = { _1296_, _1296_, _1296_ } & _0015_[15:13];
assign _0443_ = { _1294_, _1294_, _1294_ } & _0015_[47:45];
assign _0445_ = { _1299_, _1299_, _1299_ } & dscratch1_q_t0[15:13];
assign _0447_ = { _1301_, _1301_, _1301_ } & csr_depc_o_t0[15:13];
assign _0449_ = { _0769_, _0769_, _0769_ } & _0980_;
assign _0451_ = { _0258_, _0258_, _0258_ } & _0978_;
assign _0453_ = { _1303_, _1303_, _1303_ } & csr_mtval_o_t0[15:13];
assign _0455_ = { _1302_, _1302_, _1302_ } & csr_mtvec_o_t0[15:13];
assign _0994_ = { _1311_, _1311_, _1311_ } & hart_id_i_t0[15:13];
assign _0457_ = { _0778_, _0778_, _0778_ } & _0992_;
assign _0459_ = { _0264_, _0264_, _0264_ } & _0990_;
assign _0461_ = { _0259_, _0259_, _0259_ } & _0986_;
assign _0463_ = _1294_ & _0015_[48];
assign _0465_ = _0774_ & _1000_;
assign _0467_ = _1300_ & dscratch0_q_t0[16];
assign _0469_ = _1291_ & dcsr_q_t0[16];
assign _0471_ = _0775_ & _1006_;
assign _0473_ = _0260_ & _1004_;
assign _1014_ = _1303_ & csr_mtval_o_t0[16];
assign _0475_ = _1305_ & csr_mepc_o_t0[16];
assign _0477_ = _0770_ & _1014_;
assign _0479_ = _1306_ & mscratch_q_t0[16];
assign _1022_ = _1311_ & hart_id_i_t0[16];
assign _0481_ = _0771_ & _1020_;
assign _0483_ = _0253_ & _1018_;
assign _0485_ = _0261_ & _1012_;
assign _0487_ = { _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_ } & _0015_[62:54];
assign _0489_ = { _0774_, _0774_, _0774_, _0774_, _0774_, _0774_, _0774_, _0774_, _0774_ } & _1028_;
assign _0491_ = { _1300_, _1300_, _1300_, _1300_, _1300_, _1300_, _1300_, _1300_, _1300_ } & dscratch0_q_t0[30:22];
assign _0493_ = { _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_ } & dcsr_q_t0[30:22];
assign _0495_ = { _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_ } & _1034_;
assign _0497_ = { _0260_, _0260_, _0260_, _0260_, _0260_, _0260_, _0260_, _0260_, _0260_ } & _1032_;
assign _1042_ = { _1303_, _1303_, _1303_, _1303_, _1303_, _1303_, _1303_, _1303_, _1303_ } & csr_mtval_o_t0[30:22];
assign _0499_ = { _1305_, _1305_, _1305_, _1305_, _1305_, _1305_, _1305_, _1305_, _1305_ } & csr_mepc_o_t0[30:22];
assign _0501_ = { _0770_, _0770_, _0770_, _0770_, _0770_, _0770_, _0770_, _0770_, _0770_ } & _1042_;
assign _0503_ = { _1306_, _1306_, _1306_, _1306_, _1306_, _1306_, _1306_, _1306_, _1306_ } & mscratch_q_t0[30:22];
assign _1050_ = { _1311_, _1311_, _1311_, _1311_, _1311_, _1311_, _1311_, _1311_, _1311_ } & hart_id_i_t0[30:22];
assign _0505_ = { _0771_, _0771_, _0771_, _0771_, _0771_, _0771_, _0771_, _0771_, _0771_ } & _1048_;
assign _0507_ = { _0253_, _0253_, _0253_, _0253_, _0253_, _0253_, _0253_, _0253_, _0253_ } & _1046_;
assign _0509_ = { _0261_, _0261_, _0261_, _0261_, _0261_, _0261_, _0261_, _0261_, _0261_ } & _1040_;
assign _0511_ = _1294_ & _0015_[43];
assign _0513_ = _0774_ & _1058_;
assign _0515_ = _1300_ & dscratch0_q_t0[11];
assign _0517_ = _1291_ & dcsr_q_t0[11];
assign _0519_ = _0775_ & _1064_;
assign _0521_ = _0260_ & _1062_;
assign _1072_ = _1303_ & csr_mtval_o_t0[11];
assign _0523_ = _1305_ & csr_mepc_o_t0[11];
assign _0525_ = _0770_ & _1072_;
assign _0527_ = _1306_ & mscratch_q_t0[11];
assign _1080_ = _1311_ & hart_id_i_t0[11];
assign _0529_ = _1292_ & mstatus_q_t0[2];
assign _0531_ = _0771_ & _1078_;
assign _0533_ = _0253_ & _1076_;
assign _0535_ = _0261_ & _1070_;
assign _0537_ = { _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_ } & \mhpmcounter[2]_t0 ;
assign _0539_ = _1294_ & _0015_[53];
assign _0541_ = _0774_ & _1090_;
assign _0543_ = _1300_ & dscratch0_q_t0[21];
assign _0545_ = _1291_ & dcsr_q_t0[21];
assign _0547_ = _0775_ & _1096_;
assign _0549_ = _0260_ & _1094_;
assign _1104_ = _1303_ & csr_mtval_o_t0[21];
assign _0551_ = _1305_ & csr_mepc_o_t0[21];
assign _0553_ = _0770_ & _1104_;
assign _0555_ = _1306_ & mscratch_q_t0[21];
assign _1112_ = _1311_ & hart_id_i_t0[21];
assign _0557_ = _1292_ & mstatus_q_t0[0];
assign _0559_ = _0771_ & _1110_;
assign _0561_ = _0253_ & _1108_;
assign _0563_ = _0261_ & _1102_;
assign _0565_ = { _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_ } & _0107_;
assign _0567_ = { _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_ } & csr_wdata_i_t0;
assign _1122_ = _1296_ & _0015_[31];
assign _0569_ = _1294_ & _0015_[63];
assign _0571_ = _1299_ & dscratch1_q_t0[31];
assign _0573_ = _1301_ & csr_depc_o_t0[31];
assign _0575_ = _0769_ & _1126_;
assign _0577_ = _0258_ & _1124_;
assign _0579_ = _1304_ & _1244_;
assign _0581_ = _1303_ & csr_mtval_o_t0[31];
assign _0583_ = _1302_ & csr_mtvec_o_t0[31];
assign _1140_ = _1311_ & hart_id_i_t0[31];
assign _0585_ = _0778_ & _1138_;
assign _0587_ = _0264_ & _1136_;
assign _0589_ = _0259_ & _1132_;
assign _0591_ = _1297_ & cpuctrlsts_part_q_t0[7];
assign _1148_ = _1296_ & _0015_[7];
assign _0593_ = _0768_ & _1146_;
assign _0595_ = _1299_ & dscratch1_q_t0[7];
assign _0597_ = _1291_ & dcsr_q_t0[7];
assign _0599_ = _1301_ & csr_depc_o_t0[7];
assign _0601_ = _0769_ & _1152_;
assign _0603_ = _0255_ & _1150_;
assign _1162_ = _1303_ & csr_mtval_o_t0[7];
assign _0605_ = _1305_ & csr_mepc_o_t0[7];
assign _0607_ = _0770_ & _1162_;
assign _0609_ = _1306_ & mscratch_q_t0[7];
assign _1170_ = _1311_ & hart_id_i_t0[7];
assign _0611_ = _1292_ & mstatus_q_t0[4];
assign _0613_ = _0771_ & _1168_;
assign _0615_ = _0253_ & _1166_;
assign _0617_ = _0256_ & _1160_;
assign _0619_ = { _1297_, _1297_, _1297_ } & cpuctrlsts_part_q_t0[6:4];
assign _1180_ = { _1296_, _1296_, _1296_ } & _0015_[6:4];
assign _0621_ = { _0768_, _0768_, _0768_ } & _1178_;
assign _0623_ = { _1299_, _1299_, _1299_ } & dscratch1_q_t0[6:4];
assign _0625_ = { _1301_, _1301_, _1301_ } & csr_depc_o_t0[6:4];
assign _0627_ = { _0769_, _0769_, _0769_ } & _1184_;
assign _0629_ = { _0255_, _0255_, _0255_ } & _1182_;
assign _0631_ = { _1303_, _1303_, _1303_ } & csr_mtval_o_t0[6:4];
assign _0633_ = { _1305_, _1305_, _1305_ } & csr_mepc_o_t0[6:4];
assign _0635_ = { _0770_, _0770_, _0770_ } & _1192_;
assign _0637_ = { _1306_, _1306_, _1306_ } & mscratch_q_t0[6:4];
assign _0652_ = csr_save_cause_i & _0066_[1];
assign _0654_ = { nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i } & mstack_epc_q_t0;
assign _0105_[1:0] = { nmi_mode_i, nmi_mode_i } & mstack_q_t0[1:0];
assign _0105_[2] = nmi_mode_i & mstack_q_t0[2];
assign _0656_ = { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i } & _0105_;
assign _0658_ = { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i } & _0011_[4:2];
assign _0660_ = { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i } & _0086_[2:0];
assign _0662_ = csr_restore_mret_i & _0103_;
assign _0664_ = csr_restore_dret_i & _0011_[1];
assign _0666_ = csr_save_cause_i & _0011_[1];
assign _0668_ = csr_restore_mret_i & mstatus_q_t0[4];
assign _0670_ = csr_restore_dret_i & _0011_[5];
assign _0672_ = csr_save_cause_i & _0086_[3];
assign _0090_[0] = _1226_ & _0001_[6];
assign _0674_ = { debug_mode_i, debug_mode_i } & _0001_[7:6];
assign _0676_ = { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i } & { 2'h0, dummy_instr_seed_o_t0[4:0] };
assign _0678_ = { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i } & { dummy_instr_seed_o_t0[31:1], 1'h0 };
assign _0680_ = _1226_ & _0001_[7];
assign _0682_ = { debug_mode_i, debug_mode_i } & _0011_[3:2];
assign _0684_ = debug_mode_i & _0011_[4];
assign _0686_ = { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i } & dummy_instr_seed_o_t0;
assign _0688_ = { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i } & _0030_;
assign _0690_ = { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i } & debug_cause_i_t0;
assign _0692_ = { debug_csr_save_i, debug_csr_save_i } & priv_mode_id_o_t0;
assign _0694_ = { debug_csr_save_i, debug_csr_save_i } & _0001_[7:6];
assign _0696_ = { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i } & dummy_instr_seed_o_t0;
assign _0698_ = { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i } & { 2'h0, dummy_instr_seed_o_t0[4:0] };
assign _0700_ = { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i } & { dummy_instr_seed_o_t0[31:1], 1'h0 };
assign _0702_ = { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i } & _0011_[5:2];
assign _0704_ = { csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i } & pc_wb_i_t0;
assign _0706_ = { csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i } & pc_id_i_t0;
assign _0708_ = { csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i } & pc_if_i_t0;
assign _0710_ = csr_restore_dret_i & _0001_[6];
assign _0712_ = csr_save_cause_i & _0066_[0];
assign _0714_ = { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i } & _0024_;
assign _0716_ = { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i } & _0101_;
assign _0718_ = { csr_save_cause_i, csr_save_cause_i } & _0093_;
assign _0720_ = { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i } & _0049_;
assign _0722_ = { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i } & _0072_;
assign _0724_ = { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i } & { 2'h0, dummy_instr_seed_o_t0[4:0] };
assign _0726_ = { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i } & _0032_;
assign _0728_ = { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i } & _0075_;
assign _0730_ = { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i } & { dummy_instr_seed_o_t0[31:1], 1'h0 };
assign _0732_ = { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i } & _0036_;
assign _0734_ = { nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i } & mstack_cause_q_t0;
assign _1288_ = { csr_restore_mret_i, csr_restore_mret_i } & mstatus_q_t0[3:2];
assign _0736_ = { csr_restore_dret_i, csr_restore_dret_i } & dcsr_q_t0[1:0];
assign _0097_[3] = debug_mode_i & _0011_[5];
assign _0738_ = { _1292_, _1292_ } & { dummy_instr_seed_o_t0[3], dummy_instr_seed_o_t0[7] };
assign _0740_ = { _1292_, _1292_ } & _0062_;
assign _0742_ = _1291_ & dummy_instr_seed_o_t0[15];
assign _0744_ = { _1292_, _1292_ } & { dummy_instr_seed_o_t0[17], dummy_instr_seed_o_t0[21] };
assign _0746_ = { _1291_, _1291_ } & _0054_;
assign _0748_ = _1291_ & dummy_instr_seed_o_t0[2];
assign _0750_ = { _1291_, _1291_ } & dummy_instr_seed_o_t0[13:12];
assign _0752_ = { _1297_, _1297_, _1297_, _1297_, _1297_, _1297_, _1297_, _1297_ } & { dummy_instr_seed_o_t0[7:1], 1'h0 };
assign _0041_ = { _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_ } & _1238_;
assign _0039_ = { _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_ } & _1238_;
assign _0754_ = { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int } & _0018_;
assign mhpmcounterh_we_t0 = { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int } & _0041_;
assign mhpmcounter_we_t0 = { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int } & _0039_;
assign _0756_ = { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int } & { _0021_[31:9], dcsr_q_t0[8:6], _0021_[5:0] };
assign _0758_ = csr_we_int & _0052_;
assign _0760_ = { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int } & _0046_;
assign _0762_ = { csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i } & { boot_addr_i_t0[31:8], 8'h00 };
assign _0764_ = { mstatus_q[1], mstatus_q[1] } & mstatus_q_t0[3:2];
assign _0766_ = { _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_ } & minstret_next_t0;
assign _0797_ = _0290_ | _0291_;
assign csr_rdata_o_t0[6:4] = _0292_ | _0293_;
assign _0799_ = _0294_ | _0295_;
assign _0803_ = _0296_ | _0297_;
assign _0805_ = _0298_ | _0299_;
assign _0807_ = _0300_ | _0301_;
assign _0809_ = _0302_ | _0303_;
assign _0811_ = _0304_ | _0305_;
assign _0813_ = _0306_ | _0307_;
assign _0815_ = _0308_ | _0309_;
assign _0817_ = _0310_ | _0311_;
assign _0819_ = _0312_ | _0313_;
assign _0821_ = _0314_ | _0315_;
assign _0825_ = _0316_ | _0317_;
assign _0827_ = _0318_ | _0319_;
assign _0829_ = _0320_ | _0321_;
assign csr_rdata_o_t0[3] = _0322_ | _0323_;
assign _0831_ = _0324_ | _0325_;
assign _0835_ = _0326_ | _0327_;
assign _0837_ = _0328_ | _0329_;
assign _0839_ = _0330_ | _0331_;
assign _0841_ = _0332_ | _0333_;
assign _0843_ = _0334_ | _0335_;
assign _0845_ = _0336_ | _0337_;
assign _0847_ = _0338_ | _0339_;
assign _0849_ = _0340_ | _0341_;
assign _0851_ = _0342_ | _0343_;
assign _0858_ = _0344_ | _0345_;
assign _0860_ = _0346_ | _0347_;
assign csr_rdata_o_t0[2:0] = _0348_ | _0349_;
assign _0864_ = _0350_ | _0351_;
assign _0866_ = _0352_ | _0353_;
assign _0868_ = _0354_ | _0355_;
assign _0870_ = _0356_ | _0357_;
assign _0872_ = _0358_ | _0359_;
assign _0876_ = _0360_ | _0361_;
assign _0878_ = _0362_ | _0363_;
assign _0884_ = _0364_ | _0365_;
assign _0886_ = _0366_ | _0367_;
assign csr_rdata_o_t0[10:8] = _0368_ | _0369_;
assign _0888_ = _0370_ | _0371_;
assign _0892_ = _0372_ | _0373_;
assign _0894_ = _0374_ | _0375_;
assign _0896_ = _0376_ | _0377_;
assign _0898_ = _0378_ | _0379_;
assign _0900_ = _0380_ | _0381_;
assign _0904_ = _0382_ | _0383_;
assign _0906_ = _0384_ | _0385_;
assign _0908_ = _0386_ | _0387_;
assign _0914_ = _0388_ | _0389_;
assign _0916_ = _0390_ | _0391_;
assign csr_rdata_o_t0[20:18] = _0392_ | _0393_;
assign _0918_ = _0394_ | _0395_;
assign _0922_ = _0396_ | _0397_;
assign _0924_ = _0398_ | _0399_;
assign _0926_ = _0400_ | _0401_;
assign _0928_ = _0402_ | _0403_;
assign _0930_ = _0404_ | _0405_;
assign _0934_ = _0406_ | _0407_;
assign _0936_ = _0408_ | _0409_;
assign _0942_ = _0410_ | _0411_;
assign _0944_ = _0412_ | _0413_;
assign csr_rdata_o_t0[12] = _0414_ | _0415_;
assign _0946_ = _0416_ | _0417_;
assign _0950_ = _0418_ | _0419_;
assign _0952_ = _0420_ | _0421_;
assign _0954_ = _0422_ | _0423_;
assign _0956_ = _0424_ | _0425_;
assign _0958_ = _0426_ | _0427_;
assign _0962_ = _0428_ | _0429_;
assign _0964_ = _0430_ | _0431_;
assign _0966_ = _0432_ | _0433_;
assign _0970_ = _0434_ | _0435_;
assign _0972_ = _0436_ | _0437_;
assign _0974_ = _0438_ | _0439_;
assign csr_rdata_o_t0[17] = _0440_ | _0441_;
assign _0978_ = _0442_ | _0443_;
assign _0980_ = _0444_ | _0445_;
assign _0982_ = _0446_ | _0447_;
assign _0984_ = _0448_ | _0449_;
assign _0986_ = _0450_ | _0451_;
assign _0990_ = _0452_ | _0453_;
assign _0992_ = _0454_ | _0455_;
assign _0996_ = _0456_ | _0457_;
assign _0998_ = _0458_ | _0459_;
assign csr_rdata_o_t0[15:13] = _0460_ | _0461_;
assign _1000_ = _0462_ | _0463_;
assign _1004_ = _0464_ | _0465_;
assign _1006_ = _0466_ | _0467_;
assign _1008_ = _0468_ | _0469_;
assign _1010_ = _0470_ | _0471_;
assign _1012_ = _0472_ | _0473_;
assign _1016_ = _0474_ | _0475_;
assign _1018_ = _0476_ | _0477_;
assign _1020_ = _0478_ | _0479_;
assign _1024_ = _0480_ | _0481_;
assign _1026_ = _0482_ | _0483_;
assign csr_rdata_o_t0[16] = _0484_ | _0485_;
assign _1028_ = _0486_ | _0487_;
assign _1032_ = _0488_ | _0489_;
assign _1034_ = _0490_ | _0491_;
assign _1036_ = _0492_ | _0493_;
assign _1038_ = _0494_ | _0495_;
assign _1040_ = _0496_ | _0497_;
assign _1044_ = _0498_ | _0499_;
assign _1046_ = _0500_ | _0501_;
assign _1048_ = _0502_ | _0503_;
assign _1054_ = _0504_ | _0505_;
assign _1056_ = _0506_ | _0507_;
assign csr_rdata_o_t0[30:22] = _0508_ | _0509_;
assign _1058_ = _0510_ | _0511_;
assign _1062_ = _0512_ | _0513_;
assign _1064_ = _0514_ | _0515_;
assign _1066_ = _0516_ | _0517_;
assign _1068_ = _0518_ | _0519_;
assign _1070_ = _0520_ | _0521_;
assign _1074_ = _0522_ | _0523_;
assign _1076_ = _0524_ | _0525_;
assign _1078_ = _0526_ | _0527_;
assign _1082_ = _0528_ | _0529_;
assign _1084_ = _0530_ | _0531_;
assign _1086_ = _0532_ | _0533_;
assign csr_rdata_o_t0[11] = _0534_ | _0535_;
assign _1088_ = _0536_ | _0537_;
assign _1090_ = _0538_ | _0539_;
assign _1094_ = _0540_ | _0541_;
assign _1096_ = _0542_ | _0543_;
assign _1098_ = _0544_ | _0545_;
assign _1100_ = _0546_ | _0547_;
assign _1102_ = _0548_ | _0549_;
assign _1106_ = _0550_ | _0551_;
assign _1108_ = _0552_ | _0553_;
assign _1110_ = _0554_ | _0555_;
assign _1114_ = _0556_ | _0557_;
assign _1116_ = _0558_ | _0559_;
assign _1118_ = _0560_ | _0561_;
assign csr_rdata_o_t0[21] = _0562_ | _0563_;
assign _1120_ = _0564_ | _0565_;
assign dummy_instr_seed_o_t0 = _0566_ | _0567_;
assign _1124_ = _0568_ | _0569_;
assign _1126_ = _0570_ | _0571_;
assign _1128_ = _0572_ | _0573_;
assign _1130_ = _0574_ | _0575_;
assign _1132_ = _0576_ | _0577_;
assign _1134_ = _0578_ | _0579_;
assign _1136_ = _0580_ | _0581_;
assign _1138_ = _0582_ | _0583_;
assign _1142_ = _0584_ | _0585_;
assign _1144_ = _0586_ | _0587_;
assign csr_rdata_o_t0[31] = _0588_ | _0589_;
assign _1146_ = _0590_ | _0591_;
assign _1150_ = _0592_ | _0593_;
assign _1152_ = _0594_ | _0595_;
assign _1154_ = _0596_ | _0597_;
assign _1156_ = _0598_ | _0599_;
assign _1158_ = _0600_ | _0601_;
assign _1160_ = _0602_ | _0603_;
assign _1164_ = _0604_ | _0605_;
assign _1166_ = _0606_ | _0607_;
assign _1168_ = _0608_ | _0609_;
assign _1172_ = _0610_ | _0611_;
assign _1174_ = _0612_ | _0613_;
assign _1176_ = _0614_ | _0615_;
assign csr_rdata_o_t0[7] = _0616_ | _0617_;
assign _1178_ = _0618_ | _0619_;
assign _1182_ = _0620_ | _0621_;
assign _1184_ = _0622_ | _0623_;
assign _1186_ = _0624_ | _0625_;
assign _1188_ = _0626_ | _0627_;
assign _1190_ = _0628_ | _0629_;
assign _1192_ = _0630_ | _0631_;
assign _1194_ = _0632_ | _0633_;
assign _1196_ = _0634_ | _0635_;
assign _0792_ = _0636_ | _0637_;
assign cpuctrlsts_part_d_t0[7] = _0651_ | _0652_;
assign _0075_ = _0653_ | _0654_;
assign _1252_ = _0655_ | _0656_;
assign _1254_ = _0657_ | _0658_;
assign mstatus_d_t0[4:2] = _0659_ | _0660_;
assign _1256_ = _0661_ | _0662_;
assign _1258_ = _0663_ | _0664_;
assign mstatus_d_t0[1] = _0665_ | _0666_;
assign _1260_ = _0667_ | _0668_;
assign _1262_ = _0669_ | _0670_;
assign mstatus_d_t0[5] = _0671_ | _0672_;
assign _0080_ = _0673_ | _0674_;
assign _0057_ = _0675_ | _0676_;
assign _0059_ = _0677_ | _0678_;
assign _0090_[1] = _0679_ | _0680_;
assign _0097_[1:0] = _0681_ | _0682_;
assign _0097_[2] = _0683_ | _0684_;
assign _0064_ = _0685_ | _0686_;
assign _0024_ = _0687_ | _0688_;
assign _0101_ = _0689_ | _0690_;
assign _0093_ = _0691_ | _0692_;
assign _0066_ = _0693_ | _0694_;
assign _0049_ = _0695_ | _0696_;
assign _0032_ = _0697_ | _0698_;
assign _0036_ = _0699_ | _0700_;
assign _0086_ = _0701_ | _0702_;
assign _1264_ = _0703_ | _0704_;
assign _1266_ = _0705_ | _0706_;
assign _0030_ = _0707_ | _0708_;
assign _1272_ = _0709_ | _0710_;
assign cpuctrlsts_part_d_t0[6] = _0711_ | _0712_;
assign depc_d_t0 = _0713_ | _0714_;
assign dcsr_d_t0[8:6] = _0715_ | _0716_;
assign dcsr_d_t0[1:0] = _0717_ | _0718_;
assign mtval_d_t0 = _0719_ | _0720_;
assign _1276_ = _0721_ | _0722_;
assign _1278_ = _0723_ | _0724_;
assign mcause_d_t0 = _0725_ | _0726_;
assign _1282_ = _0727_ | _0728_;
assign _1284_ = _0729_ | _0730_;
assign mepc_d_t0 = _0731_ | _0732_;
assign _0072_ = _0733_ | _0734_;
assign _1290_ = _0735_ | _0736_;
assign _0046_[5:4] = _0737_ | _0738_;
assign _0046_[3:2] = _0739_ | _0740_;
assign _0021_[15] = _0741_ | _0742_;
assign _0046_[1:0] = _0743_ | _0744_;
assign _0021_[1:0] = _0745_ | _0746_;
assign _0021_[2] = _0747_ | _0748_;
assign _0021_[13:12] = _0749_ | _0750_;
assign _0018_ = _0751_ | _0752_;
assign { _0001_[7:6], cpuctrlsts_part_d_t0[5:0] } = _0753_ | _0754_;
assign { dcsr_d_t0[31:9], _0004_[8:6], dcsr_d_t0[5:2], _0004_[1:0] } = _0755_ | _0756_;
assign mtvec_en_t0 = _0757_ | _0758_;
assign { _0011_[5:1], mstatus_d_t0[0] } = _0759_ | _0760_;
assign mtvec_d_t0 = _0761_ | _0762_;
assign priv_mode_lsu_o_t0 = _0763_ | _0764_;
assign \mhpmcounter[2]_t0  = _0765_ | _0766_;
assign _0265_ = | { csr_save_cause_i, csr_restore_dret_i, csr_restore_mret_i };
assign _0266_ = | { _1352_, _1351_, _1350_, _1349_, _1348_, _1347_, _1346_, _1313_, _1312_, _1311_, _1309_, _1307_, _1306_, _1305_, _1304_, _1303_, _1302_, _1301_, _1300_, _1299_, _1298_, _1297_, _1295_, _1293_, _1292_, _1291_, _1223_, _1217_, _1216_, _1215_, _1214_, _1213_, _1212_, _1211_, _1210_, _1209_, _1208_, _1207_, _1206_, _1205_, _1204_, _1203_, _1202_, _1201_, _1200_, _1199_, _1198_ };
assign _0267_ = | { _1345_, _1344_, _1343_, _1342_, _1341_, _1340_, _1339_, _1338_, _1337_, _1336_, _1335_, _1334_, _1333_, _1332_, _1331_, _1330_, _1329_, _1328_, _1327_, _1326_, _1325_, _1324_, _1323_, _1322_, _1321_, _1320_, _1319_, _1318_, _1317_, _1316_, _1315_, _1314_ };
assign _0268_ = | { _1301_, _1300_, _1299_, _1291_ };
assign _0269_ = | { _1222_, _1250_ };
assign _0270_ = | { _1344_, _1342_, _1341_, _1340_, _1339_, _1338_, _1337_, _1336_, _1335_, _1334_, _1333_, _1332_, _1331_, _1330_, _1329_, _1328_, _1327_, _1326_, _1325_, _1324_, _1323_, _1322_, _1321_, _1320_, _1319_, _1318_, _1317_, _1316_, _1315_, _1314_ };
assign _0167_ = ~ _1346_;
assign _0243_ = ~ _1240_;
assign _0244_ = ~ mcause_q[5];
assign _0245_ = ~ csr_wdata_i;
assign _0246_ = ~ mstatus_err;
assign _0247_ = ~ _1248_;
assign _0248_ = ~ mcause_q[6];
assign _0249_ = ~ csr_rdata_o;
assign _0250_ = ~ debug_mode_entering_i;
assign _0251_ = ~ mtvec_err;
assign _0252_ = ~ cpuctrlsts_part_err;
assign _0638_ = mcause_q_t0[5] & _0248_;
assign _0641_ = csr_wdata_i_t0 & _0249_;
assign _0642_ = debug_mode_i_t0 & _0250_;
assign _0645_ = mstatus_err_t0 & _0251_;
assign _0648_ = _1249_ & _0252_;
assign _1242_ = illegal_csr_dbg_t0 & _0243_;
assign _0639_ = mcause_q_t0[6] & _0244_;
assign _0275_ = csr_rdata_o_t0 & _0245_;
assign _0643_ = debug_mode_entering_i_t0 & _0208_;
assign _0646_ = mtvec_err_t0 & _0246_;
assign _0649_ = cpuctrlsts_part_err_t0 & _0247_;
assign _0640_ = mcause_q_t0[5] & mcause_q_t0[6];
assign _0644_ = debug_mode_i_t0 & debug_mode_entering_i_t0;
assign _0647_ = mstatus_err_t0 & mtvec_err_t0;
assign _0650_ = _1249_ & cpuctrlsts_part_err_t0;
assign _0786_ = _0638_ | _0639_;
assign _0787_ = _0641_ | _0275_;
assign _0788_ = _0642_ | _0643_;
assign _0789_ = _0645_ | _0646_;
assign _0790_ = _0648_ | _0649_;
assign _1244_ = _0786_ | _0640_;
assign _1246_ = _0787_ | _0276_;
assign _1236_ = _0788_ | _0644_;
assign _1249_ = _0789_ | _0647_;
assign csr_shadow_err_o_t0 = _0790_ | _0650_;
assign _0767_ = _1311_ | _1306_;
assign _0768_ = _1294_ | _1297_;
assign _0772_ = _1299_ | _1298_;
assign _0773_ = _1346_ | _1306_;
assign _0776_ = _1305_ | _1304_;
assign _0777_ = _1292_ | _1346_;
assign _0769_ = _1300_ | _1299_;
assign _0778_ = _1306_ | _1302_;
assign _0774_ = _1296_ | _1294_;
assign _0775_ = _1301_ | _1300_;
assign _0770_ = _1304_ | _1303_;
assign _0771_ = _1307_ | _1306_;
assign _0254_ = | { _0768_, _0769_, _1309_, _1301_, _1295_, _1291_ };
assign _0256_ = | { _0768_, _0769_, _1312_, _1309_, _1301_, _1295_, _1291_ };
assign _0255_ = | { _0768_, _1309_, _1295_ };
assign _0257_ = | { _0768_, _0772_, _1309_, _1301_, _1300_, _1295_, _1291_ };
assign _0262_ = | { _1306_, _1302_, _0776_ };
assign _0263_ = | { _0774_, _0775_, _1309_, _1303_, _1299_, _1291_ };
assign _0261_ = | { _0774_, _0775_, _1312_, _1309_, _1299_, _1291_ };
assign _0258_ = | { _1309_, _1295_, _1293_ };
assign _0264_ = | { _1305_, _1304_, _1303_ };
assign _0259_ = | { _0769_, _1309_, _1301_, _1295_, _1293_, _1291_ };
assign _0260_ = | { _0774_, _1309_, _1299_ };
assign _0253_ = | { _0770_, _1305_, _1302_ };
assign _0793_ = _1313_ ? 3'h1 : 3'h0;
assign _0794_ = _0767_ ? _0791_ : _0793_;
assign _0796_ = _0253_ ? _1195_ : _0794_;
assign csr_rdata_o[6:4] = _0254_ ? _1189_ : _0796_;
assign _0798_ = _1297_ ? cpuctrlsts_part_q[3] : _0014_[35];
assign _0800_ = _1296_ ? _0014_[3] : _0016_[3];
assign _0802_ = _0768_ ? _0798_ : _0800_;
assign _0804_ = _1299_ ? dscratch1_q[3] : dscratch0_q[3];
assign _0806_ = _1291_ ? dcsr_q[3] : irq_software_i;
assign _0808_ = _1301_ ? csr_depc_o[3] : _0806_;
assign _0810_ = _0769_ ? _0804_ : _0808_;
assign _0812_ = _0255_ ? _0802_ : _0810_;
assign _0814_ = _1303_ ? csr_mtval_o[3] : mcause_q[3];
assign _0816_ = _1305_ ? csr_mepc_o[3] : csr_mtvec_o[3];
assign _0818_ = _0770_ ? _0814_ : _0816_;
assign _0820_ = _1306_ ? mscratch_q[3] : mie_q[17];
assign _0822_ = _1311_ ? hart_id_i[3] : 1'h0;
assign _0824_ = _1292_ ? mstatus_q[5] : _0822_;
assign _0826_ = _0771_ ? _0820_ : _0824_;
assign _0828_ = _0253_ ? _0818_ : _0826_;
assign csr_rdata_o[3] = _0256_ ? _0812_ : _0828_;
assign _0830_ = _1297_ ? cpuctrlsts_part_q[2:0] : _0014_[34:32];
assign _0832_ = _1296_ ? _0014_[2:0] : _0016_[2:0];
assign _0834_ = _0768_ ? _0830_ : _0832_;
assign _0836_ = _1298_ ? { mcountinhibit[2], 1'h0, mcountinhibit[0] } : dscratch1_q[2:0];
assign _0838_ = _1301_ ? csr_depc_o[2:0] : dcsr_q[2:0];
assign _0840_ = _1300_ ? dscratch0_q[2:0] : _0838_;
assign _0842_ = _0772_ ? _0836_ : _0840_;
assign _0844_ = _0255_ ? _0834_ : _0842_;
assign _0846_ = _1303_ ? csr_mtval_o[2:0] : mcause_q[2:0];
assign _0848_ = _1305_ ? csr_mepc_o[2:0] : csr_mtvec_o[2:0];
assign _0850_ = _0770_ ? _0846_ : _0848_;
assign _0852_ = _1306_ ? mscratch_q[2:0] : 3'h4;
assign _0854_ = _1313_ ? 3'h6 : 3'h0;
assign _0855_ = _1311_ ? hart_id_i[2:0] : _0854_;
assign _0857_ = _0773_ ? _0852_ : _0855_;
assign _0859_ = _0253_ ? _0850_ : _0857_;
assign csr_rdata_o[2:0] = _0257_ ? _0844_ : _0859_;
assign _0861_ = _1296_ ? _0014_[10:8] : _0016_[10:8];
assign _0863_ = _1294_ ? _0014_[42:40] : _0861_;
assign _0865_ = _1299_ ? dscratch1_q[10:8] : dscratch0_q[10:8];
assign _0867_ = _1301_ ? csr_depc_o[10:8] : dcsr_q[10:8];
assign _0869_ = _0769_ ? _0865_ : _0867_;
assign _0871_ = _0258_ ? _0863_ : _0869_;
assign _0873_ = _1303_ ? csr_mtval_o[10:8] : _1353_[5:3];
assign _0875_ = _1305_ ? csr_mepc_o[10:8] : csr_mtvec_o[10:8];
assign _0877_ = _0770_ ? _0873_ : _0875_;
assign _0879_ = _1306_ ? mscratch_q[10:8] : 3'h1;
assign _0881_ = _1311_ ? hart_id_i[10:8] : 3'h0;
assign _0883_ = _0773_ ? _0879_ : _0881_;
assign _0885_ = _0253_ ? _0877_ : _0883_;
assign csr_rdata_o[10:8] = _0259_ ? _0871_ : _0885_;
assign _0887_ = _1294_ ? _0014_[52:50] : _0014_[20:18];
assign _0889_ = _1310_ ? _0016_[20:18] : dscratch1_q[20:18];
assign _0891_ = _0774_ ? _0887_ : _0889_;
assign _0893_ = _1300_ ? dscratch0_q[20:18] : csr_depc_o[20:18];
assign _0895_ = _1291_ ? dcsr_q[20:18] : irq_fast_i[4:2];
assign _0897_ = _0775_ ? _0893_ : _0895_;
assign _0899_ = _0260_ ? _0891_ : _0897_;
assign _0901_ = _1303_ ? csr_mtval_o[20:18] : _1353_[15:13];
assign _0903_ = _1305_ ? csr_mepc_o[20:18] : csr_mtvec_o[20:18];
assign _0905_ = _0770_ ? _0901_ : _0903_;
assign _0907_ = _1306_ ? mscratch_q[20:18] : mie_q[4:2];
assign _0909_ = _1311_ ? hart_id_i[20:18] : 3'h0;
assign _0911_ = _1346_ ? 3'h4 : _0909_;
assign _0913_ = _0771_ ? _0907_ : _0911_;
assign _0915_ = _0253_ ? _0905_ : _0913_;
assign csr_rdata_o[20:18] = _0261_ ? _0899_ : _0915_;
assign _0917_ = _1294_ ? _0014_[44] : _0014_[12];
assign _0919_ = _1310_ ? _0016_[12] : dscratch1_q[12];
assign _0921_ = _0774_ ? _0917_ : _0919_;
assign _0923_ = _1300_ ? dscratch0_q[12] : csr_depc_o[12];
assign _0925_ = _1291_ ? dcsr_q[12] : csr_mtval_o[12];
assign _0927_ = _0775_ ? _0923_ : _0925_;
assign _0929_ = _0260_ ? _0921_ : _0927_;
assign _0931_ = _1304_ ? _1353_[7] : csr_mepc_o[12];
assign _0933_ = _1302_ ? csr_mtvec_o[12] : mscratch_q[12];
assign _0935_ = _0776_ ? _0931_ : _0933_;
assign _0937_ = _1346_ ? 1'h1 : mstatus_q[3];
assign _0939_ = _1311_ ? hart_id_i[12] : 1'h0;
assign _0941_ = _0777_ ? _0937_ : _0939_;
assign _0943_ = _0262_ ? _0935_ : _0941_;
assign csr_rdata_o[12] = _0263_ ? _0929_ : _0943_;
assign _0945_ = _1294_ ? _0014_[49] : _0014_[17];
assign _0947_ = _1310_ ? _0016_[17] : dscratch1_q[17];
assign _0949_ = _0774_ ? _0945_ : _0947_;
assign _0951_ = _1300_ ? dscratch0_q[17] : csr_depc_o[17];
assign _0953_ = _1291_ ? dcsr_q[17] : irq_fast_i[1];
assign _0955_ = _0775_ ? _0951_ : _0953_;
assign _0957_ = _0260_ ? _0949_ : _0955_;
assign _0959_ = _1303_ ? csr_mtval_o[17] : _1353_[12];
assign _0961_ = _1305_ ? csr_mepc_o[17] : csr_mtvec_o[17];
assign _0963_ = _0770_ ? _0959_ : _0961_;
assign _0965_ = _1306_ ? mscratch_q[17] : mie_q[1];
assign _0967_ = _1311_ ? hart_id_i[17] : 1'h0;
assign _0969_ = _1292_ ? mstatus_q[1] : _0967_;
assign _0971_ = _0771_ ? _0965_ : _0969_;
assign _0973_ = _0253_ ? _0963_ : _0971_;
assign csr_rdata_o[17] = _0261_ ? _0957_ : _0973_;
assign _0975_ = _1296_ ? _0014_[15:13] : _0016_[15:13];
assign _0977_ = _1294_ ? _0014_[47:45] : _0975_;
assign _0979_ = _1299_ ? dscratch1_q[15:13] : dscratch0_q[15:13];
assign _0981_ = _1301_ ? csr_depc_o[15:13] : dcsr_q[15:13];
assign _0983_ = _0769_ ? _0979_ : _0981_;
assign _0985_ = _0258_ ? _0977_ : _0983_;
assign _0987_ = _1304_ ? _1353_[10:8] : csr_mepc_o[15:13];
assign _0989_ = _1303_ ? csr_mtval_o[15:13] : _0987_;
assign _0991_ = _1302_ ? csr_mtvec_o[15:13] : mscratch_q[15:13];
assign _0993_ = _1311_ ? hart_id_i[15:13] : 3'h0;
assign _0995_ = _0778_ ? _0991_ : _0993_;
assign _0997_ = _0264_ ? _0989_ : _0995_;
assign csr_rdata_o[15:13] = _0259_ ? _0985_ : _0997_;
assign _0999_ = _1294_ ? _0014_[48] : _0014_[16];
assign _1001_ = _1310_ ? _0016_[16] : dscratch1_q[16];
assign _1003_ = _0774_ ? _0999_ : _1001_;
assign _1005_ = _1300_ ? dscratch0_q[16] : csr_depc_o[16];
assign _1007_ = _1291_ ? dcsr_q[16] : irq_fast_i[0];
assign _1009_ = _0775_ ? _1005_ : _1007_;
assign _1011_ = _0260_ ? _1003_ : _1009_;
assign _1013_ = _1303_ ? csr_mtval_o[16] : _1353_[11];
assign _1015_ = _1305_ ? csr_mepc_o[16] : csr_mtvec_o[16];
assign _1017_ = _0770_ ? _1013_ : _1015_;
assign _1019_ = _1306_ ? mscratch_q[16] : mie_q[0];
assign _1021_ = _1311_ ? hart_id_i[16] : 1'h0;
assign _1023_ = _0771_ ? _1019_ : _1021_;
assign _1025_ = _0253_ ? _1017_ : _1023_;
assign csr_rdata_o[16] = _0261_ ? _1011_ : _1025_;
assign _1027_ = _1294_ ? _0014_[62:54] : _0014_[30:22];
assign _1029_ = _1310_ ? _0016_[30:22] : dscratch1_q[30:22];
assign _1031_ = _0774_ ? _1027_ : _1029_;
assign _1033_ = _1300_ ? dscratch0_q[30:22] : csr_depc_o[30:22];
assign _1035_ = _1291_ ? dcsr_q[30:22] : irq_fast_i[14:6];
assign _1037_ = _0775_ ? _1033_ : _1035_;
assign _1039_ = _0260_ ? _1031_ : _1037_;
assign _1041_ = _1303_ ? csr_mtval_o[30:22] : _1353_[25:17];
assign _1043_ = _1305_ ? csr_mepc_o[30:22] : csr_mtvec_o[30:22];
assign _1045_ = _0770_ ? _1041_ : _1043_;
assign _1047_ = _1306_ ? mscratch_q[30:22] : mie_q[14:6];
assign _1049_ = _1311_ ? hart_id_i[30:22] : 9'h000;
assign _1051_ = _1346_ ? 9'h100 : _1049_;
assign _1053_ = _0771_ ? _1047_ : _1051_;
assign _1055_ = _0253_ ? _1045_ : _1053_;
assign csr_rdata_o[30:22] = _0261_ ? _1039_ : _1055_;
assign _1057_ = _1294_ ? _0014_[43] : _0014_[11];
assign _1059_ = _1310_ ? _0016_[11] : dscratch1_q[11];
assign _1061_ = _0774_ ? _1057_ : _1059_;
assign _1063_ = _1300_ ? dscratch0_q[11] : csr_depc_o[11];
assign _1065_ = _1291_ ? dcsr_q[11] : irq_external_i;
assign _1067_ = _0775_ ? _1063_ : _1065_;
assign _1069_ = _0260_ ? _1061_ : _1067_;
assign _1071_ = _1303_ ? csr_mtval_o[11] : _1353_[6];
assign _1073_ = _1305_ ? csr_mepc_o[11] : csr_mtvec_o[11];
assign _1075_ = _0770_ ? _1071_ : _1073_;
assign _1077_ = _1306_ ? mscratch_q[11] : mie_q[15];
assign _1079_ = _1311_ ? hart_id_i[11] : 1'h0;
assign _1081_ = _1292_ ? mstatus_q[2] : _1079_;
assign _1083_ = _0771_ ? _1077_ : _1081_;
assign _1085_ = _0253_ ? _1075_ : _1083_;
assign csr_rdata_o[11] = _0261_ ? _1069_ : _1085_;
assign _1087_ = _1343_ ? \mhpmcounter[2]  : \mhpmcounter[0] ;
assign _0014_ = _0270_ ? 64'h0000000000000000 : _1087_;
assign _1089_ = _1294_ ? _0014_[53] : _0014_[21];
assign _1091_ = _1310_ ? _0016_[21] : dscratch1_q[21];
assign _1093_ = _0774_ ? _1089_ : _1091_;
assign _1095_ = _1300_ ? dscratch0_q[21] : csr_depc_o[21];
assign _1097_ = _1291_ ? dcsr_q[21] : irq_fast_i[5];
assign _1099_ = _0775_ ? _1095_ : _1097_;
assign _1101_ = _0260_ ? _1093_ : _1099_;
assign _1103_ = _1303_ ? csr_mtval_o[21] : _1353_[16];
assign _1105_ = _1305_ ? csr_mepc_o[21] : csr_mtvec_o[21];
assign _1107_ = _0770_ ? _1103_ : _1105_;
assign _1109_ = _1306_ ? mscratch_q[21] : mie_q[5];
assign _1111_ = _1311_ ? hart_id_i[21] : 1'h0;
assign _1113_ = _1292_ ? mstatus_q[0] : _1111_;
assign _1115_ = _0771_ ? _1109_ : _1113_;
assign _1117_ = _0253_ ? _1107_ : _1115_;
assign csr_rdata_o[21] = _0261_ ? _1101_ : _1117_;
assign _1119_ = _1220_ ? _0106_ : _1245_;
assign dummy_instr_seed_o = _0269_ ? csr_wdata_i : _1119_;
assign _1121_ = _1296_ ? _0014_[31] : _0016_[31];
assign _1123_ = _1294_ ? _0014_[63] : _1121_;
assign _1125_ = _1299_ ? dscratch1_q[31] : dscratch0_q[31];
assign _1127_ = _1301_ ? csr_depc_o[31] : dcsr_q[31];
assign _1129_ = _0769_ ? _1125_ : _1127_;
assign _1131_ = _0258_ ? _1123_ : _1129_;
assign _1133_ = _1304_ ? _1243_ : csr_mepc_o[31];
assign _1135_ = _1303_ ? csr_mtval_o[31] : _1133_;
assign _1137_ = _1302_ ? csr_mtvec_o[31] : mscratch_q[31];
assign _1139_ = _1311_ ? hart_id_i[31] : 1'h0;
assign _1141_ = _0778_ ? _1137_ : _1139_;
assign _1143_ = _0264_ ? _1135_ : _1141_;
assign csr_rdata_o[31] = _0259_ ? _1131_ : _1143_;
assign _1145_ = _1297_ ? cpuctrlsts_part_q[7] : _0014_[39];
assign _1147_ = _1296_ ? _0014_[7] : _0016_[7];
assign _1149_ = _0768_ ? _1145_ : _1147_;
assign _1151_ = _1299_ ? dscratch1_q[7] : dscratch0_q[7];
assign _1153_ = _1291_ ? dcsr_q[7] : irq_timer_i;
assign _1155_ = _1301_ ? csr_depc_o[7] : _1153_;
assign _1157_ = _0769_ ? _1151_ : _1155_;
assign _1159_ = _0255_ ? _1149_ : _1157_;
assign _1161_ = _1303_ ? csr_mtval_o[7] : _1353_[2];
assign _1163_ = _1305_ ? csr_mepc_o[7] : csr_mtvec_o[7];
assign _1165_ = _0770_ ? _1161_ : _1163_;
assign _1167_ = _1306_ ? mscratch_q[7] : mie_q[16];
assign _1169_ = _1311_ ? hart_id_i[7] : 1'h0;
assign _1171_ = _1292_ ? mstatus_q[4] : _1169_;
assign _1173_ = _0771_ ? _1167_ : _1171_;
assign _1175_ = _0253_ ? _1165_ : _1173_;
assign csr_rdata_o[7] = _0256_ ? _1159_ : _1175_;
assign _1177_ = _1297_ ? cpuctrlsts_part_q[6:4] : _0014_[38:36];
assign _1179_ = _1296_ ? _0014_[6:4] : _0016_[6:4];
assign _1181_ = _0768_ ? _1177_ : _1179_;
assign _1183_ = _1299_ ? dscratch1_q[6:4] : dscratch0_q[6:4];
assign _1185_ = _1301_ ? csr_depc_o[6:4] : dcsr_q[6:4];
assign _1187_ = _0769_ ? _1183_ : _1185_;
assign _1189_ = _0255_ ? _1181_ : _1187_;
assign _1191_ = _1303_ ? csr_mtval_o[6:4] : { _1353_[1:0], mcause_q[4] };
assign _1193_ = _1305_ ? csr_mepc_o[6:4] : csr_mtvec_o[6:4];
assign _1195_ = _0770_ ? _1191_ : _1193_;
assign _0791_ = _1306_ ? mscratch_q[6:4] : hart_id_i[6:4];
assign _1238_ = 1'h0 >> _1232_;
assign _1197_ = csr_addr_i[11:10] == /* src = "generated/sv2v_out.v:13958.30-13958.54" */ 2'h3;
assign _1218_ = dummy_instr_seed_o[31:30] == /* src = "generated/sv2v_out.v:14127.46-14127.75" */ 2'h2;
assign _1219_ = dummy_instr_seed_o[31:30] == /* src = "generated/sv2v_out.v:14127.15-14127.44" */ 2'h3;
assign illegal_csr_priv = csr_addr_i[9:8] > /* src = "generated/sv2v_out.v:13957.28-13957.56" */ priv_mode_id_o;
assign illegal_csr_write = _1197_ && /* src = "generated/sv2v_out.v:13958.29-13958.65" */ csr_wr;
assign _1224_ = _1227_ && /* src = "generated/sv2v_out.v:14154.10-14154.66" */ _1228_;
assign _1225_ = _1229_ && /* src = "generated/sv2v_out.v:14166.10-14166.60" */ _1230_;
assign dummy_instr_seed_en_o = csr_we_int && /* src = "generated/sv2v_out.v:14824.35-14824.70" */ _1223_;
assign _1226_ = csr_mcause_i[5] || /* src = "generated/sv2v_out.v:14221.12-14221.38" */ csr_mcause_i[6];
assign _1227_ = dummy_instr_seed_o[12:11] != /* src = "generated/sv2v_out.v:14154.11-14154.35" */ 2'h3;
assign _1228_ = | /* src = "generated/sv2v_out.v:14154.41-14154.65" */ dummy_instr_seed_o[12:11];
assign _1229_ = dummy_instr_seed_o[1:0] != /* src = "generated/sv2v_out.v:14166.11-14166.32" */ 2'h3;
assign _1230_ = | /* src = "generated/sv2v_out.v:14166.38-14166.59" */ dummy_instr_seed_o[1:0];
assign _1231_ = mstatus_q[3:2] != /* src = "generated/sv2v_out.v:14236.9-14236.33" */ 2'h3;
assign _1232_ = - /* src = "generated/sv2v_out.v:0.0-0.0" */ $signed({ 27'h0000000, csr_addr_i[4:0] });
assign _1233_ = ~ /* src = "generated/sv2v_out.v:14273.47-14273.66" */ illegal_csr_insn_o;
assign _0109_ = ~ /* src = "generated/sv2v_out.v:14645.40-14645.57" */ mcountinhibit[0];
assign _1234_ = ~ /* src = "generated/sv2v_out.v:14664.46-14664.63" */ mcountinhibit[2];
assign _1235_ = ~ /* src = "generated/sv2v_out.v:14868.50-14868.89" */ _1247_;
assign _1239_ = illegal_csr | /* src = "generated/sv2v_out.v:13959.48-13959.79" */ illegal_csr_write;
assign _1240_ = _1239_ | /* src = "generated/sv2v_out.v:13959.47-13959.99" */ illegal_csr_priv;
assign _1241_ = _1240_ | /* src = "generated/sv2v_out.v:13959.46-13959.118" */ illegal_csr_dbg;
assign _1243_ = mcause_q[5] | /* src = "generated/sv2v_out.v:14014.30-14014.55" */ mcause_q[6];
assign _1245_ = csr_wdata_i | /* src = "generated/sv2v_out.v:14267.26-14267.51" */ csr_rdata_o;
assign _1247_ = debug_mode_i | /* src = "generated/sv2v_out.v:14868.52-14868.88" */ debug_mode_entering_i;
assign _1248_ = mstatus_err | /* src = "generated/sv2v_out.v:14881.31-14881.54" */ mtvec_err;
assign csr_shadow_err_o = _1248_ | /* src = "generated/sv2v_out.v:14881.29-14881.92" */ cpuctrlsts_part_err;
assign _1250_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14265.3-14271.10" */ csr_op_i;
assign _1220_ = csr_op_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14265.3-14271.10" */ 2'h3;
assign _1221_ = csr_op_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14265.3-14271.10" */ 2'h2;
assign _1222_ = csr_op_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14265.3-14271.10" */ 2'h1;
assign cpuctrlsts_part_d[7] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0065_[1] : _0000_[7];
assign _0094_ = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14240.9-14240.19|generated/sv2v_out.v:14240.5-14251.8" */ 1'h1 : _0008_;
assign _0074_ = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14240.9-14240.19|generated/sv2v_out.v:14240.5-14251.8" */ mstack_epc_q : { dummy_instr_seed_o[31:1], 1'h0 };
assign _0095_ = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14240.9-14240.19|generated/sv2v_out.v:14240.5-14251.8" */ 1'h1 : _0009_;
assign _0104_[1:0] = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14240.9-14240.19|generated/sv2v_out.v:14240.5-14251.8" */ mstack_q[1:0] : 2'h0;
assign _0104_[2] = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14240.9-14240.19|generated/sv2v_out.v:14240.5-14251.8" */ mstack_q[2] : 1'h1;
assign _0102_ = _1231_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14236.9-14236.33|generated/sv2v_out.v:14236.5-14237.26" */ 1'h0 : _0010_[1];
assign _1251_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0104_ : _0010_[4:2];
assign _1253_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0010_[4:2] : _1251_;
assign mstatus_d[4:2] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0085_[2:0] : _1253_;
assign _1255_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0102_ : _0010_[1];
assign _1257_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0010_[1] : _1255_;
assign mstatus_d[1] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0010_[1] : _1257_;
assign _1259_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ mstatus_q[4] : _0010_[5];
assign _1261_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0010_[5] : _1259_;
assign mstatus_d[5] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0085_[3] : _1261_;
assign _0082_ = cpuctrlsts_part_q[6] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14224.11-14224.31|generated/sv2v_out.v:14224.7-14227.10" */ 1'h1 : 1'h0;
assign _0089_[0] = _1226_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14221.10-14221.39|generated/sv2v_out.v:14221.6-14228.9" */ _0000_[6] : 1'h1;
assign _0070_ = _1226_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14221.10-14221.39|generated/sv2v_out.v:14221.6-14228.9" */ 1'h0 : _0082_;
assign _0098_ = cpuctrlsts_part_q[6] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14224.11-14224.31|generated/sv2v_out.v:14224.7-14227.10" */ 1'h1 : _0000_[7];
assign _0091_ = _1226_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14221.10-14221.39|generated/sv2v_out.v:14221.6-14228.9" */ _0002_ : 1'h1;
assign _0081_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14209.14-14209.27|generated/sv2v_out.v:14209.10-14229.8" */ _0002_ : _0091_;
assign _0079_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14209.14-14209.27|generated/sv2v_out.v:14209.10-14229.8" */ _0000_[7:6] : _0089_;
assign _0055_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14209.14-14209.27|generated/sv2v_out.v:14209.10-14229.8" */ 1'h0 : _0070_;
assign _0060_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14209.14-14209.27|generated/sv2v_out.v:14209.10-14229.8" */ 1'h0 : 1'h1;
assign _0056_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14209.14-14209.27|generated/sv2v_out.v:14209.10-14229.8" */ { _1219_, _1218_, dummy_instr_seed_o[4:0] } : csr_mcause_i;
assign _0083_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14209.14-14209.27|generated/sv2v_out.v:14209.10-14229.8" */ _0008_ : 1'h1;
assign _0058_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14209.14-14209.27|generated/sv2v_out.v:14209.10-14229.8" */ { dummy_instr_seed_o[31:1], 1'h0 } : _0029_;
assign _0084_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14209.14-14209.27|generated/sv2v_out.v:14209.10-14229.8" */ _0009_ : 1'h1;
assign _0089_[1] = _1226_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14221.10-14221.39|generated/sv2v_out.v:14221.6-14228.9" */ _0000_[7] : _0098_;
assign _0096_[1:0] = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14209.14-14209.27|generated/sv2v_out.v:14209.10-14229.8" */ _0010_[3:2] : priv_mode_id_o;
assign _0096_[2] = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14209.14-14209.27|generated/sv2v_out.v:14209.10-14229.8" */ _0010_[4] : mstatus_q[5];
assign _0087_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14209.14-14209.27|generated/sv2v_out.v:14209.10-14229.8" */ _0012_ : 1'h1;
assign _0063_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14209.14-14209.27|generated/sv2v_out.v:14209.10-14229.8" */ dummy_instr_seed_o : csr_mtval_i;
assign _0088_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14209.14-14209.27|generated/sv2v_out.v:14209.10-14229.8" */ _0013_ : 1'h1;
assign _0069_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ 1'h1 : _0006_;
assign _0023_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ _0029_ : { dummy_instr_seed_o[31:1], 1'h0 };
assign _0068_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ 1'h1 : _0005_;
assign _0100_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ debug_cause_i : _0003_[8:6];
assign _0092_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ priv_mode_id_o : _0003_[1:0];
assign _0067_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ _0002_ : _0081_;
assign _0065_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ _0000_[7:6] : _0079_;
assign _0044_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ 1'h0 : _0060_;
assign _0078_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ _0013_ : _0088_;
assign _0048_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ dummy_instr_seed_o : _0063_;
assign _0073_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ _0008_ : _0083_;
assign _0031_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ { _1219_, _1218_, dummy_instr_seed_o[4:0] } : _0056_;
assign _0076_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ _0009_ : _0084_;
assign _0035_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ { dummy_instr_seed_o[31:1], 1'h0 } : _0058_;
assign _0077_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ _0012_ : _0087_;
assign _0085_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ _0010_[5:2] : _0096_;
assign _0026_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14202.9-14202.25|generated/sv2v_out.v:14202.5-14229.8" */ 1'h0 : _0055_;
assign _1263_ = csr_save_wb_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14194.5-14200.12" */ pc_wb_i : pc_id_i;
assign _1265_ = csr_save_id_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14194.5-14200.12" */ pc_id_i : _1263_;
assign _0029_ = csr_save_if_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14194.5-14200.12" */ pc_if_i : _1265_;
assign _1267_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ 1'h1 : _0002_;
assign _1268_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0002_ : _1267_;
assign cpuctrlsts_part_we = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0067_ : _1268_;
assign _1269_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ 1'h0 : _0000_[6];
assign _1271_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0000_[6] : _1269_;
assign cpuctrlsts_part_d[6] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0065_[0] : _1271_;
assign mstack_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0044_ : 1'h0;
assign depc_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0069_ : _0006_;
assign depc_d = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0023_ : { dummy_instr_seed_o[31:1], 1'h0 };
assign dcsr_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0068_ : _0005_;
assign dcsr_d[8:6] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0100_ : _0003_[8:6];
assign dcsr_d[1:0] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0092_ : _0003_[1:0];
assign mtval_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0078_ : _0013_;
assign mtval_d = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0048_ : dummy_instr_seed_o;
assign _1273_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0094_ : _0008_;
assign _1274_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0008_ : _1273_;
assign mcause_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0073_ : _1274_;
assign _1275_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0071_ : { _1219_, _1218_, dummy_instr_seed_o[4:0] };
assign _1277_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ { _1219_, _1218_, dummy_instr_seed_o[4:0] } : _1275_;
assign mcause_d = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0031_ : _1277_;
assign _1279_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0095_ : _0009_;
assign _1280_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0009_ : _1279_;
assign mepc_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0076_ : _1280_;
assign _1281_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0074_ : { dummy_instr_seed_o[31:1], 1'h0 };
assign _1283_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ { dummy_instr_seed_o[31:1], 1'h0 } : _1281_;
assign mepc_d = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0035_ : _1283_;
assign _1285_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ 1'h1 : _0012_;
assign _1286_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0012_ : _1285_;
assign mstatus_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0077_ : _1286_;
assign _0071_ = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14240.9-14240.19|generated/sv2v_out.v:14240.5-14251.8" */ mstack_cause_q : { _1219_, _1218_, dummy_instr_seed_o[4:0] };
assign double_fault_seen_o = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ _0026_ : 1'h0;
assign _1287_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ mstatus_q[3:2] : 2'hx;
assign _1289_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ dcsr_q[1:0] : _1287_;
assign priv_lvl_d = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.3-14255.10" */ 2'h3 : _1289_;
assign _0096_[3] = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14209.14-14209.27|generated/sv2v_out.v:14209.10-14229.8" */ _0010_[5] : 1'h0;
assign _0020_[31:28] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 4'h4 : dcsr_q[31:28];
assign _0045_[5:4] = _1292_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ { dummy_instr_seed_o[3], dummy_instr_seed_o[7] } : mstatus_q[5:4];
assign _0045_[3:2] = _1292_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ _0061_ : mstatus_q[3:2];
assign _0020_[15] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ dummy_instr_seed_o[15] : dcsr_q[15];
assign _0020_[14] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h0 : dcsr_q[14];
assign _0020_[27:16] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 12'h000 : dcsr_q[27:16];
assign _0045_[1:0] = _1292_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ { dummy_instr_seed_o[17], dummy_instr_seed_o[21] } : mstatus_q[1:0];
assign _0020_[1:0] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ _0053_ : dcsr_q[1:0];
assign _0020_[5] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h0 : dcsr_q[5];
assign _0020_[4] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h0 : dcsr_q[4];
assign _0020_[3] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h0 : dcsr_q[3];
assign _0020_[2] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ dummy_instr_seed_o[2] : dcsr_q[2];
assign _0020_[13:12] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ dummy_instr_seed_o[13:12] : dcsr_q[13:12];
assign _0020_[11] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h0 : dcsr_q[11];
assign _0053_ = _1225_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14166.10-14166.60|generated/sv2v_out.v:14166.6-14167.28" */ 2'h0 : dummy_instr_seed_o[1:0];
assign _0020_[9] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h0 : dcsr_q[9];
assign _0061_ = _1224_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14154.10-14154.66|generated/sv2v_out.v:14154.6-14155.31" */ 2'h0 : dummy_instr_seed_o[12:11];
assign _0047_ = _1292_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h1 : 1'h0;
assign _1296_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ _1295_;
assign _0019_ = _1297_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h1 : 1'h0;
assign _0017_ = _1297_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ { dummy_instr_seed_o[7:1], 1'h0 } : cpuctrlsts_part_q;
assign _0040_ = _1294_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ _1237_ : 32'd0;
assign _0038_ = _1296_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ _1237_ : 32'd0;
assign _0034_ = _1298_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h1 : 1'h0;
assign _0028_ = _1299_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h1 : 1'h0;
assign _0027_ = _1300_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h1 : 1'h0;
assign _0025_ = _1301_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h1 : 1'h0;
assign _0022_ = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h1 : 1'h0;
assign _0020_[10] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h0 : dcsr_q[10];
assign _0051_ = _1302_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h1 : csr_mtvec_init_i;
assign _0050_ = _1303_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h1 : 1'h0;
assign _0033_ = _1304_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h1 : 1'h0;
assign _0037_ = _1305_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h1 : 1'h0;
assign _0043_ = _1306_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h1 : 1'h0;
assign _0042_ = _1307_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14150.4-14191.11" */ 1'h1 : 1'h0;
assign _0002_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0019_ : 1'h0;
assign { _0000_[7:6], cpuctrlsts_part_d[5:0] } = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0017_ : cpuctrlsts_part_q;
assign mhpmcounterh_we = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0040_ : 32'd0;
assign mhpmcounter_we = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0038_ : 32'd0;
assign mcountinhibit_we = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0034_ : 1'h0;
assign dscratch1_en = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0028_ : 1'h0;
assign dscratch0_en = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0027_ : 1'h0;
assign _0006_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0025_ : 1'h0;
assign _0005_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0022_ : 1'h0;
assign { dcsr_d[31:9], _0003_[8:6], dcsr_d[5:2], _0003_[1:0] } = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ { _0020_[31:9], dcsr_q[8:6], _0020_[5:0] } : dcsr_q;
assign mtvec_en = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0051_ : csr_mtvec_init_i;
assign _0013_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0050_ : 1'h0;
assign _0008_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0033_ : 1'h0;
assign _0009_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0037_ : 1'h0;
assign mscratch_en = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0043_ : 1'h0;
assign mie_en = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0042_ : 1'h0;
assign _0012_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0047_ : 1'h0;
assign { _0010_[5:1], mstatus_d[0] } = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14149.7-14149.17|generated/sv2v_out.v:14149.3-14191.11" */ _0045_ : mstatus_q;
assign illegal_csr = _1308_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14110.8-14110.429|generated/sv2v_out.v:14110.4-14111.24" */ 1'h1 : _0007_;
assign _0016_ = _0267_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 32'd0 : 32'hxxxxxxxx;
assign _1294_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ _1293_;
assign _1298_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h320;
assign _1313_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hf12;
assign _1310_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ _1309_;
assign _1346_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h301;
assign _1314_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1f;
assign _1315_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1e;
assign _1316_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1d;
assign _1317_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1c;
assign _1318_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1b;
assign _1319_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1a;
assign _1320_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h19;
assign _1321_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h18;
assign _1322_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h17;
assign _1323_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h16;
assign _1324_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h15;
assign _1325_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h14;
assign _1326_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h13;
assign _1327_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h12;
assign _1328_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h11;
assign _1329_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h10;
assign _1330_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0f;
assign _1331_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0e;
assign _1332_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0d;
assign _1333_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0c;
assign _1334_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0b;
assign _1335_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0a;
assign _1336_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h09;
assign _1337_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h08;
assign _1338_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h07;
assign _1339_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h06;
assign _1340_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h05;
assign _1341_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h04;
assign _1342_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h03;
assign _1343_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h02;
assign _1344_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h01;
assign _1345_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ csr_addr_i[4:0];
assign _1299_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h7b3;
assign _1300_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h7b2;
assign _1301_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h7b1;
assign _1291_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h7b0;
assign _1198_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3bf;
assign _1199_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3be;
assign _1200_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3bd;
assign _1201_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3bc;
assign _1202_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3bb;
assign _1203_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3ba;
assign _1204_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3b9;
assign _1205_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3b8;
assign _1206_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3b7;
assign _1207_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3b6;
assign _1208_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3b5;
assign _1209_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3b4;
assign _1210_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3b3;
assign _1211_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3b2;
assign _1212_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3b1;
assign _1213_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3b0;
assign _1214_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3a3;
assign _1215_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3a2;
assign _1216_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3a1;
assign _1217_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h3a0;
assign _1312_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h344;
assign _1303_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h343;
assign _1304_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h342;
assign _1305_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h341;
assign _1302_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h305;
assign _1306_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h340;
assign _1307_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h304;
assign _1292_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h300;
assign _1311_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hf14;
assign _1295_[1] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb02;
assign _1295_[10] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb0b;
assign _1295_[11] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb0c;
assign _1295_[12] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb0d;
assign _1295_[13] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb0e;
assign _1295_[14] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb0f;
assign _1295_[15] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb10;
assign _1295_[16] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb11;
assign _1295_[17] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb12;
assign _1295_[18] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb13;
assign _1295_[19] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb14;
assign _1295_[2] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb03;
assign _1295_[20] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb15;
assign _1295_[21] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb16;
assign _1295_[22] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb17;
assign _1295_[23] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb18;
assign _1295_[24] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb19;
assign _1295_[25] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb1a;
assign _1295_[26] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb1b;
assign _1295_[27] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb1c;
assign _1295_[28] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb1d;
assign _1295_[29] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb1e;
assign _1295_[3] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb04;
assign _1295_[30] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb1f;
assign _1295_[4] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb05;
assign _1295_[5] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb06;
assign _1295_[6] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb07;
assign _1295_[7] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb08;
assign _1295_[8] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb09;
assign _1295_[9] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb0a;
assign _1309_[0] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h323;
assign _1309_[1] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h324;
assign _1309_[10] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h32d;
assign _1309_[11] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h32e;
assign _1309_[12] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h32f;
assign _1309_[13] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h330;
assign _1309_[14] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h331;
assign _1309_[15] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h332;
assign _1309_[16] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h333;
assign _1309_[17] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h334;
assign _1309_[18] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h335;
assign _1309_[19] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h336;
assign _1309_[2] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h325;
assign _1309_[20] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h337;
assign _1309_[21] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h338;
assign _1309_[22] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h339;
assign _1309_[23] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h33a;
assign _1309_[24] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h33b;
assign _1309_[25] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h33c;
assign _1309_[26] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h33d;
assign _1309_[27] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h33e;
assign _1309_[28] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h33f;
assign _1309_[3] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h326;
assign _1309_[4] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h327;
assign _1309_[5] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h328;
assign _1309_[6] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h329;
assign _1309_[7] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h32a;
assign _1309_[8] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h32b;
assign _1309_[9] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h32c;
assign _0007_ = _0266_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 1'h0 : 1'h1;
assign _1223_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h7c1;
assign _1297_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h7c0;
assign _1293_[0] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb80;
assign _1293_[1] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb82;
assign _1293_[10] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb8b;
assign _1293_[11] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb8c;
assign _1293_[12] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb8d;
assign _1293_[13] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb8e;
assign _1293_[14] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb8f;
assign _1293_[15] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb90;
assign _1293_[16] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb91;
assign _1293_[17] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb92;
assign _1293_[18] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb93;
assign _1293_[19] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb94;
assign _1293_[2] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb83;
assign _1293_[20] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb95;
assign _1293_[21] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb96;
assign _1293_[22] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb97;
assign _1293_[23] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb98;
assign _1293_[24] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb99;
assign _1293_[25] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb9a;
assign _1293_[26] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb9b;
assign _1293_[27] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb9c;
assign _1293_[28] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb9d;
assign _1293_[29] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb9e;
assign _1293_[3] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb84;
assign _1293_[30] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb9f;
assign _1293_[4] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb85;
assign _1293_[5] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb86;
assign _1293_[6] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb87;
assign _1293_[7] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb88;
assign _1293_[8] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb89;
assign _1293_[9] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb8a;
assign _1295_[0] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hb00;
assign _1347_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h306;
assign _1348_[0] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h30a;
assign _1348_[1] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h31a;
assign _1349_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'h310;
assign _1350_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hf15;
assign _1351_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hf13;
assign _1352_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 12'hf11;
assign dbg_csr = _0268_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13986.3-14108.10" */ 1'h1 : 1'h0;
assign _1308_ = | /* src = "generated/sv2v_out.v:14110.8-14110.429" */ { _1217_, _1216_, _1215_, _1214_, _1213_, _1212_, _1211_, _1210_, _1209_, _1208_, _1207_, _1206_, _1205_, _1204_, _1203_, _1202_, _1201_, _1200_, _1199_, _1198_ };
assign csr_wr = | /* src = "generated/sv2v_out.v:14272.18-14272.73" */ { _1222_, _1221_, _1220_ };
assign irq_pending_o = | /* src = "generated/sv2v_out.v:14285.25-14285.32" */ irqs_o;
assign _1237_ = $signed(_1232_) < 0 ? 1'h1 << - _1232_ : 1'h1 >> _1232_;
assign _1353_ = mcause_q[6] ? /* src = "generated/sv2v_out.v:14014.58-14014.116" */ 26'h3ffffff : 26'h0000000;
assign mtvec_d = csr_mtvec_init_i ? /* src = "generated/sv2v_out.v:14131.14-14131.112" */ { boot_addr_i[31:8], 8'h01 } : { dummy_instr_seed_o[31:8], 8'h01 };
assign priv_mode_lsu_o = mstatus_q[1] ? /* src = "generated/sv2v_out.v:14263.28-14263.71" */ mstatus_q[3:2] : priv_mode_id_o;
assign \mhpmcounter[2]  = _0112_ ? /* src = "generated/sv2v_out.v:14664.27-14664.94" */ minstret_next : minstret_raw;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14642.36-14650.3" */
\$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000  mcycle_counter_i (
.clk_i(clk_i),
.counter_inc_i(_0109_),
.counter_inc_i_t0(mcountinhibit_t0[0]),
.counter_val_i(dummy_instr_seed_o),
.counter_val_i_t0(dummy_instr_seed_o_t0),
.counter_val_o(\mhpmcounter[0] ),
.counter_val_o_t0(\mhpmcounter[0]_t0 ),
.counter_we_i(mhpmcounter_we[0]),
.counter_we_i_t0(mhpmcounter_we_t0[0]),
.counterh_we_i(mhpmcounterh_we[0]),
.counterh_we_i_t0(mhpmcounterh_we_t0[0]),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14654.4-14663.3" */
\$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter  minstret_counter_i (
.clk_i(clk_i),
.counter_inc_i(_0110_),
.counter_inc_i_t0(_0111_),
.counter_val_i(dummy_instr_seed_o),
.counter_val_i_t0(dummy_instr_seed_o_t0),
.counter_val_o(minstret_raw),
.counter_val_o_t0(minstret_raw_t0),
.counter_val_upd_o(minstret_next),
.counter_val_upd_o_t0(minstret_next_t0),
.counter_we_i(mhpmcounter_we[2]),
.counter_we_i_t0(mhpmcounter_we_t0[2]),
.counterh_we_i(mhpmcounterh_we[2]),
.counterh_we_i_t0(mhpmcounterh_we_t0[2]),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14873.4-14880.3" */
\$paramod$a088b13b9337f1e1fba58a671f47d7c7701ffa49\ibex_csr  u_cpuctrlsts_part_csr (
.clk_i(clk_i),
.rd_data_o(cpuctrlsts_part_q),
.rd_data_o_t0(cpuctrlsts_part_q_t0),
.rd_error_o(cpuctrlsts_part_err),
.rd_error_o_t0(cpuctrlsts_part_err_t0),
.rst_ni(rst_ni),
.wr_data_i(cpuctrlsts_part_d),
.wr_data_i_t0(cpuctrlsts_part_d_t0),
.wr_en_i(cpuctrlsts_part_we),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14375.4-14381.3" */
\$paramod$9a435d8f6db004a67362aa9a56f32ea481a74dbe\ibex_csr  u_dcsr_csr (
.clk_i(clk_i),
.rd_data_o(dcsr_q),
.rd_data_o_t0(dcsr_q_t0),
.rst_ni(rst_ni),
.wr_data_i(dcsr_d),
.wr_data_i_t0(dcsr_d_t0),
.wr_en_i(dcsr_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14386.4-14392.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_depc_csr (
.clk_i(clk_i),
.rd_data_o(csr_depc_o),
.rd_data_o_t0(csr_depc_o_t0),
.rst_ni(rst_ni),
.wr_data_i(depc_d),
.wr_data_i_t0(depc_d_t0),
.wr_en_i(depc_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14397.4-14403.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_dscratch0_csr (
.clk_i(clk_i),
.rd_data_o(dscratch0_q),
.rd_data_o_t0(dscratch0_q_t0),
.rst_ni(rst_ni),
.wr_data_i(dummy_instr_seed_o),
.wr_data_i_t0(dummy_instr_seed_o_t0),
.wr_en_i(dscratch0_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14408.4-14414.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_dscratch1_csr (
.clk_i(clk_i),
.rd_data_o(dscratch1_q),
.rd_data_o_t0(dscratch1_q_t0),
.rst_ni(rst_ni),
.wr_data_i(dummy_instr_seed_o),
.wr_data_i_t0(dummy_instr_seed_o_t0),
.wr_en_i(dscratch1_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14340.4-14346.3" */
\$paramod$34601000fe8707ce2501f5ed778e152043201712\ibex_csr  u_mcause_csr (
.clk_i(clk_i),
.rd_data_o(mcause_q),
.rd_data_o_t0(mcause_q_t0),
.rst_ni(rst_ni),
.wr_data_i(mcause_d),
.wr_data_i_t0(mcause_d_t0),
.wr_en_i(mcause_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14303.4-14309.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_mepc_csr (
.clk_i(clk_i),
.rd_data_o(csr_mepc_o),
.rd_data_o_t0(csr_mepc_o_t0),
.rst_ni(rst_ni),
.wr_data_i(mepc_d),
.wr_data_i_t0(mepc_d_t0),
.wr_en_i(mepc_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14318.4-14324.3" */
\$paramod$e55993a14b1fbc43320d549f521b710ed37596c6\ibex_csr  u_mie_csr (
.clk_i(clk_i),
.rd_data_o(mie_q),
.rd_data_o_t0(mie_q_t0),
.rst_ni(rst_ni),
.wr_data_i({ dummy_instr_seed_o[3], dummy_instr_seed_o[7], dummy_instr_seed_o[11], dummy_instr_seed_o[30:16] }),
.wr_data_i_t0({ dummy_instr_seed_o_t0[3], dummy_instr_seed_o_t0[7], dummy_instr_seed_o_t0[11], dummy_instr_seed_o_t0[30:16] }),
.wr_en_i(mie_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14329.4-14335.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_mscratch_csr (
.clk_i(clk_i),
.rd_data_o(mscratch_q),
.rd_data_o_t0(mscratch_q_t0),
.rst_ni(rst_ni),
.wr_data_i(dummy_instr_seed_o),
.wr_data_i_t0(dummy_instr_seed_o_t0),
.wr_en_i(mscratch_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14442.4-14448.3" */
\$paramod$34601000fe8707ce2501f5ed778e152043201712\ibex_csr  u_mstack_cause_csr (
.clk_i(clk_i),
.rd_data_o(mstack_cause_q),
.rd_data_o_t0(mstack_cause_q_t0),
.rst_ni(rst_ni),
.wr_data_i(mcause_q),
.wr_data_i_t0(mcause_q_t0),
.wr_en_i(mstack_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14420.4-14426.3" */
\$paramod$410b37fbfbfa994790f1902c150d2be939cadb3b\ibex_csr  u_mstack_csr (
.clk_i(clk_i),
.rd_data_o(mstack_q),
.rd_data_o_t0(mstack_q_t0),
.rst_ni(rst_ni),
.wr_data_i(mstatus_q[4:2]),
.wr_data_i_t0(mstatus_q_t0[4:2]),
.wr_en_i(mstack_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14431.4-14437.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_mstack_epc_csr (
.clk_i(clk_i),
.rd_data_o(mstack_epc_q),
.rd_data_o_t0(mstack_epc_q_t0),
.rst_ni(rst_ni),
.wr_data_i(csr_mepc_o),
.wr_data_i_t0(csr_mepc_o_t0),
.wr_en_i(mstack_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14291.4-14298.3" */
\$paramod$5714e31d82f2b8816750797f158ebea69a089104\ibex_csr  u_mstatus_csr (
.clk_i(clk_i),
.rd_data_o(mstatus_q),
.rd_data_o_t0(mstatus_q_t0),
.rd_error_o(mstatus_err),
.rd_error_o_t0(mstatus_err_t0),
.rst_ni(rst_ni),
.wr_data_i(mstatus_d),
.wr_data_i_t0(mstatus_d_t0),
.wr_en_i(mstatus_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14351.4-14357.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_mtval_csr (
.clk_i(clk_i),
.rd_data_o(csr_mtval_o),
.rd_data_o_t0(csr_mtval_o_t0),
.rst_ni(rst_ni),
.wr_data_i(mtval_d),
.wr_data_i_t0(mtval_d_t0),
.wr_en_i(mtval_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14362.4-14369.3" */
\$paramod$4f46e25470a27719ee9ca03cee1a0827eff766f7\ibex_csr  u_mtvec_csr (
.clk_i(clk_i),
.rd_data_o(csr_mtvec_o),
.rd_data_o_t0(csr_mtvec_o_t0),
.rd_error_o(mtvec_err),
.rd_error_o_t0(mtvec_err_t0),
.rst_ni(rst_ni),
.wr_data_i(mtvec_d),
.wr_data_i_t0(mtvec_d_t0),
.wr_en_i(mtvec_en),
.wr_en_i_t0(mtvec_en_t0)
);
assign _0000_[5:0] = cpuctrlsts_part_d[5:0];
assign _0001_[5:0] = cpuctrlsts_part_d_t0[5:0];
assign { _0003_[31:9], _0003_[5:2] } = { dcsr_d[31:9], dcsr_d[5:2] };
assign { _0004_[31:9], _0004_[5:2] } = { dcsr_d_t0[31:9], dcsr_d_t0[5:2] };
assign _0010_[0] = mstatus_d[0];
assign _0011_[0] = mstatus_d_t0[0];
assign _0020_[8:6] = dcsr_q[8:6];
assign _0021_[8:6] = dcsr_q_t0[8:6];
assign csr_mstatus_mie_o = mstatus_q[5];
assign csr_mstatus_mie_o_t0 = mstatus_q_t0[5];
assign csr_mstatus_tw_o = mstatus_q[0];
assign csr_mstatus_tw_o_t0 = mstatus_q_t0[0];
assign csr_pmp_addr_o = 136'h0000000000000000000000000000000000;
assign csr_pmp_addr_o_t0 = 136'h0000000000000000000000000000000000;
assign csr_pmp_cfg_o = 24'h000000;
assign csr_pmp_cfg_o_t0 = 24'h000000;
assign csr_pmp_mseccfg_o = 3'h0;
assign csr_pmp_mseccfg_o_t0 = 3'h0;
assign data_ind_timing_o = cpuctrlsts_part_q[1];
assign data_ind_timing_o_t0 = cpuctrlsts_part_q_t0[1];
assign debug_ebreakm_o = dcsr_q[15];
assign debug_ebreakm_o_t0 = dcsr_q_t0[15];
assign debug_ebreaku_o = dcsr_q[12];
assign debug_ebreaku_o_t0 = dcsr_q_t0[12];
assign debug_single_step_o = dcsr_q[2];
assign debug_single_step_o_t0 = dcsr_q_t0[2];
assign double_fault_seen_o_t0 = 1'h0;
assign dummy_instr_en_o = cpuctrlsts_part_q[2];
assign dummy_instr_en_o_t0 = cpuctrlsts_part_q_t0[2];
assign dummy_instr_mask_o = cpuctrlsts_part_q[5:3];
assign dummy_instr_mask_o_t0 = cpuctrlsts_part_q_t0[5:3];
assign dummy_instr_seed_en_o_t0 = 1'h0;
assign irq_pending_o_t0 = 1'h0;
assign { mcountinhibit[31:3], mcountinhibit[1] } = 30'h00000000;
assign { mcountinhibit_t0[31:3], mcountinhibit_t0[1] } = 30'h00000000;
assign trigger_match_o = 1'h0;
assign trigger_match_o_t0 = 1'h0;
endmodule

module \$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter (clk_i, rst_ni, counter_inc_i, counterh_we_i, counter_we_i, counter_val_i, counter_val_o, counter_val_upd_o, counter_inc_i_t0, counter_val_i_t0, counter_val_o_t0, counter_val_upd_o_t0, counter_we_i_t0, counterh_we_i_t0);
/* src = "generated/sv2v_out.v:13636.2-13650.5" */
wire [63:0] _00_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13636.2-13650.5" */
wire [63:0] _01_;
wire [63:0] _02_;
wire _03_;
wire _04_;
wire [63:0] _05_;
wire [31:0] _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire [63:0] _12_;
wire [31:0] _13_;
wire [31:0] _14_;
wire [31:0] _15_;
wire [31:0] _16_;
wire [63:0] _17_;
wire [63:0] _18_;
wire [63:0] _19_;
wire [31:0] _20_;
wire [31:0] _21_;
wire [63:0] _22_;
wire [63:0] _23_;
wire [63:0] _24_;
/* src = "generated/sv2v_out.v:13622.13-13622.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:13634.27-13634.36" */
wire [63:0] counter_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13634.27-13634.36" */
wire [63:0] counter_d_t0;
/* src = "generated/sv2v_out.v:13624.13-13624.26" */
input counter_inc_i;
wire counter_inc_i;
/* cellift = 32'd1 */
input counter_inc_i_t0;
wire counter_inc_i_t0;
/* src = "generated/sv2v_out.v:13632.13-13632.25" */
wire [63:0] counter_load;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13632.13-13632.25" */
wire [63:0] counter_load_t0;
/* src = "generated/sv2v_out.v:13627.20-13627.33" */
input [31:0] counter_val_i;
wire [31:0] counter_val_i;
/* cellift = 32'd1 */
input [31:0] counter_val_i_t0;
wire [31:0] counter_val_i_t0;
/* src = "generated/sv2v_out.v:13628.21-13628.34" */
output [63:0] counter_val_o;
reg [63:0] counter_val_o;
/* cellift = 32'd1 */
output [63:0] counter_val_o_t0;
reg [63:0] counter_val_o_t0;
/* src = "generated/sv2v_out.v:13629.21-13629.38" */
output [63:0] counter_val_upd_o;
wire [63:0] counter_val_upd_o;
/* cellift = 32'd1 */
output [63:0] counter_val_upd_o_t0;
wire [63:0] counter_val_upd_o_t0;
/* src = "generated/sv2v_out.v:13626.13-13626.25" */
input counter_we_i;
wire counter_we_i;
/* cellift = 32'd1 */
input counter_we_i_t0;
wire counter_we_i_t0;
/* src = "generated/sv2v_out.v:13625.13-13625.26" */
input counterh_we_i;
wire counterh_we_i;
/* cellift = 32'd1 */
input counterh_we_i_t0;
wire counterh_we_i_t0;
/* src = "generated/sv2v_out.v:13623.13-13623.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:13633.6-13633.8" */
wire we;
assign counter_val_upd_o = counter_val_o + /* src = "generated/sv2v_out.v:13635.23-13635.86" */ 64'h0000000000000001;
assign _02_ = ~ counter_val_o_t0;
assign _12_ = counter_val_o & _02_;
assign _23_ = _12_ + 64'h0000000000000001;
assign _19_ = counter_val_o | counter_val_o_t0;
assign _24_ = _19_ + 64'h0000000000000001;
assign _22_ = _23_ ^ _24_;
assign counter_val_upd_o_t0 = _22_ | counter_val_o_t0;
assign _03_ = ~ _10_;
assign _04_ = ~ _11_;
assign _13_ = { _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_ } & counter_d_t0[63:32];
assign _15_ = { _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_ } & counter_d_t0[31:0];
assign _14_ = { _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_ } & counter_val_o_t0[63:32];
assign _16_ = { _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_ } & counter_val_o_t0[31:0];
assign _20_ = _13_ | _14_;
assign _21_ = _15_ | _16_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter  */
/* PC_TAINT_INFO STATE_NAME counter_val_o_t0[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o_t0[63:32] <= 32'd0;
else counter_val_o_t0[63:32] <= _20_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter  */
/* PC_TAINT_INFO STATE_NAME counter_val_o_t0[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o_t0[31:0] <= 32'd0;
else counter_val_o_t0[31:0] <= _21_;
/* src = "generated/sv2v_out.v:13652.2-13656.27" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter  */
/* PC_TAINT_INFO STATE_NAME counter_val_o[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o[63:32] <= 32'd0;
else if (_10_) counter_val_o[63:32] <= counter_d[63:32];
/* src = "generated/sv2v_out.v:13652.2-13656.27" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter  */
/* PC_TAINT_INFO STATE_NAME counter_val_o[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o[31:0] <= 32'd0;
else if (_11_) counter_val_o[31:0] <= counter_d[31:0];
assign _05_ = ~ { we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we };
assign _06_ = ~ { counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i };
assign _17_ = _05_ & _01_;
assign counter_load_t0[31:0] = _06_ & counter_val_i_t0;
assign _01_ = { counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i } & counter_val_upd_o_t0;
assign _18_ = { we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we } & counter_load_t0;
assign counter_load_t0[63:32] = { counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i } & counter_val_i_t0;
assign counter_d_t0 = _17_ | _18_;
assign _07_ = | { we, counter_inc_i };
assign _08_ = { we, counterh_we_i } != 2'h2;
assign _09_ = { we, counterh_we_i } != 2'h3;
assign _10_ = & { _08_, _07_ };
assign _11_ = & { _07_, _09_ };
assign we = counter_we_i | /* src = "generated/sv2v_out.v:13637.8-13637.36" */ counterh_we_i;
assign _00_ = counter_inc_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13646.12-13646.25|generated/sv2v_out.v:13646.8-13649.44" */ counter_val_upd_o : 64'hxxxxxxxxxxxxxxxx;
assign counter_d = we ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13644.7-13644.9|generated/sv2v_out.v:13644.3-13649.44" */ counter_load : _00_;
assign counter_load[63:32] = counterh_we_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13640.7-13640.20|generated/sv2v_out.v:13640.3-13643.6" */ counter_val_i : 32'hxxxxxxxx;
assign counter_load[31:0] = counterh_we_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13640.7-13640.20|generated/sv2v_out.v:13640.3-13643.6" */ 32'hxxxxxxxx : counter_val_i;
endmodule

module \$paramod$e55993a14b1fbc43320d549f521b710ed37596c6\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _0_;
wire [17:0] _1_;
wire [17:0] _2_;
wire [17:0] _3_;
/* src = "generated/sv2v_out.v:14894.13-14894.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14898.28-14898.37" */
output [17:0] rd_data_o;
reg [17:0] rd_data_o;
/* cellift = 32'd1 */
output [17:0] rd_data_o_t0;
reg [17:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14899.14-14899.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14895.13-14895.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14896.27-14896.36" */
input [17:0] wr_data_i;
wire [17:0] wr_data_i;
/* cellift = 32'd1 */
input [17:0] wr_data_i_t0;
wire [17:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14897.13-14897.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _0_ = ~ wr_en_i;
assign _1_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _2_ = { _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_ } & rd_data_o_t0;
assign _3_ = _1_ | _2_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$e55993a14b1fbc43320d549f521b710ed37596c6\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 18'h00000;
else rd_data_o_t0 <= _3_;
/* src = "generated/sv2v_out.v:14901.2-14905.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$e55993a14b1fbc43320d549f521b710ed37596c6\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 18'h00000;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage (clk_i, rst_ni, ctrl_busy_o, illegal_insn_o, instr_valid_i, instr_rdata_i, instr_rdata_alu_i, instr_rdata_c_i, instr_is_compressed_i, instr_bp_taken_i, instr_req_o, instr_first_cycle_id_o, instr_valid_clear_o, id_in_ready_o, instr_exec_i, icache_inval_o, branch_decision_i, pc_set_o, pc_mux_o, nt_branch_mispredict_o, nt_branch_addr_o
, exc_pc_mux_o, exc_cause_o, illegal_c_insn_i, instr_fetch_err_i, instr_fetch_err_plus2_i, pc_id_i, ex_valid_i, lsu_resp_valid_i, alu_operator_ex_o, alu_operand_a_ex_o, alu_operand_b_ex_o, imd_val_we_ex_i, imd_val_d_ex_i, imd_val_q_ex_o, bt_a_operand_o, bt_b_operand_o, mult_en_ex_o, div_en_ex_o, mult_sel_ex_o, div_sel_ex_o, multdiv_operator_ex_o
, multdiv_signed_mode_ex_o, multdiv_operand_a_ex_o, multdiv_operand_b_ex_o, multdiv_ready_id_o, csr_access_o, csr_op_o, csr_op_en_o, csr_save_if_o, csr_save_id_o, csr_save_wb_o, csr_restore_mret_id_o, csr_restore_dret_id_o, csr_save_cause_o, csr_mtval_o, priv_mode_i, csr_mstatus_tw_i, illegal_csr_insn_i, data_ind_timing_i, lsu_req_o, lsu_we_o, lsu_type_o
, lsu_sign_ext_o, lsu_wdata_o, lsu_req_done_i, lsu_addr_incr_req_i, lsu_addr_last_i, csr_mstatus_mie_i, irq_pending_i, irqs_i, irq_nm_i, nmi_mode_o, lsu_load_err_i, lsu_load_resp_intg_err_i, lsu_store_err_i, lsu_store_resp_intg_err_i, expecting_load_resp_o, expecting_store_resp_o, debug_mode_o, debug_mode_entering_o, debug_cause_o, debug_csr_save_o, debug_req_i
, debug_single_step_i, debug_ebreakm_i, debug_ebreaku_i, trigger_match_i, result_ex_i, csr_rdata_i, rf_raddr_a_o, rf_rdata_a_i, rf_raddr_b_o, rf_rdata_b_i, rf_ren_a_o, rf_ren_b_o, rf_waddr_id_o, rf_wdata_id_o, rf_we_id_o, rf_rd_a_wb_match_o, rf_rd_b_wb_match_o, rf_waddr_wb_i, rf_wdata_fwd_wb_i, rf_write_wb_i, en_wb_o
, instr_type_wb_o, instr_perf_count_id_o, ready_wb_i, outstanding_load_wb_i, outstanding_store_wb_i, perf_jump_o, perf_branch_o, perf_tbranch_o, perf_dside_wait_o, perf_mul_wait_o, perf_div_wait_o, instr_id_done_o, ready_wb_i_t0, priv_mode_i_t0, perf_tbranch_o_t0, perf_jump_o_t0, pc_set_o_t0, pc_mux_o_t0, debug_ebreaku_i_t0, debug_ebreakm_i_t0, debug_csr_save_o_t0
, debug_cause_o_t0, ctrl_busy_o_t0, csr_save_wb_o_t0, csr_save_if_o_t0, csr_save_id_o_t0, csr_save_cause_o_t0, csr_restore_mret_id_o_t0, csr_restore_dret_id_o_t0, csr_mtval_o_t0, csr_mstatus_mie_i_t0, instr_req_o_t0, instr_rdata_i_t0, rf_ren_b_o_t0, rf_ren_a_o_t0, rf_raddr_b_o_t0, rf_raddr_a_o_t0, instr_rdata_alu_i_t0, illegal_insn_o_t0, illegal_c_insn_i_t0, icache_inval_o_t0, csr_op_o_t0
, csr_access_o_t0, perf_branch_o_t0, perf_div_wait_o_t0, perf_dside_wait_o_t0, perf_mul_wait_o_t0, result_ex_i_t0, trigger_match_i_t0, pc_id_i_t0, nt_branch_mispredict_o_t0, nmi_mode_o_t0, lsu_addr_last_i_t0, irqs_i_t0, irq_pending_i_t0, instr_valid_i_t0, instr_valid_clear_o_t0, instr_is_compressed_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_i_t0, instr_exec_i_t0, instr_bp_taken_i_t0, id_in_ready_o_t0
, rf_write_wb_i_t0, exc_pc_mux_o_t0, exc_cause_o_t0, debug_single_step_i_t0, debug_req_i_t0, debug_mode_o_t0, debug_mode_entering_o_t0, rf_rd_a_wb_match_o_t0, rf_rd_b_wb_match_o_t0, rf_rdata_a_i_t0, rf_rdata_b_i_t0, rf_waddr_id_o_t0, rf_waddr_wb_i_t0, rf_wdata_fwd_wb_i_t0, rf_wdata_id_o_t0, rf_we_id_o_t0, multdiv_signed_mode_ex_o_t0, nt_branch_addr_o_t0, outstanding_load_wb_i_t0, outstanding_store_wb_i_t0, alu_operand_a_ex_o_t0
, alu_operand_b_ex_o_t0, alu_operator_ex_o_t0, branch_decision_i_t0, bt_a_operand_o_t0, bt_b_operand_o_t0, csr_mstatus_tw_i_t0, csr_op_en_o_t0, csr_rdata_i_t0, data_ind_timing_i_t0, div_en_ex_o_t0, div_sel_ex_o_t0, en_wb_o_t0, ex_valid_i_t0, expecting_load_resp_o_t0, expecting_store_resp_o_t0, illegal_csr_insn_i_t0, imd_val_d_ex_i_t0, imd_val_q_ex_o_t0, imd_val_we_ex_i_t0, instr_first_cycle_id_o_t0, instr_id_done_o_t0
, instr_perf_count_id_o_t0, instr_rdata_c_i_t0, instr_type_wb_o_t0, irq_nm_i_t0, lsu_addr_incr_req_i_t0, lsu_load_err_i_t0, lsu_load_resp_intg_err_i_t0, lsu_req_done_i_t0, lsu_req_o_t0, lsu_resp_valid_i_t0, lsu_sign_ext_o_t0, lsu_store_err_i_t0, lsu_store_resp_intg_err_i_t0, lsu_type_o_t0, lsu_wdata_o_t0, lsu_we_o_t0, mult_en_ex_o_t0, mult_sel_ex_o_t0, multdiv_operand_a_ex_o_t0, multdiv_operand_b_ex_o_t0, multdiv_operator_ex_o_t0
, multdiv_ready_id_o_t0);
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0001_;
/* src = "generated/sv2v_out.v:17501.2-17510.5" */
wire _0002_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0003_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0004_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0005_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0007_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0008_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0009_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0010_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0011_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0012_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0013_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0014_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0015_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0016_;
/* src = "generated/sv2v_out.v:17501.2-17510.5" */
wire _0017_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0018_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0019_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0020_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0021_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0022_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0023_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0024_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0025_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0026_;
/* src = "generated/sv2v_out.v:17501.2-17510.5" */
wire _0027_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0028_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0029_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0030_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0031_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0032_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0033_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0034_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0035_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0036_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0037_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0038_;
/* src = "generated/sv2v_out.v:17655.2-17714.5" */
wire _0039_;
/* src = "generated/sv2v_out.v:17321.22-17321.56" */
wire _0040_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17321.22-17321.56" */
wire _0041_;
/* src = "generated/sv2v_out.v:17321.21-17321.75" */
wire _0042_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17321.21-17321.75" */
wire _0043_;
/* src = "generated/sv2v_out.v:17436.23-17436.50" */
wire _0044_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17436.23-17436.50" */
wire _0045_;
/* src = "generated/sv2v_out.v:17512.73-17512.104" */
wire _0046_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17512.73-17512.104" */
wire _0047_;
/* src = "generated/sv2v_out.v:17587.38-17587.68" */
wire _0048_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17587.38-17587.68" */
wire _0049_;
/* src = "generated/sv2v_out.v:17595.24-17595.54" */
wire _0050_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17595.24-17595.54" */
wire _0051_;
/* src = "generated/sv2v_out.v:17703.19-17703.41" */
wire _0052_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17703.19-17703.41" */
wire _0053_;
/* src = "generated/sv2v_out.v:17704.10-17704.38" */
wire _0054_;
/* src = "generated/sv2v_out.v:17717.23-17717.44" */
wire _0055_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17717.23-17717.44" */
wire _0056_;
/* src = "generated/sv2v_out.v:17754.40-17754.93" */
wire _0057_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17754.40-17754.93" */
wire _0058_;
/* src = "generated/sv2v_out.v:17762.37-17762.64" */
wire _0059_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17762.37-17762.64" */
wire _0060_;
/* src = "generated/sv2v_out.v:17762.36-17762.86" */
wire _0061_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17762.36-17762.86" */
wire _0062_;
/* src = "generated/sv2v_out.v:17782.32-17782.61" */
wire _0063_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17782.32-17782.61" */
wire _0064_;
/* src = "generated/sv2v_out.v:17786.36-17786.64" */
wire _0065_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17786.36-17786.64" */
wire _0066_;
/* src = "generated/sv2v_out.v:17786.35-17786.85" */
wire _0067_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17786.35-17786.85" */
wire _0068_;
/* src = "generated/sv2v_out.v:17786.34-17786.108" */
wire _0069_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17786.34-17786.108" */
wire _0070_;
wire _0071_;
wire _0072_;
wire _0073_;
wire [31:0] _0074_;
wire [31:0] _0075_;
wire [31:0] _0076_;
wire [31:0] _0077_;
wire [31:0] _0078_;
wire _0079_;
wire [31:0] _0080_;
wire [31:0] _0081_;
wire [31:0] _0082_;
wire [31:0] _0083_;
wire _0084_;
wire _0085_;
wire _0086_;
wire _0087_;
wire _0088_;
wire _0089_;
wire [31:0] _0090_;
wire [31:0] _0091_;
wire _0092_;
wire _0093_;
wire _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire _0109_;
wire _0110_;
wire _0111_;
wire _0112_;
wire _0113_;
wire _0114_;
wire _0115_;
wire _0116_;
wire _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire _0139_;
wire _0140_;
wire _0141_;
wire _0142_;
wire _0143_;
wire _0144_;
wire _0145_;
wire _0146_;
wire _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
wire _0152_;
wire _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire _0186_;
wire _0187_;
wire _0188_;
wire _0189_;
wire _0190_;
wire _0191_;
wire _0192_;
wire _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire _0199_;
wire _0200_;
wire _0201_;
wire _0202_;
wire _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire [33:0] _0219_;
wire [33:0] _0220_;
wire _0221_;
wire [33:0] _0222_;
wire [33:0] _0223_;
wire [31:0] _0224_;
wire [31:0] _0225_;
wire [31:0] _0226_;
wire [31:0] _0227_;
wire [31:0] _0228_;
wire [31:0] _0229_;
wire [31:0] _0230_;
wire [31:0] _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire [31:0] _0235_;
wire [31:0] _0236_;
wire [31:0] _0237_;
wire [31:0] _0238_;
wire [31:0] _0239_;
wire [31:0] _0240_;
wire [31:0] _0241_;
wire [31:0] _0242_;
wire _0243_;
wire _0244_;
wire _0245_;
wire _0246_;
wire _0247_;
wire _0248_;
wire _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire _0271_;
wire _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire _0276_;
wire _0277_;
wire _0278_;
wire _0279_;
wire _0280_;
wire _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire _0285_;
wire _0286_;
wire _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire _0294_;
wire _0295_;
wire _0296_;
wire [31:0] _0297_;
wire [31:0] _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire _0324_;
wire _0325_;
wire _0326_;
wire _0327_;
wire _0328_;
wire _0329_;
wire _0330_;
wire _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire [33:0] _0335_;
wire [33:0] _0336_;
wire _0337_;
wire _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire _0344_;
wire _0345_;
wire _0346_;
wire _0347_;
wire _0348_;
wire _0349_;
wire _0350_;
wire [31:0] _0351_;
/* cellift = 32'd1 */
wire [31:0] _0352_;
wire [31:0] _0353_;
/* cellift = 32'd1 */
wire [31:0] _0354_;
wire [31:0] _0355_;
/* cellift = 32'd1 */
wire [31:0] _0356_;
wire [31:0] _0357_;
/* cellift = 32'd1 */
wire [31:0] _0358_;
wire [31:0] _0359_;
/* cellift = 32'd1 */
wire [31:0] _0360_;
wire [31:0] _0361_;
/* cellift = 32'd1 */
wire [31:0] _0362_;
wire [31:0] _0363_;
/* cellift = 32'd1 */
wire [31:0] _0364_;
/* src = "generated/sv2v_out.v:17503.34-17503.50" */
wire _0365_;
/* src = "generated/sv2v_out.v:17503.56-17503.72" */
wire _0366_;
/* src = "generated/sv2v_out.v:17504.11-17504.42" */
wire _0367_;
/* src = "generated/sv2v_out.v:17504.48-17504.79" */
wire _0368_;
/* src = "generated/sv2v_out.v:17504.86-17504.117" */
wire _0369_;
/* src = "generated/sv2v_out.v:17504.124-17504.153" */
wire _0370_;
/* src = "generated/sv2v_out.v:17508.11-17508.42" */
wire _0371_;
/* src = "generated/sv2v_out.v:17508.48-17508.79" */
wire _0372_;
/* src = "generated/sv2v_out.v:17508.86-17508.117" */
wire _0373_;
/* src = "generated/sv2v_out.v:17508.124-17508.155" */
wire _0374_;
/* src = "generated/sv2v_out.v:17503.7-17503.74" */
wire _0375_;
/* src = "generated/sv2v_out.v:17507.12-17507.55" */
wire _0376_;
/* src = "generated/sv2v_out.v:17503.33-17503.73" */
wire _0377_;
/* src = "generated/sv2v_out.v:17504.10-17504.80" */
wire _0378_;
/* src = "generated/sv2v_out.v:17504.9-17504.118" */
wire _0379_;
/* src = "generated/sv2v_out.v:17504.8-17504.154" */
wire _0380_;
/* src = "generated/sv2v_out.v:17508.10-17508.80" */
wire _0381_;
/* src = "generated/sv2v_out.v:17508.9-17508.118" */
wire _0382_;
/* src = "generated/sv2v_out.v:17508.8-17508.156" */
wire _0383_;
/* src = "generated/sv2v_out.v:17682.20-17682.80" */
wire _0384_;
/* src = "generated/sv2v_out.v:17507.38-17507.54" */
wire _0385_;
/* src = "generated/sv2v_out.v:17512.31-17512.51" */
wire _0386_;
/* src = "generated/sv2v_out.v:17321.38-17321.56" */
wire _0387_;
/* src = "generated/sv2v_out.v:17321.60-17321.75" */
wire _0388_;
/* src = "generated/sv2v_out.v:17511.45-17511.58" */
wire _0389_;
/* src = "generated/sv2v_out.v:17619.95-17619.115" */
wire _0390_;
/* src = "generated/sv2v_out.v:17717.23-17717.32" */
wire _0391_;
/* src = "generated/sv2v_out.v:17717.35-17717.44" */
wire _0392_;
/* src = "generated/sv2v_out.v:17754.55-17754.72" */
wire _0393_;
/* src = "generated/sv2v_out.v:17762.90-17762.97" */
wire _0394_;
/* src = "generated/sv2v_out.v:17786.36-17786.46" */
wire _0395_;
/* src = "generated/sv2v_out.v:17786.49-17786.64" */
wire _0396_;
/* src = "generated/sv2v_out.v:17512.56-17512.105" */
wire _0397_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17512.56-17512.105" */
wire _0398_;
/* src = "generated/sv2v_out.v:17513.45-17513.82" */
wire _0399_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17513.45-17513.82" */
wire _0400_;
/* src = "generated/sv2v_out.v:17513.44-17513.103" */
wire _0401_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17513.44-17513.103" */
wire _0402_;
/* src = "generated/sv2v_out.v:17513.43-17513.125" */
wire _0403_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17513.43-17513.125" */
wire _0404_;
/* src = "generated/sv2v_out.v:17619.36-17619.65" */
wire _0405_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17619.36-17619.65" */
wire _0406_;
/* src = "generated/sv2v_out.v:17619.35-17619.91" */
wire _0407_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17619.35-17619.91" */
wire _0408_;
/* src = "generated/sv2v_out.v:17683.23-17683.81" */
wire _0409_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17683.23-17683.81" */
wire _0410_;
/* src = "generated/sv2v_out.v:17716.23-17716.64" */
wire _0411_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17716.23-17716.64" */
wire _0412_;
/* src = "generated/sv2v_out.v:17716.22-17716.78" */
wire _0413_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17716.22-17716.78" */
wire _0414_;
/* src = "generated/sv2v_out.v:17716.21-17716.94" */
wire _0415_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17716.21-17716.94" */
wire _0416_;
/* src = "generated/sv2v_out.v:17754.55-17754.92" */
wire _0417_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17754.55-17754.92" */
wire _0418_;
wire _0419_;
wire _0420_;
wire _0421_;
wire _0422_;
wire _0423_;
wire _0424_;
wire _0425_;
wire _0426_;
wire _0427_;
wire _0428_;
wire _0429_;
wire _0430_;
wire _0431_;
wire _0432_;
/* cellift = 32'd1 */
wire _0433_;
wire _0434_;
/* cellift = 32'd1 */
wire _0435_;
wire _0436_;
/* cellift = 32'd1 */
wire _0437_;
wire _0438_;
/* cellift = 32'd1 */
wire _0439_;
wire _0440_;
wire _0441_;
wire _0442_;
wire _0443_;
/* cellift = 32'd1 */
wire _0444_;
wire _0445_;
/* cellift = 32'd1 */
wire _0446_;
wire _0447_;
wire _0448_;
/* cellift = 32'd1 */
wire _0449_;
wire _0450_;
/* cellift = 32'd1 */
wire _0451_;
wire _0452_;
/* cellift = 32'd1 */
wire _0453_;
wire _0454_;
wire _0455_;
wire _0456_;
wire _0457_;
wire _0458_;
/* src = "generated/sv2v_out.v:17416.21-17416.72" */
wire [31:0] _0459_;
/* src = "generated/sv2v_out.v:17682.20-17682.94" */
wire _0460_;
/* src = "generated/sv2v_out.v:17332.7-17332.25" */
wire alu_multicycle_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17332.7-17332.25" */
/* unused_bits = "0" */
wire alu_multicycle_dec_t0;
/* src = "generated/sv2v_out.v:17328.13-17328.29" */
wire [1:0] alu_op_a_mux_sel;
/* src = "generated/sv2v_out.v:17329.13-17329.33" */
wire [1:0] alu_op_a_mux_sel_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17329.13-17329.33" */
/* unused_bits = "0 1" */
wire [1:0] alu_op_a_mux_sel_dec_t0;
/* src = "generated/sv2v_out.v:17330.7-17330.23" */
wire alu_op_b_mux_sel;
/* src = "generated/sv2v_out.v:17331.7-17331.27" */
wire alu_op_b_mux_sel_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17331.7-17331.27" */
/* unused_bits = "0" */
wire alu_op_b_mux_sel_dec_t0;
/* src = "generated/sv2v_out.v:17182.21-17182.39" */
output [31:0] alu_operand_a_ex_o;
wire [31:0] alu_operand_a_ex_o;
/* cellift = 32'd1 */
output [31:0] alu_operand_a_ex_o_t0;
wire [31:0] alu_operand_a_ex_o_t0;
/* src = "generated/sv2v_out.v:17183.21-17183.39" */
output [31:0] alu_operand_b_ex_o;
wire [31:0] alu_operand_b_ex_o;
/* cellift = 32'd1 */
output [31:0] alu_operand_b_ex_o_t0;
wire [31:0] alu_operand_b_ex_o_t0;
/* src = "generated/sv2v_out.v:17181.20-17181.37" */
output [6:0] alu_operator_ex_o;
wire [6:0] alu_operator_ex_o;
/* cellift = 32'd1 */
output [6:0] alu_operator_ex_o_t0;
wire [6:0] alu_operator_ex_o_t0;
/* src = "generated/sv2v_out.v:17168.13-17168.30" */
input branch_decision_i;
wire branch_decision_i;
/* cellift = 32'd1 */
input branch_decision_i_t0;
wire branch_decision_i_t0;
/* src = "generated/sv2v_out.v:17279.7-17279.20" */
wire branch_in_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17279.7-17279.20" */
wire branch_in_dec_t0;
/* src = "generated/sv2v_out.v:17284.7-17284.29" */
wire branch_jump_set_done_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17284.7-17284.29" */
wire branch_jump_set_done_d_t0;
/* src = "generated/sv2v_out.v:17283.6-17283.28" */
reg branch_jump_set_done_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17283.6-17283.28" */
reg branch_jump_set_done_q_t0;
/* src = "generated/sv2v_out.v:17280.7-17280.17" */
wire branch_set;
/* src = "generated/sv2v_out.v:17281.7-17281.21" */
reg branch_set_raw;
/* src = "generated/sv2v_out.v:17282.6-17282.22" */
wire branch_set_raw_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17282.6-17282.22" */
wire branch_set_raw_d_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17281.7-17281.21" */
reg branch_set_raw_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17280.7-17280.17" */
wire branch_set_t0;
/* src = "generated/sv2v_out.v:17286.7-17286.19" */
wire branch_taken;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17286.7-17286.19" */
wire branch_taken_t0;
/* src = "generated/sv2v_out.v:17335.13-17335.25" */
/* unused_bits = "0 1" */
wire [1:0] bt_a_mux_sel;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17335.13-17335.25" */
/* unused_bits = "0 1" */
wire [1:0] bt_a_mux_sel_t0;
/* src = "generated/sv2v_out.v:17187.20-17187.34" */
output [31:0] bt_a_operand_o;
wire [31:0] bt_a_operand_o;
/* cellift = 32'd1 */
output [31:0] bt_a_operand_o_t0;
wire [31:0] bt_a_operand_o_t0;
/* src = "generated/sv2v_out.v:17336.13-17336.25" */
/* unused_bits = "0 1 2" */
wire [2:0] bt_b_mux_sel;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17336.13-17336.25" */
/* unused_bits = "0 1 2" */
wire [2:0] bt_b_mux_sel_t0;
/* src = "generated/sv2v_out.v:17188.20-17188.34" */
output [31:0] bt_b_operand_o;
wire [31:0] bt_b_operand_o;
/* cellift = 32'd1 */
output [31:0] bt_b_operand_o_t0;
wire [31:0] bt_b_operand_o_t0;
/* src = "generated/sv2v_out.v:17152.13-17152.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:17295.7-17295.21" */
wire controller_run;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17295.7-17295.21" */
wire controller_run_t0;
/* src = "generated/sv2v_out.v:17198.14-17198.26" */
output csr_access_o;
wire csr_access_o;
/* cellift = 32'd1 */
output csr_access_o_t0;
wire csr_access_o_t0;
/* src = "generated/sv2v_out.v:17220.13-17220.30" */
input csr_mstatus_mie_i;
wire csr_mstatus_mie_i;
/* cellift = 32'd1 */
input csr_mstatus_mie_i_t0;
wire csr_mstatus_mie_i_t0;
/* src = "generated/sv2v_out.v:17209.13-17209.29" */
input csr_mstatus_tw_i;
wire csr_mstatus_tw_i;
/* cellift = 32'd1 */
input csr_mstatus_tw_i_t0;
wire csr_mstatus_tw_i_t0;
/* src = "generated/sv2v_out.v:17207.21-17207.32" */
output [31:0] csr_mtval_o;
wire [31:0] csr_mtval_o;
/* cellift = 32'd1 */
output [31:0] csr_mtval_o_t0;
wire [31:0] csr_mtval_o_t0;
/* src = "generated/sv2v_out.v:17200.14-17200.25" */
output csr_op_en_o;
wire csr_op_en_o;
/* cellift = 32'd1 */
output csr_op_en_o_t0;
wire csr_op_en_o_t0;
/* src = "generated/sv2v_out.v:17199.20-17199.28" */
output [1:0] csr_op_o;
wire [1:0] csr_op_o;
/* cellift = 32'd1 */
output [1:0] csr_op_o_t0;
wire [1:0] csr_op_o_t0;
/* src = "generated/sv2v_out.v:17353.6-17353.20" */
wire csr_pipe_flush;
/* src = "generated/sv2v_out.v:17241.20-17241.31" */
input [31:0] csr_rdata_i;
wire [31:0] csr_rdata_i;
/* cellift = 32'd1 */
input [31:0] csr_rdata_i_t0;
wire [31:0] csr_rdata_i_t0;
/* src = "generated/sv2v_out.v:17205.14-17205.35" */
output csr_restore_dret_id_o;
wire csr_restore_dret_id_o;
/* cellift = 32'd1 */
output csr_restore_dret_id_o_t0;
wire csr_restore_dret_id_o_t0;
/* src = "generated/sv2v_out.v:17204.14-17204.35" */
output csr_restore_mret_id_o;
wire csr_restore_mret_id_o;
/* cellift = 32'd1 */
output csr_restore_mret_id_o_t0;
wire csr_restore_mret_id_o_t0;
/* src = "generated/sv2v_out.v:17206.14-17206.30" */
output csr_save_cause_o;
wire csr_save_cause_o;
/* cellift = 32'd1 */
output csr_save_cause_o_t0;
wire csr_save_cause_o_t0;
/* src = "generated/sv2v_out.v:17202.14-17202.27" */
output csr_save_id_o;
wire csr_save_id_o;
/* cellift = 32'd1 */
output csr_save_id_o_t0;
wire csr_save_id_o_t0;
/* src = "generated/sv2v_out.v:17201.14-17201.27" */
output csr_save_if_o;
wire csr_save_if_o;
/* cellift = 32'd1 */
output csr_save_if_o_t0;
wire csr_save_if_o_t0;
/* src = "generated/sv2v_out.v:17203.14-17203.27" */
output csr_save_wb_o;
wire csr_save_wb_o;
/* cellift = 32'd1 */
output csr_save_wb_o_t0;
wire csr_save_wb_o_t0;
/* src = "generated/sv2v_out.v:17154.14-17154.25" */
output ctrl_busy_o;
wire ctrl_busy_o;
/* cellift = 32'd1 */
output ctrl_busy_o_t0;
wire ctrl_busy_o_t0;
/* src = "generated/sv2v_out.v:17211.13-17211.30" */
input data_ind_timing_i;
wire data_ind_timing_i;
/* cellift = 32'd1 */
input data_ind_timing_i_t0;
wire data_ind_timing_i_t0;
/* src = "generated/sv2v_out.v:17233.20-17233.33" */
output [2:0] debug_cause_o;
wire [2:0] debug_cause_o;
/* cellift = 32'd1 */
output [2:0] debug_cause_o_t0;
wire [2:0] debug_cause_o_t0;
/* src = "generated/sv2v_out.v:17234.14-17234.30" */
output debug_csr_save_o;
wire debug_csr_save_o;
/* cellift = 32'd1 */
output debug_csr_save_o_t0;
wire debug_csr_save_o_t0;
/* src = "generated/sv2v_out.v:17237.13-17237.28" */
input debug_ebreakm_i;
wire debug_ebreakm_i;
/* cellift = 32'd1 */
input debug_ebreakm_i_t0;
wire debug_ebreakm_i_t0;
/* src = "generated/sv2v_out.v:17238.13-17238.28" */
input debug_ebreaku_i;
wire debug_ebreaku_i;
/* cellift = 32'd1 */
input debug_ebreaku_i_t0;
wire debug_ebreaku_i_t0;
/* src = "generated/sv2v_out.v:17232.14-17232.35" */
output debug_mode_entering_o;
wire debug_mode_entering_o;
/* cellift = 32'd1 */
output debug_mode_entering_o_t0;
wire debug_mode_entering_o_t0;
/* src = "generated/sv2v_out.v:17231.14-17231.26" */
output debug_mode_o;
wire debug_mode_o;
/* cellift = 32'd1 */
output debug_mode_o_t0;
wire debug_mode_o_t0;
/* src = "generated/sv2v_out.v:17235.13-17235.24" */
input debug_req_i;
wire debug_req_i;
/* cellift = 32'd1 */
input debug_req_i_t0;
wire debug_req_i_t0;
/* src = "generated/sv2v_out.v:17236.13-17236.32" */
input debug_single_step_i;
wire debug_single_step_i;
/* cellift = 32'd1 */
input debug_single_step_i_t0;
wire debug_single_step_i_t0;
/* src = "generated/sv2v_out.v:17343.7-17343.17" */
wire div_en_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17343.7-17343.17" */
wire div_en_dec_t0;
/* src = "generated/sv2v_out.v:17190.14-17190.25" */
output div_en_ex_o;
wire div_en_ex_o;
/* cellift = 32'd1 */
output div_en_ex_o_t0;
wire div_en_ex_o_t0;
/* src = "generated/sv2v_out.v:17192.14-17192.26" */
output div_sel_ex_o;
wire div_sel_ex_o;
/* cellift = 32'd1 */
output div_sel_ex_o_t0;
wire div_sel_ex_o_t0;
/* src = "generated/sv2v_out.v:17274.7-17274.20" */
wire dret_insn_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17274.7-17274.20" */
wire dret_insn_dec_t0;
/* src = "generated/sv2v_out.v:17272.7-17272.16" */
wire ebrk_insn;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17272.7-17272.16" */
wire ebrk_insn_t0;
/* src = "generated/sv2v_out.v:17275.7-17275.21" */
wire ecall_insn_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17275.7-17275.21" */
wire ecall_insn_dec_t0;
/* src = "generated/sv2v_out.v:17256.14-17256.21" */
output en_wb_o;
wire en_wb_o;
/* cellift = 32'd1 */
output en_wb_o_t0;
wire en_wb_o_t0;
/* src = "generated/sv2v_out.v:17179.13-17179.23" */
input ex_valid_i;
wire ex_valid_i;
/* cellift = 32'd1 */
input ex_valid_i_t0;
wire ex_valid_i_t0;
/* src = "generated/sv2v_out.v:17174.20-17174.31" */
output [6:0] exc_cause_o;
wire [6:0] exc_cause_o;
/* cellift = 32'd1 */
output [6:0] exc_cause_o_t0;
wire [6:0] exc_cause_o_t0;
/* src = "generated/sv2v_out.v:17173.20-17173.32" */
output [1:0] exc_pc_mux_o;
wire [1:0] exc_pc_mux_o;
/* cellift = 32'd1 */
output [1:0] exc_pc_mux_o_t0;
wire [1:0] exc_pc_mux_o_t0;
/* src = "generated/sv2v_out.v:17229.14-17229.35" */
output expecting_load_resp_o;
wire expecting_load_resp_o;
/* cellift = 32'd1 */
output expecting_load_resp_o_t0;
wire expecting_load_resp_o_t0;
/* src = "generated/sv2v_out.v:17230.14-17230.36" */
output expecting_store_resp_o;
wire expecting_store_resp_o;
/* cellift = 32'd1 */
output expecting_store_resp_o_t0;
wire expecting_store_resp_o_t0;
/* src = "generated/sv2v_out.v:17303.7-17303.15" */
wire flush_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17303.7-17303.15" */
wire flush_id_t0;
/* src = "generated/sv2v_out.v:17629.8-17629.22" */
reg \g_sec_branch_taken.branch_taken_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17629.8-17629.22" */
reg \g_sec_branch_taken.branch_taken_q_t0 ;
/* src = "generated/sv2v_out.v:17771.9-17771.28" */
/* unused_bits = "0" */
wire \gen_no_stall_mem.unused_id_exception ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17771.9-17771.28" */
/* unused_bits = "0" */
wire \gen_no_stall_mem.unused_id_exception_t0 ;
/* src = "generated/sv2v_out.v:17769.9-17769.28" */
/* unused_bits = "0" */
wire \gen_no_stall_mem.unused_wb_exception ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17769.9-17769.28" */
/* unused_bits = "0" */
wire \gen_no_stall_mem.unused_wb_exception_t0 ;
/* src = "generated/sv2v_out.v:17167.14-17167.28" */
output icache_inval_o;
wire icache_inval_o;
/* cellift = 32'd1 */
output icache_inval_o_t0;
wire icache_inval_o_t0;
/* src = "generated/sv2v_out.v:17648.6-17648.14" */
wire id_fsm_d;
/* src = "generated/sv2v_out.v:17647.6-17647.14" */
reg id_fsm_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17647.6-17647.14" */
reg id_fsm_q_t0;
/* src = "generated/sv2v_out.v:17165.14-17165.27" */
output id_in_ready_o;
wire id_in_ready_o;
/* cellift = 32'd1 */
output id_in_ready_o_t0;
wire id_in_ready_o_t0;
/* src = "generated/sv2v_out.v:17175.13-17175.29" */
input illegal_c_insn_i;
wire illegal_c_insn_i;
/* cellift = 32'd1 */
input illegal_c_insn_i_t0;
wire illegal_c_insn_i_t0;
/* src = "generated/sv2v_out.v:17210.13-17210.31" */
input illegal_csr_insn_i;
wire illegal_csr_insn_i;
/* cellift = 32'd1 */
input illegal_csr_insn_i_t0;
wire illegal_csr_insn_i_t0;
/* src = "generated/sv2v_out.v:17270.7-17270.24" */
wire illegal_dret_insn;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17270.7-17270.24" */
wire illegal_dret_insn_t0;
/* src = "generated/sv2v_out.v:17269.7-17269.23" */
wire illegal_insn_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17269.7-17269.23" */
wire illegal_insn_dec_t0;
/* src = "generated/sv2v_out.v:17155.14-17155.28" */
output illegal_insn_o;
wire illegal_insn_o;
/* cellift = 32'd1 */
output illegal_insn_o_t0;
wire illegal_insn_o_t0;
/* src = "generated/sv2v_out.v:17271.7-17271.25" */
wire illegal_umode_insn;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17271.7-17271.25" */
wire illegal_umode_insn_t0;
/* src = "generated/sv2v_out.v:17185.20-17185.34" */
input [67:0] imd_val_d_ex_i;
wire [67:0] imd_val_d_ex_i;
/* cellift = 32'd1 */
input [67:0] imd_val_d_ex_i_t0;
wire [67:0] imd_val_d_ex_i_t0;
/* src = "generated/sv2v_out.v:17186.21-17186.35" */
output [67:0] imd_val_q_ex_o;
reg [67:0] imd_val_q_ex_o;
/* cellift = 32'd1 */
output [67:0] imd_val_q_ex_o_t0;
reg [67:0] imd_val_q_ex_o_t0;
/* src = "generated/sv2v_out.v:17184.19-17184.34" */
input [1:0] imd_val_we_ex_i;
wire [1:0] imd_val_we_ex_i;
/* cellift = 32'd1 */
input [1:0] imd_val_we_ex_i_t0;
wire [1:0] imd_val_we_ex_i_t0;
/* src = "generated/sv2v_out.v:17312.14-17312.19" */
wire [31:0] imm_a;
/* src = "generated/sv2v_out.v:17337.7-17337.20" */
wire imm_a_mux_sel;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17337.7-17337.20" */
/* unused_bits = "0" */
wire imm_a_mux_sel_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17312.14-17312.19" */
wire [31:0] imm_a_t0;
/* src = "generated/sv2v_out.v:17313.13-17313.18" */
wire [31:0] imm_b;
/* src = "generated/sv2v_out.v:17338.13-17338.26" */
wire [2:0] imm_b_mux_sel;
/* src = "generated/sv2v_out.v:17339.13-17339.30" */
wire [2:0] imm_b_mux_sel_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17339.13-17339.30" */
/* unused_bits = "0 1 2" */
wire [2:0] imm_b_mux_sel_dec_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17313.13-17313.18" */
wire [31:0] imm_b_t0;
/* src = "generated/sv2v_out.v:17308.14-17308.24" */
wire [31:0] imm_b_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17308.14-17308.24" */
wire [31:0] imm_b_type_t0;
/* src = "generated/sv2v_out.v:17306.14-17306.24" */
wire [31:0] imm_i_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17306.14-17306.24" */
wire [31:0] imm_i_type_t0;
/* src = "generated/sv2v_out.v:17310.14-17310.24" */
wire [31:0] imm_j_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17310.14-17310.24" */
wire [31:0] imm_j_type_t0;
/* src = "generated/sv2v_out.v:17307.14-17307.24" */
wire [31:0] imm_s_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17307.14-17307.24" */
wire [31:0] imm_s_type_t0;
/* src = "generated/sv2v_out.v:17309.14-17309.24" */
wire [31:0] imm_u_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17309.14-17309.24" */
wire [31:0] imm_u_type_t0;
/* src = "generated/sv2v_out.v:17161.13-17161.29" */
input instr_bp_taken_i;
wire instr_bp_taken_i;
/* cellift = 32'd1 */
input instr_bp_taken_i_t0;
wire instr_bp_taken_i_t0;
/* src = "generated/sv2v_out.v:17166.13-17166.25" */
input instr_exec_i;
wire instr_exec_i;
/* cellift = 32'd1 */
input instr_exec_i_t0;
wire instr_exec_i_t0;
/* src = "generated/sv2v_out.v:17293.7-17293.22" */
wire instr_executing;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17293.7-17293.22" */
wire instr_executing_t0;
/* src = "generated/sv2v_out.v:17176.13-17176.30" */
input instr_fetch_err_i;
wire instr_fetch_err_i;
/* cellift = 32'd1 */
input instr_fetch_err_i_t0;
wire instr_fetch_err_i_t0;
/* src = "generated/sv2v_out.v:17177.13-17177.36" */
input instr_fetch_err_plus2_i;
wire instr_fetch_err_plus2_i;
/* cellift = 32'd1 */
input instr_fetch_err_plus2_i_t0;
wire instr_fetch_err_plus2_i_t0;
/* src = "generated/sv2v_out.v:17163.14-17163.36" */
output instr_first_cycle_id_o;
wire instr_first_cycle_id_o;
/* cellift = 32'd1 */
output instr_first_cycle_id_o_t0;
wire instr_first_cycle_id_o_t0;
/* src = "generated/sv2v_out.v:17268.14-17268.29" */
output instr_id_done_o;
wire instr_id_done_o;
/* cellift = 32'd1 */
output instr_id_done_o_t0;
wire instr_id_done_o_t0;
/* src = "generated/sv2v_out.v:17160.13-17160.34" */
input instr_is_compressed_i;
wire instr_is_compressed_i;
/* cellift = 32'd1 */
input instr_is_compressed_i_t0;
wire instr_is_compressed_i_t0;
/* src = "generated/sv2v_out.v:17258.14-17258.35" */
output instr_perf_count_id_o;
wire instr_perf_count_id_o;
/* cellift = 32'd1 */
output instr_perf_count_id_o_t0;
wire instr_perf_count_id_o_t0;
/* src = "generated/sv2v_out.v:17158.20-17158.37" */
input [31:0] instr_rdata_alu_i;
wire [31:0] instr_rdata_alu_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_alu_i_t0;
wire [31:0] instr_rdata_alu_i_t0;
/* src = "generated/sv2v_out.v:17159.20-17159.35" */
input [15:0] instr_rdata_c_i;
wire [15:0] instr_rdata_c_i;
/* cellift = 32'd1 */
input [15:0] instr_rdata_c_i_t0;
wire [15:0] instr_rdata_c_i_t0;
/* src = "generated/sv2v_out.v:17157.20-17157.33" */
input [31:0] instr_rdata_i;
wire [31:0] instr_rdata_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_i_t0;
wire [31:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:17162.14-17162.25" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:17257.20-17257.35" */
output [1:0] instr_type_wb_o;
wire [1:0] instr_type_wb_o;
/* cellift = 32'd1 */
output [1:0] instr_type_wb_o_t0;
wire [1:0] instr_type_wb_o_t0;
/* src = "generated/sv2v_out.v:17164.14-17164.33" */
output instr_valid_clear_o;
wire instr_valid_clear_o;
/* cellift = 32'd1 */
output instr_valid_clear_o_t0;
wire instr_valid_clear_o_t0;
/* src = "generated/sv2v_out.v:17156.13-17156.26" */
input instr_valid_i;
wire instr_valid_i;
/* cellift = 32'd1 */
input instr_valid_i_t0;
wire instr_valid_i_t0;
/* src = "generated/sv2v_out.v:17223.13-17223.21" */
input irq_nm_i;
wire irq_nm_i;
/* cellift = 32'd1 */
input irq_nm_i_t0;
wire irq_nm_i_t0;
/* src = "generated/sv2v_out.v:17221.13-17221.26" */
input irq_pending_i;
wire irq_pending_i;
/* cellift = 32'd1 */
input irq_pending_i_t0;
wire irq_pending_i_t0;
/* src = "generated/sv2v_out.v:17222.20-17222.26" */
input [17:0] irqs_i;
wire [17:0] irqs_i;
/* cellift = 32'd1 */
input [17:0] irqs_i_t0;
wire [17:0] irqs_i_t0;
/* src = "generated/sv2v_out.v:17287.7-17287.18" */
wire jump_in_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17287.7-17287.18" */
wire jump_in_dec_t0;
/* src = "generated/sv2v_out.v:17289.7-17289.15" */
wire jump_set;
/* src = "generated/sv2v_out.v:17288.7-17288.19" */
wire jump_set_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17288.7-17288.19" */
wire jump_set_dec_t0;
/* src = "generated/sv2v_out.v:17290.6-17290.18" */
wire jump_set_raw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17290.6-17290.18" */
wire jump_set_raw_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17289.7-17289.15" */
wire jump_set_t0;
/* src = "generated/sv2v_out.v:17218.13-17218.32" */
input lsu_addr_incr_req_i;
wire lsu_addr_incr_req_i;
/* cellift = 32'd1 */
input lsu_addr_incr_req_i_t0;
wire lsu_addr_incr_req_i_t0;
/* src = "generated/sv2v_out.v:17219.20-17219.35" */
input [31:0] lsu_addr_last_i;
wire [31:0] lsu_addr_last_i;
/* cellift = 32'd1 */
input [31:0] lsu_addr_last_i_t0;
wire [31:0] lsu_addr_last_i_t0;
/* src = "generated/sv2v_out.v:17225.13-17225.27" */
input lsu_load_err_i;
wire lsu_load_err_i;
/* cellift = 32'd1 */
input lsu_load_err_i_t0;
wire lsu_load_err_i_t0;
/* src = "generated/sv2v_out.v:17226.13-17226.37" */
input lsu_load_resp_intg_err_i;
wire lsu_load_resp_intg_err_i;
/* cellift = 32'd1 */
input lsu_load_resp_intg_err_i_t0;
wire lsu_load_resp_intg_err_i_t0;
/* src = "generated/sv2v_out.v:17351.7-17351.18" */
wire lsu_req_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17351.7-17351.18" */
wire lsu_req_dec_t0;
/* src = "generated/sv2v_out.v:17217.13-17217.27" */
input lsu_req_done_i;
wire lsu_req_done_i;
/* cellift = 32'd1 */
input lsu_req_done_i_t0;
wire lsu_req_done_i_t0;
/* src = "generated/sv2v_out.v:17212.14-17212.23" */
output lsu_req_o;
wire lsu_req_o;
/* cellift = 32'd1 */
output lsu_req_o_t0;
wire lsu_req_o_t0;
/* src = "generated/sv2v_out.v:17180.13-17180.29" */
input lsu_resp_valid_i;
wire lsu_resp_valid_i;
/* cellift = 32'd1 */
input lsu_resp_valid_i_t0;
wire lsu_resp_valid_i_t0;
/* src = "generated/sv2v_out.v:17215.14-17215.28" */
output lsu_sign_ext_o;
wire lsu_sign_ext_o;
/* cellift = 32'd1 */
output lsu_sign_ext_o_t0;
wire lsu_sign_ext_o_t0;
/* src = "generated/sv2v_out.v:17227.13-17227.28" */
input lsu_store_err_i;
wire lsu_store_err_i;
/* cellift = 32'd1 */
input lsu_store_err_i_t0;
wire lsu_store_err_i_t0;
/* src = "generated/sv2v_out.v:17228.13-17228.38" */
input lsu_store_resp_intg_err_i;
wire lsu_store_resp_intg_err_i;
/* cellift = 32'd1 */
input lsu_store_resp_intg_err_i_t0;
wire lsu_store_resp_intg_err_i_t0;
/* src = "generated/sv2v_out.v:17214.20-17214.30" */
output [1:0] lsu_type_o;
wire [1:0] lsu_type_o;
/* cellift = 32'd1 */
output [1:0] lsu_type_o_t0;
wire [1:0] lsu_type_o_t0;
/* src = "generated/sv2v_out.v:17216.21-17216.32" */
output [31:0] lsu_wdata_o;
wire [31:0] lsu_wdata_o;
/* cellift = 32'd1 */
output [31:0] lsu_wdata_o_t0;
wire [31:0] lsu_wdata_o_t0;
/* src = "generated/sv2v_out.v:17213.14-17213.22" */
output lsu_we_o;
wire lsu_we_o;
/* cellift = 32'd1 */
output lsu_we_o_t0;
wire lsu_we_o_t0;
/* src = "generated/sv2v_out.v:17305.7-17305.24" */
wire mem_resp_intg_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17305.7-17305.24" */
wire mem_resp_intg_err_t0;
/* src = "generated/sv2v_out.v:17273.7-17273.20" */
wire mret_insn_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17273.7-17273.20" */
wire mret_insn_dec_t0;
/* src = "generated/sv2v_out.v:17341.7-17341.18" */
wire mult_en_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17341.7-17341.18" */
wire mult_en_dec_t0;
/* src = "generated/sv2v_out.v:17189.14-17189.26" */
output mult_en_ex_o;
wire mult_en_ex_o;
/* cellift = 32'd1 */
output mult_en_ex_o_t0;
wire mult_en_ex_o_t0;
/* src = "generated/sv2v_out.v:17191.14-17191.27" */
output mult_sel_ex_o;
wire mult_sel_ex_o;
/* cellift = 32'd1 */
output mult_sel_ex_o_t0;
wire mult_sel_ex_o_t0;
/* src = "generated/sv2v_out.v:17344.7-17344.21" */
wire multdiv_en_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17344.7-17344.21" */
wire multdiv_en_dec_t0;
/* src = "generated/sv2v_out.v:17195.21-17195.43" */
output [31:0] multdiv_operand_a_ex_o;
wire [31:0] multdiv_operand_a_ex_o;
/* cellift = 32'd1 */
output [31:0] multdiv_operand_a_ex_o_t0;
wire [31:0] multdiv_operand_a_ex_o_t0;
/* src = "generated/sv2v_out.v:17196.21-17196.43" */
output [31:0] multdiv_operand_b_ex_o;
wire [31:0] multdiv_operand_b_ex_o;
/* cellift = 32'd1 */
output [31:0] multdiv_operand_b_ex_o_t0;
wire [31:0] multdiv_operand_b_ex_o_t0;
/* src = "generated/sv2v_out.v:17193.20-17193.41" */
output [1:0] multdiv_operator_ex_o;
wire [1:0] multdiv_operator_ex_o;
/* cellift = 32'd1 */
output [1:0] multdiv_operator_ex_o_t0;
wire [1:0] multdiv_operator_ex_o_t0;
/* src = "generated/sv2v_out.v:17197.14-17197.32" */
output multdiv_ready_id_o;
wire multdiv_ready_id_o;
/* cellift = 32'd1 */
output multdiv_ready_id_o_t0;
wire multdiv_ready_id_o_t0;
/* src = "generated/sv2v_out.v:17194.20-17194.44" */
output [1:0] multdiv_signed_mode_ex_o;
wire [1:0] multdiv_signed_mode_ex_o;
/* cellift = 32'd1 */
output [1:0] multdiv_signed_mode_ex_o_t0;
wire [1:0] multdiv_signed_mode_ex_o_t0;
/* src = "generated/sv2v_out.v:17304.7-17304.22" */
wire multicycle_done;
/* src = "generated/sv2v_out.v:17224.14-17224.24" */
output nmi_mode_o;
wire nmi_mode_o;
/* cellift = 32'd1 */
output nmi_mode_o_t0;
wire nmi_mode_o_t0;
/* src = "generated/sv2v_out.v:17172.21-17172.37" */
output [31:0] nt_branch_addr_o;
wire [31:0] nt_branch_addr_o;
/* cellift = 32'd1 */
output [31:0] nt_branch_addr_o_t0;
wire [31:0] nt_branch_addr_o_t0;
/* src = "generated/sv2v_out.v:17171.14-17171.36" */
output nt_branch_mispredict_o;
wire nt_branch_mispredict_o;
/* cellift = 32'd1 */
output nt_branch_mispredict_o_t0;
wire nt_branch_mispredict_o_t0;
/* src = "generated/sv2v_out.v:17260.13-17260.34" */
input outstanding_load_wb_i;
wire outstanding_load_wb_i;
/* cellift = 32'd1 */
input outstanding_load_wb_i_t0;
wire outstanding_load_wb_i_t0;
/* src = "generated/sv2v_out.v:17261.13-17261.35" */
input outstanding_store_wb_i;
wire outstanding_store_wb_i;
/* cellift = 32'd1 */
input outstanding_store_wb_i_t0;
wire outstanding_store_wb_i_t0;
/* src = "generated/sv2v_out.v:17178.20-17178.27" */
input [31:0] pc_id_i;
wire [31:0] pc_id_i;
/* cellift = 32'd1 */
input [31:0] pc_id_i_t0;
wire [31:0] pc_id_i_t0;
/* src = "generated/sv2v_out.v:17170.20-17170.28" */
output [2:0] pc_mux_o;
wire [2:0] pc_mux_o;
/* cellift = 32'd1 */
output [2:0] pc_mux_o_t0;
wire [2:0] pc_mux_o_t0;
/* src = "generated/sv2v_out.v:17169.14-17169.22" */
output pc_set_o;
wire pc_set_o;
/* cellift = 32'd1 */
output pc_set_o_t0;
wire pc_set_o_t0;
/* src = "generated/sv2v_out.v:17263.13-17263.26" */
output perf_branch_o;
wire perf_branch_o;
/* cellift = 32'd1 */
output perf_branch_o_t0;
wire perf_branch_o_t0;
/* src = "generated/sv2v_out.v:17267.14-17267.29" */
output perf_div_wait_o;
wire perf_div_wait_o;
/* cellift = 32'd1 */
output perf_div_wait_o_t0;
wire perf_div_wait_o_t0;
/* src = "generated/sv2v_out.v:17265.14-17265.31" */
output perf_dside_wait_o;
wire perf_dside_wait_o;
/* cellift = 32'd1 */
output perf_dside_wait_o_t0;
wire perf_dside_wait_o_t0;
/* src = "generated/sv2v_out.v:17262.14-17262.25" */
output perf_jump_o;
wire perf_jump_o;
/* cellift = 32'd1 */
output perf_jump_o_t0;
wire perf_jump_o_t0;
/* src = "generated/sv2v_out.v:17266.14-17266.29" */
output perf_mul_wait_o;
wire perf_mul_wait_o;
/* cellift = 32'd1 */
output perf_mul_wait_o_t0;
wire perf_mul_wait_o_t0;
/* src = "generated/sv2v_out.v:17264.14-17264.28" */
output perf_tbranch_o;
wire perf_tbranch_o;
/* cellift = 32'd1 */
output perf_tbranch_o_t0;
wire perf_tbranch_o_t0;
/* src = "generated/sv2v_out.v:17208.19-17208.30" */
input [1:0] priv_mode_i;
wire [1:0] priv_mode_i;
/* cellift = 32'd1 */
input [1:0] priv_mode_i_t0;
wire [1:0] priv_mode_i_t0;
/* src = "generated/sv2v_out.v:17259.13-17259.23" */
input ready_wb_i;
wire ready_wb_i;
/* cellift = 32'd1 */
input ready_wb_i_t0;
wire ready_wb_i_t0;
/* src = "generated/sv2v_out.v:17240.20-17240.31" */
input [31:0] result_ex_i;
wire [31:0] result_ex_i;
/* cellift = 32'd1 */
input [31:0] result_ex_i_t0;
wire [31:0] result_ex_i_t0;
/* src = "generated/sv2v_out.v:17242.20-17242.32" */
output [4:0] rf_raddr_a_o;
wire [4:0] rf_raddr_a_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_a_o_t0;
wire [4:0] rf_raddr_a_o_t0;
/* src = "generated/sv2v_out.v:17244.20-17244.32" */
output [4:0] rf_raddr_b_o;
wire [4:0] rf_raddr_b_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_b_o_t0;
wire [4:0] rf_raddr_b_o_t0;
/* src = "generated/sv2v_out.v:17251.14-17251.32" */
output rf_rd_a_wb_match_o;
wire rf_rd_a_wb_match_o;
/* cellift = 32'd1 */
output rf_rd_a_wb_match_o_t0;
wire rf_rd_a_wb_match_o_t0;
/* src = "generated/sv2v_out.v:17252.14-17252.32" */
output rf_rd_b_wb_match_o;
wire rf_rd_b_wb_match_o;
/* cellift = 32'd1 */
output rf_rd_b_wb_match_o_t0;
wire rf_rd_b_wb_match_o_t0;
/* src = "generated/sv2v_out.v:17243.20-17243.32" */
input [31:0] rf_rdata_a_i;
wire [31:0] rf_rdata_a_i;
/* cellift = 32'd1 */
input [31:0] rf_rdata_a_i_t0;
wire [31:0] rf_rdata_a_i_t0;
/* src = "generated/sv2v_out.v:17245.20-17245.32" */
input [31:0] rf_rdata_b_i;
wire [31:0] rf_rdata_b_i;
/* cellift = 32'd1 */
input [31:0] rf_rdata_b_i_t0;
wire [31:0] rf_rdata_b_i_t0;
/* src = "generated/sv2v_out.v:17319.7-17319.19" */
wire rf_ren_a_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17319.7-17319.19" */
wire rf_ren_a_dec_t0;
/* src = "generated/sv2v_out.v:17246.14-17246.24" */
output rf_ren_a_o;
wire rf_ren_a_o;
/* cellift = 32'd1 */
output rf_ren_a_o_t0;
wire rf_ren_a_o_t0;
/* src = "generated/sv2v_out.v:17320.7-17320.19" */
wire rf_ren_b_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17320.7-17320.19" */
wire rf_ren_b_dec_t0;
/* src = "generated/sv2v_out.v:17247.14-17247.24" */
output rf_ren_b_o;
wire rf_ren_b_o;
/* cellift = 32'd1 */
output rf_ren_b_o_t0;
wire rf_ren_b_o_t0;
/* src = "generated/sv2v_out.v:17248.20-17248.33" */
output [4:0] rf_waddr_id_o;
wire [4:0] rf_waddr_id_o;
/* cellift = 32'd1 */
output [4:0] rf_waddr_id_o_t0;
wire [4:0] rf_waddr_id_o_t0;
/* src = "generated/sv2v_out.v:17253.19-17253.32" */
input [4:0] rf_waddr_wb_i;
wire [4:0] rf_waddr_wb_i;
/* cellift = 32'd1 */
input [4:0] rf_waddr_wb_i_t0;
wire [4:0] rf_waddr_wb_i_t0;
/* src = "generated/sv2v_out.v:17254.20-17254.37" */
input [31:0] rf_wdata_fwd_wb_i;
wire [31:0] rf_wdata_fwd_wb_i;
/* cellift = 32'd1 */
input [31:0] rf_wdata_fwd_wb_i_t0;
wire [31:0] rf_wdata_fwd_wb_i_t0;
/* src = "generated/sv2v_out.v:17249.20-17249.33" */
output [31:0] rf_wdata_id_o;
wire [31:0] rf_wdata_id_o;
/* cellift = 32'd1 */
output [31:0] rf_wdata_id_o_t0;
wire [31:0] rf_wdata_id_o_t0;
/* src = "generated/sv2v_out.v:17314.7-17314.19" */
wire rf_wdata_sel;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17314.7-17314.19" */
/* unused_bits = "0" */
wire rf_wdata_sel_t0;
/* src = "generated/sv2v_out.v:17315.7-17315.16" */
wire rf_we_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17315.7-17315.16" */
wire rf_we_dec_t0;
/* src = "generated/sv2v_out.v:17250.14-17250.24" */
output rf_we_id_o;
wire rf_we_id_o;
/* cellift = 32'd1 */
output rf_we_id_o_t0;
wire rf_we_id_o_t0;
/* src = "generated/sv2v_out.v:17316.6-17316.15" */
wire rf_we_raw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17316.6-17316.15" */
wire rf_we_raw_t0;
/* src = "generated/sv2v_out.v:17255.13-17255.26" */
input rf_write_wb_i;
wire rf_write_wb_i;
/* cellift = 32'd1 */
input rf_write_wb_i_t0;
wire rf_write_wb_i_t0;
/* src = "generated/sv2v_out.v:17153.13-17153.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:17333.6-17333.15" */
wire stall_alu;
/* src = "generated/sv2v_out.v:17299.6-17299.18" */
wire stall_branch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17299.6-17299.18" */
wire stall_branch_t0;
/* src = "generated/sv2v_out.v:17301.7-17301.15" */
wire stall_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17301.7-17301.15" */
wire stall_id_t0;
/* src = "generated/sv2v_out.v:17300.6-17300.16" */
wire stall_jump;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17300.6-17300.16" */
wire stall_jump_t0;
/* src = "generated/sv2v_out.v:17297.7-17297.16" */
wire stall_mem;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17297.7-17297.16" */
wire stall_mem_t0;
/* src = "generated/sv2v_out.v:17298.6-17298.19" */
wire stall_multdiv;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17298.6-17298.19" */
wire stall_multdiv_t0;
/* src = "generated/sv2v_out.v:17239.13-17239.28" */
input trigger_match_i;
wire trigger_match_i;
/* cellift = 32'd1 */
input trigger_match_i_t0;
wire trigger_match_i_t0;
/* src = "generated/sv2v_out.v:17276.7-17276.19" */
wire wfi_insn_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17276.7-17276.19" */
wire wfi_insn_dec_t0;
/* src = "generated/sv2v_out.v:17311.14-17311.27" */
wire [31:0] zimm_rs1_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17311.14-17311.27" */
wire [31:0] zimm_rs1_type_t0;
assign rf_ren_a_o = _0042_ & /* src = "generated/sv2v_out.v:17321.20-17321.91" */ rf_ren_a_dec;
assign _0042_ = _0040_ & /* src = "generated/sv2v_out.v:17322.21-17322.75" */ _0388_;
assign rf_ren_b_o = _0042_ & /* src = "generated/sv2v_out.v:17322.20-17322.91" */ rf_ren_b_dec;
assign _0044_ = rf_we_raw & /* src = "generated/sv2v_out.v:17436.23-17436.50" */ instr_executing;
assign rf_we_id_o = _0044_ & /* src = "generated/sv2v_out.v:17436.22-17436.73" */ _0105_;
assign illegal_dret_insn = dret_insn_dec & /* src = "generated/sv2v_out.v:17511.29-17511.58" */ _0389_;
assign _0046_ = csr_mstatus_tw_i & /* src = "generated/sv2v_out.v:17512.73-17512.104" */ wfi_insn_dec;
assign illegal_umode_insn = _0386_ & /* src = "generated/sv2v_out.v:17512.30-17512.106" */ _0397_;
assign illegal_insn_o = instr_valid_i & /* src = "generated/sv2v_out.v:17513.26-17513.126" */ _0403_;
assign _0048_ = instr_first_cycle_id_o & /* src = "generated/sv2v_out.v:17587.38-17587.68" */ lsu_req_dec;
assign _0050_ = csr_access_o & /* src = "generated/sv2v_out.v:17595.24-17595.54" */ instr_executing;
assign csr_op_en_o = _0050_ & /* src = "generated/sv2v_out.v:17595.23-17595.73" */ en_wb_o;
assign branch_jump_set_done_d = _0407_ & /* src = "generated/sv2v_out.v:17619.34-17619.115" */ _0390_;
assign jump_set = jump_set_raw & /* src = "generated/sv2v_out.v:17625.20-17625.58" */ _0111_;
assign branch_set = branch_set_raw & /* src = "generated/sv2v_out.v:17626.22-17626.62" */ _0111_;
assign _0052_ = rf_we_dec & /* src = "generated/sv2v_out.v:17703.19-17703.41" */ ex_valid_i;
assign _0054_ = multicycle_done & /* src = "generated/sv2v_out.v:17704.10-17704.38" */ ready_wb_i;
assign _0055_ = _0391_ & /* src = "generated/sv2v_out.v:17717.23-17717.44" */ _0392_;
assign en_wb_o = _0055_ & /* src = "generated/sv2v_out.v:17717.22-17717.63" */ instr_executing;
assign instr_first_cycle_id_o = instr_valid_i & /* src = "generated/sv2v_out.v:17718.29-17718.63" */ _0079_;
assign _0057_ = lsu_req_dec & /* src = "generated/sv2v_out.v:17754.40-17754.93" */ _0417_;
assign stall_mem = instr_valid_i & /* src = "generated/sv2v_out.v:17754.23-17754.94" */ _0057_;
assign _0040_ = instr_valid_i & /* src = "generated/sv2v_out.v:17756.35-17756.69" */ _0387_;
assign instr_executing = _0040_ & /* src = "generated/sv2v_out.v:17756.34-17756.87" */ controller_run;
assign expecting_load_resp_o = _0061_ & /* src = "generated/sv2v_out.v:17762.35-17762.97" */ _0394_;
assign _0059_ = instr_valid_i & /* src = "generated/sv2v_out.v:17763.38-17763.65" */ lsu_req_dec;
assign _0061_ = _0059_ & /* src = "generated/sv2v_out.v:17763.37-17763.87" */ _0118_;
assign expecting_store_resp_o = _0061_ & /* src = "generated/sv2v_out.v:17763.36-17763.97" */ lsu_we_o;
assign _0063_ = instr_executing & /* src = "generated/sv2v_out.v:17782.32-17782.61" */ lsu_req_dec;
assign perf_dside_wait_o = _0063_ & /* src = "generated/sv2v_out.v:17782.31-17782.82" */ _0393_;
assign _0065_ = _0395_ & /* src = "generated/sv2v_out.v:17786.36-17786.64" */ _0396_;
assign _0067_ = _0065_ & /* src = "generated/sv2v_out.v:17786.35-17786.85" */ _0093_;
assign _0069_ = _0067_ & /* src = "generated/sv2v_out.v:17786.34-17786.108" */ _0105_;
assign instr_perf_count_id_o = _0069_ & /* src = "generated/sv2v_out.v:17786.33-17786.130" */ _0387_;
assign perf_mul_wait_o = stall_multdiv & /* src = "generated/sv2v_out.v:17788.27-17788.54" */ mult_en_dec;
assign perf_div_wait_o = stall_multdiv & /* src = "generated/sv2v_out.v:17789.27-17789.53" */ div_en_dec;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME \g_sec_branch_taken.branch_taken_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_sec_branch_taken.branch_taken_q_t0  <= 1'h0;
else \g_sec_branch_taken.branch_taken_q_t0  <= branch_decision_i_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME branch_set_raw_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_set_raw_t0 <= 1'h0;
else branch_set_raw_t0 <= branch_set_raw_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME branch_jump_set_done_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_jump_set_done_q_t0 <= 1'h0;
else branch_jump_set_done_q_t0 <= branch_jump_set_done_d_t0;
assign _0071_ = ~ imd_val_we_ex_i[1];
assign _0073_ = ~ imd_val_we_ex_i[0];
assign _0219_ = { imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1] } & imd_val_d_ex_i_t0[33:0];
assign _0222_ = { imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0] } & imd_val_d_ex_i_t0[67:34];
assign _0220_ = { _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_ } & imd_val_q_ex_o_t0[33:0];
assign _0221_ = _0072_ & id_fsm_q_t0;
assign _0223_ = { _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_, _0073_ } & imd_val_q_ex_o_t0[67:34];
assign _0335_ = _0219_ | _0220_;
assign _0336_ = _0222_ | _0223_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME imd_val_q_ex_o_t0[33:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) imd_val_q_ex_o_t0[33:0] <= 34'h000000000;
else imd_val_q_ex_o_t0[33:0] <= _0335_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME id_fsm_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) id_fsm_q_t0 <= 1'h0;
else id_fsm_q_t0 <= _0221_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME imd_val_q_ex_o_t0[67:34] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) imd_val_q_ex_o_t0[67:34] <= 34'h000000000;
else imd_val_q_ex_o_t0[67:34] <= _0336_;
assign _0120_ = _0043_ & rf_ren_a_dec;
assign _0123_ = _0041_ & _0388_;
assign _0126_ = _0043_ & rf_ren_b_dec;
assign _0129_ = rf_we_raw_t0 & instr_executing;
assign _0132_ = _0045_ & _0105_;
assign _0135_ = dret_insn_dec_t0 & _0389_;
assign _0138_ = csr_mstatus_tw_i_t0 & wfi_insn_dec;
assign _0141_ = instr_valid_i_t0 & _0403_;
assign _0144_ = instr_first_cycle_id_o_t0 & lsu_req_dec;
assign _0147_ = csr_access_o_t0 & instr_executing;
assign _0150_ = _0051_ & en_wb_o;
assign _0153_ = _0408_ & _0390_;
assign _0156_ = jump_set_raw_t0 & _0111_;
assign _0159_ = branch_set_raw_t0 & _0111_;
assign _0029_ = rf_we_dec_t0 & ex_valid_i;
assign _0164_ = stall_id_t0 & _0392_;
assign _0167_ = _0056_ & instr_executing;
assign _0170_ = instr_valid_i_t0 & _0079_;
assign _0173_ = lsu_req_dec_t0 & _0417_;
assign _0176_ = instr_valid_i_t0 & _0057_;
assign _0179_ = instr_valid_i_t0 & _0387_;
assign _0182_ = _0041_ & controller_run;
assign _0185_ = _0062_ & _0394_;
assign _0188_ = instr_valid_i_t0 & lsu_req_dec;
assign _0191_ = _0060_ & _0118_;
assign _0194_ = _0062_ & lsu_we_o;
assign _0195_ = instr_executing_t0 & lsu_req_dec;
assign _0198_ = _0064_ & _0393_;
assign _0201_ = ebrk_insn_t0 & _0396_;
assign _0204_ = _0066_ & _0093_;
assign _0207_ = _0068_ & _0105_;
assign _0210_ = _0070_ & _0387_;
assign _0213_ = stall_multdiv_t0 & mult_en_dec;
assign _0216_ = stall_multdiv_t0 & div_en_dec;
assign _0121_ = rf_ren_a_dec_t0 & _0042_;
assign _0124_ = illegal_insn_o_t0 & _0040_;
assign _0127_ = rf_ren_b_dec_t0 & _0042_;
assign _0130_ = instr_executing_t0 & rf_we_raw;
assign _0133_ = illegal_csr_insn_i_t0 & _0044_;
assign _0136_ = debug_mode_o_t0 & dret_insn_dec;
assign _0139_ = wfi_insn_dec_t0 & csr_mstatus_tw_i;
assign illegal_umode_insn_t0 = _0398_ & _0386_;
assign _0142_ = _0404_ & instr_valid_i;
assign _0145_ = lsu_req_dec_t0 & instr_first_cycle_id_o;
assign _0148_ = instr_executing_t0 & csr_access_o;
assign _0151_ = en_wb_o_t0 & _0050_;
assign _0154_ = instr_valid_clear_o_t0 & _0407_;
assign _0157_ = branch_jump_set_done_q_t0 & jump_set_raw;
assign _0160_ = branch_jump_set_done_q_t0 & branch_set_raw;
assign _0162_ = ex_valid_i_t0 & rf_we_dec;
assign _0165_ = flush_id_t0 & _0391_;
assign _0168_ = instr_executing_t0 & _0055_;
assign _0171_ = id_fsm_q_t0 & instr_valid_i;
assign _0174_ = _0418_ & lsu_req_dec;
assign _0177_ = _0058_ & instr_valid_i;
assign _0180_ = instr_fetch_err_i_t0 & instr_valid_i;
assign _0183_ = controller_run_t0 & _0040_;
assign _0186_ = lsu_we_o_t0 & _0061_;
assign _0189_ = lsu_req_dec_t0 & instr_valid_i;
assign _0192_ = instr_first_cycle_id_o_t0 & _0059_;
assign _0196_ = lsu_req_dec_t0 & instr_executing;
assign _0199_ = lsu_resp_valid_i_t0 & _0063_;
assign _0202_ = ecall_insn_dec_t0 & _0395_;
assign _0205_ = illegal_insn_dec_t0 & _0065_;
assign _0208_ = illegal_csr_insn_i_t0 & _0067_;
assign _0211_ = instr_fetch_err_i_t0 & _0069_;
assign _0214_ = mult_en_dec_t0 & stall_multdiv;
assign _0217_ = div_en_dec_t0 & stall_multdiv;
assign _0122_ = _0043_ & rf_ren_a_dec_t0;
assign _0125_ = _0041_ & illegal_insn_o_t0;
assign _0128_ = _0043_ & rf_ren_b_dec_t0;
assign _0131_ = rf_we_raw_t0 & instr_executing_t0;
assign _0134_ = _0045_ & illegal_csr_insn_i_t0;
assign _0137_ = dret_insn_dec_t0 & debug_mode_o_t0;
assign _0140_ = csr_mstatus_tw_i_t0 & wfi_insn_dec_t0;
assign _0143_ = instr_valid_i_t0 & _0404_;
assign _0146_ = instr_first_cycle_id_o_t0 & lsu_req_dec_t0;
assign _0149_ = csr_access_o_t0 & instr_executing_t0;
assign _0152_ = _0051_ & en_wb_o_t0;
assign _0155_ = _0408_ & instr_valid_clear_o_t0;
assign _0158_ = jump_set_raw_t0 & branch_jump_set_done_q_t0;
assign _0161_ = branch_set_raw_t0 & branch_jump_set_done_q_t0;
assign _0163_ = rf_we_dec_t0 & ex_valid_i_t0;
assign _0166_ = stall_id_t0 & flush_id_t0;
assign _0169_ = _0056_ & instr_executing_t0;
assign _0172_ = instr_valid_i_t0 & id_fsm_q_t0;
assign _0175_ = lsu_req_dec_t0 & _0418_;
assign _0178_ = instr_valid_i_t0 & _0058_;
assign _0181_ = instr_valid_i_t0 & instr_fetch_err_i_t0;
assign _0184_ = _0041_ & controller_run_t0;
assign _0187_ = _0062_ & lsu_we_o_t0;
assign _0190_ = instr_valid_i_t0 & lsu_req_dec_t0;
assign _0193_ = _0060_ & instr_first_cycle_id_o_t0;
assign _0197_ = instr_executing_t0 & lsu_req_dec_t0;
assign _0200_ = _0064_ & lsu_resp_valid_i_t0;
assign _0203_ = ebrk_insn_t0 & ecall_insn_dec_t0;
assign _0206_ = _0066_ & illegal_insn_dec_t0;
assign _0209_ = _0068_ & illegal_csr_insn_i_t0;
assign _0212_ = _0070_ & instr_fetch_err_i_t0;
assign _0215_ = stall_multdiv_t0 & mult_en_dec_t0;
assign _0218_ = stall_multdiv_t0 & div_en_dec_t0;
assign _0301_ = _0120_ | _0121_;
assign _0302_ = _0123_ | _0124_;
assign _0303_ = _0126_ | _0127_;
assign _0304_ = _0129_ | _0130_;
assign _0305_ = _0132_ | _0133_;
assign _0306_ = _0135_ | _0136_;
assign _0307_ = _0138_ | _0139_;
assign _0308_ = _0141_ | _0142_;
assign _0309_ = _0144_ | _0145_;
assign _0310_ = _0147_ | _0148_;
assign _0311_ = _0150_ | _0151_;
assign _0312_ = _0153_ | _0154_;
assign _0313_ = _0156_ | _0157_;
assign _0314_ = _0159_ | _0160_;
assign _0315_ = _0029_ | _0162_;
assign _0316_ = _0164_ | _0165_;
assign _0317_ = _0167_ | _0168_;
assign _0318_ = _0170_ | _0171_;
assign _0319_ = _0173_ | _0174_;
assign _0320_ = _0176_ | _0177_;
assign _0321_ = _0179_ | _0180_;
assign _0322_ = _0182_ | _0183_;
assign _0323_ = _0185_ | _0186_;
assign _0324_ = _0188_ | _0189_;
assign _0325_ = _0191_ | _0192_;
assign _0326_ = _0194_ | _0186_;
assign _0327_ = _0195_ | _0196_;
assign _0328_ = _0198_ | _0199_;
assign _0329_ = _0201_ | _0202_;
assign _0330_ = _0204_ | _0205_;
assign _0331_ = _0207_ | _0208_;
assign _0332_ = _0210_ | _0211_;
assign _0333_ = _0213_ | _0214_;
assign _0334_ = _0216_ | _0217_;
assign rf_ren_a_o_t0 = _0301_ | _0122_;
assign _0043_ = _0302_ | _0125_;
assign rf_ren_b_o_t0 = _0303_ | _0128_;
assign _0045_ = _0304_ | _0131_;
assign rf_we_id_o_t0 = _0305_ | _0134_;
assign illegal_dret_insn_t0 = _0306_ | _0137_;
assign _0047_ = _0307_ | _0140_;
assign illegal_insn_o_t0 = _0308_ | _0143_;
assign _0049_ = _0309_ | _0146_;
assign _0051_ = _0310_ | _0149_;
assign csr_op_en_o_t0 = _0311_ | _0152_;
assign branch_jump_set_done_d_t0 = _0312_ | _0155_;
assign jump_set_t0 = _0313_ | _0158_;
assign branch_set_t0 = _0314_ | _0161_;
assign _0053_ = _0315_ | _0163_;
assign _0056_ = _0316_ | _0166_;
assign en_wb_o_t0 = _0317_ | _0169_;
assign instr_first_cycle_id_o_t0 = _0318_ | _0172_;
assign _0058_ = _0319_ | _0175_;
assign stall_mem_t0 = _0320_ | _0178_;
assign _0041_ = _0321_ | _0181_;
assign instr_executing_t0 = _0322_ | _0184_;
assign expecting_load_resp_o_t0 = _0323_ | _0187_;
assign _0060_ = _0324_ | _0190_;
assign _0062_ = _0325_ | _0193_;
assign expecting_store_resp_o_t0 = _0326_ | _0187_;
assign _0064_ = _0327_ | _0197_;
assign perf_dside_wait_o_t0 = _0328_ | _0200_;
assign _0066_ = _0329_ | _0203_;
assign _0068_ = _0330_ | _0206_;
assign _0070_ = _0331_ | _0209_;
assign instr_perf_count_id_o_t0 = _0332_ | _0212_;
assign perf_mul_wait_o_t0 = _0333_ | _0215_;
assign perf_div_wait_o_t0 = _0334_ | _0218_;
/* src = "generated/sv2v_out.v:17427.4-17432.7" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME imd_val_q_ex_o[33:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) imd_val_q_ex_o[33:0] <= 34'h000000000;
else if (imd_val_we_ex_i[1]) imd_val_q_ex_o[33:0] <= imd_val_d_ex_i[33:0];
/* src = "generated/sv2v_out.v:17649.2-17654.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME id_fsm_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) id_fsm_q <= 1'h0;
else if (instr_executing) id_fsm_q <= id_fsm_d;
/* src = "generated/sv2v_out.v:17427.4-17432.7" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME imd_val_q_ex_o[67:34] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) imd_val_q_ex_o[67:34] <= 34'h000000000;
else if (imd_val_we_ex_i[0]) imd_val_q_ex_o[67:34] <= imd_val_d_ex_i[67:34];
assign _0074_ = ~ { _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_ };
assign _0075_ = ~ { _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_, _0419_ };
assign _0076_ = ~ { _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_ };
assign _0077_ = ~ { _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_ };
assign _0078_ = ~ { _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_ };
assign _0079_ = ~ id_fsm_q;
assign _0080_ = ~ { rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel };
assign _0081_ = ~ { _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_ };
assign _0082_ = ~ { _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_ };
assign _0083_ = ~ { _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_ };
assign _0084_ = ~ _0054_;
assign _0085_ = ~ multdiv_en_dec;
assign _0086_ = ~ alu_multicycle_dec;
assign _0087_ = ~ jump_in_dec;
assign _0088_ = ~ branch_in_dec;
assign _0089_ = ~ lsu_req_dec;
assign _0072_ = ~ instr_executing;
assign _0090_ = ~ { imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel };
assign _0091_ = ~ { alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel };
assign _0224_ = _0074_ & imm_u_type_t0;
assign _0354_ = _0075_ & _0352_;
assign _0226_ = _0076_ & imm_s_type_t0;
assign _0228_ = _0077_ & _0358_;
assign _0230_ = _0078_ & _0360_;
assign _0232_ = _0079_ & _0023_;
assign _0001_ = _0079_ & _0016_;
assign _0004_ = _0079_ & _0020_;
assign _0235_ = _0080_ & result_ex_i_t0;
assign _0237_ = _0081_ & pc_id_i_t0;
assign _0239_ = _0082_ & rf_rdata_a_i_t0;
assign _0241_ = _0083_ & _0364_;
assign _0033_ = _0084_ & jump_in_dec_t0;
assign _0031_ = _0084_ & branch_in_dec_t0;
assign _0038_ = _0084_ & multdiv_en_dec_t0;
assign _0285_ = _0085_ & rf_we_dec_t0;
assign _0433_ = _0086_ & rf_we_dec_t0;
assign _0287_ = _0087_ & _0433_;
assign _0289_ = _0088_ & _0435_;
assign _0291_ = _0085_ & _0437_;
assign _0293_ = _0089_ & _0439_;
assign _0446_ = _0085_ & _0444_;
assign _0016_ = _0089_ & _0446_;
assign _0451_ = _0088_ & _0449_;
assign _0453_ = _0085_ & _0451_;
assign _0020_ = _0089_ & _0453_;
assign _0295_ = _0072_ & rf_we_dec_t0;
assign imm_a_t0 = _0090_ & zimm_rs1_type_t0;
assign _0297_ = _0091_ & rf_rdata_b_i_t0;
assign _0225_ = { _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_ } & imm_j_type_t0;
assign _0227_ = { _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_ } & imm_b_type_t0;
assign _0358_ = { _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_, _0424_ } & imm_i_type_t0;
assign _0229_ = { _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_ } & _0356_;
assign _0231_ = { _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_ } & _0354_;
assign _0233_ = id_fsm_q & _0036_;
assign _0012_ = id_fsm_q & _0033_;
assign _0234_ = id_fsm_q & _0031_;
assign _0014_ = id_fsm_q & _0038_;
assign _0236_ = { rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel } & csr_rdata_i_t0;
assign _0238_ = { _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_ } & imm_a_t0;
assign _0240_ = { _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_ } & lsu_addr_last_i_t0;
assign _0242_ = { _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_ } & _0362_;
assign _0286_ = multdiv_en_dec & _0053_;
assign _0288_ = jump_in_dec & rf_we_dec_t0;
assign _0290_ = branch_in_dec & rf_we_dec_t0;
assign _0292_ = multdiv_en_dec & _0029_;
assign _0294_ = lsu_req_dec & rf_we_dec_t0;
assign _0444_ = branch_in_dec & _0410_;
assign _0449_ = jump_in_dec & jump_set_dec_t0;
assign _0296_ = instr_executing & _0007_;
assign stall_jump_t0 = instr_executing & _0012_;
assign stall_branch_t0 = instr_executing & _0010_;
assign stall_multdiv_t0 = instr_executing & _0014_;
assign jump_set_raw_t0 = instr_executing & _0004_;
assign branch_set_raw_d_t0 = instr_executing & _0001_;
assign _0298_ = { alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel } & imm_b_t0;
assign lsu_req_o_t0 = instr_executing & _0049_;
assign mult_en_ex_o_t0 = instr_executing & mult_en_dec_t0;
assign div_en_ex_o_t0 = instr_executing & div_en_dec_t0;
assign _0352_ = _0224_ | _0225_;
assign _0356_ = _0226_ | _0227_;
assign _0360_ = _0228_ | _0229_;
assign imm_b_t0 = _0230_ | _0231_;
assign _0007_ = _0232_ | _0233_;
assign _0010_ = _0001_ | _0234_;
assign rf_wdata_id_o_t0 = _0235_ | _0236_;
assign _0362_ = _0237_ | _0238_;
assign _0364_ = _0239_ | _0240_;
assign alu_operand_a_ex_o_t0 = _0241_ | _0242_;
assign _0036_ = _0285_ | _0286_;
assign _0435_ = _0287_ | _0288_;
assign _0437_ = _0289_ | _0290_;
assign _0439_ = _0291_ | _0292_;
assign _0023_ = _0293_ | _0294_;
assign rf_we_raw_t0 = _0295_ | _0296_;
assign alu_operand_b_ex_o_t0 = _0297_ | _0298_;
assign _0092_ = ~ mret_insn_dec;
assign _0093_ = ~ illegal_insn_dec;
assign _0094_ = ~ _0399_;
assign _0095_ = ~ _0401_;
assign _0096_ = ~ lsu_load_resp_intg_err_i;
assign _0097_ = ~ mult_en_dec;
assign _0098_ = ~ branch_set_raw;
assign _0099_ = ~ _0405_;
assign _0100_ = ~ branch_decision_i;
assign _0101_ = ~ stall_mem;
assign _0102_ = ~ _0411_;
assign _0103_ = ~ _0413_;
assign _0104_ = ~ _0046_;
assign _0105_ = ~ illegal_csr_insn_i;
assign _0106_ = ~ illegal_dret_insn;
assign _0107_ = ~ illegal_umode_insn;
assign _0108_ = ~ lsu_store_resp_intg_err_i;
assign _0109_ = ~ div_en_dec;
assign _0110_ = ~ jump_set_raw;
assign _0111_ = ~ branch_jump_set_done_q;
assign _0112_ = ~ \g_sec_branch_taken.branch_taken_q ;
assign _0113_ = ~ data_ind_timing_i;
assign _0114_ = ~ stall_multdiv;
assign _0115_ = ~ stall_jump;
assign _0116_ = ~ stall_branch;
assign _0117_ = ~ stall_alu;
assign _0118_ = ~ instr_first_cycle_id_o;
assign _0243_ = mret_insn_dec_t0 & _0104_;
assign _0246_ = illegal_insn_dec_t0 & _0105_;
assign _0249_ = _0400_ & _0106_;
assign _0252_ = _0402_ & _0107_;
assign _0255_ = lsu_load_resp_intg_err_i_t0 & _0108_;
assign _0258_ = mult_en_dec_t0 & _0109_;
assign _0261_ = branch_set_raw_t0 & _0110_;
assign _0264_ = _0406_ & _0111_;
assign _0267_ = data_ind_timing_i_t0 & _0112_;
assign _0270_ = branch_decision_i_t0 & _0113_;
assign _0273_ = stall_mem_t0 & _0114_;
assign _0276_ = _0412_ & _0115_;
assign _0279_ = _0414_ & _0116_;
assign stall_id_t0 = _0416_ & _0117_;
assign _0282_ = lsu_resp_valid_i_t0 & _0118_;
assign _0244_ = _0047_ & _0092_;
assign _0247_ = illegal_csr_insn_i_t0 & _0093_;
assign _0250_ = illegal_dret_insn_t0 & _0094_;
assign _0253_ = illegal_umode_insn_t0 & _0095_;
assign _0256_ = lsu_store_resp_intg_err_i_t0 & _0096_;
assign _0259_ = div_en_dec_t0 & _0097_;
assign _0262_ = jump_set_raw_t0 & _0098_;
assign _0265_ = branch_jump_set_done_q_t0 & _0099_;
assign _0268_ = \g_sec_branch_taken.branch_taken_q_t0  & data_ind_timing_i;
assign _0271_ = data_ind_timing_i_t0 & _0100_;
assign _0274_ = stall_multdiv_t0 & _0101_;
assign _0277_ = stall_jump_t0 & _0102_;
assign _0280_ = stall_branch_t0 & _0103_;
assign _0283_ = instr_first_cycle_id_o_t0 & lsu_resp_valid_i;
assign _0245_ = mret_insn_dec_t0 & _0047_;
assign _0248_ = illegal_insn_dec_t0 & illegal_csr_insn_i_t0;
assign _0251_ = _0400_ & illegal_dret_insn_t0;
assign _0254_ = _0402_ & illegal_umode_insn_t0;
assign _0257_ = lsu_load_resp_intg_err_i_t0 & lsu_store_resp_intg_err_i_t0;
assign _0260_ = mult_en_dec_t0 & div_en_dec_t0;
assign _0263_ = branch_set_raw_t0 & jump_set_raw_t0;
assign _0266_ = _0406_ & branch_jump_set_done_q_t0;
assign _0269_ = data_ind_timing_i_t0 & \g_sec_branch_taken.branch_taken_q_t0 ;
assign _0272_ = branch_decision_i_t0 & data_ind_timing_i_t0;
assign _0275_ = stall_mem_t0 & stall_multdiv_t0;
assign _0278_ = _0412_ & stall_jump_t0;
assign _0281_ = _0414_ & stall_branch_t0;
assign _0284_ = lsu_resp_valid_i_t0 & instr_first_cycle_id_o_t0;
assign _0337_ = _0243_ | _0244_;
assign _0338_ = _0246_ | _0247_;
assign _0339_ = _0249_ | _0250_;
assign _0340_ = _0252_ | _0253_;
assign _0341_ = _0255_ | _0256_;
assign _0342_ = _0258_ | _0259_;
assign _0343_ = _0261_ | _0262_;
assign _0344_ = _0264_ | _0265_;
assign _0345_ = _0267_ | _0268_;
assign _0346_ = _0270_ | _0271_;
assign _0347_ = _0273_ | _0274_;
assign _0348_ = _0276_ | _0277_;
assign _0349_ = _0279_ | _0280_;
assign _0350_ = _0282_ | _0283_;
assign _0398_ = _0337_ | _0245_;
assign _0400_ = _0338_ | _0248_;
assign _0402_ = _0339_ | _0251_;
assign _0404_ = _0340_ | _0254_;
assign mem_resp_intg_err_t0 = _0341_ | _0257_;
assign multdiv_en_dec_t0 = _0342_ | _0260_;
assign _0406_ = _0343_ | _0263_;
assign _0408_ = _0344_ | _0266_;
assign branch_taken_t0 = _0345_ | _0269_;
assign _0410_ = _0346_ | _0272_;
assign _0412_ = _0347_ | _0275_;
assign _0414_ = _0348_ | _0278_;
assign _0416_ = _0349_ | _0281_;
assign _0418_ = _0350_ | _0284_;
assign _0299_ = _0423_ | _0422_;
assign _0300_ = _0457_ | _0456_;
assign _0119_ = | { _0421_, _0420_, _0419_ };
assign _0351_ = _0420_ ? imm_j_type : imm_u_type;
assign _0353_ = _0419_ ? _0459_ : _0351_;
assign _0355_ = _0422_ ? imm_b_type : imm_s_type;
assign _0357_ = _0424_ ? imm_i_type : 32'd4;
assign _0359_ = _0299_ ? _0355_ : _0357_;
assign imm_b = _0119_ ? _0353_ : _0359_;
assign id_fsm_d = id_fsm_q ? _0039_ : _0018_;
assign _0008_ = id_fsm_q ? 1'h0 : _0024_;
assign _0006_ = id_fsm_q ? _0035_ : _0022_;
assign _0011_ = id_fsm_q ? _0032_ : _0025_;
assign _0009_ = id_fsm_q ? _0030_ : _0015_;
assign _0013_ = id_fsm_q ? _0037_ : _0026_;
assign _0003_ = id_fsm_q ? 1'h0 : _0019_;
assign _0000_ = id_fsm_q ? 1'h0 : _0015_;
assign _0005_ = id_fsm_q ? 1'h0 : _0021_;
assign rf_wdata_id_o = rf_wdata_sel ? csr_rdata_i : result_ex_i;
assign _0361_ = _0456_ ? imm_a : pc_id_i;
assign _0363_ = _0458_ ? lsu_addr_last_i : rf_rdata_a_i;
assign alu_operand_a_ex_o = _0300_ ? _0361_ : _0363_;
assign _0365_ = csr_op_o == /* src = "generated/sv2v_out.v:17503.34-17503.50" */ 2'h1;
assign _0366_ = csr_op_o == /* src = "generated/sv2v_out.v:17503.56-17503.72" */ 2'h2;
assign _0367_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17504.11-17504.42" */ 12'h300;
assign _0368_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17504.48-17504.79" */ 12'h304;
assign _0369_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17504.86-17504.117" */ 12'h747;
assign _0370_ = instr_rdata_i[31:25] == /* src = "generated/sv2v_out.v:17504.124-17504.153" */ 7'h1d;
assign _0371_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17508.11-17508.42" */ 12'h7b0;
assign _0372_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17508.48-17508.79" */ 12'h7b1;
assign _0373_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17508.86-17508.117" */ 12'h7b2;
assign _0374_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17508.124-17508.155" */ 12'h7b3;
assign _0375_ = csr_op_en_o && /* src = "generated/sv2v_out.v:17503.7-17503.74" */ _0377_;
assign _0376_ = csr_op_en_o && /* src = "generated/sv2v_out.v:17507.12-17507.55" */ _0385_;
assign _0377_ = _0365_ || /* src = "generated/sv2v_out.v:17503.33-17503.73" */ _0366_;
assign _0378_ = _0367_ || /* src = "generated/sv2v_out.v:17504.10-17504.80" */ _0368_;
assign _0379_ = _0378_ || /* src = "generated/sv2v_out.v:17504.9-17504.118" */ _0369_;
assign _0380_ = _0379_ || /* src = "generated/sv2v_out.v:17504.8-17504.154" */ _0370_;
assign _0381_ = _0371_ || /* src = "generated/sv2v_out.v:17508.10-17508.80" */ _0372_;
assign _0382_ = _0381_ || /* src = "generated/sv2v_out.v:17508.9-17508.118" */ _0373_;
assign _0383_ = _0382_ || /* src = "generated/sv2v_out.v:17508.8-17508.156" */ _0374_;
assign _0384_ = data_ind_timing_i || /* src = "generated/sv2v_out.v:17682.20-17682.80" */ branch_decision_i;
assign _0385_ = | /* src = "generated/sv2v_out.v:17507.38-17507.54" */ csr_op_o;
assign _0386_ = priv_mode_i != /* src = "generated/sv2v_out.v:17512.31-17512.51" */ 2'h3;
assign _0388_ = ~ /* src = "generated/sv2v_out.v:17322.60-17322.75" */ illegal_insn_o;
assign _0389_ = ~ /* src = "generated/sv2v_out.v:17511.45-17511.58" */ debug_mode_o;
assign _0390_ = ~ /* src = "generated/sv2v_out.v:17619.95-17619.115" */ instr_valid_clear_o;
assign _0391_ = ~ /* src = "generated/sv2v_out.v:17717.23-17717.32" */ stall_id;
assign _0392_ = ~ /* src = "generated/sv2v_out.v:17717.35-17717.44" */ flush_id;
assign _0387_ = ~ /* src = "generated/sv2v_out.v:17756.51-17756.69" */ instr_fetch_err_i;
assign _0394_ = ~ /* src = "generated/sv2v_out.v:17762.90-17762.97" */ lsu_we_o;
assign _0393_ = ~ /* src = "generated/sv2v_out.v:17782.65-17782.82" */ lsu_resp_valid_i;
assign _0395_ = ~ /* src = "generated/sv2v_out.v:17786.36-17786.46" */ ebrk_insn;
assign _0396_ = ~ /* src = "generated/sv2v_out.v:17786.49-17786.64" */ ecall_insn_dec;
assign _0397_ = mret_insn_dec | /* src = "generated/sv2v_out.v:17512.56-17512.105" */ _0046_;
assign _0399_ = illegal_insn_dec | /* src = "generated/sv2v_out.v:17513.45-17513.82" */ illegal_csr_insn_i;
assign _0401_ = _0399_ | /* src = "generated/sv2v_out.v:17513.44-17513.103" */ illegal_dret_insn;
assign _0403_ = _0401_ | /* src = "generated/sv2v_out.v:17513.43-17513.125" */ illegal_umode_insn;
assign mem_resp_intg_err = lsu_load_resp_intg_err_i | /* src = "generated/sv2v_out.v:17514.29-17514.81" */ lsu_store_resp_intg_err_i;
assign multdiv_en_dec = mult_en_dec | /* src = "generated/sv2v_out.v:17586.26-17586.50" */ div_en_dec;
assign _0405_ = branch_set_raw | /* src = "generated/sv2v_out.v:17619.36-17619.65" */ jump_set_raw;
assign _0407_ = _0405_ | /* src = "generated/sv2v_out.v:17619.35-17619.91" */ branch_jump_set_done_q;
assign branch_taken = _0113_ | /* src = "generated/sv2v_out.v:17635.26-17635.61" */ \g_sec_branch_taken.branch_taken_q ;
assign _0409_ = branch_decision_i | /* src = "generated/sv2v_out.v:17684.27-17684.64" */ data_ind_timing_i;
assign _0411_ = stall_mem | /* src = "generated/sv2v_out.v:17716.23-17716.64" */ stall_multdiv;
assign _0413_ = _0411_ | /* src = "generated/sv2v_out.v:17716.22-17716.78" */ stall_jump;
assign _0415_ = _0413_ | /* src = "generated/sv2v_out.v:17716.21-17716.94" */ stall_branch;
assign stall_id = _0415_ | /* src = "generated/sv2v_out.v:17716.20-17716.107" */ stall_alu;
assign _0417_ = _0393_ | /* src = "generated/sv2v_out.v:17754.55-17754.92" */ instr_first_cycle_id_o;
/* src = "generated/sv2v_out.v:17630.4-17634.42" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME \g_sec_branch_taken.branch_taken_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_sec_branch_taken.branch_taken_q  <= 1'h0;
else \g_sec_branch_taken.branch_taken_q  <= branch_decision_i;
/* src = "generated/sv2v_out.v:17611.4-17615.43" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME branch_set_raw */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_set_raw <= 1'h0;
else branch_set_raw <= branch_set_raw_d;
/* src = "generated/sv2v_out.v:17620.2-17624.53" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME branch_jump_set_done_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_jump_set_done_q <= 1'h0;
else branch_jump_set_done_q <= branch_jump_set_done_d;
assign _0419_ = imm_b_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17410.5-17419.12" */ 3'h5;
assign _0420_ = imm_b_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17410.5-17419.12" */ 3'h4;
assign _0421_ = imm_b_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17410.5-17419.12" */ 3'h3;
assign _0422_ = imm_b_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17410.5-17419.12" */ 3'h2;
assign _0423_ = imm_b_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17410.5-17419.12" */ 3'h1;
assign _0424_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17410.5-17419.12" */ imm_b_mux_sel;
assign _0039_ = _0054_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17704.10-17704.38|generated/sv2v_out.v:17704.6-17710.9" */ 1'h0 : 1'h1;
assign _0032_ = _0054_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17704.10-17704.38|generated/sv2v_out.v:17704.6-17710.9" */ 1'h0 : jump_in_dec;
assign _0030_ = _0054_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17704.10-17704.38|generated/sv2v_out.v:17704.6-17710.9" */ 1'h0 : branch_in_dec;
assign _0037_ = _0054_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17704.10-17704.38|generated/sv2v_out.v:17704.6-17710.9" */ 1'h0 : multdiv_en_dec;
assign _0035_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17702.10-17702.24|generated/sv2v_out.v:17702.6-17703.42" */ _0052_ : rf_we_dec;
assign _0028_ = ex_valid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17676.12-17676.23|generated/sv2v_out.v:17676.8-17680.11" */ rf_we_dec : 1'h0;
assign _0034_ = ex_valid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17676.12-17676.23|generated/sv2v_out.v:17676.8-17680.11" */ 1'h0 : 1'h1;
assign _0425_ = alu_multicycle_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h1 : 1'h0;
assign _0426_ = jump_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h1 : _0425_;
assign _0427_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ _0460_ : _0426_;
assign _0428_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ _0034_ : _0427_;
assign _0018_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h1 : _0428_;
assign _0429_ = jump_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h0 : _0425_;
assign _0430_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h0 : _0429_;
assign _0431_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h0 : _0430_;
assign _0024_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h0 : _0431_;
assign _0432_ = alu_multicycle_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h0 : rf_we_dec;
assign _0434_ = jump_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ rf_we_dec : _0432_;
assign _0436_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ rf_we_dec : _0434_;
assign _0438_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ _0028_ : _0436_;
assign _0022_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ rf_we_dec : _0438_;
assign _0440_ = jump_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h1 : 1'h0;
assign _0441_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h0 : _0440_;
assign _0442_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h0 : _0441_;
assign _0025_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h0 : _0442_;
assign _0443_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ _0409_ : 1'h0;
assign _0445_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h0 : _0443_;
assign _0015_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h0 : _0445_;
assign _0447_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ _0034_ : 1'h0;
assign _0026_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h0 : _0447_;
assign _0448_ = jump_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ jump_set_dec : 1'h0;
assign _0450_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h0 : _0448_;
assign _0452_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h0 : _0450_;
assign _0019_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h0 : _0452_;
assign _0454_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h1 : 1'h0;
assign _0455_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h0 : _0454_;
assign _0021_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17669.6-17700.13" */ 1'h0 : _0455_;
assign stall_alu = instr_executing ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17666.7-17666.27|generated/sv2v_out.v:17666.3-17713.11" */ _0008_ : 1'h0;
assign rf_we_raw = instr_executing ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17666.7-17666.27|generated/sv2v_out.v:17666.3-17713.11" */ _0006_ : rf_we_dec;
assign stall_jump = instr_executing ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17666.7-17666.27|generated/sv2v_out.v:17666.3-17713.11" */ _0011_ : 1'h0;
assign stall_branch = instr_executing ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17666.7-17666.27|generated/sv2v_out.v:17666.3-17713.11" */ _0009_ : 1'h0;
assign stall_multdiv = instr_executing ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17666.7-17666.27|generated/sv2v_out.v:17666.3-17713.11" */ _0013_ : 1'h0;
assign jump_set_raw = instr_executing ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17666.7-17666.27|generated/sv2v_out.v:17666.3-17713.11" */ _0003_ : 1'h0;
assign branch_set_raw_d = instr_executing ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17666.7-17666.27|generated/sv2v_out.v:17666.3-17713.11" */ _0000_ : 1'h0;
assign perf_branch_o = instr_executing ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17666.7-17666.27|generated/sv2v_out.v:17666.3-17713.11" */ _0005_ : 1'h0;
assign _0027_ = _0383_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17508.8-17508.156|generated/sv2v_out.v:17508.4-17509.27" */ 1'h1 : 1'h0;
assign _0017_ = _0376_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17507.12-17507.55|generated/sv2v_out.v:17507.8-17509.27" */ _0027_ : 1'h0;
assign _0002_ = _0380_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17504.8-17504.154|generated/sv2v_out.v:17504.4-17505.27" */ 1'h1 : 1'h0;
assign csr_pipe_flush = _0375_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17503.7-17503.74|generated/sv2v_out.v:17503.3-17509.27" */ _0002_ : _0017_;
assign _0456_ = alu_op_a_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17361.3-17367.10" */ 2'h3;
assign _0457_ = alu_op_a_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17361.3-17367.10" */ 2'h2;
assign _0458_ = alu_op_a_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17361.3-17367.10" */ 2'h1;
assign alu_op_a_mux_sel = lsu_addr_incr_req_i ? /* src = "generated/sv2v_out.v:17356.29-17356.78" */ 2'h1 : alu_op_a_mux_sel_dec;
assign alu_op_b_mux_sel = lsu_addr_incr_req_i ? /* src = "generated/sv2v_out.v:17357.29-17357.78" */ 1'h1 : alu_op_b_mux_sel_dec;
assign imm_b_mux_sel = lsu_addr_incr_req_i ? /* src = "generated/sv2v_out.v:17358.26-17358.72" */ 3'h6 : imm_b_mux_sel_dec;
assign imm_a = imm_a_mux_sel ? /* src = "generated/sv2v_out.v:17359.18-17359.70" */ 32'd0 : zimm_rs1_type;
assign _0459_ = instr_is_compressed_i ? /* src = "generated/sv2v_out.v:17416.21-17416.72" */ 32'd2 : 32'd4;
assign alu_operand_b_ex_o = alu_op_b_mux_sel ? /* src = "generated/sv2v_out.v:17423.26-17423.75" */ imm_b : rf_rdata_b_i;
assign lsu_req_o = instr_executing ? /* src = "generated/sv2v_out.v:17587.20-17587.75" */ _0048_ : 1'h0;
assign mult_en_ex_o = instr_executing ? /* src = "generated/sv2v_out.v:17588.23-17588.59" */ mult_en_dec : 1'h0;
assign div_en_ex_o = instr_executing ? /* src = "generated/sv2v_out.v:17589.22-17589.57" */ div_en_dec : 1'h0;
assign _0460_ = _0384_ ? /* src = "generated/sv2v_out.v:17682.20-17682.94" */ 1'h1 : 1'h0;
assign multicycle_done = lsu_req_dec ? /* src = "generated/sv2v_out.v:17752.30-17752.73" */ lsu_resp_valid_i : ex_valid_i;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:17519.4-17585.3" */
\$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  controller_i (
.branch_not_set_i(1'h0),
.branch_not_set_i_t0(1'h0),
.branch_set_i(branch_set),
.branch_set_i_t0(branch_set_t0),
.clk_i(clk_i),
.controller_run_o(controller_run),
.controller_run_o_t0(controller_run_t0),
.csr_mstatus_mie_i(csr_mstatus_mie_i),
.csr_mstatus_mie_i_t0(csr_mstatus_mie_i_t0),
.csr_mtval_o(csr_mtval_o),
.csr_mtval_o_t0(csr_mtval_o_t0),
.csr_pipe_flush_i(csr_pipe_flush),
.csr_pipe_flush_i_t0(1'h0),
.csr_restore_dret_id_o(csr_restore_dret_id_o),
.csr_restore_dret_id_o_t0(csr_restore_dret_id_o_t0),
.csr_restore_mret_id_o(csr_restore_mret_id_o),
.csr_restore_mret_id_o_t0(csr_restore_mret_id_o_t0),
.csr_save_cause_o(csr_save_cause_o),
.csr_save_cause_o_t0(csr_save_cause_o_t0),
.csr_save_id_o(csr_save_id_o),
.csr_save_id_o_t0(csr_save_id_o_t0),
.csr_save_if_o(csr_save_if_o),
.csr_save_if_o_t0(csr_save_if_o_t0),
.csr_save_wb_o(csr_save_wb_o),
.csr_save_wb_o_t0(csr_save_wb_o_t0),
.ctrl_busy_o(ctrl_busy_o),
.ctrl_busy_o_t0(ctrl_busy_o_t0),
.debug_cause_o(debug_cause_o),
.debug_cause_o_t0(debug_cause_o_t0),
.debug_csr_save_o(debug_csr_save_o),
.debug_csr_save_o_t0(debug_csr_save_o_t0),
.debug_ebreakm_i(debug_ebreakm_i),
.debug_ebreakm_i_t0(debug_ebreakm_i_t0),
.debug_ebreaku_i(debug_ebreaku_i),
.debug_ebreaku_i_t0(debug_ebreaku_i_t0),
.debug_mode_entering_o(debug_mode_entering_o),
.debug_mode_entering_o_t0(debug_mode_entering_o_t0),
.debug_mode_o(debug_mode_o),
.debug_mode_o_t0(debug_mode_o_t0),
.debug_req_i(debug_req_i),
.debug_req_i_t0(debug_req_i_t0),
.debug_single_step_i(debug_single_step_i),
.debug_single_step_i_t0(debug_single_step_i_t0),
.dret_insn_i(dret_insn_dec),
.dret_insn_i_t0(dret_insn_dec_t0),
.ebrk_insn_i(ebrk_insn),
.ebrk_insn_i_t0(ebrk_insn_t0),
.ecall_insn_i(ecall_insn_dec),
.ecall_insn_i_t0(ecall_insn_dec_t0),
.exc_cause_o(exc_cause_o),
.exc_cause_o_t0(exc_cause_o_t0),
.exc_pc_mux_o(exc_pc_mux_o),
.exc_pc_mux_o_t0(exc_pc_mux_o_t0),
.flush_id_o(flush_id),
.flush_id_o_t0(flush_id_t0),
.id_exception_o(\gen_no_stall_mem.unused_id_exception ),
.id_exception_o_t0(\gen_no_stall_mem.unused_id_exception_t0 ),
.id_in_ready_o(id_in_ready_o),
.id_in_ready_o_t0(id_in_ready_o_t0),
.illegal_insn_i(illegal_insn_o),
.illegal_insn_i_t0(illegal_insn_o_t0),
.instr_bp_taken_i(instr_bp_taken_i),
.instr_bp_taken_i_t0(instr_bp_taken_i_t0),
.instr_compressed_i(instr_rdata_c_i),
.instr_compressed_i_t0(instr_rdata_c_i_t0),
.instr_exec_i(instr_exec_i),
.instr_exec_i_t0(instr_exec_i_t0),
.instr_fetch_err_i(instr_fetch_err_i),
.instr_fetch_err_i_t0(instr_fetch_err_i_t0),
.instr_fetch_err_plus2_i(instr_fetch_err_plus2_i),
.instr_fetch_err_plus2_i_t0(instr_fetch_err_plus2_i_t0),
.instr_i(instr_rdata_i),
.instr_i_t0(instr_rdata_i_t0),
.instr_is_compressed_i(instr_is_compressed_i),
.instr_is_compressed_i_t0(instr_is_compressed_i_t0),
.instr_req_o(instr_req_o),
.instr_req_o_t0(instr_req_o_t0),
.instr_valid_clear_o(instr_valid_clear_o),
.instr_valid_clear_o_t0(instr_valid_clear_o_t0),
.instr_valid_i(instr_valid_i),
.instr_valid_i_t0(instr_valid_i_t0),
.irq_nm_ext_i(irq_nm_i),
.irq_nm_ext_i_t0(irq_nm_i_t0),
.irq_pending_i(irq_pending_i),
.irq_pending_i_t0(irq_pending_i_t0),
.irqs_i(irqs_i),
.irqs_i_t0(irqs_i_t0),
.jump_set_i(jump_set),
.jump_set_i_t0(jump_set_t0),
.load_err_i(lsu_load_err_i),
.load_err_i_t0(lsu_load_err_i_t0),
.lsu_addr_last_i(lsu_addr_last_i),
.lsu_addr_last_i_t0(lsu_addr_last_i_t0),
.mem_resp_intg_err_i(mem_resp_intg_err),
.mem_resp_intg_err_i_t0(mem_resp_intg_err_t0),
.mret_insn_i(mret_insn_dec),
.mret_insn_i_t0(mret_insn_dec_t0),
.nmi_mode_o(nmi_mode_o),
.nmi_mode_o_t0(nmi_mode_o_t0),
.nt_branch_mispredict_o(nt_branch_mispredict_o),
.nt_branch_mispredict_o_t0(nt_branch_mispredict_o_t0),
.pc_id_i(pc_id_i),
.pc_id_i_t0(pc_id_i_t0),
.pc_mux_o(pc_mux_o),
.pc_mux_o_t0(pc_mux_o_t0),
.pc_set_o(pc_set_o),
.pc_set_o_t0(pc_set_o_t0),
.perf_jump_o(perf_jump_o),
.perf_jump_o_t0(perf_jump_o_t0),
.perf_tbranch_o(perf_tbranch_o),
.perf_tbranch_o_t0(perf_tbranch_o_t0),
.priv_mode_i(priv_mode_i),
.priv_mode_i_t0(priv_mode_i_t0),
.ready_wb_i(ready_wb_i),
.ready_wb_i_t0(ready_wb_i_t0),
.rst_ni(rst_ni),
.stall_id_i(stall_id),
.stall_id_i_t0(stall_id_t0),
.stall_wb_i(1'h0),
.stall_wb_i_t0(1'h0),
.store_err_i(lsu_store_err_i),
.store_err_i_t0(lsu_store_err_i_t0),
.trigger_match_i(trigger_match_i),
.trigger_match_i_t0(trigger_match_i_t0),
.wb_exception_o(\gen_no_stall_mem.unused_wb_exception ),
.wb_exception_o_t0(\gen_no_stall_mem.unused_wb_exception_t0 ),
.wfi_insn_i(wfi_insn_dec),
.wfi_insn_i_t0(wfi_insn_dec_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:17449.4-17500.3" */
\$paramod$5ffe4cc9ba21eb548f33468a0c4a93d38de3dae5\ibex_decoder  decoder_i (
.alu_multicycle_o(alu_multicycle_dec),
.alu_multicycle_o_t0(alu_multicycle_dec_t0),
.alu_op_a_mux_sel_o(alu_op_a_mux_sel_dec),
.alu_op_a_mux_sel_o_t0(alu_op_a_mux_sel_dec_t0),
.alu_op_b_mux_sel_o(alu_op_b_mux_sel_dec),
.alu_op_b_mux_sel_o_t0(alu_op_b_mux_sel_dec_t0),
.alu_operator_o(alu_operator_ex_o),
.alu_operator_o_t0(alu_operator_ex_o_t0),
.branch_in_dec_o(branch_in_dec),
.branch_in_dec_o_t0(branch_in_dec_t0),
.branch_taken_i(branch_taken),
.branch_taken_i_t0(branch_taken_t0),
.bt_a_mux_sel_o(bt_a_mux_sel),
.bt_a_mux_sel_o_t0(bt_a_mux_sel_t0),
.bt_b_mux_sel_o(bt_b_mux_sel),
.bt_b_mux_sel_o_t0(bt_b_mux_sel_t0),
.clk_i(clk_i),
.csr_access_o(csr_access_o),
.csr_access_o_t0(csr_access_o_t0),
.csr_op_o(csr_op_o),
.csr_op_o_t0(csr_op_o_t0),
.data_req_o(lsu_req_dec),
.data_req_o_t0(lsu_req_dec_t0),
.data_sign_extension_o(lsu_sign_ext_o),
.data_sign_extension_o_t0(lsu_sign_ext_o_t0),
.data_type_o(lsu_type_o),
.data_type_o_t0(lsu_type_o_t0),
.data_we_o(lsu_we_o),
.data_we_o_t0(lsu_we_o_t0),
.div_en_o(div_en_dec),
.div_en_o_t0(div_en_dec_t0),
.div_sel_o(div_sel_ex_o),
.div_sel_o_t0(div_sel_ex_o_t0),
.dret_insn_o(dret_insn_dec),
.dret_insn_o_t0(dret_insn_dec_t0),
.ebrk_insn_o(ebrk_insn),
.ebrk_insn_o_t0(ebrk_insn_t0),
.ecall_insn_o(ecall_insn_dec),
.ecall_insn_o_t0(ecall_insn_dec_t0),
.icache_inval_o(icache_inval_o),
.icache_inval_o_t0(icache_inval_o_t0),
.illegal_c_insn_i(illegal_c_insn_i),
.illegal_c_insn_i_t0(illegal_c_insn_i_t0),
.illegal_insn_o(illegal_insn_dec),
.illegal_insn_o_t0(illegal_insn_dec_t0),
.imm_a_mux_sel_o(imm_a_mux_sel),
.imm_a_mux_sel_o_t0(imm_a_mux_sel_t0),
.imm_b_mux_sel_o(imm_b_mux_sel_dec),
.imm_b_mux_sel_o_t0(imm_b_mux_sel_dec_t0),
.imm_b_type_o(imm_b_type),
.imm_b_type_o_t0(imm_b_type_t0),
.imm_i_type_o(imm_i_type),
.imm_i_type_o_t0(imm_i_type_t0),
.imm_j_type_o(imm_j_type),
.imm_j_type_o_t0(imm_j_type_t0),
.imm_s_type_o(imm_s_type),
.imm_s_type_o_t0(imm_s_type_t0),
.imm_u_type_o(imm_u_type),
.imm_u_type_o_t0(imm_u_type_t0),
.instr_first_cycle_i(instr_first_cycle_id_o),
.instr_first_cycle_i_t0(instr_first_cycle_id_o_t0),
.instr_rdata_alu_i(instr_rdata_alu_i),
.instr_rdata_alu_i_t0(instr_rdata_alu_i_t0),
.instr_rdata_i(instr_rdata_i),
.instr_rdata_i_t0(instr_rdata_i_t0),
.jump_in_dec_o(jump_in_dec),
.jump_in_dec_o_t0(jump_in_dec_t0),
.jump_set_o(jump_set_dec),
.jump_set_o_t0(jump_set_dec_t0),
.mret_insn_o(mret_insn_dec),
.mret_insn_o_t0(mret_insn_dec_t0),
.mult_en_o(mult_en_dec),
.mult_en_o_t0(mult_en_dec_t0),
.mult_sel_o(mult_sel_ex_o),
.mult_sel_o_t0(mult_sel_ex_o_t0),
.multdiv_operator_o(multdiv_operator_ex_o),
.multdiv_operator_o_t0(multdiv_operator_ex_o_t0),
.multdiv_signed_mode_o(multdiv_signed_mode_ex_o),
.multdiv_signed_mode_o_t0(multdiv_signed_mode_ex_o_t0),
.rf_raddr_a_o(rf_raddr_a_o),
.rf_raddr_a_o_t0(rf_raddr_a_o_t0),
.rf_raddr_b_o(rf_raddr_b_o),
.rf_raddr_b_o_t0(rf_raddr_b_o_t0),
.rf_ren_a_o(rf_ren_a_dec),
.rf_ren_a_o_t0(rf_ren_a_dec_t0),
.rf_ren_b_o(rf_ren_b_dec),
.rf_ren_b_o_t0(rf_ren_b_dec_t0),
.rf_waddr_o(rf_waddr_id_o),
.rf_waddr_o_t0(rf_waddr_id_o_t0),
.rf_wdata_sel_o(rf_wdata_sel),
.rf_wdata_sel_o_t0(rf_wdata_sel_t0),
.rf_we_o(rf_we_dec),
.rf_we_o_t0(rf_we_dec_t0),
.rst_ni(rst_ni),
.wfi_insn_o(wfi_insn_dec),
.wfi_insn_o_t0(wfi_insn_dec_t0),
.zimm_rs1_type_o(zimm_rs1_type),
.zimm_rs1_type_o_t0(zimm_rs1_type_t0)
);
assign bt_a_operand_o = 32'd0;
assign bt_a_operand_o_t0 = 32'd0;
assign bt_b_operand_o = 32'd0;
assign bt_b_operand_o_t0 = 32'd0;
assign instr_id_done_o = en_wb_o;
assign instr_id_done_o_t0 = en_wb_o_t0;
assign instr_type_wb_o = 2'h2;
assign instr_type_wb_o_t0 = 2'h0;
assign lsu_wdata_o = rf_rdata_b_i;
assign lsu_wdata_o_t0 = rf_rdata_b_i_t0;
assign multdiv_operand_a_ex_o = rf_rdata_a_i;
assign multdiv_operand_a_ex_o_t0 = rf_rdata_a_i_t0;
assign multdiv_operand_b_ex_o = rf_rdata_b_i;
assign multdiv_operand_b_ex_o_t0 = rf_rdata_b_i_t0;
assign multdiv_ready_id_o = ready_wb_i;
assign multdiv_ready_id_o_t0 = ready_wb_i_t0;
assign nt_branch_addr_o = 32'd0;
assign nt_branch_addr_o_t0 = 32'd0;
assign perf_branch_o_t0 = 1'h0;
assign rf_rd_a_wb_match_o = 1'h0;
assign rf_rd_a_wb_match_o_t0 = 1'h0;
assign rf_rd_b_wb_match_o = 1'h0;
assign rf_rd_b_wb_match_o_t0 = 1'h0;
endmodule

module \$paramod\ibex_alu\RV32B=s32'00000000000000000000000000000000 (operator_i, operand_a_i, operand_b_i, instr_first_cycle_i, multdiv_operand_a_i, multdiv_operand_b_i, multdiv_sel_i, imd_val_q_i, imd_val_d_o, imd_val_we_o, adder_result_o, adder_result_ext_o, result_o, comparison_result_o, is_equal_result_o, instr_first_cycle_i_t0, imd_val_d_o_t0, imd_val_q_i_t0, imd_val_we_o_t0, operator_i_t0, adder_result_ext_o_t0
, adder_result_o_t0, comparison_result_o_t0, is_equal_result_o_t0, multdiv_operand_a_i_t0, multdiv_operand_b_i_t0, multdiv_sel_i_t0, operand_a_i_t0, operand_b_i_t0, result_o_t0);
/* src = "generated/sv2v_out.v:11397.52-11397.83" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11397.52-11397.83" */
wire _001_;
wire [33:0] _002_;
wire [33:0] _003_;
wire [31:0] _004_;
wire [31:0] _005_;
wire [31:0] _006_;
wire _007_;
wire [31:0] _008_;
wire [31:0] _009_;
wire _010_;
wire [32:0] _011_;
wire [32:0] _012_;
wire [31:0] _013_;
wire [31:0] _014_;
wire [31:0] _015_;
wire _016_;
wire [33:0] _017_;
wire [33:0] _018_;
wire [31:0] _019_;
wire [31:0] _020_;
wire [31:0] _021_;
wire [31:0] _022_;
wire [31:0] _023_;
wire [31:0] _024_;
wire [31:0] _025_;
wire [31:0] _026_;
wire [31:0] _027_;
wire _028_;
wire _029_;
wire [31:0] _030_;
wire [31:0] _031_;
wire [31:0] _032_;
wire [31:0] _033_;
wire [31:0] _034_;
wire [31:0] _035_;
wire _036_;
wire _037_;
wire [32:0] _038_;
wire [32:0] _039_;
wire [32:0] _040_;
wire [32:0] _041_;
wire [32:0] _042_;
wire [32:0] _043_;
wire [31:0] _044_;
wire [31:0] _045_;
wire [31:0] _046_;
wire [31:0] _047_;
wire _048_;
wire _049_;
wire [33:0] _050_;
wire [33:0] _051_;
wire [33:0] _052_;
wire [31:0] _053_;
wire [31:0] _054_;
wire [33:0] _055_;
wire [33:0] _056_;
wire [33:0] _057_;
wire [31:0] _058_;
/* cellift = 32'd1 */
wire [31:0] _059_;
wire [31:0] _060_;
/* cellift = 32'd1 */
wire [31:0] _061_;
wire [31:0] _062_;
/* cellift = 32'd1 */
wire [31:0] _063_;
wire _064_;
/* cellift = 32'd1 */
wire _065_;
wire _066_;
/* src = "generated/sv2v_out.v:11318.23-11318.47" */
wire _067_;
/* src = "generated/sv2v_out.v:11426.23-11426.41" */
wire _068_;
/* src = "generated/sv2v_out.v:11426.46-11426.64" */
wire _069_;
/* src = "generated/sv2v_out.v:11427.24-11427.42" */
wire _070_;
/* src = "generated/sv2v_out.v:11427.47-11427.65" */
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
/* src = "generated/sv2v_out.v:11325.24-11325.33" */
wire _088_;
/* src = "generated/sv2v_out.v:11327.59-11327.76" */
wire _089_;
wire [7:0] _090_;
wire _091_;
wire [4:0] _092_;
wire _093_;
wire [4:0] _094_;
wire _095_;
wire [5:0] _096_;
wire _097_;
wire [31:0] _098_;
/* cellift = 32'd1 */
wire [31:0] _099_;
wire [5:0] _100_;
wire _101_;
wire [3:0] _102_;
wire _103_;
wire _104_;
wire [32:0] _105_;
/* cellift = 32'd1 */
wire [32:0] _106_;
/* src = "generated/sv2v_out.v:11364.27-11364.48" */
/* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] _107_;
/* src = "generated/sv2v_out.v:11317.8-11317.41" */
wire _108_;
/* src = "generated/sv2v_out.v:11320.23-11320.51" */
wire _109_;
/* src = "generated/sv2v_out.v:11265.13-11265.23" */
wire [32:0] adder_in_a;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11265.13-11265.23" */
wire [32:0] adder_in_a_t0;
/* src = "generated/sv2v_out.v:11266.13-11266.23" */
wire [32:0] adder_in_b;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11266.13-11266.23" */
wire [32:0] adder_in_b_t0;
/* src = "generated/sv2v_out.v:11264.6-11264.23" */
wire adder_op_b_negate;
/* src = "generated/sv2v_out.v:11249.21-11249.39" */
output [33:0] adder_result_ext_o;
wire [33:0] adder_result_ext_o;
/* cellift = 32'd1 */
output [33:0] adder_result_ext_o_t0;
wire [33:0] adder_result_ext_o_t0;
/* src = "generated/sv2v_out.v:11248.21-11248.35" */
output [31:0] adder_result_o;
wire [31:0] adder_result_o;
/* cellift = 32'd1 */
output [31:0] adder_result_o_t0;
wire [31:0] adder_result_o_t0;
/* src = "generated/sv2v_out.v:11409.7-11409.18" */
wire bwlogic_and;
/* src = "generated/sv2v_out.v:11412.14-11412.32" */
wire [31:0] bwlogic_and_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11412.14-11412.32" */
wire [31:0] bwlogic_and_result_t0;
/* src = "generated/sv2v_out.v:11408.7-11408.17" */
wire bwlogic_or;
/* src = "generated/sv2v_out.v:11411.14-11411.31" */
wire [31:0] bwlogic_or_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11411.14-11411.31" */
wire [31:0] bwlogic_or_result_t0;
/* src = "generated/sv2v_out.v:11414.13-11414.27" */
wire [31:0] bwlogic_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11414.13-11414.27" */
wire [31:0] bwlogic_result_t0;
/* src = "generated/sv2v_out.v:11413.14-11413.32" */
wire [31:0] bwlogic_xor_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11413.14-11413.32" */
wire [31:0] bwlogic_xor_result_t0;
/* src = "generated/sv2v_out.v:11308.6-11308.16" */
wire cmp_signed;
/* src = "generated/sv2v_out.v:11251.14-11251.33" */
output comparison_result_o;
wire comparison_result_o;
/* cellift = 32'd1 */
output comparison_result_o_t0;
wire comparison_result_o_t0;
/* src = "generated/sv2v_out.v:11246.20-11246.31" */
output [63:0] imd_val_d_o;
wire [63:0] imd_val_d_o;
/* cellift = 32'd1 */
output [63:0] imd_val_d_o_t0;
wire [63:0] imd_val_d_o_t0;
/* src = "generated/sv2v_out.v:11245.20-11245.31" */
input [63:0] imd_val_q_i;
wire [63:0] imd_val_q_i;
/* cellift = 32'd1 */
input [63:0] imd_val_q_i_t0;
wire [63:0] imd_val_q_i_t0;
/* src = "generated/sv2v_out.v:11247.19-11247.31" */
output [1:0] imd_val_we_o;
wire [1:0] imd_val_we_o;
/* cellift = 32'd1 */
output [1:0] imd_val_we_o_t0;
wire [1:0] imd_val_we_o_t0;
/* src = "generated/sv2v_out.v:11241.13-11241.32" */
input instr_first_cycle_i;
wire instr_first_cycle_i;
/* cellift = 32'd1 */
input instr_first_cycle_i_t0;
wire instr_first_cycle_i_t0;
/* src = "generated/sv2v_out.v:11252.14-11252.31" */
output is_equal_result_o;
wire is_equal_result_o;
/* cellift = 32'd1 */
output is_equal_result_o_t0;
wire is_equal_result_o_t0;
/* src = "generated/sv2v_out.v:11307.6-11307.22" */
wire is_greater_equal;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11307.6-11307.22" */
wire is_greater_equal_t0;
/* src = "generated/sv2v_out.v:11242.20-11242.39" */
input [32:0] multdiv_operand_a_i;
wire [32:0] multdiv_operand_a_i;
/* cellift = 32'd1 */
input [32:0] multdiv_operand_a_i_t0;
wire [32:0] multdiv_operand_a_i_t0;
/* src = "generated/sv2v_out.v:11243.20-11243.39" */
input [32:0] multdiv_operand_b_i;
wire [32:0] multdiv_operand_b_i;
/* cellift = 32'd1 */
input [32:0] multdiv_operand_b_i_t0;
wire [32:0] multdiv_operand_b_i_t0;
/* src = "generated/sv2v_out.v:11244.13-11244.26" */
input multdiv_sel_i;
wire multdiv_sel_i;
/* cellift = 32'd1 */
input multdiv_sel_i_t0;
wire multdiv_sel_i_t0;
/* src = "generated/sv2v_out.v:11239.20-11239.31" */
input [31:0] operand_a_i;
wire [31:0] operand_a_i;
/* cellift = 32'd1 */
input [31:0] operand_a_i_t0;
wire [31:0] operand_a_i_t0;
/* src = "generated/sv2v_out.v:11240.20-11240.31" */
input [31:0] operand_b_i;
wire [31:0] operand_b_i;
/* cellift = 32'd1 */
input [31:0] operand_b_i_t0;
wire [31:0] operand_b_i_t0;
/* src = "generated/sv2v_out.v:11254.14-11254.27" */
wire [32:0] operand_b_neg;
/* src = "generated/sv2v_out.v:11238.19-11238.29" */
input [6:0] operator_i;
wire [6:0] operator_i;
/* cellift = 32'd1 */
input [6:0] operator_i_t0;
wire [6:0] operator_i_t0;
/* src = "generated/sv2v_out.v:11250.20-11250.28" */
output [31:0] result_o;
wire [31:0] result_o;
/* cellift = 32'd1 */
output [31:0] result_o_t0;
wire [31:0] result_o_t0;
/* src = "generated/sv2v_out.v:11336.12-11336.21" */
wire [5:0] shift_amt;
/* src = "generated/sv2v_out.v:11337.13-11337.28" */
/* unused_bits = "5" */
wire [5:0] shift_amt_compl;
/* src = "generated/sv2v_out.v:11333.7-11333.18" */
wire shift_arith;
/* src = "generated/sv2v_out.v:11331.6-11331.16" */
wire shift_left;
/* src = "generated/sv2v_out.v:11338.13-11338.26" */
wire [31:0] shift_operand;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11338.13-11338.26" */
wire [31:0] shift_operand_t0;
/* src = "generated/sv2v_out.v:11342.13-11342.25" */
wire [31:0] shift_result;
/* src = "generated/sv2v_out.v:11340.13-11340.29" */
/* unused_bits = "32" */
wire [32:0] shift_result_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11340.13-11340.29" */
/* unused_bits = "32" */
wire [32:0] shift_result_ext_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11342.13-11342.25" */
wire [31:0] shift_result_t0;
assign adder_result_ext_o = { 1'h0, adder_in_a } + /* src = "generated/sv2v_out.v:11303.30-11303.75" */ { 1'h0, adder_in_b };
assign _000_ = shift_arith & /* src = "generated/sv2v_out.v:11397.52-11397.83" */ shift_operand[31];
assign bwlogic_and_result = operand_a_i & /* src = "generated/sv2v_out.v:11424.30-11424.61" */ operand_b_i;
assign _002_ = ~ { 1'h0, adder_in_a_t0 };
assign _003_ = ~ { 1'h0, adder_in_b_t0 };
assign _017_ = { 1'h0, adder_in_a } & _002_;
assign _018_ = { 1'h0, adder_in_b } & _003_;
assign _056_ = _017_ + _018_;
assign _050_ = { 1'h0, adder_in_a } | { 1'h0, adder_in_a_t0 };
assign _051_ = { 1'h0, adder_in_b } | { 1'h0, adder_in_b_t0 };
assign _057_ = _050_ + _051_;
assign _055_ = _056_ ^ _057_;
assign _052_ = _055_ | { 1'h0, adder_in_a_t0 };
assign adder_result_ext_o_t0 = _052_ | { 1'h0, adder_in_b_t0 };
assign _019_ = operand_a_i_t0 & operand_b_i;
assign _001_ = shift_operand_t0[31] & shift_arith;
assign _020_ = operand_b_i_t0 & operand_a_i;
assign _021_ = operand_a_i_t0 & operand_b_i_t0;
assign _053_ = _019_ | _020_;
assign bwlogic_and_result_t0 = _053_ | _021_;
assign _004_ = ~ { _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_ };
assign _005_ = ~ { _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_ };
assign _006_ = ~ { _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_ };
assign _008_ = ~ { bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and };
assign _009_ = ~ { bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or };
assign _010_ = ~ _108_;
assign _011_ = ~ { adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate };
assign _012_ = ~ { multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i };
assign _013_ = ~ { shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left };
assign _022_ = _004_ & shift_result_t0;
assign _024_ = _005_ & _061_;
assign _026_ = _006_ & _063_;
assign _028_ = _007_ & is_greater_equal_t0;
assign _032_ = _008_ & bwlogic_xor_result_t0;
assign _034_ = _009_ & _099_;
assign _036_ = _010_ & adder_result_ext_o_t0[32];
assign _038_ = _011_ & { operand_b_i_t0, 1'h0 };
assign _040_ = _012_ & _106_;
assign _042_ = _012_ & { operand_a_i_t0, 1'h0 };
assign _044_ = _013_ & operand_a_i_t0;
assign _046_ = _013_ & shift_result_ext_t0[31:0];
assign _023_ = { _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_ } & { 31'h00000000, comparison_result_o_t0 };
assign _061_ = { _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_ } & bwlogic_result_t0;
assign _025_ = { _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_ } & adder_result_ext_o_t0[32:1];
assign _027_ = { _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_ } & _059_;
assign _029_ = _101_ & is_greater_equal_t0;
assign comparison_result_o_t0 = _049_ & _065_;
assign _033_ = { bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and } & bwlogic_and_result_t0;
assign _035_ = { bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or } & bwlogic_or_result_t0;
assign _037_ = _108_ & operand_a_i_t0[31];
assign _039_ = { adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate } & { operand_b_i_t0, 1'h0 };
assign _041_ = { multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i } & multdiv_operand_b_i_t0;
assign _043_ = { multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i } & multdiv_operand_a_i_t0;
assign _045_ = { shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left } & { operand_a_i_t0[0], operand_a_i_t0[1], operand_a_i_t0[2], operand_a_i_t0[3], operand_a_i_t0[4], operand_a_i_t0[5], operand_a_i_t0[6], operand_a_i_t0[7], operand_a_i_t0[8], operand_a_i_t0[9], operand_a_i_t0[10], operand_a_i_t0[11], operand_a_i_t0[12], operand_a_i_t0[13], operand_a_i_t0[14], operand_a_i_t0[15], operand_a_i_t0[16], operand_a_i_t0[17], operand_a_i_t0[18], operand_a_i_t0[19], operand_a_i_t0[20], operand_a_i_t0[21], operand_a_i_t0[22], operand_a_i_t0[23], operand_a_i_t0[24], operand_a_i_t0[25], operand_a_i_t0[26], operand_a_i_t0[27], operand_a_i_t0[28], operand_a_i_t0[29], operand_a_i_t0[30], operand_a_i_t0[31] };
assign _047_ = { shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left } & { shift_result_ext_t0[0], shift_result_ext_t0[1], shift_result_ext_t0[2], shift_result_ext_t0[3], shift_result_ext_t0[4], shift_result_ext_t0[5], shift_result_ext_t0[6], shift_result_ext_t0[7], shift_result_ext_t0[8], shift_result_ext_t0[9], shift_result_ext_t0[10], shift_result_ext_t0[11], shift_result_ext_t0[12], shift_result_ext_t0[13], shift_result_ext_t0[14], shift_result_ext_t0[15], shift_result_ext_t0[16], shift_result_ext_t0[17], shift_result_ext_t0[18], shift_result_ext_t0[19], shift_result_ext_t0[20], shift_result_ext_t0[21], shift_result_ext_t0[22], shift_result_ext_t0[23], shift_result_ext_t0[24], shift_result_ext_t0[25], shift_result_ext_t0[26], shift_result_ext_t0[27], shift_result_ext_t0[28], shift_result_ext_t0[29], shift_result_ext_t0[30], shift_result_ext_t0[31] };
assign _059_ = _022_ | _023_;
assign _063_ = _024_ | _025_;
assign result_o_t0 = _026_ | _027_;
assign _065_ = _028_ | _029_;
assign _099_ = _032_ | _033_;
assign bwlogic_result_t0 = _034_ | _035_;
assign is_greater_equal_t0 = _036_ | _037_;
assign _106_ = _038_ | _039_;
assign adder_in_b_t0 = _040_ | _041_;
assign adder_in_a_t0 = _042_ | _043_;
assign shift_operand_t0 = _044_ | _045_;
assign shift_result_t0 = _046_ | _047_;
assign operand_b_neg = ~ { operand_b_i, 1'h0 };
assign _014_ = ~ operand_a_i;
assign _007_ = ~ _101_;
assign _015_ = ~ operand_b_i;
assign _030_ = operand_a_i_t0 & _015_;
assign _031_ = operand_b_i_t0 & _014_;
assign _054_ = _030_ | _031_;
assign bwlogic_or_result_t0 = _054_ | _021_;
assign _048_ = _093_ | _091_;
assign _049_ = _103_ | _101_;
assign _058_ = _091_ ? { 31'h00000000, comparison_result_o } : shift_result;
assign _060_ = _097_ ? bwlogic_result : 32'd0;
assign _062_ = _095_ ? adder_result_ext_o[32:1] : _060_;
assign result_o = _048_ ? _058_ : _062_;
assign _064_ = _101_ ? _089_ : is_greater_equal;
assign _066_ = _090_[1] ? _088_ : is_equal_result_o;
assign comparison_result_o = _049_ ? _064_ : _066_;
assign shift_result_ext_t0 = { _001_, shift_operand_t0 } >>> shift_amt[4:0];
assign bwlogic_xor_result_t0 = operand_a_i_t0 | operand_b_i_t0;
assign is_equal_result_o = ! /* src = "generated/sv2v_out.v:11314.20-11314.72" */ adder_result_ext_o[32:1];
assign _067_ = ~ /* src = "generated/sv2v_out.v:11318.23-11318.47" */ adder_result_ext_o[32];
assign _016_ = operator_i[5] ? _073_ : _072_;
assign _072_ = operator_i[4] ? _075_ : _074_;
assign _073_ = operator_i[4] ? 1'h0 : _076_;
assign _074_ = operator_i[3] ? 1'h0 : _077_;
assign _075_ = operator_i[3] ? _078_ : 1'h0;
assign _076_ = operator_i[3] ? _080_ : _079_;
assign _077_ = operator_i[2] ? 1'h0 : _081_;
assign _078_ = operator_i[2] ? 1'h1 : _082_;
assign _079_ = operator_i[2] ? 1'h0 : _083_;
assign _080_ = operator_i[2] ? _085_ : _084_;
assign _081_ = operator_i[1] ? 1'h0 : _086_;
assign _084_ = operator_i[1] ? _086_ : 1'h0;
assign _085_ = operator_i[1] ? 1'h0 : _087_;
assign _082_ = operator_i[1] ? 1'h1 : _086_;
assign _083_ = operator_i[1] ? _087_ : 1'h1;
assign _086_ = operator_i[0] ? 1'h1 : 1'h0;
assign _087_ = operator_i[0] ? 1'h0 : 1'h1;
assign _088_ = ~ /* src = "generated/sv2v_out.v:11325.24-11325.33" */ is_equal_result_o;
assign _089_ = ~ /* src = "generated/sv2v_out.v:11327.59-11327.76" */ is_greater_equal;
assign bwlogic_or_result = operand_a_i | /* src = "generated/sv2v_out.v:11423.29-11423.60" */ operand_b_i;
assign bwlogic_or = _068_ | /* src = "generated/sv2v_out.v:11426.22-11426.65" */ _069_;
assign bwlogic_and = _070_ | /* src = "generated/sv2v_out.v:11427.23-11427.66" */ _071_;
assign _091_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ _090_;
assign _090_[0] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h1d;
assign _093_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ { _092_[4:3], _092_[1:0], shift_arith };
assign _092_[1] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h09;
assign shift_arith = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h08;
assign _092_[3] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h0c;
assign _092_[4] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h0b;
assign _095_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ _094_;
assign _094_[0] = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ operator_i;
assign _094_[1] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h01;
assign _094_[2] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h16;
assign _094_[3] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h17;
assign _094_[4] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h18;
assign _097_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ { _096_[1:0], _071_, _070_, _069_, _068_ };
assign _096_[0] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h02;
assign _096_[1] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h05;
assign _068_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h03;
assign _069_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h06;
assign _070_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h04;
assign _071_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h07;
assign _098_ = bwlogic_and ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11429.3-11433.10" */ bwlogic_and_result : bwlogic_xor_result;
assign bwlogic_result = bwlogic_or ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11429.3-11433.10" */ bwlogic_or_result : _098_;
assign shift_left = _092_[0] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11372.3-11381.10" */ 1'h1 : 1'h0;
assign _092_[0] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11372.3-11381.10" */ 7'h0a;
assign _101_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ { _100_[3:2], _090_[7:4] };
assign _090_[4] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h19;
assign _090_[5] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h1a;
assign _100_[2] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h1f;
assign _100_[3] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h20;
assign _090_[6] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h2b;
assign _090_[7] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h2c;
assign _103_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ { _102_[3:2], _090_[3:2] };
assign _090_[3] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h1c;
assign _102_[2] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h21;
assign _102_[3] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h22;
assign _090_[1] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h1e;
assign is_greater_equal = _108_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:11317.7-11317.50|generated/sv2v_out.v:11317.3-11320.52" */ _109_ : _067_;
assign cmp_signed = _104_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11310.3-11313.10" */ 1'h1 : 1'h0;
assign _104_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11310.3-11313.10" */ { _102_[2], _100_[2], _090_[6], _090_[4], _090_[2] };
assign _090_[2] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11310.3-11313.10" */ 7'h1b;
assign _105_ = adder_op_b_negate ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11298.3-11302.10" */ operand_b_neg : { operand_b_i, 1'h0 };
assign adder_in_b = multdiv_sel_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11298.3-11302.10" */ multdiv_operand_b_i : _105_;
assign adder_in_a = multdiv_sel_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11289.3-11295.10" */ multdiv_operand_a_i : { operand_a_i, 1'h1 };
assign adder_op_b_negate = operator_i[6] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:11273.3-11286.10" */ 1'h0 : _016_;
assign shift_result_ext = $signed({ _000_, shift_operand }) >>> /* src = "generated/sv2v_out.v:11397.29-11397.120" */ shift_amt[4:0];
assign { _107_[31:6], shift_amt_compl } = 32'd32 - /* src = "generated/sv2v_out.v:11364.27-11364.48" */ operand_b_i[4:0];
assign shift_amt[4:0] = instr_first_cycle_i ? /* src = "generated/sv2v_out.v:11369.22-11369.195" */ operand_b_i[4:0] : shift_amt_compl[4:0];
assign shift_operand = shift_left ? /* src = "generated/sv2v_out.v:11390.21-11390.61" */ { operand_a_i[0], operand_a_i[1], operand_a_i[2], operand_a_i[3], operand_a_i[4], operand_a_i[5], operand_a_i[6], operand_a_i[7], operand_a_i[8], operand_a_i[9], operand_a_i[10], operand_a_i[11], operand_a_i[12], operand_a_i[13], operand_a_i[14], operand_a_i[15], operand_a_i[16], operand_a_i[17], operand_a_i[18], operand_a_i[19], operand_a_i[20], operand_a_i[21], operand_a_i[22], operand_a_i[23], operand_a_i[24], operand_a_i[25], operand_a_i[26], operand_a_i[27], operand_a_i[28], operand_a_i[29], operand_a_i[30], operand_a_i[31] } : operand_a_i;
assign shift_result = shift_left ? /* src = "generated/sv2v_out.v:11406.19-11406.63" */ { shift_result_ext[0], shift_result_ext[1], shift_result_ext[2], shift_result_ext[3], shift_result_ext[4], shift_result_ext[5], shift_result_ext[6], shift_result_ext[7], shift_result_ext[8], shift_result_ext[9], shift_result_ext[10], shift_result_ext[11], shift_result_ext[12], shift_result_ext[13], shift_result_ext[14], shift_result_ext[15], shift_result_ext[16], shift_result_ext[17], shift_result_ext[18], shift_result_ext[19], shift_result_ext[20], shift_result_ext[21], shift_result_ext[22], shift_result_ext[23], shift_result_ext[24], shift_result_ext[25], shift_result_ext[26], shift_result_ext[27], shift_result_ext[28], shift_result_ext[29], shift_result_ext[30], shift_result_ext[31] } : shift_result_ext[31:0];
assign _108_ = operand_a_i[31] ^ /* src = "generated/sv2v_out.v:11317.8-11317.41" */ operand_b_i[31];
assign _109_ = operand_a_i[31] ^ /* src = "generated/sv2v_out.v:11320.23-11320.51" */ cmp_signed;
assign bwlogic_xor_result = operand_a_i ^ /* src = "generated/sv2v_out.v:11425.30-11425.61" */ operand_b_i;
assign _092_[2] = shift_arith;
assign _096_[5:2] = { _071_, _070_, _069_, _068_ };
assign { _100_[5:4], _100_[1:0] } = _090_[7:4];
assign _102_[1:0] = _090_[3:2];
assign _107_[5:0] = shift_amt_compl;
assign adder_result_o = adder_result_ext_o[32:1];
assign adder_result_o_t0 = adder_result_ext_o_t0[32:1];
assign imd_val_d_o = 64'h0000000000000000;
assign imd_val_d_o_t0 = 64'h0000000000000000;
assign imd_val_we_o = 2'h0;
assign imd_val_we_o_t0 = 2'h0;
assign is_equal_result_o_t0 = 1'h0;
assign shift_amt[5] = 1'h0;
endmodule

module \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1 (clk_i, rst_ni, ctrl_busy_o, illegal_insn_i, ecall_insn_i, mret_insn_i, dret_insn_i, wfi_insn_i, ebrk_insn_i, csr_pipe_flush_i, instr_valid_i, instr_i, instr_compressed_i, instr_is_compressed_i, instr_bp_taken_i, instr_fetch_err_i, instr_fetch_err_plus2_i, pc_id_i, instr_valid_clear_o, id_in_ready_o, controller_run_o
, instr_exec_i, instr_req_o, pc_set_o, pc_mux_o, nt_branch_mispredict_o, exc_pc_mux_o, exc_cause_o, lsu_addr_last_i, load_err_i, store_err_i, mem_resp_intg_err_i, wb_exception_o, id_exception_o, branch_set_i, branch_not_set_i, jump_set_i, csr_mstatus_mie_i, irq_pending_i, irqs_i, irq_nm_ext_i, nmi_mode_o
, debug_req_i, debug_cause_o, debug_csr_save_o, debug_mode_o, debug_mode_entering_o, debug_single_step_i, debug_ebreakm_i, debug_ebreaku_i, trigger_match_i, csr_save_if_o, csr_save_id_o, csr_save_wb_o, csr_restore_mret_id_o, csr_restore_dret_id_o, csr_save_cause_o, csr_mtval_o, priv_mode_i, stall_id_i, stall_wb_i, flush_id_o, ready_wb_i
, perf_jump_o, perf_tbranch_o, stall_wb_i_t0, stall_id_i_t0, ready_wb_i_t0, priv_mode_i_t0, perf_tbranch_o_t0, perf_jump_o_t0, pc_set_o_t0, pc_mux_o_t0, debug_ebreaku_i_t0, debug_ebreakm_i_t0, debug_csr_save_o_t0, debug_cause_o_t0, ctrl_busy_o_t0, csr_save_wb_o_t0, csr_save_if_o_t0, csr_save_id_o_t0, csr_save_cause_o_t0, csr_restore_mret_id_o_t0, csr_restore_dret_id_o_t0
, csr_pipe_flush_i_t0, csr_mtval_o_t0, csr_mstatus_mie_i_t0, controller_run_o_t0, branch_set_i_t0, branch_not_set_i_t0, instr_req_o_t0, wfi_insn_i_t0, wb_exception_o_t0, trigger_match_i_t0, store_err_i_t0, pc_id_i_t0, nt_branch_mispredict_o_t0, nmi_mode_o_t0, mret_insn_i_t0, mem_resp_intg_err_i_t0, lsu_addr_last_i_t0, load_err_i_t0, jump_set_i_t0, irqs_i_t0, irq_pending_i_t0
, irq_nm_ext_i_t0, instr_valid_i_t0, instr_valid_clear_o_t0, instr_is_compressed_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_i_t0, instr_exec_i_t0, instr_compressed_i_t0, instr_bp_taken_i_t0, illegal_insn_i_t0, id_in_ready_o_t0, id_exception_o_t0, flush_id_o_t0, exc_pc_mux_o_t0, exc_cause_o_t0, ecall_insn_i_t0, ebrk_insn_i_t0, dret_insn_i_t0, debug_single_step_i_t0, debug_req_i_t0, debug_mode_o_t0
, debug_mode_entering_o_t0, instr_i_t0);
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _000_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _001_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _002_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _003_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _004_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _005_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _006_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _007_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _008_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _009_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _010_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _011_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _012_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _013_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _014_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _015_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _016_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _017_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _018_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _019_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _020_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _021_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _022_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _023_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _024_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _025_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _026_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [1:0] _027_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _028_;
/* src = "generated/sv2v_out.v:12399.4-12411.7" */
wire _029_;
/* src = "generated/sv2v_out.v:12399.4-12411.7" */
wire _030_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _031_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _032_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _033_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _034_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _035_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [2:0] _036_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _037_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _038_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _039_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _040_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _041_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _042_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _043_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _044_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _045_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _046_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _047_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _048_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _049_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _050_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _051_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _052_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _053_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _054_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _055_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _056_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _057_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _058_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [2:0] _059_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _060_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _061_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _062_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _063_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _064_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _065_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _066_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _067_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _068_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _069_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _070_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _071_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _072_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _073_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _074_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [2:0] _075_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _076_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _077_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _078_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _079_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _080_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _081_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _082_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _083_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _084_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _085_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _086_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _087_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _088_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _089_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _090_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _091_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _092_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _093_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _094_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _095_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _096_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _097_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _098_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _099_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _100_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _101_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _102_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _103_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _104_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _105_;
/* src = "generated/sv2v_out.v:12638.49-12638.64" */
wire [31:0] _106_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12638.49-12638.64" */
wire [31:0] _107_;
/* src = "generated/sv2v_out.v:12404.10-12404.38" */
wire _108_;
/* src = "generated/sv2v_out.v:12412.46-12412.108" */
wire _109_;
/* src = "generated/sv2v_out.v:12434.45-12434.80" */
wire _110_;
/* src = "generated/sv2v_out.v:12436.55-12436.86" */
wire _111_;
/* src = "generated/sv2v_out.v:12440.24-12440.60" */
wire _112_;
/* src = "generated/sv2v_out.v:12440.23-12440.75" */
wire _113_;
/* src = "generated/sv2v_out.v:12440.90-12440.117" */
wire _114_;
/* src = "generated/sv2v_out.v:12451.52-12451.86" */
wire _115_;
/* src = "generated/sv2v_out.v:12578.11-12578.37" */
wire _116_;
/* src = "generated/sv2v_out.v:12697.26-12697.43" */
wire _117_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12697.26-12697.43" */
wire _118_;
wire [31:0] _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire [31:0] _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire [31:0] _130_;
wire [31:0] _131_;
wire [31:0] _132_;
wire [31:0] _133_;
wire [31:0] _134_;
wire _135_;
wire _136_;
wire _137_;
wire [31:0] _138_;
wire [31:0] _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire [31:0] _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire [31:0] _177_;
wire [31:0] _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire [31:0] _183_;
wire [31:0] _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire [31:0] _197_;
wire [31:0] _198_;
wire [31:0] _199_;
wire [31:0] _200_;
wire [31:0] _201_;
wire [31:0] _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire [31:0] _207_;
wire [31:0] _208_;
wire [31:0] _209_;
wire [31:0] _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire [31:0] _216_;
wire _217_;
wire _218_;
wire _219_;
wire [31:0] _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire [31:0] _225_;
wire [31:0] _226_;
wire [31:0] _227_;
wire [3:0] _228_;
wire [3:0] _229_;
wire [3:0] _230_;
wire [3:0] _231_;
wire [3:0] _232_;
wire [3:0] _233_;
wire [3:0] _234_;
wire _235_;
wire _236_;
wire _237_;
wire [2:0] _238_;
wire [2:0] _239_;
wire _240_;
wire _241_;
wire _242_;
/* cellift = 32'd1 */
wire _243_;
wire _244_;
wire _245_;
wire [31:0] _246_;
/* cellift = 32'd1 */
wire [31:0] _247_;
wire _248_;
wire _249_;
wire [6:0] _250_;
wire [1:0] _251_;
wire _252_;
/* src = "generated/sv2v_out.v:12437.30-12437.50" */
wire _253_;
/* src = "generated/sv2v_out.v:12437.72-12437.92" */
wire _254_;
/* src = "generated/sv2v_out.v:12557.9-12557.69" */
wire _255_;
/* src = "generated/sv2v_out.v:12559.10-12559.32" */
wire _256_;
/* src = "generated/sv2v_out.v:12559.9-12559.51" */
wire _257_;
/* src = "generated/sv2v_out.v:12576.10-12576.31" */
wire _258_;
/* src = "generated/sv2v_out.v:12610.9-12610.43" */
wire _259_;
/* src = "generated/sv2v_out.v:12682.38-12682.73" */
wire _260_;
/* src = "generated/sv2v_out.v:12682.9-12682.74" */
wire _261_;
/* src = "generated/sv2v_out.v:12404.25-12404.38" */
wire _262_;
/* src = "generated/sv2v_out.v:12559.10-12559.16" */
wire _263_;
/* src = "generated/sv2v_out.v:12559.20-12559.32" */
wire _264_;
/* src = "generated/sv2v_out.v:12559.37-12559.51" */
wire _265_;
/* src = "generated/sv2v_out.v:12576.20-12576.31" */
wire _266_;
/* src = "generated/sv2v_out.v:12610.30-12610.43" */
wire _267_;
/* src = "generated/sv2v_out.v:12682.36-12682.74" */
wire _268_;
/* src = "generated/sv2v_out.v:12524.12-12524.35" */
wire _269_;
/* src = "generated/sv2v_out.v:12524.11-12524.51" */
wire _270_;
/* src = "generated/sv2v_out.v:12524.10-12524.68" */
wire _271_;
/* src = "generated/sv2v_out.v:12524.9-12524.92" */
wire _272_;
/* src = "generated/sv2v_out.v:12549.9-12549.35" */
wire _273_;
/* src = "generated/sv2v_out.v:12557.10-12557.40" */
wire _274_;
/* src = "generated/sv2v_out.v:12557.46-12557.68" */
wire _275_;
/* src = "generated/sv2v_out.v:12623.10-12623.34" */
wire _276_;
/* src = "generated/sv2v_out.v:12623.9-12623.49" */
wire _277_;
/* src = "generated/sv2v_out.v:12335.44-12335.63" */
wire _278_;
/* src = "generated/sv2v_out.v:12582.15-12582.52" */
wire _279_;
/* src = "generated/sv2v_out.v:12342.41-12342.52" */
wire _280_;
/* src = "generated/sv2v_out.v:12398.39-12398.50" */
wire _281_;
/* src = "generated/sv2v_out.v:12412.80-12412.108" */
wire _282_;
/* src = "generated/sv2v_out.v:12440.40-12440.60" */
wire _283_;
/* src = "generated/sv2v_out.v:12697.35-12697.43" */
wire _284_;
/* src = "generated/sv2v_out.v:12698.31-12698.51" */
wire _285_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12698.31-12698.51" */
wire _286_;
/* src = "generated/sv2v_out.v:12336.24-12336.46" */
wire _287_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12336.24-12336.46" */
wire _288_;
/* src = "generated/sv2v_out.v:12336.23-12336.64" */
wire _289_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12336.23-12336.64" */
wire _290_;
/* src = "generated/sv2v_out.v:12336.22-12336.83" */
wire _291_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12336.22-12336.83" */
wire _292_;
/* src = "generated/sv2v_out.v:12340.35-12340.56" */
wire _293_;
/* src = "generated/sv2v_out.v:12340.34-12340.69" */
wire _294_;
/* src = "generated/sv2v_out.v:12435.36-12435.66" */
wire _295_;
/* src = "generated/sv2v_out.v:12440.80-12440.118" */
wire _296_;
/* src = "generated/sv2v_out.v:12646.12-12646.44" */
wire _297_;
wire _298_;
wire [31:0] _299_;
/* cellift = 32'd1 */
wire [31:0] _300_;
wire [31:0] _301_;
/* cellift = 32'd1 */
wire [31:0] _302_;
wire [31:0] _303_;
/* cellift = 32'd1 */
wire [31:0] _304_;
wire [31:0] _305_;
/* cellift = 32'd1 */
wire [31:0] _306_;
wire [31:0] _307_;
/* cellift = 32'd1 */
wire [31:0] _308_;
wire [6:0] _309_;
wire [6:0] _310_;
wire [6:0] _311_;
wire [6:0] _312_;
wire [6:0] _313_;
wire [3:0] _314_;
wire [3:0] _315_;
wire [3:0] _316_;
wire _317_;
wire _318_;
wire _319_;
wire _320_;
wire _321_;
wire _322_;
wire _323_;
wire _324_;
wire _325_;
wire _326_;
wire _327_;
wire _328_;
/* src = "generated/sv2v_out.v:12437.72-12437.117" */
wire _329_;
/* src = "generated/sv2v_out.v:12451.119-12451.149" */
wire [2:0] _330_;
/* src = "generated/sv2v_out.v:12451.97-12451.150" */
wire [2:0] _331_;
/* src = "generated/sv2v_out.v:12451.52-12451.151" */
wire [2:0] _332_;
/* src = "generated/sv2v_out.v:12577.22-12577.87" */
wire [6:0] _333_;
/* src = "generated/sv2v_out.v:12626.22-12626.48" */
wire [1:0] _334_;
/* src = "generated/sv2v_out.v:12638.23-12638.74" */
wire [31:0] _335_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12638.23-12638.74" */
wire [31:0] _336_;
/* src = "generated/sv2v_out.v:12642.23-12642.99" */
wire [31:0] _337_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12642.23-12642.99" */
wire [31:0] _338_;
/* src = "generated/sv2v_out.v:12644.39-12644.119" */
wire [6:0] _339_;
/* src = "generated/sv2v_out.v:12244.13-12244.29" */
input branch_not_set_i;
wire branch_not_set_i;
/* cellift = 32'd1 */
input branch_not_set_i_t0;
wire branch_not_set_i_t0;
/* src = "generated/sv2v_out.v:12243.13-12243.25" */
input branch_set_i;
wire branch_set_i;
/* cellift = 32'd1 */
input branch_set_i_t0;
wire branch_set_i_t0;
/* src = "generated/sv2v_out.v:12209.13-12209.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:12229.13-12229.29" */
output controller_run_o;
wire controller_run_o;
/* cellift = 32'd1 */
output controller_run_o_t0;
wire controller_run_o_t0;
/* src = "generated/sv2v_out.v:12246.13-12246.30" */
input csr_mstatus_mie_i;
wire csr_mstatus_mie_i;
/* cellift = 32'd1 */
input csr_mstatus_mie_i_t0;
wire csr_mstatus_mie_i_t0;
/* src = "generated/sv2v_out.v:12266.20-12266.31" */
output [31:0] csr_mtval_o;
wire [31:0] csr_mtval_o;
/* cellift = 32'd1 */
output [31:0] csr_mtval_o_t0;
wire [31:0] csr_mtval_o_t0;
/* src = "generated/sv2v_out.v:12324.7-12324.21" */
wire csr_pipe_flush;
/* src = "generated/sv2v_out.v:12218.13-12218.29" */
input csr_pipe_flush_i;
wire csr_pipe_flush_i;
/* cellift = 32'd1 */
input csr_pipe_flush_i_t0;
wire csr_pipe_flush_i_t0;
/* src = "generated/sv2v_out.v:12264.13-12264.34" */
output csr_restore_dret_id_o;
wire csr_restore_dret_id_o;
/* cellift = 32'd1 */
output csr_restore_dret_id_o_t0;
wire csr_restore_dret_id_o_t0;
/* src = "generated/sv2v_out.v:12263.13-12263.34" */
output csr_restore_mret_id_o;
wire csr_restore_mret_id_o;
/* cellift = 32'd1 */
output csr_restore_mret_id_o_t0;
wire csr_restore_mret_id_o_t0;
/* src = "generated/sv2v_out.v:12265.13-12265.29" */
output csr_save_cause_o;
wire csr_save_cause_o;
/* cellift = 32'd1 */
output csr_save_cause_o_t0;
wire csr_save_cause_o_t0;
/* src = "generated/sv2v_out.v:12261.13-12261.26" */
output csr_save_id_o;
wire csr_save_id_o;
/* cellift = 32'd1 */
output csr_save_id_o_t0;
wire csr_save_id_o_t0;
/* src = "generated/sv2v_out.v:12260.13-12260.26" */
output csr_save_if_o;
wire csr_save_if_o;
/* cellift = 32'd1 */
output csr_save_if_o_t0;
wire csr_save_if_o_t0;
/* src = "generated/sv2v_out.v:12262.13-12262.26" */
output csr_save_wb_o;
wire csr_save_wb_o;
/* cellift = 32'd1 */
output csr_save_wb_o_t0;
wire csr_save_wb_o_t0;
/* src = "generated/sv2v_out.v:12211.13-12211.24" */
output ctrl_busy_o;
wire ctrl_busy_o;
/* cellift = 32'd1 */
output ctrl_busy_o_t0;
wire ctrl_busy_o_t0;
/* src = "generated/sv2v_out.v:12274.12-12274.23" */
reg [3:0] ctrl_fsm_cs;
/* src = "generated/sv2v_out.v:12275.12-12275.23" */
wire [3:0] ctrl_fsm_ns;
/* src = "generated/sv2v_out.v:12280.13-12280.26" */
wire [2:0] debug_cause_d;
/* src = "generated/sv2v_out.v:12252.20-12252.33" */
output [2:0] debug_cause_o;
reg [2:0] debug_cause_o;
/* cellift = 32'd1 */
output [2:0] debug_cause_o_t0;
wire [2:0] debug_cause_o_t0;
/* src = "generated/sv2v_out.v:12253.13-12253.29" */
output debug_csr_save_o;
wire debug_csr_save_o;
/* cellift = 32'd1 */
output debug_csr_save_o_t0;
wire debug_csr_save_o_t0;
/* src = "generated/sv2v_out.v:12257.13-12257.28" */
input debug_ebreakm_i;
wire debug_ebreakm_i;
/* cellift = 32'd1 */
input debug_ebreakm_i_t0;
wire debug_ebreakm_i_t0;
/* src = "generated/sv2v_out.v:12258.13-12258.28" */
input debug_ebreaku_i;
wire debug_ebreaku_i;
/* cellift = 32'd1 */
input debug_ebreaku_i_t0;
wire debug_ebreaku_i_t0;
/* src = "generated/sv2v_out.v:12279.6-12279.18" */
wire debug_mode_d;
/* src = "generated/sv2v_out.v:12255.13-12255.34" */
output debug_mode_entering_o;
wire debug_mode_entering_o;
/* cellift = 32'd1 */
output debug_mode_entering_o_t0;
wire debug_mode_entering_o_t0;
/* src = "generated/sv2v_out.v:12254.14-12254.26" */
output debug_mode_o;
reg debug_mode_o;
/* cellift = 32'd1 */
output debug_mode_o_t0;
reg debug_mode_o_t0;
/* src = "generated/sv2v_out.v:12251.13-12251.24" */
input debug_req_i;
wire debug_req_i;
/* cellift = 32'd1 */
input debug_req_i_t0;
wire debug_req_i_t0;
/* src = "generated/sv2v_out.v:12256.13-12256.32" */
input debug_single_step_i;
wire debug_single_step_i;
/* cellift = 32'd1 */
input debug_single_step_i_t0;
wire debug_single_step_i_t0;
/* src = "generated/sv2v_out.v:12304.7-12304.23" */
wire do_single_step_d;
/* src = "generated/sv2v_out.v:12305.6-12305.22" */
reg do_single_step_q;
/* src = "generated/sv2v_out.v:12321.7-12321.16" */
wire dret_insn;
/* src = "generated/sv2v_out.v:12215.13-12215.24" */
input dret_insn_i;
wire dret_insn_i;
/* cellift = 32'd1 */
input dret_insn_i_t0;
wire dret_insn_i_t0;
/* src = "generated/sv2v_out.v:12309.7-12309.24" */
wire ebreak_into_debug;
/* src = "generated/sv2v_out.v:12323.7-12323.16" */
wire ebrk_insn;
/* src = "generated/sv2v_out.v:12217.13-12217.24" */
input ebrk_insn_i;
wire ebrk_insn_i;
/* cellift = 32'd1 */
input ebrk_insn_i_t0;
wire ebrk_insn_i_t0;
/* src = "generated/sv2v_out.v:12293.6-12293.20" */
wire ebrk_insn_prio;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12323.7-12323.16" */
wire ebrk_insn_t0;
/* src = "generated/sv2v_out.v:12319.7-12319.17" */
wire ecall_insn;
/* src = "generated/sv2v_out.v:12213.13-12213.25" */
input ecall_insn_i;
wire ecall_insn_i;
/* cellift = 32'd1 */
input ecall_insn_i_t0;
wire ecall_insn_i_t0;
/* src = "generated/sv2v_out.v:12292.6-12292.21" */
wire ecall_insn_prio;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12319.7-12319.17" */
wire ecall_insn_t0;
/* src = "generated/sv2v_out.v:12308.7-12308.23" */
wire enter_debug_mode;
/* src = "generated/sv2v_out.v:12306.7-12306.30" */
wire enter_debug_mode_prio_d;
/* src = "generated/sv2v_out.v:12307.6-12307.29" */
reg enter_debug_mode_prio_q;
/* src = "generated/sv2v_out.v:12236.19-12236.30" */
output [6:0] exc_cause_o;
wire [6:0] exc_cause_o;
/* cellift = 32'd1 */
output [6:0] exc_cause_o_t0;
wire [6:0] exc_cause_o_t0;
/* src = "generated/sv2v_out.v:12235.19-12235.31" */
output [1:0] exc_pc_mux_o;
wire [1:0] exc_pc_mux_o;
/* cellift = 32'd1 */
output [1:0] exc_pc_mux_o_t0;
wire [1:0] exc_pc_mux_o_t0;
/* src = "generated/sv2v_out.v:12300.7-12300.18" */
wire exc_req_lsu;
/* src = "generated/sv2v_out.v:12286.6-12286.15" */
reg exc_req_q;
/* src = "generated/sv2v_out.v:12270.14-12270.24" */
output flush_id_o;
wire flush_id_o;
/* cellift = 32'd1 */
output flush_id_o_t0;
wire flush_id_o_t0;
/* src = "generated/sv2v_out.v:12397.9-12397.21" */
wire \g_intg_irq_int.entering_nmi ;
/* src = "generated/sv2v_out.v:12393.15-12393.39" */
reg [31:0] \g_intg_irq_int.mem_resp_intg_err_addr_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12393.15-12393.39" */
reg [31:0] \g_intg_irq_int.mem_resp_intg_err_addr_q_t0 ;
/* src = "generated/sv2v_out.v:12396.8-12396.35" */
wire \g_intg_irq_int.mem_resp_intg_err_irq_clear ;
/* src = "generated/sv2v_out.v:12392.9-12392.40" */
wire \g_intg_irq_int.mem_resp_intg_err_irq_pending_d ;
/* src = "generated/sv2v_out.v:12391.8-12391.39" */
reg \g_intg_irq_int.mem_resp_intg_err_irq_pending_q ;
/* src = "generated/sv2v_out.v:12395.8-12395.33" */
wire \g_intg_irq_int.mem_resp_intg_err_irq_set ;
/* src = "generated/sv2v_out.v:12297.6-12297.13" */
wire halt_if;
/* src = "generated/sv2v_out.v:12311.7-12311.17" */
wire handle_irq;
/* src = "generated/sv2v_out.v:12242.14-12242.28" */
output id_exception_o;
wire id_exception_o;
/* cellift = 32'd1 */
output id_exception_o_t0;
wire id_exception_o_t0;
/* src = "generated/sv2v_out.v:12228.14-12228.27" */
output id_in_ready_o;
wire id_in_ready_o;
/* cellift = 32'd1 */
output id_in_ready_o_t0;
wire id_in_ready_o_t0;
/* src = "generated/sv2v_out.v:12312.7-12312.20" */
wire id_wb_pending;
/* src = "generated/sv2v_out.v:12289.7-12289.21" */
wire illegal_insn_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12289.7-12289.21" */
wire illegal_insn_d_t0;
/* src = "generated/sv2v_out.v:12212.13-12212.27" */
input illegal_insn_i;
wire illegal_insn_i;
/* cellift = 32'd1 */
input illegal_insn_i_t0;
wire illegal_insn_i_t0;
/* src = "generated/sv2v_out.v:12291.6-12291.23" */
wire illegal_insn_prio;
/* src = "generated/sv2v_out.v:12288.6-12288.20" */
reg illegal_insn_q;
/* src = "generated/sv2v_out.v:12223.13-12223.29" */
input instr_bp_taken_i;
wire instr_bp_taken_i;
/* cellift = 32'd1 */
input instr_bp_taken_i_t0;
wire instr_bp_taken_i_t0;
/* src = "generated/sv2v_out.v:12221.20-12221.38" */
input [15:0] instr_compressed_i;
wire [15:0] instr_compressed_i;
/* cellift = 32'd1 */
input [15:0] instr_compressed_i_t0;
wire [15:0] instr_compressed_i_t0;
/* src = "generated/sv2v_out.v:12230.13-12230.25" */
input instr_exec_i;
wire instr_exec_i;
/* cellift = 32'd1 */
input instr_exec_i_t0;
wire instr_exec_i_t0;
/* src = "generated/sv2v_out.v:12325.7-12325.22" */
wire instr_fetch_err;
/* src = "generated/sv2v_out.v:12224.13-12224.30" */
input instr_fetch_err_i;
wire instr_fetch_err_i;
/* cellift = 32'd1 */
input instr_fetch_err_i_t0;
wire instr_fetch_err_i_t0;
/* src = "generated/sv2v_out.v:12225.13-12225.36" */
input instr_fetch_err_plus2_i;
wire instr_fetch_err_plus2_i;
/* cellift = 32'd1 */
input instr_fetch_err_plus2_i_t0;
wire instr_fetch_err_plus2_i_t0;
/* src = "generated/sv2v_out.v:12290.6-12290.26" */
wire instr_fetch_err_prio;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12325.7-12325.22" */
wire instr_fetch_err_t0;
/* src = "generated/sv2v_out.v:12220.20-12220.27" */
input [31:0] instr_i;
wire [31:0] instr_i;
/* cellift = 32'd1 */
input [31:0] instr_i_t0;
wire [31:0] instr_i_t0;
/* src = "generated/sv2v_out.v:12222.13-12222.34" */
input instr_is_compressed_i;
wire instr_is_compressed_i;
/* cellift = 32'd1 */
input instr_is_compressed_i_t0;
wire instr_is_compressed_i_t0;
/* src = "generated/sv2v_out.v:12231.13-12231.24" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:12227.14-12227.33" */
output instr_valid_clear_o;
wire instr_valid_clear_o;
/* cellift = 32'd1 */
output instr_valid_clear_o_t0;
wire instr_valid_clear_o_t0;
/* src = "generated/sv2v_out.v:12219.13-12219.26" */
input instr_valid_i;
wire instr_valid_i;
/* cellift = 32'd1 */
input instr_valid_i_t0;
wire instr_valid_i_t0;
/* src = "generated/sv2v_out.v:12310.7-12310.18" */
wire irq_enabled;
/* src = "generated/sv2v_out.v:12313.7-12313.13" */
wire irq_nm;
/* src = "generated/sv2v_out.v:12249.13-12249.25" */
input irq_nm_ext_i;
wire irq_nm_ext_i;
/* cellift = 32'd1 */
input irq_nm_ext_i_t0;
wire irq_nm_ext_i_t0;
/* src = "generated/sv2v_out.v:12314.7-12314.17" */
wire irq_nm_int;
/* src = "generated/sv2v_out.v:12247.13-12247.26" */
input irq_pending_i;
wire irq_pending_i;
/* cellift = 32'd1 */
input irq_pending_i_t0;
wire irq_pending_i_t0;
/* src = "generated/sv2v_out.v:12248.20-12248.26" */
input [17:0] irqs_i;
wire [17:0] irqs_i;
/* cellift = 32'd1 */
input [17:0] irqs_i_t0;
wire [17:0] irqs_i_t0;
/* src = "generated/sv2v_out.v:12245.13-12245.23" */
input jump_set_i;
wire jump_set_i;
/* cellift = 32'd1 */
input jump_set_i_t0;
wire jump_set_i_t0;
/* src = "generated/sv2v_out.v:12238.13-12238.23" */
input load_err_i;
wire load_err_i;
/* cellift = 32'd1 */
input load_err_i_t0;
wire load_err_i_t0;
/* src = "generated/sv2v_out.v:12295.6-12295.19" */
wire load_err_prio;
/* src = "generated/sv2v_out.v:12282.6-12282.16" */
reg load_err_q;
/* src = "generated/sv2v_out.v:12237.20-12237.35" */
input [31:0] lsu_addr_last_i;
wire [31:0] lsu_addr_last_i;
/* cellift = 32'd1 */
input [31:0] lsu_addr_last_i_t0;
wire [31:0] lsu_addr_last_i_t0;
/* src = "generated/sv2v_out.v:12240.13-12240.32" */
input mem_resp_intg_err_i;
wire mem_resp_intg_err_i;
/* cellift = 32'd1 */
input mem_resp_intg_err_i_t0;
wire mem_resp_intg_err_i_t0;
/* src = "generated/sv2v_out.v:12317.12-12317.19" */
wire [3:0] mfip_id;
/* src = "generated/sv2v_out.v:12320.7-12320.16" */
wire mret_insn;
/* src = "generated/sv2v_out.v:12214.13-12214.24" */
input mret_insn_i;
wire mret_insn_i;
/* cellift = 32'd1 */
input mret_insn_i_t0;
wire mret_insn_i_t0;
/* src = "generated/sv2v_out.v:12277.6-12277.16" */
wire nmi_mode_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12277.6-12277.16" */
wire nmi_mode_d_t0;
/* src = "generated/sv2v_out.v:12250.14-12250.24" */
output nmi_mode_o;
reg nmi_mode_o;
/* cellift = 32'd1 */
output nmi_mode_o_t0;
reg nmi_mode_o_t0;
/* src = "generated/sv2v_out.v:12234.13-12234.35" */
output nt_branch_mispredict_o;
wire nt_branch_mispredict_o;
/* cellift = 32'd1 */
output nt_branch_mispredict_o_t0;
wire nt_branch_mispredict_o_t0;
/* src = "generated/sv2v_out.v:12226.20-12226.27" */
input [31:0] pc_id_i;
wire [31:0] pc_id_i;
/* cellift = 32'd1 */
input [31:0] pc_id_i_t0;
wire [31:0] pc_id_i_t0;
/* src = "generated/sv2v_out.v:12233.19-12233.27" */
output [2:0] pc_mux_o;
wire [2:0] pc_mux_o;
/* cellift = 32'd1 */
output [2:0] pc_mux_o_t0;
wire [2:0] pc_mux_o_t0;
/* src = "generated/sv2v_out.v:12232.13-12232.21" */
output pc_set_o;
wire pc_set_o;
/* cellift = 32'd1 */
output pc_set_o_t0;
wire pc_set_o_t0;
/* src = "generated/sv2v_out.v:12272.13-12272.24" */
output perf_jump_o;
wire perf_jump_o;
/* cellift = 32'd1 */
output perf_jump_o_t0;
wire perf_jump_o_t0;
/* src = "generated/sv2v_out.v:12273.13-12273.27" */
output perf_tbranch_o;
wire perf_tbranch_o;
/* cellift = 32'd1 */
output perf_tbranch_o_t0;
wire perf_tbranch_o_t0;
/* src = "generated/sv2v_out.v:12267.19-12267.30" */
input [1:0] priv_mode_i;
wire [1:0] priv_mode_i;
/* cellift = 32'd1 */
input [1:0] priv_mode_i_t0;
wire [1:0] priv_mode_i_t0;
/* src = "generated/sv2v_out.v:12271.13-12271.23" */
input ready_wb_i;
wire ready_wb_i;
/* cellift = 32'd1 */
input ready_wb_i_t0;
wire ready_wb_i_t0;
/* src = "generated/sv2v_out.v:12298.6-12298.15" */
wire retain_id;
/* src = "generated/sv2v_out.v:12210.13-12210.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:12301.7-12301.18" */
wire special_req;
/* src = "generated/sv2v_out.v:12303.7-12303.29" */
wire special_req_flush_only;
/* src = "generated/sv2v_out.v:12302.7-12302.28" */
wire special_req_pc_change;
/* src = "generated/sv2v_out.v:12296.7-12296.12" */
wire stall;
/* src = "generated/sv2v_out.v:12268.13-12268.23" */
input stall_id_i;
wire stall_id_i;
/* cellift = 32'd1 */
input stall_id_i_t0;
wire stall_id_i_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12296.7-12296.12" */
wire stall_t0;
/* src = "generated/sv2v_out.v:12269.13-12269.23" */
input stall_wb_i;
wire stall_wb_i;
/* cellift = 32'd1 */
input stall_wb_i_t0;
wire stall_wb_i_t0;
/* src = "generated/sv2v_out.v:12239.13-12239.24" */
input store_err_i;
wire store_err_i;
/* cellift = 32'd1 */
input store_err_i_t0;
wire store_err_i_t0;
/* src = "generated/sv2v_out.v:12294.6-12294.20" */
wire store_err_prio;
/* src = "generated/sv2v_out.v:12284.6-12284.17" */
reg store_err_q;
/* src = "generated/sv2v_out.v:12259.13-12259.28" */
input trigger_match_i;
wire trigger_match_i;
/* cellift = 32'd1 */
input trigger_match_i_t0;
wire trigger_match_i_t0;
/* src = "generated/sv2v_out.v:12241.14-12241.28" */
output wb_exception_o;
wire wb_exception_o;
/* cellift = 32'd1 */
output wb_exception_o_t0;
wire wb_exception_o_t0;
/* src = "generated/sv2v_out.v:12322.7-12322.15" */
wire wfi_insn;
/* src = "generated/sv2v_out.v:12216.13-12216.23" */
input wfi_insn_i;
wire wfi_insn_i;
/* cellift = 32'd1 */
input wfi_insn_i_t0;
wire wfi_insn_i_t0;
assign _106_ = pc_id_i + /* src = "generated/sv2v_out.v:12638.49-12638.64" */ 32'd2;
assign ecall_insn = ecall_insn_i & /* src = "generated/sv2v_out.v:12328.22-12328.50" */ instr_valid_i;
assign mret_insn = mret_insn_i & /* src = "generated/sv2v_out.v:12329.21-12329.48" */ instr_valid_i;
assign dret_insn = dret_insn_i & /* src = "generated/sv2v_out.v:12330.21-12330.48" */ instr_valid_i;
assign wfi_insn = wfi_insn_i & /* src = "generated/sv2v_out.v:12331.20-12331.46" */ instr_valid_i;
assign ebrk_insn = ebrk_insn_i & /* src = "generated/sv2v_out.v:12332.21-12332.48" */ instr_valid_i;
assign csr_pipe_flush = csr_pipe_flush_i & /* src = "generated/sv2v_out.v:12333.26-12333.58" */ instr_valid_i;
assign instr_fetch_err = instr_fetch_err_i & /* src = "generated/sv2v_out.v:12334.27-12334.60" */ instr_valid_i;
assign illegal_insn_d = illegal_insn_i & /* src = "generated/sv2v_out.v:12335.26-12335.64" */ _278_;
assign id_exception_o = _291_ & /* src = "generated/sv2v_out.v:12336.21-12336.108" */ _278_;
assign \g_intg_irq_int.entering_nmi  = nmi_mode_d & /* src = "generated/sv2v_out.v:12398.26-12398.50" */ _281_;
assign _108_ = \g_intg_irq_int.entering_nmi  & /* src = "generated/sv2v_out.v:12404.10-12404.38" */ _262_;
assign _109_ = \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  & /* src = "generated/sv2v_out.v:12412.46-12412.108" */ _282_;
assign _110_ = _142_ & /* src = "generated/sv2v_out.v:12434.45-12434.80" */ debug_single_step_i;
assign enter_debug_mode_prio_d = _295_ & /* src = "generated/sv2v_out.v:12435.35-12435.83" */ _142_;
assign _111_ = trigger_match_i & /* src = "generated/sv2v_out.v:12436.55-12436.86" */ _142_;
assign _112_ = _142_ & /* src = "generated/sv2v_out.v:12440.24-12440.60" */ _283_;
assign _113_ = _112_ & /* src = "generated/sv2v_out.v:12440.23-12440.75" */ _281_;
assign _114_ = irq_pending_i & /* src = "generated/sv2v_out.v:12440.90-12440.117" */ irq_enabled;
assign handle_irq = _113_ & /* src = "generated/sv2v_out.v:12440.22-12440.119" */ _296_;
assign _115_ = ebrk_insn_prio & /* src = "generated/sv2v_out.v:12451.52-12451.86" */ ebreak_into_debug;
assign _116_ = irq_nm_int & /* src = "generated/sv2v_out.v:12578.11-12578.37" */ _262_;
assign _117_ = _144_ & /* src = "generated/sv2v_out.v:12697.26-12697.43" */ _284_;
assign id_in_ready_o = _117_ & /* src = "generated/sv2v_out.v:12697.25-12697.57" */ _148_;
assign _119_ = ~ pc_id_i_t0;
assign _166_ = pc_id_i & _119_;
assign _226_ = _166_ + 32'd2;
assign _216_ = pc_id_i | pc_id_i_t0;
assign _227_ = _216_ + 32'd2;
assign _225_ = _226_ ^ _227_;
assign _107_ = _225_ | pc_id_i_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME nmi_mode_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) nmi_mode_o_t0 <= 1'h0;
else nmi_mode_o_t0 <= nmi_mode_d_t0;
assign _120_ = ~ _158_;
assign _121_ = ~ _160_;
assign _177_ = { _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_, _160_ } & lsu_addr_last_i_t0;
assign _176_ = _120_ & debug_mode_o_t0;
assign _178_ = { _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_, _121_ } & \g_intg_irq_int.mem_resp_intg_err_addr_q_t0 ;
assign _220_ = _177_ | _178_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME debug_mode_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) debug_mode_o_t0 <= 1'h0;
else debug_mode_o_t0 <= _176_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_intg_irq_int.mem_resp_intg_err_addr_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_intg_irq_int.mem_resp_intg_err_addr_q_t0  <= 32'd0;
else \g_intg_irq_int.mem_resp_intg_err_addr_q_t0  <= _220_;
assign _167_ = ecall_insn_i_t0 & instr_valid_i;
assign _170_ = ebrk_insn_i_t0 & instr_valid_i;
assign _173_ = instr_fetch_err_i_t0 & instr_valid_i;
assign illegal_insn_d_t0 = illegal_insn_i_t0 & _278_;
assign id_exception_o_t0 = _292_ & _278_;
assign _118_ = stall_t0 & _284_;
assign id_in_ready_o_t0 = _118_ & _148_;
assign _168_ = instr_valid_i_t0 & ecall_insn_i;
assign _171_ = instr_valid_i_t0 & ebrk_insn_i;
assign _174_ = instr_valid_i_t0 & instr_fetch_err_i;
assign _169_ = ecall_insn_i_t0 & instr_valid_i_t0;
assign _172_ = ebrk_insn_i_t0 & instr_valid_i_t0;
assign _175_ = instr_fetch_err_i_t0 & instr_valid_i_t0;
assign _217_ = _167_ | _168_;
assign _218_ = _170_ | _171_;
assign _219_ = _173_ | _174_;
assign ecall_insn_t0 = _217_ | _169_;
assign ebrk_insn_t0 = _218_ | _172_;
assign instr_fetch_err_t0 = _219_ | _175_;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME debug_mode_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) debug_mode_o <= 1'h0;
else if (_158_) debug_mode_o <= debug_mode_d;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME ctrl_fsm_cs */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) ctrl_fsm_cs <= 4'h0;
else if (_159_) ctrl_fsm_cs <= ctrl_fsm_ns;
/* src = "generated/sv2v_out.v:12413.4-12421.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_intg_irq_int.mem_resp_intg_err_addr_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_intg_irq_int.mem_resp_intg_err_addr_q  <= 32'd0;
else if (_160_) \g_intg_irq_int.mem_resp_intg_err_addr_q  <= lsu_addr_last_i;
assign _124_ = ~ { _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_ };
assign _123_ = ~ _321_;
assign _125_ = ~ \g_intg_irq_int.mem_resp_intg_err_irq_pending_q ;
assign _126_ = ~ ebrk_insn;
assign _127_ = ~ ecall_insn;
assign _128_ = ~ instr_fetch_err;
assign _129_ = ~ mret_insn;
assign _130_ = ~ { store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio };
assign _131_ = ~ { ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio };
assign _132_ = ~ { ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio };
assign _133_ = ~ { illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio };
assign _134_ = ~ { instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio };
assign _135_ = ~ _277_;
assign _136_ = ~ _258_;
assign _137_ = ~ handle_irq;
assign _122_ = ~ _298_;
assign _138_ = ~ { instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i };
assign _139_ = ~ { instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i };
assign _179_ = _123_ & nmi_mode_o_t0;
assign _181_ = _122_ & _243_;
assign _183_ = _124_ & _247_;
assign _086_ = _129_ & nmi_mode_o_t0;
assign _197_ = _130_ & _300_;
assign _304_ = _131_ & _302_;
assign _306_ = _132_ & _304_;
assign _199_ = _133_ & _306_;
assign _201_ = _134_ & _308_;
assign _203_ = _135_ & _086_;
assign _058_ = _136_ & nmi_mode_o_t0;
assign _205_ = _137_ & nmi_mode_o_t0;
assign _207_ = _138_ & pc_id_i_t0;
assign _209_ = _139_ & instr_i_t0;
assign _180_ = _321_ & _035_;
assign _182_ = _298_ & _074_;
assign _247_ = { _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_, _321_ } & _016_;
assign _184_ = { _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_, _298_ } & _079_;
assign _300_ = { load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio } & lsu_addr_last_i_t0;
assign _198_ = { store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio } & lsu_addr_last_i_t0;
assign _200_ = { illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio } & _338_;
assign _202_ = { instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio } & _336_;
assign _079_ = { _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_ } & _089_;
assign _204_ = _277_ & nmi_mode_o_t0;
assign _062_ = { _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_, _116_ } & \g_intg_irq_int.mem_resp_intg_err_addr_q_t0 ;
assign _045_ = { _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_, _258_ } & _062_;
assign _206_ = handle_irq & _058_;
assign _016_ = { handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq } & _045_;
assign _039_ = _273_ & jump_set_i_t0;
assign _041_ = _273_ & branch_set_i_t0;
assign perf_tbranch_o_t0 = _322_ & _041_;
assign perf_jump_o_t0 = _322_ & _039_;
assign _208_ = { instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i } & _107_;
assign _210_ = { instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i } & { 16'h0000, instr_compressed_i_t0 };
assign _243_ = _179_ | _180_;
assign nmi_mode_d_t0 = _181_ | _182_;
assign csr_mtval_o_t0 = _183_ | _184_;
assign _302_ = _197_ | _198_;
assign _308_ = _199_ | _200_;
assign _089_ = _201_ | _202_;
assign _074_ = _203_ | _204_;
assign _035_ = _205_ | _206_;
assign _336_ = _207_ | _208_;
assign _338_ = _209_ | _210_;
assign _152_ = { _298_, _277_, dret_insn, mret_insn } != 4'h8;
assign _153_ = { _298_, _277_, mret_insn } != 3'h5;
assign _154_ = { _298_, _277_ } != 2'h3;
assign _155_ = | { _150_, _298_ };
assign _156_ = { _323_, id_in_ready_o, handle_irq, enter_debug_mode } != 4'h8;
assign _157_ = { _324_, _272_ } != 2'h2;
assign _158_ = & { _155_, _154_, _153_, _152_ };
assign _159_ = & { _156_, _157_ };
assign _160_ = & { _125_, mem_resp_intg_err_i };
assign _161_ = | { _328_, _327_, _325_, _320_ };
assign _162_ = | { _325_, _321_, _320_ };
assign _163_ = | { _326_, _324_, _298_ };
assign _164_ = | { _327_, _325_, _323_, _322_, _321_, _320_, _298_ };
assign _165_ = | { _326_, _325_, _324_, _320_ };
assign _140_ = ~ _287_;
assign _141_ = ~ _289_;
assign _142_ = ~ debug_mode_o;
assign _143_ = ~ stall_id_i;
assign _144_ = ~ stall;
assign _146_ = ~ illegal_insn_d;
assign _147_ = ~ stall_wb_i;
assign _148_ = ~ retain_id;
assign _149_ = ~ flush_id_o;
assign _185_ = ecall_insn_t0 & _126_;
assign _188_ = _288_ & _146_;
assign _191_ = _290_ & _128_;
assign _194_ = stall_id_i_t0 & _147_;
assign _286_ = stall_t0 & _148_;
assign instr_valid_clear_o_t0 = _286_ & _149_;
assign _186_ = ebrk_insn_t0 & _127_;
assign _189_ = illegal_insn_d_t0 & _140_;
assign _192_ = instr_fetch_err_t0 & _141_;
assign _195_ = stall_wb_i_t0 & _143_;
assign _187_ = ecall_insn_t0 & ebrk_insn_t0;
assign _190_ = _288_ & illegal_insn_d_t0;
assign _193_ = _290_ & instr_fetch_err_t0;
assign _196_ = stall_id_i_t0 & stall_wb_i_t0;
assign _221_ = _185_ | _186_;
assign _222_ = _188_ | _189_;
assign _223_ = _191_ | _192_;
assign _224_ = _194_ | _195_;
assign _288_ = _221_ | _187_;
assign _290_ = _222_ | _190_;
assign _292_ = _223_ | _193_;
assign stall_t0 = _224_ | _196_;
assign _150_ = | { _325_, _320_ };
assign _212_ = _326_ | _324_;
assign _213_ = _161_ | _298_;
assign _211_ = _162_ | _298_;
assign _214_ = _322_ | _163_;
assign _215_ = _320_ | _298_;
assign _151_ = | { _323_, _322_, _211_ };
assign _228_ = _298_ ? _012_ : 4'h5;
assign _229_ = _322_ ? _100_ : _080_;
assign _230_ = _211_ ? _228_ : _229_;
assign _231_ = _324_ ? _022_ : 4'h3;
assign _232_ = _328_ ? 4'h1 : 4'h0;
assign _233_ = _327_ ? 4'h4 : _232_;
assign _234_ = _212_ ? _231_ : _233_;
assign ctrl_fsm_ns = _151_ ? _230_ : _234_;
assign _235_ = _298_ ? _076_ : 1'h1;
assign _236_ = _322_ ? _037_ : 1'h0;
assign _237_ = _321_ ? _019_ : _236_;
assign pc_set_o = _213_ ? _235_ : _237_;
assign _238_ = _298_ ? _036_ : 3'h2;
assign _239_ = _322_ ? 3'h1 : 3'h0;
assign pc_mux_o = _211_ ? _238_ : _239_;
assign _240_ = _163_ ? 1'h1 : _082_;
assign _241_ = _323_ ? _054_ : 1'h0;
assign _013_ = _214_ ? _240_ : _241_;
assign debug_mode_d = _298_ ? _023_ : 1'h1;
assign _242_ = _321_ ? _034_ : nmi_mode_o;
assign nmi_mode_d = _298_ ? _073_ : _242_;
assign _244_ = _165_ ? 1'h1 : 1'h0;
assign flush_id_o = _298_ ? _028_ : _244_;
assign _245_ = _325_ ? 1'h1 : 1'h0;
assign debug_csr_save_o = _320_ ? _020_ : _245_;
assign _246_ = _321_ ? _015_ : 32'd0;
assign csr_mtval_o = _298_ ? _078_ : _246_;
assign _248_ = _298_ ? _064_ : _020_;
assign csr_save_if_o = _325_ ? 1'h1 : _249_;
assign csr_save_cause_o = _215_ ? _248_ : csr_save_if_o;
assign _249_ = _321_ ? _019_ : 1'h0;
assign _250_ = _321_ ? _026_ : 7'h00;
assign exc_cause_o = _298_ ? _096_ : _250_;
assign _251_ = _150_ ? 2'h2 : 2'h1;
assign exc_pc_mux_o = _298_ ? _027_ : _251_;
assign _252_ = _326_ ? 1'h0 : 1'h1;
assign ctrl_busy_o = _324_ ? _021_ : _252_;
assign _254_ = ! /* src = "generated/sv2v_out.v:12439.44-12439.64" */ priv_mode_i;
assign _253_ = priv_mode_i == /* src = "generated/sv2v_out.v:12644.39-12644.59" */ 2'h3;
assign _255_ = _274_ && /* src = "generated/sv2v_out.v:12557.9-12557.69" */ _275_;
assign _256_ = _263_ && /* src = "generated/sv2v_out.v:12559.10-12559.32" */ _264_;
assign _257_ = _256_ && /* src = "generated/sv2v_out.v:12559.9-12559.51" */ _265_;
assign _258_ = irq_nm && /* src = "generated/sv2v_out.v:12576.10-12576.31" */ _266_;
assign _259_ = ebreak_into_debug && /* src = "generated/sv2v_out.v:12610.9-12610.43" */ _267_;
assign _260_ = ebrk_insn_prio && /* src = "generated/sv2v_out.v:12682.38-12682.73" */ ebreak_into_debug;
assign _261_ = enter_debug_mode_prio_q && /* src = "generated/sv2v_out.v:12682.9-12682.74" */ _268_;
assign _262_ = ! /* src = "generated/sv2v_out.v:12404.25-12404.38" */ irq_nm_ext_i;
assign _263_ = ! /* src = "generated/sv2v_out.v:12559.10-12559.16" */ stall;
assign _264_ = ! /* src = "generated/sv2v_out.v:12559.20-12559.32" */ special_req;
assign _265_ = ! /* src = "generated/sv2v_out.v:12559.37-12559.51" */ id_wb_pending;
assign _266_ = ! /* src = "generated/sv2v_out.v:12576.20-12576.31" */ nmi_mode_o;
assign _267_ = ! /* src = "generated/sv2v_out.v:12610.30-12610.43" */ debug_mode_o;
assign _268_ = ! /* src = "generated/sv2v_out.v:12682.36-12682.74" */ _260_;
assign _269_ = irq_nm || /* src = "generated/sv2v_out.v:12524.12-12524.35" */ irq_pending_i;
assign _270_ = _269_ || /* src = "generated/sv2v_out.v:12524.11-12524.51" */ debug_req_i;
assign _271_ = _270_ || /* src = "generated/sv2v_out.v:12524.10-12524.68" */ debug_mode_o;
assign _272_ = _271_ || /* src = "generated/sv2v_out.v:12524.9-12524.92" */ debug_single_step_i;
assign _273_ = branch_set_i || /* src = "generated/sv2v_out.v:12549.9-12549.35" */ jump_set_i;
assign _274_ = enter_debug_mode || /* src = "generated/sv2v_out.v:12557.10-12557.40" */ handle_irq;
assign _275_ = stall || /* src = "generated/sv2v_out.v:12557.46-12557.68" */ id_wb_pending;
assign _276_ = exc_req_q || /* src = "generated/sv2v_out.v:12623.10-12623.34" */ store_err_q;
assign _277_ = _276_ || /* src = "generated/sv2v_out.v:12623.9-12623.49" */ load_err_q;
assign _278_ = ctrl_fsm_cs != /* src = "generated/sv2v_out.v:12336.88-12336.107" */ 4'h6;
assign _279_ = | /* src = "generated/sv2v_out.v:12582.15-12582.52" */ irqs_i[14:0];
assign _280_ = ~ /* src = "generated/sv2v_out.v:12342.41-12342.52" */ ready_wb_i;
assign _281_ = ~ /* src = "generated/sv2v_out.v:12398.39-12398.50" */ nmi_mode_o;
assign _282_ = ~ /* src = "generated/sv2v_out.v:12412.80-12412.108" */ \g_intg_irq_int.mem_resp_intg_err_irq_clear ;
assign _283_ = ~ /* src = "generated/sv2v_out.v:12440.40-12440.60" */ debug_single_step_i;
assign _284_ = ~ /* src = "generated/sv2v_out.v:12697.35-12697.43" */ halt_if;
assign _285_ = ~ /* src = "generated/sv2v_out.v:12698.31-12698.51" */ _145_;
assign _287_ = ecall_insn | /* src = "generated/sv2v_out.v:12336.24-12336.46" */ ebrk_insn;
assign _289_ = _287_ | /* src = "generated/sv2v_out.v:12336.23-12336.64" */ illegal_insn_d;
assign _291_ = _289_ | /* src = "generated/sv2v_out.v:12336.22-12336.83" */ instr_fetch_err;
assign exc_req_lsu = store_err_i | /* src = "generated/sv2v_out.v:12337.23-12337.47" */ load_err_i;
assign special_req_flush_only = wfi_insn | /* src = "generated/sv2v_out.v:12339.34-12339.59" */ csr_pipe_flush;
assign _293_ = mret_insn | /* src = "generated/sv2v_out.v:12340.35-12340.56" */ dret_insn;
assign _294_ = _293_ | /* src = "generated/sv2v_out.v:12340.34-12340.69" */ id_exception_o;
assign special_req_pc_change = _294_ | /* src = "generated/sv2v_out.v:12340.33-12340.84" */ exc_req_lsu;
assign special_req = special_req_pc_change | /* src = "generated/sv2v_out.v:12341.23-12341.69" */ special_req_flush_only;
assign id_wb_pending = instr_valid_i | /* src = "generated/sv2v_out.v:12342.25-12342.52" */ _280_;
assign \g_intg_irq_int.mem_resp_intg_err_irq_pending_d  = _109_ | /* src = "generated/sv2v_out.v:12412.45-12412.137" */ \g_intg_irq_int.mem_resp_intg_err_irq_set ;
assign irq_nm_int = \g_intg_irq_int.mem_resp_intg_err_irq_set  | /* src = "generated/sv2v_out.v:12422.24-12422.83" */ \g_intg_irq_int.mem_resp_intg_err_irq_pending_q ;
assign _295_ = debug_req_i | /* src = "generated/sv2v_out.v:12435.36-12435.66" */ do_single_step_d;
assign enter_debug_mode = enter_debug_mode_prio_d | /* src = "generated/sv2v_out.v:12436.28-12436.87" */ _111_;
assign irq_nm = irq_nm_ext_i | /* src = "generated/sv2v_out.v:12438.18-12438.43" */ irq_nm_int;
assign irq_enabled = csr_mstatus_mie_i | /* src = "generated/sv2v_out.v:12439.23-12439.65" */ _254_;
assign _296_ = irq_nm | /* src = "generated/sv2v_out.v:12440.80-12440.118" */ _114_;
assign _297_ = debug_mode_o | /* src = "generated/sv2v_out.v:12646.12-12646.44" */ ebreak_into_debug;
assign stall = stall_id_i | /* src = "generated/sv2v_out.v:12696.17-12696.40" */ stall_wb_i;
assign _145_ = stall | /* src = "generated/sv2v_out.v:12698.33-12698.50" */ retain_id;
assign instr_valid_clear_o = _285_ | /* src = "generated/sv2v_out.v:12698.31-12698.62" */ flush_id_o;
/* src = "generated/sv2v_out.v:12413.4-12421.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  <= 1'h0;
else \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  <= \g_intg_irq_int.mem_resp_intg_err_irq_pending_d ;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME nmi_mode_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) nmi_mode_o <= 1'h0;
else nmi_mode_o <= nmi_mode_d;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME load_err_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) load_err_q <= 1'h0;
else load_err_q <= load_err_i;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME store_err_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) store_err_q <= 1'h0;
else store_err_q <= store_err_i;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME exc_req_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) exc_req_q <= 1'h0;
else exc_req_q <= id_exception_o;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME illegal_insn_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) illegal_insn_q <= 1'h0;
else illegal_insn_q <= illegal_insn_d;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME do_single_step_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) do_single_step_q <= 1'h0;
else do_single_step_q <= do_single_step_d;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME enter_debug_mode_prio_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) enter_debug_mode_prio_q <= 1'h0;
else enter_debug_mode_prio_q <= enter_debug_mode_prio_d;
/* src = "generated/sv2v_out.v:12452.2-12456.35" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME debug_cause_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) debug_cause_o <= 3'h0;
else debug_cause_o <= debug_cause_d;
assign _030_ = mem_resp_intg_err_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12407.14-12407.33|generated/sv2v_out.v:12407.10-12410.8" */ 1'h1 : 1'h0;
assign _029_ = _108_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12404.10-12404.38|generated/sv2v_out.v:12404.6-12405.42" */ 1'h1 : 1'h0;
assign \g_intg_irq_int.mem_resp_intg_err_irq_clear  = \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12403.9-12403.40|generated/sv2v_out.v:12403.5-12410.8" */ _029_ : 1'h0;
assign \g_intg_irq_int.mem_resp_intg_err_irq_set  = \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12403.9-12403.40|generated/sv2v_out.v:12403.5-12410.8" */ 1'h0 : _030_;
assign _093_ = load_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12385.14-12385.24|generated/sv2v_out.v:12385.10-12386.27" */ 1'h1 : 1'h0;
assign _087_ = store_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12383.14-12383.25|generated/sv2v_out.v:12383.10-12386.27" */ 1'h1 : 1'h0;
assign _083_ = store_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12383.14-12383.25|generated/sv2v_out.v:12383.10-12386.27" */ 1'h0 : _093_;
assign _067_ = ebrk_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12381.14-12381.23|generated/sv2v_out.v:12381.10-12386.27" */ 1'h1 : 1'h0;
assign _071_ = ebrk_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12381.14-12381.23|generated/sv2v_out.v:12381.10-12386.27" */ 1'h0 : _083_;
assign _077_ = ebrk_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12381.14-12381.23|generated/sv2v_out.v:12381.10-12386.27" */ 1'h0 : _087_;
assign _051_ = ecall_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12379.14-12379.24|generated/sv2v_out.v:12379.10-12386.27" */ 1'h1 : 1'h0;
assign _055_ = ecall_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12379.14-12379.24|generated/sv2v_out.v:12379.10-12386.27" */ 1'h0 : _071_;
assign _060_ = ecall_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12379.14-12379.24|generated/sv2v_out.v:12379.10-12386.27" */ 1'h0 : _077_;
assign _050_ = ecall_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12379.14-12379.24|generated/sv2v_out.v:12379.10-12386.27" */ 1'h0 : _067_;
assign _031_ = illegal_insn_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12377.14-12377.28|generated/sv2v_out.v:12377.10-12386.27" */ 1'h1 : 1'h0;
assign _032_ = illegal_insn_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12377.14-12377.28|generated/sv2v_out.v:12377.10-12386.27" */ 1'h0 : _055_;
assign _043_ = illegal_insn_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12377.14-12377.28|generated/sv2v_out.v:12377.10-12386.27" */ 1'h0 : _060_;
assign _024_ = illegal_insn_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12377.14-12377.28|generated/sv2v_out.v:12377.10-12386.27" */ 1'h0 : _050_;
assign _025_ = illegal_insn_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12377.14-12377.28|generated/sv2v_out.v:12377.10-12386.27" */ 1'h0 : _051_;
assign instr_fetch_err_prio = instr_fetch_err ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12375.9-12375.24|generated/sv2v_out.v:12375.5-12386.27" */ 1'h1 : 1'h0;
assign load_err_prio = instr_fetch_err ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12375.9-12375.24|generated/sv2v_out.v:12375.5-12386.27" */ 1'h0 : _032_;
assign store_err_prio = instr_fetch_err ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12375.9-12375.24|generated/sv2v_out.v:12375.5-12386.27" */ 1'h0 : _043_;
assign ebrk_insn_prio = instr_fetch_err ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12375.9-12375.24|generated/sv2v_out.v:12375.5-12386.27" */ 1'h0 : _024_;
assign ecall_insn_prio = instr_fetch_err ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12375.9-12375.24|generated/sv2v_out.v:12375.5-12386.27" */ 1'h0 : _025_;
assign illegal_insn_prio = instr_fetch_err ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12375.9-12375.24|generated/sv2v_out.v:12375.5-12386.27" */ 1'h0 : _031_;
assign halt_if = instr_exec_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12690.7-12690.20|generated/sv2v_out.v:12690.3-12691.19" */ _013_ : 1'h1;
assign _012_ = _261_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12682.9-12682.74|generated/sv2v_out.v:12682.5-12683.25" */ 4'h8 : _002_;
assign _011_ = wfi_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12680.14-12680.22|generated/sv2v_out.v:12680.10-12681.25" */ 4'h2 : 4'h5;
assign _066_ = dret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12674.14-12674.23|generated/sv2v_out.v:12674.10-12681.25" */ 1'h0 : 1'hx;
assign _063_ = dret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12674.14-12674.23|generated/sv2v_out.v:12674.10-12681.25" */ 1'h1 : 1'h0;
assign _075_ = dret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12674.14-12674.23|generated/sv2v_out.v:12674.10-12681.25" */ 3'h4 : 3'h0;
assign _010_ = dret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12674.14-12674.23|generated/sv2v_out.v:12674.10-12681.25" */ 4'h5 : _011_;
assign _085_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12667.14-12667.23|generated/sv2v_out.v:12667.10-12681.25" */ 1'h0 : nmi_mode_o;
assign _047_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12667.14-12667.23|generated/sv2v_out.v:12667.10-12681.25" */ 1'h1 : 1'h0;
assign _099_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12667.14-12667.23|generated/sv2v_out.v:12667.10-12681.25" */ 1'h1 : _063_;
assign _059_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12667.14-12667.23|generated/sv2v_out.v:12667.10-12681.25" */ 3'h3 : _075_;
assign _049_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12667.14-12667.23|generated/sv2v_out.v:12667.10-12681.25" */ 1'hx : _066_;
assign _008_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12667.14-12667.23|generated/sv2v_out.v:12667.10-12681.25" */ 4'h5 : _010_;
assign _046_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12667.14-12667.23|generated/sv2v_out.v:12667.10-12681.25" */ 1'h0 : _063_;
assign _006_ = _297_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12646.12-12646.44|generated/sv2v_out.v:12646.8-12654.51" */ 4'h9 : 4'h5;
assign _069_ = _297_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12646.12-12646.44|generated/sv2v_out.v:12646.8-12654.51" */ 1'h0 : 1'h1;
assign _104_ = _297_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12646.12-12646.44|generated/sv2v_out.v:12646.8-12654.51" */ 7'h00 : 7'h03;
assign _299_ = load_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ lsu_addr_last_i : 32'd0;
assign _301_ = store_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ lsu_addr_last_i : _299_;
assign _303_ = ebrk_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 32'd0 : _301_;
assign _305_ = ecall_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 32'd0 : _303_;
assign _307_ = illegal_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ _337_ : _305_;
assign _088_ = instr_fetch_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ _335_ : _307_;
assign _309_ = load_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 7'h05 : 7'h00;
assign _310_ = store_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 7'h07 : _309_;
assign _311_ = ebrk_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ _104_ : _310_;
assign _312_ = ecall_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ _339_ : _311_;
assign _313_ = illegal_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 7'h02 : _312_;
assign _101_ = instr_fetch_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 7'h01 : _313_;
assign _314_ = ebrk_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ _006_ : 4'h5;
assign _315_ = ecall_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 4'h5 : _314_;
assign _316_ = illegal_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 4'h5 : _315_;
assign _004_ = instr_fetch_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 4'h5 : _316_;
assign _318_ = ecall_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 1'h1 : _317_;
assign _319_ = illegal_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 1'h1 : _318_;
assign _053_ = instr_fetch_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 1'h1 : _319_;
assign _317_ = ebrk_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ _069_ : 1'h1;
assign _002_ = _277_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ _004_ : _008_;
assign _028_ = _277_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ _053_ : 1'h1;
assign _078_ = _277_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ _088_ : 32'd0;
assign _064_ = _277_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ _053_ : 1'h0;
assign _096_ = _277_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ _101_ : 7'h00;
assign _076_ = _277_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ _053_ : _099_;
assign _027_ = _277_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ _334_ : 2'h1;
assign _036_ = _277_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ 3'h2 : _059_;
assign _023_ = _277_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ 1'hx : _049_;
assign _073_ = _277_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ nmi_mode_o : _085_;
assign _017_ = _277_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ 1'h0 : _046_;
assign _018_ = _277_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ 1'h0 : _047_;
assign _020_ = _259_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12610.9-12610.43|generated/sv2v_out.v:12610.5-12614.8" */ 1'h1 : 1'h0;
assign _091_ = irqs_i[17] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12586.15-12586.25|generated/sv2v_out.v:12586.11-12589.48" */ 7'h23 : 7'h27;
assign _081_ = irqs_i[15] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12584.15-12584.25|generated/sv2v_out.v:12584.11-12589.48" */ 7'h2b : _091_;
assign _068_ = _279_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12582.15-12582.52|generated/sv2v_out.v:12582.11-12589.48" */ { 3'h3, mfip_id } : _081_;
assign _061_ = _116_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12578.11-12578.37|generated/sv2v_out.v:12578.7-12579.39" */ \g_intg_irq_int.mem_resp_intg_err_addr_q  : 32'd0;
assign _057_ = _258_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12576.10-12576.31|generated/sv2v_out.v:12576.6-12589.48" */ 1'h1 : nmi_mode_o;
assign _044_ = _258_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12576.10-12576.31|generated/sv2v_out.v:12576.6-12589.48" */ _061_ : 32'd0;
assign _052_ = _258_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12576.10-12576.31|generated/sv2v_out.v:12576.6-12589.48" */ _333_ : _068_;
assign _034_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12572.9-12572.19|generated/sv2v_out.v:12572.5-12590.8" */ _057_ : nmi_mode_o;
assign _015_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12572.9-12572.19|generated/sv2v_out.v:12572.5-12590.8" */ _044_ : 32'd0;
assign _026_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12572.9-12572.19|generated/sv2v_out.v:12572.5-12590.8" */ _052_ : 7'h00;
assign _019_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12572.9-12572.19|generated/sv2v_out.v:12572.5-12590.8" */ 1'h1 : 1'h0;
assign _097_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12564.15-12564.25|generated/sv2v_out.v:12564.11-12567.9" */ 1'h1 : _070_;
assign _000_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12564.15-12564.25|generated/sv2v_out.v:12564.11-12567.9" */ 4'h7 : _090_;
assign _092_ = enter_debug_mode ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12560.10-12560.26|generated/sv2v_out.v:12560.6-12567.9" */ 1'h1 : _097_;
assign _103_ = enter_debug_mode ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12560.10-12560.26|generated/sv2v_out.v:12560.6-12567.9" */ 4'h8 : _000_;
assign _082_ = _257_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12559.9-12559.51|generated/sv2v_out.v:12559.5-12567.9" */ _092_ : _070_;
assign _100_ = _257_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12559.9-12559.51|generated/sv2v_out.v:12559.5-12567.9" */ _103_ : _090_;
assign _070_ = _255_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12557.9-12557.69|generated/sv2v_out.v:12557.5-12558.21" */ 1'h1 : 1'h0;
assign _038_ = _273_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12549.9-12549.35|generated/sv2v_out.v:12549.5-12553.8" */ jump_set_i : 1'h0;
assign _040_ = _273_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12549.9-12549.35|generated/sv2v_out.v:12549.5-12553.8" */ branch_set_i : 1'h0;
assign _037_ = _273_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12549.9-12549.35|generated/sv2v_out.v:12549.5-12553.8" */ 1'h1 : 1'h0;
assign _095_ = ready_wb_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12546.10-12546.37|generated/sv2v_out.v:12546.6-12547.26" */ 4'h6 : ctrl_fsm_cs;
assign _090_ = special_req ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12544.9-12544.20|generated/sv2v_out.v:12544.5-12548.8" */ _095_ : ctrl_fsm_cs;
assign _042_ = special_req ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12544.9-12544.20|generated/sv2v_out.v:12544.5-12548.8" */ 1'h1 : 1'h0;
assign _054_ = enter_debug_mode ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12536.9-12536.25|generated/sv2v_out.v:12536.5-12539.8" */ 1'h1 : _019_;
assign _080_ = enter_debug_mode ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12536.9-12536.25|generated/sv2v_out.v:12536.5-12539.8" */ 4'h8 : _065_;
assign _065_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12532.9-12532.19|generated/sv2v_out.v:12532.5-12535.8" */ 4'h7 : _048_;
assign _048_ = id_in_ready_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12530.9-12530.22|generated/sv2v_out.v:12530.5-12531.25" */ 4'h5 : 4'hx;
assign _022_ = _272_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12524.9-12524.92|generated/sv2v_out.v:12524.5-12527.25" */ 4'h4 : 4'hx;
assign _021_ = _272_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12524.9-12524.92|generated/sv2v_out.v:12524.5-12527.25" */ 1'h1 : 1'h0;
assign _328_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ ctrl_fsm_cs;
assign instr_req_o = _164_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 1'h1 : 1'h0;
assign _327_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h1;
assign retain_id = _322_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ _042_ : 1'h0;
assign _323_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h4;
assign _321_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h7;
assign controller_run_o = _322_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 1'h1 : 1'h0;
assign _298_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h6;
assign _325_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h8;
assign _324_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h3;
assign _326_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h2;
assign perf_tbranch_o = _322_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ _040_ : 1'h0;
assign perf_jump_o = _322_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ _038_ : 1'h0;
assign _322_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h5;
assign _320_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h9;
assign debug_mode_entering_o = _150_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 1'h1 : 1'h0;
assign csr_restore_dret_id_o = _298_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ _017_ : 1'h0;
assign csr_restore_mret_id_o = _298_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ _018_ : 1'h0;
assign csr_save_id_o = _320_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ _020_ : 1'h0;
assign mfip_id = irqs_i[0] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h0 : _009_;
assign _009_ = irqs_i[1] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h1 : _007_;
assign _007_ = irqs_i[2] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h2 : _005_;
assign _005_ = irqs_i[3] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h3 : _003_;
assign _003_ = irqs_i[4] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h4 : _001_;
assign _001_ = irqs_i[5] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h5 : _105_;
assign _105_ = irqs_i[6] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h6 : _102_;
assign _102_ = irqs_i[7] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h7 : _098_;
assign _098_ = irqs_i[8] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h8 : _094_;
assign _094_ = irqs_i[9] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h9 : _084_;
assign _084_ = irqs_i[10] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'ha : _072_;
assign _072_ = irqs_i[11] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'hb : _056_;
assign _056_ = irqs_i[12] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'hc : _033_;
assign _033_ = irqs_i[13] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'hd : _014_;
assign _014_ = irqs_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'he : 4'h0;
assign do_single_step_d = instr_valid_i ? /* src = "generated/sv2v_out.v:12434.29-12434.99" */ _110_ : do_single_step_q;
assign _329_ = _254_ ? /* src = "generated/sv2v_out.v:12437.72-12437.117" */ debug_ebreaku_i : 1'h0;
assign ebreak_into_debug = _253_ ? /* src = "generated/sv2v_out.v:12437.30-12437.118" */ debug_ebreakm_i : _329_;
assign _330_ = do_single_step_d ? /* src = "generated/sv2v_out.v:12451.119-12451.149" */ 3'h4 : 3'h0;
assign _331_ = debug_req_i ? /* src = "generated/sv2v_out.v:12451.97-12451.150" */ 3'h3 : _330_;
assign _332_ = _115_ ? /* src = "generated/sv2v_out.v:12451.52-12451.151" */ 3'h1 : _331_;
assign debug_cause_d = trigger_match_i ? /* src = "generated/sv2v_out.v:12451.26-12451.152" */ 3'h2 : _332_;
assign _333_ = irq_nm_ext_i ? /* src = "generated/sv2v_out.v:12577.22-12577.87" */ 7'h3f : 7'h40;
assign _334_ = debug_mode_o ? /* src = "generated/sv2v_out.v:12626.22-12626.48" */ 2'h3 : 2'h0;
assign _335_ = instr_fetch_err_plus2_i ? /* src = "generated/sv2v_out.v:12638.23-12638.74" */ _106_ : pc_id_i;
assign _337_ = instr_is_compressed_i ? /* src = "generated/sv2v_out.v:12642.23-12642.99" */ { 16'h0000, instr_compressed_i } : instr_i;
assign _339_ = _253_ ? /* src = "generated/sv2v_out.v:12644.39-12644.119" */ 7'h0b : 7'h08;
assign controller_run_o_t0 = 1'h0;
assign csr_restore_dret_id_o_t0 = 1'h0;
assign csr_restore_mret_id_o_t0 = 1'h0;
assign csr_save_cause_o_t0 = 1'h0;
assign csr_save_id_o_t0 = 1'h0;
assign csr_save_if_o_t0 = 1'h0;
assign csr_save_wb_o = 1'h0;
assign csr_save_wb_o_t0 = 1'h0;
assign ctrl_busy_o_t0 = 1'h0;
assign debug_cause_o_t0 = 3'h0;
assign debug_csr_save_o_t0 = 1'h0;
assign debug_mode_entering_o_t0 = 1'h0;
assign exc_cause_o_t0 = 7'h00;
assign exc_pc_mux_o_t0 = 2'h0;
assign flush_id_o_t0 = 1'h0;
assign instr_req_o_t0 = 1'h0;
assign nt_branch_mispredict_o = 1'h0;
assign nt_branch_mispredict_o_t0 = 1'h0;
assign pc_mux_o_t0 = 3'h0;
assign pc_set_o_t0 = 1'h0;
assign wb_exception_o = 1'h0;
assign wb_exception_o_t0 = 1'h0;
endmodule

module \$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000 (clk_i, rst_ni, counter_inc_i, counterh_we_i, counter_we_i, counter_val_i, counter_val_o, counter_val_upd_o, counter_inc_i_t0, counter_val_i_t0, counter_val_o_t0, counter_val_upd_o_t0, counter_we_i_t0, counterh_we_i_t0);
/* src = "generated/sv2v_out.v:13636.2-13650.5" */
wire [63:0] _00_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13636.2-13650.5" */
wire [63:0] _01_;
wire [63:0] _02_;
wire _03_;
wire _04_;
wire [63:0] _05_;
wire [31:0] _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire [63:0] _12_;
wire [31:0] _13_;
wire [31:0] _14_;
wire [31:0] _15_;
wire [31:0] _16_;
wire [63:0] _17_;
wire [63:0] _18_;
wire [63:0] _19_;
wire [31:0] _20_;
wire [31:0] _21_;
wire [63:0] _22_;
wire [63:0] _23_;
wire [63:0] _24_;
/* src = "generated/sv2v_out.v:13622.13-13622.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:13634.27-13634.36" */
wire [63:0] counter_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13634.27-13634.36" */
wire [63:0] counter_d_t0;
/* src = "generated/sv2v_out.v:13624.13-13624.26" */
input counter_inc_i;
wire counter_inc_i;
/* cellift = 32'd1 */
input counter_inc_i_t0;
wire counter_inc_i_t0;
/* src = "generated/sv2v_out.v:13632.13-13632.25" */
wire [63:0] counter_load;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13632.13-13632.25" */
wire [63:0] counter_load_t0;
/* src = "generated/sv2v_out.v:13631.28-13631.39" */
wire [63:0] counter_upd;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13631.28-13631.39" */
wire [63:0] counter_upd_t0;
/* src = "generated/sv2v_out.v:13627.20-13627.33" */
input [31:0] counter_val_i;
wire [31:0] counter_val_i;
/* cellift = 32'd1 */
input [31:0] counter_val_i_t0;
wire [31:0] counter_val_i_t0;
/* src = "generated/sv2v_out.v:13628.21-13628.34" */
output [63:0] counter_val_o;
reg [63:0] counter_val_o;
/* cellift = 32'd1 */
output [63:0] counter_val_o_t0;
reg [63:0] counter_val_o_t0;
/* src = "generated/sv2v_out.v:13629.21-13629.38" */
output [63:0] counter_val_upd_o;
wire [63:0] counter_val_upd_o;
/* cellift = 32'd1 */
output [63:0] counter_val_upd_o_t0;
wire [63:0] counter_val_upd_o_t0;
/* src = "generated/sv2v_out.v:13626.13-13626.25" */
input counter_we_i;
wire counter_we_i;
/* cellift = 32'd1 */
input counter_we_i_t0;
wire counter_we_i_t0;
/* src = "generated/sv2v_out.v:13625.13-13625.26" */
input counterh_we_i;
wire counterh_we_i;
/* cellift = 32'd1 */
input counterh_we_i_t0;
wire counterh_we_i_t0;
/* src = "generated/sv2v_out.v:13623.13-13623.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:13633.6-13633.8" */
wire we;
assign counter_upd = counter_val_o + /* src = "generated/sv2v_out.v:13635.23-13635.86" */ 64'h0000000000000001;
assign _02_ = ~ counter_val_o_t0;
assign _12_ = counter_val_o & _02_;
assign _23_ = _12_ + 64'h0000000000000001;
assign _19_ = counter_val_o | counter_val_o_t0;
assign _24_ = _19_ + 64'h0000000000000001;
assign _22_ = _23_ ^ _24_;
assign counter_upd_t0 = _22_ | counter_val_o_t0;
assign _03_ = ~ _10_;
assign _04_ = ~ _11_;
assign _13_ = { _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_ } & counter_d_t0[63:32];
assign _15_ = { _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_ } & counter_d_t0[31:0];
assign _14_ = { _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_ } & counter_val_o_t0[63:32];
assign _16_ = { _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_ } & counter_val_o_t0[31:0];
assign _20_ = _13_ | _14_;
assign _21_ = _15_ | _16_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000  */
/* PC_TAINT_INFO STATE_NAME counter_val_o_t0[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o_t0[63:32] <= 32'd0;
else counter_val_o_t0[63:32] <= _20_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000  */
/* PC_TAINT_INFO STATE_NAME counter_val_o_t0[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o_t0[31:0] <= 32'd0;
else counter_val_o_t0[31:0] <= _21_;
/* src = "generated/sv2v_out.v:13652.2-13656.27" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000  */
/* PC_TAINT_INFO STATE_NAME counter_val_o[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o[63:32] <= 32'd0;
else if (_10_) counter_val_o[63:32] <= counter_d[63:32];
/* src = "generated/sv2v_out.v:13652.2-13656.27" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000  */
/* PC_TAINT_INFO STATE_NAME counter_val_o[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o[31:0] <= 32'd0;
else if (_11_) counter_val_o[31:0] <= counter_d[31:0];
assign _05_ = ~ { we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we };
assign _06_ = ~ { counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i };
assign _17_ = _05_ & _01_;
assign counter_load_t0[31:0] = _06_ & counter_val_i_t0;
assign _01_ = { counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i } & counter_upd_t0;
assign _18_ = { we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we } & counter_load_t0;
assign counter_load_t0[63:32] = { counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i } & counter_val_i_t0;
assign counter_d_t0 = _17_ | _18_;
assign _07_ = | { we, counter_inc_i };
assign _08_ = { we, counterh_we_i } != 2'h2;
assign _09_ = { we, counterh_we_i } != 2'h3;
assign _10_ = & { _07_, _08_ };
assign _11_ = & { _07_, _09_ };
assign we = counter_we_i | /* src = "generated/sv2v_out.v:13637.8-13637.36" */ counterh_we_i;
assign _00_ = counter_inc_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13646.12-13646.25|generated/sv2v_out.v:13646.8-13649.44" */ counter_upd : 64'hxxxxxxxxxxxxxxxx;
assign counter_d = we ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13644.7-13644.9|generated/sv2v_out.v:13644.3-13649.44" */ counter_load : _00_;
assign counter_load[63:32] = counterh_we_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13640.7-13640.20|generated/sv2v_out.v:13640.3-13643.6" */ counter_val_i : 32'hxxxxxxxx;
assign counter_load[31:0] = counterh_we_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13640.7-13640.20|generated/sv2v_out.v:13640.3-13643.6" */ 32'hxxxxxxxx : counter_val_i;
assign counter_val_upd_o = 64'h0000000000000000;
assign counter_val_upd_o_t0 = 64'h0000000000000000;
endmodule

module \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1 (clk_i, rst_ni, clear_i, busy_o, in_valid_i, in_addr_i, in_rdata_i, in_err_i, out_valid_o, out_ready_i, out_addr_o, out_rdata_o, out_err_o, out_err_plus2_o, out_valid_o_t0, out_ready_i_t0, out_rdata_o_t0, out_err_plus2_o_t0, out_err_o_t0, out_addr_o_t0, in_valid_i_t0
, in_rdata_i_t0, in_err_i_t0, in_addr_i_t0, clear_i_t0, busy_o_t0);
/* src = "generated/sv2v_out.v:16150.2-16165.6" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16150.2-16165.6" */
wire _001_;
/* src = "generated/sv2v_out.v:16145.40-16145.75" */
wire _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16145.40-16145.75" */
wire _003_;
/* src = "generated/sv2v_out.v:16145.91-16145.112" */
wire _004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16145.91-16145.112" */
wire _005_;
/* src = "generated/sv2v_out.v:16145.117-16145.168" */
wire _006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16145.117-16145.168" */
wire _007_;
/* src = "generated/sv2v_out.v:16146.35-16146.55" */
wire _008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16146.35-16146.55" */
wire _009_;
/* src = "generated/sv2v_out.v:16146.59-16146.80" */
wire _010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16146.59-16146.80" */
wire _011_;
/* src = "generated/sv2v_out.v:16146.58-16146.93" */
wire _012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16146.58-16146.93" */
wire _013_;
/* src = "generated/sv2v_out.v:16147.48-16147.71" */
wire _014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16147.48-16147.71" */
wire _015_;
/* src = "generated/sv2v_out.v:16166.36-16166.61" */
wire _016_;
/* src = "generated/sv2v_out.v:16197.30-16197.63" */
wire _017_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16197.30-16197.63" */
wire _018_;
/* src = "generated/sv2v_out.v:16197.30-16197.63" */
wire _019_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16197.30-16197.63" */
wire _020_;
/* src = "generated/sv2v_out.v:16200.26-16200.56" */
wire _021_;
/* src = "generated/sv2v_out.v:16200.61-16200.108" */
wire _022_;
/* src = "generated/sv2v_out.v:16200.26-16200.56" */
wire _023_;
/* src = "generated/sv2v_out.v:16200.61-16200.108" */
wire _024_;
wire [30:0] _025_;
wire [30:0] _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire [31:0] _033_;
wire [31:0] _034_;
wire [31:0] _035_;
wire _036_;
wire [30:0] _037_;
wire _038_;
wire [31:0] _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire [30:0] _049_;
wire [30:0] _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire [31:0] _098_;
wire [31:0] _099_;
wire _100_;
wire _101_;
wire [31:0] _102_;
wire [31:0] _103_;
wire _104_;
wire _105_;
wire [31:0] _106_;
wire [31:0] _107_;
wire [30:0] _108_;
wire [30:0] _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire [31:0] _136_;
wire [31:0] _137_;
wire [31:0] _138_;
wire [31:0] _139_;
wire _140_;
wire [31:0] _141_;
wire [31:0] _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire [30:0] _148_;
wire [30:0] _149_;
wire _150_;
wire _151_;
wire [31:0] _152_;
wire [31:0] _153_;
wire [31:0] _154_;
wire [31:0] _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire [30:0] _160_;
wire [30:0] _161_;
wire [30:0] _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire [31:0] _179_;
wire _180_;
wire [31:0] _181_;
wire _182_;
wire [31:0] _183_;
wire [30:0] _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire [30:0] _192_;
wire [30:0] _193_;
wire [30:0] _194_;
/* src = "generated/sv2v_out.v:16148.36-16148.57" */
wire _195_;
/* src = "generated/sv2v_out.v:16149.34-16149.53" */
wire _196_;
/* src = "generated/sv2v_out.v:16148.61-16148.65" */
wire _197_;
/* src = "generated/sv2v_out.v:16168.56-16168.70" */
wire _198_;
/* src = "generated/sv2v_out.v:16187.51-16187.73" */
wire _199_;
/* src = "generated/sv2v_out.v:16145.39-16145.87" */
wire _200_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16145.39-16145.87" */
wire _201_;
/* src = "generated/sv2v_out.v:16145.129-16145.167" */
wire _202_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16145.129-16145.167" */
wire _203_;
/* src = "generated/sv2v_out.v:16145.90-16145.169" */
wire _204_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16145.90-16145.169" */
wire _205_;
/* src = "generated/sv2v_out.v:16187.51-16187.89" */
wire _206_;
/* src = "generated/sv2v_out.v:16135.7-16135.20" */
wire addr_incr_two;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16135.7-16135.20" */
wire addr_incr_two_t0;
/* src = "generated/sv2v_out.v:16133.7-16133.28" */
wire aligned_is_compressed;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16133.7-16133.28" */
wire aligned_is_compressed_t0;
/* src = "generated/sv2v_out.v:16103.31-16103.37" */
output [1:0] busy_o;
wire [1:0] busy_o;
/* cellift = 32'd1 */
output [1:0] busy_o_t0;
wire [1:0] busy_o_t0;
/* src = "generated/sv2v_out.v:16102.13-16102.20" */
input clear_i;
wire clear_i;
/* cellift = 32'd1 */
input clear_i_t0;
wire clear_i_t0;
/* src = "generated/sv2v_out.v:16100.13-16100.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:16124.21-16124.29" */
wire [2:0] entry_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16124.21-16124.29" */
/* unused_bits = "0 1" */
wire [2:0] entry_en_t0;
/* src = "generated/sv2v_out.v:16128.7-16128.10" */
wire err;
/* src = "generated/sv2v_out.v:16117.21-16117.26" */
wire [2:0] err_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16117.21-16117.26" */
wire [2:0] err_d_t0;
/* src = "generated/sv2v_out.v:16130.7-16130.16" */
wire err_plus2;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16130.7-16130.16" */
wire err_plus2_t0;
/* src = "generated/sv2v_out.v:16118.20-16118.25" */
reg [2:0] err_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16118.20-16118.25" */
reg [2:0] err_q_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16128.7-16128.10" */
wire err_t0;
/* src = "generated/sv2v_out.v:16129.7-16129.20" */
wire err_unaligned;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16129.7-16129.20" */
wire err_unaligned_t0;
/* src = "generated/sv2v_out.v:16105.20-16105.29" */
input [31:0] in_addr_i;
wire [31:0] in_addr_i;
/* cellift = 32'd1 */
input [31:0] in_addr_i_t0;
wire [31:0] in_addr_i_t0;
/* src = "generated/sv2v_out.v:16107.13-16107.21" */
input in_err_i;
wire in_err_i;
/* cellift = 32'd1 */
input in_err_i_t0;
wire in_err_i_t0;
/* src = "generated/sv2v_out.v:16106.20-16106.30" */
input [31:0] in_rdata_i;
wire [31:0] in_rdata_i;
/* cellift = 32'd1 */
input [31:0] in_rdata_i_t0;
wire [31:0] in_rdata_i_t0;
/* src = "generated/sv2v_out.v:16104.13-16104.23" */
input in_valid_i;
wire in_valid_i;
/* cellift = 32'd1 */
input in_valid_i_t0;
wire in_valid_i_t0;
/* src = "generated/sv2v_out.v:16137.14-16137.26" */
wire [31:1] instr_addr_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16137.14-16137.26" */
wire [31:1] instr_addr_d_t0;
/* src = "generated/sv2v_out.v:16139.7-16139.20" */
wire instr_addr_en;
/* src = "generated/sv2v_out.v:16136.14-16136.29" */
wire [31:1] instr_addr_next;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16136.14-16136.29" */
wire [31:1] instr_addr_next_t0;
/* src = "generated/sv2v_out.v:16138.13-16138.25" */
reg [31:1] instr_addr_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16138.13-16138.25" */
reg [31:1] instr_addr_q_t0;
/* src = "generated/sv2v_out.v:16121.21-16121.38" */
wire [2:0] lowest_free_entry;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16121.21-16121.38" */
wire [2:0] lowest_free_entry_t0;
/* src = "generated/sv2v_out.v:16110.21-16110.31" */
output [31:0] out_addr_o;
wire [31:0] out_addr_o;
/* cellift = 32'd1 */
output [31:0] out_addr_o_t0;
wire [31:0] out_addr_o_t0;
/* src = "generated/sv2v_out.v:16112.13-16112.22" */
output out_err_o;
wire out_err_o;
/* cellift = 32'd1 */
output out_err_o_t0;
wire out_err_o_t0;
/* src = "generated/sv2v_out.v:16113.13-16113.28" */
output out_err_plus2_o;
wire out_err_plus2_o;
/* cellift = 32'd1 */
output out_err_plus2_o_t0;
wire out_err_plus2_o_t0;
/* src = "generated/sv2v_out.v:16111.20-16111.31" */
output [31:0] out_rdata_o;
wire [31:0] out_rdata_o;
/* cellift = 32'd1 */
output [31:0] out_rdata_o_t0;
wire [31:0] out_rdata_o_t0;
/* src = "generated/sv2v_out.v:16109.13-16109.24" */
input out_ready_i;
wire out_ready_i;
/* cellift = 32'd1 */
input out_ready_i_t0;
wire out_ready_i_t0;
/* src = "generated/sv2v_out.v:16108.13-16108.24" */
output out_valid_o;
wire out_valid_o;
/* cellift = 32'd1 */
output out_valid_o_t0;
wire out_valid_o_t0;
/* src = "generated/sv2v_out.v:16125.7-16125.15" */
wire pop_fifo;
/* src = "generated/sv2v_out.v:16126.14-16126.19" */
wire [31:0] rdata;
/* src = "generated/sv2v_out.v:16115.28-16115.35" */
wire [95:0] rdata_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16115.28-16115.35" */
wire [95:0] rdata_d_t0;
/* src = "generated/sv2v_out.v:16116.27-16116.34" */
reg [95:0] rdata_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16116.27-16116.34" */
reg [95:0] rdata_q_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16126.14-16126.19" */
wire [31:0] rdata_t0;
/* src = "generated/sv2v_out.v:16127.14-16127.29" */
wire [31:0] rdata_unaligned;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16127.14-16127.29" */
wire [31:0] rdata_unaligned_t0;
/* src = "generated/sv2v_out.v:16101.13-16101.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:16134.7-16134.30" */
wire unaligned_is_compressed;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16134.7-16134.30" */
wire unaligned_is_compressed_t0;
/* src = "generated/sv2v_out.v:16131.7-16131.12" */
wire valid;
/* src = "generated/sv2v_out.v:16119.21-16119.28" */
wire [2:0] valid_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16119.21-16119.28" */
wire [2:0] valid_d_t0;
/* src = "generated/sv2v_out.v:16123.21-16123.33" */
wire [2:0] valid_popped;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16123.21-16123.33" */
wire [2:0] valid_popped_t0;
/* src = "generated/sv2v_out.v:16122.21-16122.33" */
wire [2:0] valid_pushed;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16122.21-16122.33" */
wire [2:0] valid_pushed_t0;
/* src = "generated/sv2v_out.v:16120.20-16120.27" */
reg [2:0] valid_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16120.20-16120.27" */
reg [2:0] valid_q_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16131.7-16131.12" */
wire valid_t0;
/* src = "generated/sv2v_out.v:16132.7-16132.22" */
wire valid_unaligned;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16132.7-16132.22" */
wire valid_unaligned_t0;
assign instr_addr_next = instr_addr_q + /* src = "generated/sv2v_out.v:16168.27-16168.86" */ { 29'h00000000, _198_, addr_incr_two };
assign _002_ = err_q[1] & /* src = "generated/sv2v_out.v:16145.40-16145.75" */ _031_;
assign _004_ = valid_q[0] & /* src = "generated/sv2v_out.v:16145.91-16145.112" */ err_q[0];
assign _006_ = in_err_i & /* src = "generated/sv2v_out.v:16145.117-16145.168" */ _202_;
assign _008_ = err_q[1] & /* src = "generated/sv2v_out.v:16146.35-16146.55" */ _047_;
assign _010_ = in_err_i & /* src = "generated/sv2v_out.v:16146.59-16146.80" */ valid_q[0];
assign _012_ = _010_ & /* src = "generated/sv2v_out.v:16146.58-16146.93" */ _047_;
assign _014_ = valid_q[0] & /* src = "generated/sv2v_out.v:16147.48-16147.71" */ in_valid_i;
assign unaligned_is_compressed = _195_ & /* src = "generated/sv2v_out.v:16148.35-16148.65" */ _197_;
assign aligned_is_compressed = _196_ & /* src = "generated/sv2v_out.v:16149.33-16149.61" */ _197_;
assign _016_ = out_ready_i & /* src = "generated/sv2v_out.v:16187.21-16187.46" */ out_valid_o;
assign pop_fifo = _016_ & /* src = "generated/sv2v_out.v:16187.20-16187.90" */ _206_;
assign lowest_free_entry[1] = _036_ & /* src = "generated/sv2v_out.v:16195.35-16195.63" */ valid_q[0];
assign valid_d[0] = valid_popped[0] & /* src = "generated/sv2v_out.v:16199.24-16199.50" */ _043_;
assign valid_d[1] = valid_popped[1] & /* src = "generated/sv2v_out.v:16199.24-16199.50" */ _043_;
assign _021_ = valid_pushed[1] & /* src = "generated/sv2v_out.v:16200.26-16200.56" */ pop_fifo;
assign _017_ = in_valid_i & /* src = "generated/sv2v_out.v:16200.62-16200.95" */ lowest_free_entry[0];
assign _022_ = _017_ & /* src = "generated/sv2v_out.v:16200.61-16200.108" */ _038_;
assign _023_ = valid_pushed[2] & /* src = "generated/sv2v_out.v:16200.26-16200.56" */ pop_fifo;
assign _019_ = in_valid_i & /* src = "generated/sv2v_out.v:16200.62-16200.95" */ lowest_free_entry[1];
assign _024_ = _019_ & /* src = "generated/sv2v_out.v:16200.61-16200.108" */ _038_;
assign lowest_free_entry[2] = _040_ & /* src = "generated/sv2v_out.v:16205.40-16205.80" */ valid_q[1];
assign valid_d[2] = valid_popped[2] & /* src = "generated/sv2v_out.v:16208.30-16208.64" */ _043_;
assign entry_en[2] = in_valid_i & /* src = "generated/sv2v_out.v:16209.31-16209.72" */ lowest_free_entry[2];
assign _025_ = ~ instr_addr_q_t0;
assign _026_ = ~ { 29'h00000000, addr_incr_two_t0, addr_incr_two_t0 };
assign _049_ = instr_addr_q & _025_;
assign _050_ = { 29'h00000000, _198_, addr_incr_two } & _026_;
assign _193_ = _049_ + _050_;
assign _160_ = instr_addr_q | instr_addr_q_t0;
assign _161_ = { 29'h00000000, _198_, addr_incr_two } | { 29'h00000000, addr_incr_two_t0, addr_incr_two_t0 };
assign _194_ = _160_ + _161_;
assign _192_ = _193_ ^ _194_;
assign _162_ = _192_ | instr_addr_q_t0;
assign instr_addr_next_t0 = _162_ | { 29'h00000000, addr_incr_two_t0, addr_incr_two_t0 };
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME valid_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) valid_q_t0 <= 3'h0;
else valid_q_t0 <= valid_d_t0;
assign _027_ = ~ entry_en[2];
assign _028_ = ~ entry_en[1];
assign _029_ = ~ entry_en[0];
assign _030_ = ~ instr_addr_en;
assign _096_ = entry_en[2] & in_err_i_t0;
assign _098_ = { entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2] } & in_rdata_i_t0;
assign _100_ = entry_en[1] & err_d_t0[1];
assign _102_ = { entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1] } & rdata_d_t0[63:32];
assign _104_ = entry_en[0] & err_d_t0[0];
assign _106_ = { entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0] } & rdata_d_t0[31:0];
assign _108_ = { instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en } & instr_addr_d_t0;
assign _097_ = _027_ & err_q_t0[2];
assign _099_ = { _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_ } & rdata_q_t0[95:64];
assign _101_ = _028_ & err_q_t0[1];
assign _103_ = { _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_ } & rdata_q_t0[63:32];
assign _105_ = _029_ & err_q_t0[0];
assign _107_ = { _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_ } & rdata_q_t0[31:0];
assign _109_ = { _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_ } & instr_addr_q_t0;
assign _178_ = _096_ | _097_;
assign _179_ = _098_ | _099_;
assign _180_ = _100_ | _101_;
assign _181_ = _102_ | _103_;
assign _182_ = _104_ | _105_;
assign _183_ = _106_ | _107_;
assign _184_ = _108_ | _109_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q_t0[2] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q_t0[2] <= 1'h0;
else err_q_t0[2] <= _178_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q_t0[95:64] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q_t0[95:64] <= 32'd0;
else rdata_q_t0[95:64] <= _179_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q_t0[1] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q_t0[1] <= 1'h0;
else err_q_t0[1] <= _180_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q_t0[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q_t0[63:32] <= 32'd0;
else rdata_q_t0[63:32] <= _181_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q_t0[0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q_t0[0] <= 1'h0;
else err_q_t0[0] <= _182_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q_t0[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q_t0[31:0] <= 32'd0;
else rdata_q_t0[31:0] <= _183_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME instr_addr_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_addr_q_t0 <= 31'h00000000;
else instr_addr_q_t0 <= _184_;
assign _051_ = err_q_t0[1] & _031_;
assign _054_ = valid_q_t0[0] & err_q[0];
assign _057_ = in_err_i_t0 & _202_;
assign _060_ = err_q_t0[1] & _047_;
assign _063_ = in_err_i_t0 & valid_q[0];
assign _066_ = _011_ & _047_;
assign _069_ = valid_q_t0[0] & in_valid_i;
assign _072_ = valid_q_t0[1] & valid_q[0];
assign _075_ = valid_popped_t0[0] & _043_;
assign _078_ = valid_popped_t0[1] & _043_;
assign _081_ = valid_pushed_t0[1] & pop_fifo;
assign _082_ = in_valid_i_t0 & lowest_free_entry[0];
assign _083_ = valid_pushed_t0[2] & pop_fifo;
assign _084_ = in_valid_i_t0 & lowest_free_entry[1];
assign _087_ = valid_q_t0[2] & valid_q[1];
assign _090_ = valid_popped_t0[2] & _043_;
assign _093_ = in_valid_i_t0 & lowest_free_entry[2];
assign _052_ = unaligned_is_compressed_t0 & err_q[1];
assign _055_ = err_q_t0[0] & valid_q[0];
assign _058_ = _203_ & in_err_i;
assign _061_ = err_q_t0[0] & err_q[1];
assign _064_ = valid_q_t0[0] & in_err_i;
assign _067_ = err_q_t0[0] & _010_;
assign _070_ = in_valid_i_t0 & valid_q[0];
assign unaligned_is_compressed_t0 = err_t0 & _195_;
assign aligned_is_compressed_t0 = err_t0 & _196_;
assign _073_ = valid_q_t0[0] & _036_;
assign _076_ = clear_i_t0 & valid_popped[0];
assign _079_ = clear_i_t0 & valid_popped[1];
assign _085_ = lowest_free_entry_t0[1] & in_valid_i;
assign _088_ = valid_q_t0[1] & _040_;
assign _091_ = clear_i_t0 & valid_popped[2];
assign _094_ = lowest_free_entry_t0[2] & in_valid_i;
assign _053_ = err_q_t0[1] & unaligned_is_compressed_t0;
assign _056_ = valid_q_t0[0] & err_q_t0[0];
assign _059_ = in_err_i_t0 & _203_;
assign _062_ = err_q_t0[1] & err_q_t0[0];
assign _065_ = in_err_i_t0 & valid_q_t0[0];
assign _068_ = _011_ & err_q_t0[0];
assign _071_ = valid_q_t0[0] & in_valid_i_t0;
assign _074_ = valid_q_t0[1] & valid_q_t0[0];
assign _077_ = valid_popped_t0[0] & clear_i_t0;
assign _080_ = valid_popped_t0[1] & clear_i_t0;
assign _086_ = in_valid_i_t0 & lowest_free_entry_t0[1];
assign _089_ = valid_q_t0[2] & valid_q_t0[1];
assign _092_ = valid_popped_t0[2] & clear_i_t0;
assign _095_ = in_valid_i_t0 & lowest_free_entry_t0[2];
assign _163_ = _051_ | _052_;
assign _164_ = _054_ | _055_;
assign _165_ = _057_ | _058_;
assign _166_ = _060_ | _061_;
assign _167_ = _063_ | _064_;
assign _168_ = _066_ | _067_;
assign _169_ = _069_ | _070_;
assign _170_ = _072_ | _073_;
assign _171_ = _075_ | _076_;
assign _172_ = _078_ | _079_;
assign _173_ = _082_ | _069_;
assign _174_ = _084_ | _085_;
assign _175_ = _087_ | _088_;
assign _176_ = _090_ | _091_;
assign _177_ = _093_ | _094_;
assign _003_ = _163_ | _053_;
assign _005_ = _164_ | _056_;
assign _007_ = _165_ | _059_;
assign _009_ = _166_ | _062_;
assign _011_ = _167_ | _065_;
assign _013_ = _168_ | _068_;
assign _015_ = _169_ | _071_;
assign lowest_free_entry_t0[1] = _170_ | _074_;
assign valid_d_t0[0] = _171_ | _077_;
assign valid_d_t0[1] = _172_ | _080_;
assign _018_ = _173_ | _071_;
assign _020_ = _174_ | _086_;
assign lowest_free_entry_t0[2] = _175_ | _089_;
assign valid_d_t0[2] = _176_ | _092_;
assign entry_en_t0[2] = _177_ | _095_;
/* src = "generated/sv2v_out.v:16220.5-16228.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q[2] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q[2] <= 1'h0;
else if (entry_en[2]) err_q[2] <= in_err_i;
/* src = "generated/sv2v_out.v:16220.5-16228.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q[95:64] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q[95:64] <= 32'd0;
else if (entry_en[2]) rdata_q[95:64] <= in_rdata_i;
/* src = "generated/sv2v_out.v:16220.5-16228.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q[1] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q[1] <= 1'h0;
else if (entry_en[1]) err_q[1] <= err_d[1];
/* src = "generated/sv2v_out.v:16220.5-16228.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q[63:32] <= 32'd0;
else if (entry_en[1]) rdata_q[63:32] <= rdata_d[63:32];
/* src = "generated/sv2v_out.v:16220.5-16228.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q[0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q[0] <= 1'h0;
else if (entry_en[0]) err_q[0] <= err_d[0];
/* src = "generated/sv2v_out.v:16220.5-16228.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q[31:0] <= 32'd0;
else if (entry_en[0]) rdata_q[31:0] <= rdata_d[31:0];
/* src = "generated/sv2v_out.v:16172.4-16176.35" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME instr_addr_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_addr_q <= 31'h00000000;
else if (instr_addr_en) instr_addr_q <= instr_addr_d;
assign _031_ = ~ unaligned_is_compressed;
assign _032_ = ~ instr_addr_q[1];
assign _033_ = ~ { instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1] };
assign _034_ = ~ { valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0] };
assign lowest_free_entry[0] = ~ valid_q[0];
assign _035_ = ~ { valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1] };
assign _036_ = ~ valid_q[1];
assign _037_ = ~ { clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i };
assign _038_ = ~ pop_fifo;
assign _039_ = ~ { valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2] };
assign _040_ = ~ valid_q[2];
assign _130_ = _031_ & valid_unaligned_t0;
assign _132_ = _032_ & valid_t0;
assign _134_ = _032_ & err_t0;
assign _136_ = _033_ & rdata_t0;
assign _138_ = _034_ & in_rdata_i_t0;
assign _140_ = lowest_free_entry[0] & in_err_i_t0;
assign _141_ = _035_ & { in_rdata_i_t0[15:0], rdata_t0[31:16] };
assign _143_ = _036_ & _205_;
assign _145_ = _036_ & _013_;
assign valid_unaligned_t0 = _036_ & _015_;
assign _120_ = _032_ & aligned_is_compressed_t0;
assign _148_ = _037_ & instr_addr_next_t0;
assign _150_ = _038_ & valid_pushed_t0[0];
assign _151_ = _038_ & valid_pushed_t0[1];
assign _152_ = _035_ & in_rdata_i_t0;
assign _154_ = _039_ & in_rdata_i_t0;
assign _156_ = _036_ & in_err_i_t0;
assign _158_ = _040_ & in_err_i_t0;
assign valid_popped_t0[2] = _038_ & valid_pushed_t0[2];
assign _131_ = unaligned_is_compressed & valid_t0;
assign _133_ = instr_addr_q[1] & _001_;
assign out_err_plus2_o_t0 = instr_addr_q[1] & err_plus2_t0;
assign _135_ = instr_addr_q[1] & err_unaligned_t0;
assign _137_ = { instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1] } & rdata_unaligned_t0;
assign _139_ = { valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0] } & rdata_q_t0[31:0];
assign _142_ = { valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1] } & { rdata_q_t0[47:32], rdata_t0[31:16] };
assign _144_ = valid_q[1] & _201_;
assign _146_ = valid_q[1] & _009_;
assign _147_ = instr_addr_q[1] & unaligned_is_compressed_t0;
assign _149_ = { clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i } & in_addr_i_t0[31:1];
assign _153_ = { valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1] } & rdata_q_t0[63:32];
assign _155_ = { valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2] } & rdata_q_t0[95:64];
assign _157_ = valid_q[1] & err_q_t0[1];
assign _159_ = valid_q[2] & err_q_t0[2];
assign _001_ = _130_ | _131_;
assign out_valid_o_t0 = _132_ | _133_;
assign out_err_o_t0 = _134_ | _135_;
assign out_rdata_o_t0 = _136_ | _137_;
assign rdata_t0 = _138_ | _139_;
assign err_t0 = _140_ | _055_;
assign rdata_unaligned_t0 = _141_ | _142_;
assign err_unaligned_t0 = _143_ | _144_;
assign err_plus2_t0 = _145_ | _146_;
assign addr_incr_two_t0 = _120_ | _147_;
assign instr_addr_d_t0 = _148_ | _149_;
assign valid_popped_t0[0] = _150_ | _081_;
assign valid_popped_t0[1] = _151_ | _083_;
assign rdata_d_t0[31:0] = _152_ | _153_;
assign rdata_d_t0[63:32] = _154_ | _155_;
assign err_d_t0[0] = _156_ | _157_;
assign err_d_t0[1] = _158_ | _159_;
assign _041_ = ~ _002_;
assign _042_ = ~ _004_;
assign _043_ = ~ clear_i;
assign _044_ = ~ _017_;
assign _045_ = ~ _019_;
assign _046_ = ~ in_valid_i;
assign _047_ = ~ err_q[0];
assign _048_ = ~ _006_;
assign _110_ = valid_q_t0[0] & _046_;
assign _111_ = _003_ & _047_;
assign _114_ = valid_q_t0[0] & unaligned_is_compressed;
assign _117_ = _005_ & _048_;
assign _121_ = _018_ & lowest_free_entry[0];
assign _124_ = _020_ & _036_;
assign _127_ = valid_q_t0[2] & _027_;
assign _112_ = err_q_t0[0] & _041_;
assign _115_ = unaligned_is_compressed_t0 & valid_q[0];
assign _118_ = _007_ & _042_;
assign _122_ = valid_q_t0[0] & _044_;
assign _125_ = valid_q_t0[1] & _045_;
assign _128_ = entry_en_t0[2] & _040_;
assign _113_ = _003_ & err_q_t0[0];
assign _116_ = valid_q_t0[0] & unaligned_is_compressed_t0;
assign _119_ = _005_ & _007_;
assign _123_ = _018_ & valid_q_t0[0];
assign _126_ = _020_ & valid_q_t0[1];
assign _129_ = valid_q_t0[2] & entry_en_t0[2];
assign _185_ = _110_ | _082_;
assign _186_ = _111_ | _112_;
assign _187_ = _114_ | _115_;
assign _188_ = _117_ | _118_;
assign _189_ = _121_ | _122_;
assign _190_ = _124_ | _125_;
assign _191_ = _127_ | _128_;
assign valid_t0 = _185_ | _071_;
assign _201_ = _186_ | _113_;
assign _203_ = _187_ | _116_;
assign _205_ = _188_ | _119_;
assign valid_pushed_t0[0] = _189_ | _123_;
assign valid_pushed_t0[1] = _190_ | _126_;
assign valid_pushed_t0[2] = _191_ | _129_;
assign _195_ = rdata[17:16] != /* src = "generated/sv2v_out.v:16148.36-16148.57" */ 2'h3;
assign _196_ = rdata[1:0] != /* src = "generated/sv2v_out.v:16149.34-16149.53" */ 2'h3;
assign _197_ = ~ /* src = "generated/sv2v_out.v:16149.57-16149.61" */ err;
assign _198_ = ~ /* src = "generated/sv2v_out.v:16168.56-16168.70" */ addr_incr_two;
assign _199_ = ~ /* src = "generated/sv2v_out.v:16187.51-16187.73" */ aligned_is_compressed;
assign valid = valid_q[0] | /* src = "generated/sv2v_out.v:16143.17-16143.40" */ in_valid_i;
assign _200_ = _002_ | /* src = "generated/sv2v_out.v:16145.39-16145.87" */ err_q[0];
assign _202_ = lowest_free_entry[0] | /* src = "generated/sv2v_out.v:16145.129-16145.167" */ _031_;
assign _204_ = _004_ | /* src = "generated/sv2v_out.v:16145.90-16145.169" */ _006_;
assign instr_addr_en = clear_i | /* src = "generated/sv2v_out.v:16166.25-16166.62" */ _016_;
assign _206_ = _199_ | /* src = "generated/sv2v_out.v:16187.51-16187.89" */ instr_addr_q[1];
assign valid_pushed[0] = _017_ | /* src = "generated/sv2v_out.v:16197.29-16197.77" */ valid_q[0];
assign valid_pushed[1] = _019_ | /* src = "generated/sv2v_out.v:16197.29-16197.77" */ valid_q[1];
assign entry_en[0] = _021_ | /* src = "generated/sv2v_out.v:16200.25-16200.109" */ _022_;
assign entry_en[1] = _023_ | /* src = "generated/sv2v_out.v:16200.25-16200.109" */ _024_;
assign valid_pushed[2] = valid_q[2] | /* src = "generated/sv2v_out.v:16206.35-16206.99" */ entry_en[2];
/* src = "generated/sv2v_out.v:16212.2-16216.23" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME valid_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) valid_q <= 3'h0;
else valid_q <= valid_d;
assign _000_ = unaligned_is_compressed ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:16155.8-16155.31|generated/sv2v_out.v:16155.4-16158.35" */ valid : valid_unaligned;
assign out_valid_o = instr_addr_q[1] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:16151.7-16151.20|generated/sv2v_out.v:16151.3-16165.6" */ _000_ : valid;
assign out_err_plus2_o = instr_addr_q[1] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:16151.7-16151.20|generated/sv2v_out.v:16151.3-16165.6" */ err_plus2 : 1'h0;
assign out_err_o = instr_addr_q[1] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:16151.7-16151.20|generated/sv2v_out.v:16151.3-16165.6" */ err_unaligned : err;
assign out_rdata_o = instr_addr_q[1] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:16151.7-16151.20|generated/sv2v_out.v:16151.3-16165.6" */ rdata_unaligned : rdata;
assign rdata = valid_q[0] ? /* src = "generated/sv2v_out.v:16141.18-16141.58" */ rdata_q[31:0] : in_rdata_i;
assign err = valid_q[0] ? /* src = "generated/sv2v_out.v:16142.16-16142.48" */ err_q[0] : in_err_i;
assign rdata_unaligned = valid_q[1] ? /* src = "generated/sv2v_out.v:16144.28-16144.107" */ { rdata_q[47:32], rdata[31:16] } : { in_rdata_i[15:0], rdata[31:16] };
assign err_unaligned = valid_q[1] ? /* src = "generated/sv2v_out.v:16145.26-16145.169" */ _200_ : _204_;
assign err_plus2 = valid_q[1] ? /* src = "generated/sv2v_out.v:16146.22-16146.93" */ _008_ : _012_;
assign valid_unaligned = valid_q[1] ? /* src = "generated/sv2v_out.v:16147.28-16147.71" */ 1'h1 : _014_;
assign addr_incr_two = instr_addr_q[1] ? /* src = "generated/sv2v_out.v:16167.26-16167.91" */ unaligned_is_compressed : aligned_is_compressed;
assign instr_addr_d = clear_i ? /* src = "generated/sv2v_out.v:16169.25-16169.68" */ in_addr_i[31:1] : instr_addr_next;
assign valid_popped[0] = pop_fifo ? /* src = "generated/sv2v_out.v:16198.30-16198.78" */ valid_pushed[1] : valid_pushed[0];
assign valid_popped[1] = pop_fifo ? /* src = "generated/sv2v_out.v:16198.30-16198.78" */ valid_pushed[2] : valid_pushed[1];
assign rdata_d[31:0] = valid_q[1] ? /* src = "generated/sv2v_out.v:16201.34-16201.89" */ rdata_q[63:32] : in_rdata_i;
assign rdata_d[63:32] = valid_q[2] ? /* src = "generated/sv2v_out.v:16201.34-16201.89" */ rdata_q[95:64] : in_rdata_i;
assign err_d[0] = valid_q[1] ? /* src = "generated/sv2v_out.v:16202.23-16202.63" */ err_q[1] : in_err_i;
assign err_d[1] = valid_q[2] ? /* src = "generated/sv2v_out.v:16202.23-16202.63" */ err_q[2] : in_err_i;
assign valid_popped[2] = pop_fifo ? /* src = "generated/sv2v_out.v:16207.36-16207.77" */ 1'h0 : valid_pushed[2];
assign busy_o = valid_q[2:1];
assign busy_o_t0 = valid_q_t0[2:1];
assign err_d[2] = in_err_i;
assign err_d_t0[2] = in_err_i_t0;
assign lowest_free_entry_t0[0] = valid_q_t0[0];
assign out_addr_o = { instr_addr_q, 1'h0 };
assign out_addr_o_t0 = { instr_addr_q_t0, 1'h0 };
assign rdata_d[95:64] = in_rdata_i;
assign rdata_d_t0[95:64] = in_rdata_i_t0;
endmodule

module \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111 (clk_i, rst_ni, data_req_o, data_gnt_i, data_rvalid_i, data_bus_err_i, data_pmp_err_i, data_addr_o, data_we_o, data_be_o, data_wdata_o, data_rdata_i, lsu_we_i, lsu_type_i, lsu_wdata_i, lsu_sign_ext_i, lsu_rdata_o, lsu_rdata_valid_o, lsu_req_i, adder_result_ex_i, addr_incr_req_o
, addr_last_o, lsu_req_done_o, lsu_resp_valid_o, load_err_o, load_resp_intg_err_o, store_err_o, store_resp_intg_err_o, busy_o, perf_load_o, perf_store_o, data_we_o_t0, data_req_o_t0, store_resp_intg_err_o_t0, store_err_o_t0, perf_store_o_t0, perf_load_o_t0, lsu_we_i_t0, lsu_wdata_i_t0, lsu_type_i_t0, lsu_sign_ext_i_t0, lsu_resp_valid_o_t0
, lsu_req_i_t0, lsu_req_done_o_t0, lsu_rdata_valid_o_t0, lsu_rdata_o_t0, data_rdata_i_t0, data_pmp_err_i_t0, data_gnt_i_t0, data_bus_err_i_t0, data_be_o_t0, data_addr_o_t0, addr_last_o_t0, addr_incr_req_o_t0, adder_result_ex_i_t0, load_resp_intg_err_o_t0, load_err_o_t0, data_rvalid_i_t0, data_wdata_o_t0, busy_o_t0);
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _000_;
/* src = "generated/sv2v_out.v:18438.2-18477.10" */
wire [3:0] _001_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _002_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _003_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire [2:0] _004_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _005_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _007_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _008_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _009_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _010_;
/* src = "generated/sv2v_out.v:18542.2-18565.10" */
wire [31:0] _011_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18542.2-18565.10" */
wire [31:0] _012_;
/* src = "generated/sv2v_out.v:18518.2-18541.10" */
wire [31:0] _013_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18518.2-18541.10" */
wire [31:0] _014_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _015_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _016_;
/* src = "generated/sv2v_out.v:18438.2-18477.10" */
wire [3:0] _017_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _018_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire [2:0] _019_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _021_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _022_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _023_;
/* src = "generated/sv2v_out.v:18542.2-18565.10" */
wire [31:0] _024_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18542.2-18565.10" */
wire [31:0] _025_;
/* src = "generated/sv2v_out.v:18518.2-18541.10" */
wire [31:0] _026_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18518.2-18541.10" */
wire [31:0] _027_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _028_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _029_;
/* src = "generated/sv2v_out.v:18438.2-18477.10" */
wire [3:0] _030_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _031_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire [2:0] _032_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _033_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _034_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _035_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _036_;
/* src = "generated/sv2v_out.v:18542.2-18565.10" */
wire [31:0] _037_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18542.2-18565.10" */
wire [31:0] _038_;
/* src = "generated/sv2v_out.v:18518.2-18541.10" */
wire [31:0] _039_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18518.2-18541.10" */
wire [31:0] _040_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _041_;
/* src = "generated/sv2v_out.v:18438.2-18477.10" */
wire [3:0] _042_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _043_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _044_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire [2:0] _045_;
/* src = "generated/sv2v_out.v:18542.2-18565.10" */
wire [31:0] _046_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18542.2-18565.10" */
wire [31:0] _047_;
/* src = "generated/sv2v_out.v:18518.2-18541.10" */
wire [31:0] _048_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18518.2-18541.10" */
wire [31:0] _049_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _050_;
/* src = "generated/sv2v_out.v:18438.2-18477.10" */
wire [3:0] _051_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _052_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire [2:0] _053_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _054_;
/* src = "generated/sv2v_out.v:18438.2-18477.10" */
wire [3:0] _055_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire _056_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire [2:0] _057_;
/* src = "generated/sv2v_out.v:18592.2-18670.5" */
wire [2:0] _058_;
/* src = "generated/sv2v_out.v:18640.20-18640.62" */
wire _059_;
/* src = "generated/sv2v_out.v:18687.32-18687.67" */
wire _060_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18687.32-18687.67" */
wire _061_;
/* src = "generated/sv2v_out.v:18687.31-18687.87" */
wire _062_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18687.31-18687.87" */
wire _063_;
/* src = "generated/sv2v_out.v:18687.30-18687.101" */
wire _064_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18687.30-18687.101" */
wire _065_;
/* src = "generated/sv2v_out.v:18705.23-18705.51" */
wire _066_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18705.23-18705.51" */
wire _067_;
/* src = "generated/sv2v_out.v:18706.24-18706.51" */
wire _068_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18706.24-18706.51" */
wire _069_;
/* src = "generated/sv2v_out.v:18707.33-18707.62" */
wire _070_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18707.33-18707.62" */
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire [31:0] _082_;
wire [31:0] _083_;
wire [31:0] _084_;
wire [31:0] _085_;
wire [31:0] _086_;
wire [31:0] _087_;
wire [31:0] _088_;
wire [31:0] _089_;
wire _090_;
wire _091_;
wire [31:0] _092_;
wire [31:0] _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire [23:0] _143_;
wire [23:0] _144_;
wire [31:0] _145_;
wire [31:0] _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire [31:0] _153_;
wire [31:0] _154_;
wire [31:0] _155_;
wire [31:0] _156_;
wire [31:0] _157_;
wire [31:0] _158_;
wire [31:0] _159_;
wire [31:0] _160_;
wire [31:0] _161_;
wire [31:0] _162_;
wire [31:0] _163_;
wire [31:0] _164_;
wire [31:0] _165_;
wire [31:0] _166_;
wire [31:0] _167_;
wire [31:0] _168_;
wire [31:0] _169_;
wire [31:0] _170_;
wire [31:0] _171_;
wire [31:0] _172_;
wire [31:0] _173_;
wire [31:0] _174_;
wire [31:0] _175_;
wire [31:0] _176_;
wire [31:0] _177_;
wire [31:0] _178_;
wire [31:0] _179_;
wire [31:0] _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire [31:0] _193_;
wire [31:0] _194_;
wire [31:0] _195_;
wire [31:0] _196_;
wire [31:0] _197_;
wire [31:0] _198_;
wire [31:0] _199_;
wire [31:0] _200_;
wire [31:0] _201_;
wire [31:0] _202_;
wire [31:0] _203_;
wire [31:0] _204_;
wire [31:0] _205_;
wire [31:0] _206_;
wire [31:0] _207_;
wire [31:0] _208_;
wire [31:0] _209_;
wire [31:0] _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire [23:0] _226_;
wire [31:0] _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire [2:0] _232_;
wire [2:0] _233_;
wire [2:0] _234_;
wire [2:0] _235_;
wire _236_;
/* cellift = 32'd1 */
wire _237_;
wire _238_;
/* cellift = 32'd1 */
wire _239_;
wire _240_;
/* cellift = 32'd1 */
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
/* cellift = 32'd1 */
wire _250_;
wire [31:0] _251_;
/* cellift = 32'd1 */
wire [31:0] _252_;
wire [31:0] _253_;
/* cellift = 32'd1 */
wire [31:0] _254_;
wire [31:0] _255_;
/* cellift = 32'd1 */
wire [31:0] _256_;
wire [31:0] _257_;
/* cellift = 32'd1 */
wire [31:0] _258_;
wire [31:0] _259_;
/* cellift = 32'd1 */
wire [31:0] _260_;
wire [31:0] _261_;
/* cellift = 32'd1 */
wire [31:0] _262_;
wire [31:0] _263_;
/* cellift = 32'd1 */
wire [31:0] _264_;
wire [31:0] _265_;
/* cellift = 32'd1 */
wire [31:0] _266_;
wire [31:0] _267_;
/* cellift = 32'd1 */
wire [31:0] _268_;
wire [3:0] _269_;
wire [3:0] _270_;
wire [3:0] _271_;
wire [3:0] _272_;
wire [3:0] _273_;
wire [3:0] _274_;
wire [3:0] _275_;
wire [3:0] _276_;
/* src = "generated/sv2v_out.v:18591.37-18591.56" */
wire _277_;
/* src = "generated/sv2v_out.v:18591.90-18591.109" */
wire _278_;
/* src = "generated/sv2v_out.v:18591.115-18591.135" */
wire _279_;
/* src = "generated/sv2v_out.v:18671.63-18671.80" */
wire _280_;
/* src = "generated/sv2v_out.v:18686.59-18686.76" */
wire _281_;
/* src = "generated/sv2v_out.v:18591.36-18591.83" */
wire _282_;
/* src = "generated/sv2v_out.v:18591.89-18591.136" */
wire _283_;
/* src = "generated/sv2v_out.v:18625.9-18625.32" */
wire _284_;
/* src = "generated/sv2v_out.v:18635.9-18635.35" */
wire _285_;
/* src = "generated/sv2v_out.v:18591.62-18591.82" */
wire _286_;
/* src = "generated/sv2v_out.v:18611.20-18611.29" */
wire _287_;
/* src = "generated/sv2v_out.v:18638.21-18638.31" */
wire _288_;
/* src = "generated/sv2v_out.v:18640.33-18640.62" */
wire _289_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18640.33-18640.62" */
wire _290_;
/* src = "generated/sv2v_out.v:18687.71-18687.87" */
wire _291_;
/* src = "generated/sv2v_out.v:18687.105-18687.119" */
wire _292_;
/* src = "generated/sv2v_out.v:18637.18-18637.44" */
wire _293_;
/* src = "generated/sv2v_out.v:18671.27-18671.58" */
wire _294_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18671.27-18671.58" */
wire _295_;
/* src = "generated/sv2v_out.v:18685.28-18685.54" */
wire _296_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18685.28-18685.54" */
wire _297_;
/* src = "generated/sv2v_out.v:18686.29-18686.54" */
wire _298_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18686.29-18686.54" */
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire [1:0] _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire [1:0] _312_;
wire _313_;
/* src = "generated/sv2v_out.v:18617.20-18617.57" */
wire [2:0] _314_;
/* src = "generated/sv2v_out.v:18620.20-18620.57" */
wire [2:0] _315_;
/* src = "generated/sv2v_out.v:18639.19-18639.43" */
wire [2:0] _316_;
/* src = "generated/sv2v_out.v:18394.20-18394.37" */
input [31:0] adder_result_ex_i;
wire [31:0] adder_result_ex_i;
/* cellift = 32'd1 */
input [31:0] adder_result_ex_i_t0;
wire [31:0] adder_result_ex_i_t0;
/* src = "generated/sv2v_out.v:18395.13-18395.28" */
output addr_incr_req_o;
wire addr_incr_req_o;
/* cellift = 32'd1 */
output addr_incr_req_o_t0;
wire addr_incr_req_o_t0;
/* src = "generated/sv2v_out.v:18409.14-18409.25" */
wire [31:0] addr_last_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18409.14-18409.25" */
wire [31:0] addr_last_d_t0;
/* src = "generated/sv2v_out.v:18396.21-18396.32" */
output [31:0] addr_last_o;
reg [31:0] addr_last_o;
/* cellift = 32'd1 */
output [31:0] addr_last_o_t0;
reg [31:0] addr_last_o_t0;
/* src = "generated/sv2v_out.v:18410.6-18410.17" */
wire addr_update;
/* src = "generated/sv2v_out.v:18403.14-18403.20" */
output busy_o;
wire busy_o;
/* cellift = 32'd1 */
output busy_o_t0;
wire busy_o_t0;
/* src = "generated/sv2v_out.v:18375.13-18375.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:18411.6-18411.17" */
wire ctrl_update;
/* src = "generated/sv2v_out.v:18382.21-18382.32" */
output [31:0] data_addr_o;
wire [31:0] data_addr_o;
/* cellift = 32'd1 */
output [31:0] data_addr_o_t0;
wire [31:0] data_addr_o_t0;
/* src = "generated/sv2v_out.v:18384.20-18384.29" */
output [3:0] data_be_o;
wire [3:0] data_be_o;
/* cellift = 32'd1 */
output [3:0] data_be_o_t0;
wire [3:0] data_be_o_t0;
/* src = "generated/sv2v_out.v:18380.13-18380.27" */
input data_bus_err_i;
wire data_bus_err_i;
/* cellift = 32'd1 */
input data_bus_err_i_t0;
wire data_bus_err_i_t0;
/* src = "generated/sv2v_out.v:18378.13-18378.23" */
input data_gnt_i;
wire data_gnt_i;
/* cellift = 32'd1 */
input data_gnt_i_t0;
wire data_gnt_i_t0;
/* src = "generated/sv2v_out.v:18432.7-18432.20" */
wire data_intg_err;
/* src = "generated/sv2v_out.v:18433.7-18433.22" */
wire data_or_pmp_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18433.7-18433.22" */
wire data_or_pmp_err_t0;
/* src = "generated/sv2v_out.v:18381.13-18381.27" */
input data_pmp_err_i;
wire data_pmp_err_i;
/* cellift = 32'd1 */
input data_pmp_err_i_t0;
wire data_pmp_err_i_t0;
/* src = "generated/sv2v_out.v:18386.34-18386.46" */
input [38:0] data_rdata_i;
wire [38:0] data_rdata_i;
/* cellift = 32'd1 */
input [38:0] data_rdata_i_t0;
wire [38:0] data_rdata_i_t0;
/* src = "generated/sv2v_out.v:18377.13-18377.23" */
output data_req_o;
wire data_req_o;
/* cellift = 32'd1 */
output data_req_o_t0;
wire data_req_o_t0;
/* src = "generated/sv2v_out.v:18379.13-18379.26" */
input data_rvalid_i;
wire data_rvalid_i;
/* cellift = 32'd1 */
input data_rvalid_i_t0;
wire data_rvalid_i_t0;
/* src = "generated/sv2v_out.v:18416.6-18416.21" */
reg data_sign_ext_q;
/* src = "generated/sv2v_out.v:18415.12-18415.23" */
reg [1:0] data_type_q;
/* src = "generated/sv2v_out.v:18420.13-18420.23" */
wire [31:0] data_wdata;
/* src = "generated/sv2v_out.v:18385.35-18385.47" */
output [38:0] data_wdata_o;
wire [38:0] data_wdata_o;
/* cellift = 32'd1 */
output [38:0] data_wdata_o_t0;
wire [38:0] data_wdata_o_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18420.13-18420.23" */
wire [31:0] data_wdata_t0;
/* src = "generated/sv2v_out.v:18383.14-18383.23" */
output data_we_o;
wire data_we_o;
/* cellift = 32'd1 */
output data_we_o_t0;
wire data_we_o_t0;
/* src = "generated/sv2v_out.v:18417.6-18417.15" */
reg data_we_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18417.6-18417.15" */
reg data_we_q_t0;
/* src = "generated/sv2v_out.v:18576.30-18576.44" */
wire [38:0] \g_mem_rdata_ecc.data_rdata_buf ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18576.30-18576.44" */
wire [38:0] \g_mem_rdata_ecc.data_rdata_buf_t0 ;
/* src = "generated/sv2v_out.v:18575.15-18575.22" */
wire [1:0] \g_mem_rdata_ecc.ecc_err ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18575.15-18575.22" */
/* unused_bits = "0 1" */
wire [1:0] \g_mem_rdata_ecc.ecc_err_t0 ;
/* src = "generated/sv2v_out.v:18427.6-18427.25" */
wire handle_misaligned_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18427.6-18427.25" */
wire handle_misaligned_d_t0;
/* src = "generated/sv2v_out.v:18426.6-18426.25" */
reg handle_misaligned_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18426.6-18426.25" */
reg handle_misaligned_q_t0;
/* src = "generated/sv2v_out.v:18399.14-18399.24" */
output load_err_o;
wire load_err_o;
/* cellift = 32'd1 */
output load_err_o_t0;
wire load_err_o_t0;
/* src = "generated/sv2v_out.v:18400.14-18400.34" */
output load_resp_intg_err_o;
wire load_resp_intg_err_o;
/* cellift = 32'd1 */
output load_resp_intg_err_o_t0;
wire load_resp_intg_err_o_t0;
/* src = "generated/sv2v_out.v:18434.12-18434.21" */
reg [2:0] ls_fsm_cs;
/* src = "generated/sv2v_out.v:18435.12-18435.21" */
wire [2:0] ls_fsm_ns;
/* src = "generated/sv2v_out.v:18431.6-18431.15" */
wire lsu_err_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18431.6-18431.15" */
wire lsu_err_d_t0;
/* src = "generated/sv2v_out.v:18430.6-18430.15" */
reg lsu_err_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18430.6-18430.15" */
reg lsu_err_q_t0;
/* src = "generated/sv2v_out.v:18391.21-18391.32" */
output [31:0] lsu_rdata_o;
wire [31:0] lsu_rdata_o;
/* cellift = 32'd1 */
output [31:0] lsu_rdata_o_t0;
wire [31:0] lsu_rdata_o_t0;
/* src = "generated/sv2v_out.v:18392.14-18392.31" */
output lsu_rdata_valid_o;
wire lsu_rdata_valid_o;
/* cellift = 32'd1 */
output lsu_rdata_valid_o_t0;
wire lsu_rdata_valid_o_t0;
/* src = "generated/sv2v_out.v:18397.14-18397.28" */
output lsu_req_done_o;
wire lsu_req_done_o;
/* cellift = 32'd1 */
output lsu_req_done_o_t0;
wire lsu_req_done_o_t0;
/* src = "generated/sv2v_out.v:18393.13-18393.22" */
input lsu_req_i;
wire lsu_req_i;
/* cellift = 32'd1 */
input lsu_req_i_t0;
wire lsu_req_i_t0;
/* src = "generated/sv2v_out.v:18398.14-18398.30" */
output lsu_resp_valid_o;
wire lsu_resp_valid_o;
/* cellift = 32'd1 */
output lsu_resp_valid_o_t0;
wire lsu_resp_valid_o_t0;
/* src = "generated/sv2v_out.v:18390.13-18390.27" */
input lsu_sign_ext_i;
wire lsu_sign_ext_i;
/* cellift = 32'd1 */
input lsu_sign_ext_i_t0;
wire lsu_sign_ext_i_t0;
/* src = "generated/sv2v_out.v:18388.19-18388.29" */
input [1:0] lsu_type_i;
wire [1:0] lsu_type_i;
/* cellift = 32'd1 */
input [1:0] lsu_type_i_t0;
wire [1:0] lsu_type_i_t0;
/* src = "generated/sv2v_out.v:18389.20-18389.31" */
input [31:0] lsu_wdata_i;
wire [31:0] lsu_wdata_i;
/* cellift = 32'd1 */
input [31:0] lsu_wdata_i_t0;
wire [31:0] lsu_wdata_i_t0;
/* src = "generated/sv2v_out.v:18387.13-18387.21" */
input lsu_we_i;
wire lsu_we_i;
/* cellift = 32'd1 */
input lsu_we_i_t0;
wire lsu_we_i_t0;
/* src = "generated/sv2v_out.v:18404.13-18404.24" */
output perf_load_o;
wire perf_load_o;
/* cellift = 32'd1 */
output perf_load_o_t0;
wire perf_load_o_t0;
/* src = "generated/sv2v_out.v:18405.13-18405.25" */
output perf_store_o;
wire perf_store_o;
/* cellift = 32'd1 */
output perf_store_o_t0;
wire perf_store_o_t0;
/* src = "generated/sv2v_out.v:18429.6-18429.15" */
wire pmp_err_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18429.6-18429.15" */
wire pmp_err_d_t0;
/* src = "generated/sv2v_out.v:18428.6-18428.15" */
reg pmp_err_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18428.6-18428.15" */
reg pmp_err_q_t0;
/* src = "generated/sv2v_out.v:18424.13-18424.24" */
wire [31:0] rdata_b_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18424.13-18424.24" */
wire [31:0] rdata_b_ext_t0;
/* src = "generated/sv2v_out.v:18423.13-18423.24" */
wire [31:0] rdata_h_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18423.13-18423.24" */
wire [31:0] rdata_h_ext_t0;
/* src = "generated/sv2v_out.v:18414.12-18414.26" */
reg [1:0] rdata_offset_q;
/* src = "generated/sv2v_out.v:18413.13-18413.20" */
reg [31:8] rdata_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18413.13-18413.20" */
reg [31:8] rdata_q_t0;
/* src = "generated/sv2v_out.v:18412.6-18412.18" */
wire rdata_update;
/* src = "generated/sv2v_out.v:18422.13-18422.24" */
wire [31:0] rdata_w_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18422.13-18422.24" */
wire [31:0] rdata_w_ext_t0;
/* src = "generated/sv2v_out.v:18376.13-18376.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:18425.7-18425.30" */
wire split_misaligned_access;
/* src = "generated/sv2v_out.v:18401.14-18401.25" */
output store_err_o;
wire store_err_o;
/* cellift = 32'd1 */
output store_err_o_t0;
wire store_err_o_t0;
/* src = "generated/sv2v_out.v:18402.14-18402.35" */
output store_resp_intg_err_o;
wire store_resp_intg_err_o;
/* cellift = 32'd1 */
output store_resp_intg_err_o_t0;
wire store_resp_intg_err_o_t0;
assign _059_ = data_gnt_i & /* src = "generated/sv2v_out.v:18640.20-18640.62" */ _289_;
assign lsu_req_done_o = _294_ & /* src = "generated/sv2v_out.v:18671.26-18671.81" */ _280_;
assign lsu_resp_valid_o = _298_ & /* src = "generated/sv2v_out.v:18686.28-18686.77" */ _281_;
assign _060_ = _281_ & /* src = "generated/sv2v_out.v:18687.32-18687.67" */ data_rvalid_i;
assign _062_ = _060_ & /* src = "generated/sv2v_out.v:18687.31-18687.87" */ _291_;
assign _064_ = _062_ & /* src = "generated/sv2v_out.v:18687.30-18687.101" */ _288_;
assign lsu_rdata_valid_o = _064_ & /* src = "generated/sv2v_out.v:18687.29-18687.119" */ _292_;
assign _066_ = data_or_pmp_err & /* src = "generated/sv2v_out.v:18705.23-18705.51" */ _288_;
assign load_err_o = _066_ & /* src = "generated/sv2v_out.v:18705.22-18705.71" */ lsu_resp_valid_o;
assign _068_ = data_or_pmp_err & /* src = "generated/sv2v_out.v:18706.24-18706.51" */ data_we_q;
assign store_err_o = _068_ & /* src = "generated/sv2v_out.v:18706.23-18706.71" */ lsu_resp_valid_o;
assign load_resp_intg_err_o = _070_ & /* src = "generated/sv2v_out.v:18707.32-18707.76" */ _288_;
assign _070_ = data_intg_err & /* src = "generated/sv2v_out.v:18708.34-18708.63" */ data_rvalid_i;
assign store_resp_intg_err_o = _070_ & /* src = "generated/sv2v_out.v:18708.33-18708.76" */ data_we_q;
assign _072_ = ~ _110_;
assign _073_ = ~ ctrl_update;
assign _074_ = ~ _111_;
assign _075_ = ~ _112_;
assign _076_ = ~ rdata_update;
assign _077_ = ~ addr_update;
assign _135_ = _110_ & handle_misaligned_d_t0;
assign _137_ = ctrl_update & lsu_we_i_t0;
assign _139_ = _111_ & pmp_err_d_t0;
assign _141_ = _112_ & lsu_err_d_t0;
assign _143_ = { rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update } & data_rdata_i_t0[31:8];
assign _145_ = { addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update } & addr_last_d_t0;
assign _136_ = _072_ & handle_misaligned_q_t0;
assign _138_ = _073_ & data_we_q_t0;
assign _140_ = _074_ & pmp_err_q_t0;
assign _142_ = _075_ & lsu_err_q_t0;
assign _144_ = { _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_ } & rdata_q_t0;
assign _146_ = { _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_ } & addr_last_o_t0;
assign _222_ = _135_ | _136_;
assign _223_ = _137_ | _138_;
assign _224_ = _139_ | _140_;
assign _225_ = _141_ | _142_;
assign _226_ = _143_ | _144_;
assign _227_ = _145_ | _146_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME handle_misaligned_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) handle_misaligned_q_t0 <= 1'h0;
else handle_misaligned_q_t0 <= _222_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME data_we_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) data_we_q_t0 <= 1'h0;
else data_we_q_t0 <= _223_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME pmp_err_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) pmp_err_q_t0 <= 1'h0;
else pmp_err_q_t0 <= _224_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME lsu_err_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) lsu_err_q_t0 <= 1'h0;
else lsu_err_q_t0 <= _225_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME rdata_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q_t0 <= 24'h000000;
else rdata_q_t0 <= _226_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME addr_last_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) addr_last_o_t0 <= 32'd0;
else addr_last_o_t0 <= _227_;
assign lsu_req_done_o_t0 = _295_ & _280_;
assign lsu_resp_valid_o_t0 = _299_ & _281_;
assign _115_ = _061_ & _291_;
assign _118_ = _063_ & _288_;
assign lsu_rdata_valid_o_t0 = _065_ & _292_;
assign _121_ = data_or_pmp_err_t0 & _288_;
assign _124_ = _067_ & lsu_resp_valid_o;
assign _127_ = data_or_pmp_err_t0 & data_we_q;
assign _128_ = _069_ & lsu_resp_valid_o;
assign _131_ = _071_ & _288_;
assign _134_ = _071_ & data_we_q;
assign _061_ = data_rvalid_i_t0 & _281_;
assign _116_ = data_or_pmp_err_t0 & _060_;
assign _119_ = data_we_q_t0 & _062_;
assign _125_ = lsu_resp_valid_o_t0 & _066_;
assign _122_ = data_we_q_t0 & data_or_pmp_err;
assign _129_ = lsu_resp_valid_o_t0 & _068_;
assign _071_ = data_rvalid_i_t0 & data_intg_err;
assign _132_ = data_we_q_t0 & _070_;
assign _117_ = _061_ & data_or_pmp_err_t0;
assign _120_ = _063_ & data_we_q_t0;
assign _126_ = _067_ & lsu_resp_valid_o_t0;
assign _123_ = data_or_pmp_err_t0 & data_we_q_t0;
assign _130_ = _069_ & lsu_resp_valid_o_t0;
assign _133_ = _071_ & data_we_q_t0;
assign _214_ = _115_ | _116_;
assign _215_ = _118_ | _119_;
assign _216_ = _121_ | _122_;
assign _217_ = _124_ | _125_;
assign _218_ = _127_ | _122_;
assign _219_ = _128_ | _129_;
assign _220_ = _131_ | _132_;
assign _221_ = _134_ | _132_;
assign _063_ = _214_ | _117_;
assign _065_ = _215_ | _120_;
assign _067_ = _216_ | _123_;
assign load_err_o_t0 = _217_ | _126_;
assign _069_ = _218_ | _123_;
assign store_err_o_t0 = _219_ | _130_;
assign load_resp_intg_err_o_t0 = _220_ | _133_;
assign store_resp_intg_err_o_t0 = _221_ | _133_;
/* src = "generated/sv2v_out.v:18672.2-18684.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME handle_misaligned_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) handle_misaligned_q <= 1'h0;
else if (_110_) handle_misaligned_q <= handle_misaligned_d;
/* src = "generated/sv2v_out.v:18491.2-18503.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME data_we_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) data_we_q <= 1'h0;
else if (ctrl_update) data_we_q <= lsu_we_i;
/* src = "generated/sv2v_out.v:18672.2-18684.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME pmp_err_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) pmp_err_q <= 1'h0;
else if (_111_) pmp_err_q <= pmp_err_d;
/* src = "generated/sv2v_out.v:18672.2-18684.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME lsu_err_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) lsu_err_q <= 1'h0;
else if (_112_) lsu_err_q <= lsu_err_d;
/* src = "generated/sv2v_out.v:18486.2-18490.34" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME rdata_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q <= 24'h000000;
else if (rdata_update) rdata_q <= data_rdata_i[31:8];
/* src = "generated/sv2v_out.v:18505.2-18509.31" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME addr_last_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) addr_last_o <= 32'd0;
else if (addr_update) addr_last_o <= addr_last_d;
/* src = "generated/sv2v_out.v:18491.2-18503.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME rdata_offset_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_offset_q <= 2'h0;
else if (ctrl_update) rdata_offset_q <= adder_result_ex_i[1:0];
/* src = "generated/sv2v_out.v:18491.2-18503.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME data_type_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) data_type_q <= 2'h0;
else if (ctrl_update) data_type_q <= lsu_type_i;
/* src = "generated/sv2v_out.v:18491.2-18503.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME data_sign_ext_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) data_sign_ext_q <= 1'h0;
else if (ctrl_update) data_sign_ext_q <= lsu_sign_ext_i;
assign _078_ = ~ _302_;
assign _079_ = ~ _300_;
assign _080_ = ~ _301_;
assign _081_ = ~ _099_;
assign _082_ = ~ { _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_ };
assign _083_ = ~ { _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_ };
assign _084_ = ~ { _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_ };
assign _085_ = ~ { _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_ };
assign _086_ = ~ { _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_ };
assign _087_ = ~ { _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_ };
assign _088_ = ~ { _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_ };
assign _089_ = ~ { _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_ };
assign _090_ = ~ data_rvalid_i;
assign _091_ = ~ data_gnt_i;
assign _092_ = ~ { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q };
assign _093_ = ~ { addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o };
assign _147_ = _079_ & _237_;
assign _149_ = _078_ & _010_;
assign _151_ = _079_ & _239_;
assign _241_ = _080_ & _044_;
assign addr_incr_req_o_t0 = _081_ & _250_;
assign _153_ = _082_ & rdata_w_ext_t0;
assign _155_ = _083_ & _252_;
assign _157_ = _084_ & _038_;
assign _159_ = _085_ & _012_;
assign _161_ = _086_ & _256_;
assign _163_ = _084_ & _040_;
assign _165_ = _085_ & _014_;
assign _167_ = _086_ & _260_;
assign _169_ = _084_ & { data_rdata_i_t0[15:0], rdata_q_t0[31:16] };
assign _171_ = _085_ & data_rdata_i_t0[31:0];
assign _173_ = _086_ & _264_;
assign _175_ = _087_ & { lsu_wdata_i_t0[15:0], lsu_wdata_i_t0[31:16] };
assign _177_ = _088_ & lsu_wdata_i_t0;
assign _179_ = _089_ & _268_;
assign _193_ = _092_ & { 24'h000000, data_rdata_i_t0[31:24] };
assign _195_ = _092_ & { 24'h000000, data_rdata_i_t0[23:16] };
assign _197_ = _092_ & { 24'h000000, data_rdata_i_t0[15:8] };
assign _199_ = _092_ & { 24'h000000, data_rdata_i_t0[7:0] };
assign _201_ = _092_ & { 16'h0000, data_rdata_i_t0[7:0], rdata_q_t0[31:24] };
assign _203_ = _092_ & { 16'h0000, data_rdata_i_t0[31:16] };
assign _205_ = _092_ & { 16'h0000, data_rdata_i_t0[23:8] };
assign _207_ = _092_ & { 16'h0000, data_rdata_i_t0[15:0] };
assign _209_ = _093_ & adder_result_ex_i_t0;
assign _237_ = _302_ & _021_;
assign _148_ = _300_ & _034_;
assign _150_ = _302_ & _023_;
assign _152_ = _300_ & _036_;
assign handle_misaligned_d_t0 = _211_ & _241_;
assign _250_ = _301_ & handle_misaligned_q_t0;
assign _154_ = { _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_ } & rdata_h_ext_t0;
assign _156_ = { _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_ } & rdata_b_ext_t0;
assign _158_ = { _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_ } & _047_;
assign _160_ = { _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_ } & _025_;
assign _162_ = { _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_ } & _254_;
assign _164_ = { _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_ } & _049_;
assign _166_ = { _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_ } & _027_;
assign _168_ = { _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_ } & _258_;
assign _170_ = { _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_ } & { data_rdata_i_t0[23:0], rdata_q_t0[31:24] };
assign _172_ = { _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_ } & { data_rdata_i_t0[7:0], rdata_q_t0 };
assign _174_ = { _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_ } & _262_;
assign _176_ = { _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_ } & { lsu_wdata_i_t0[7:0], lsu_wdata_i_t0[31:8] };
assign _178_ = { _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_ } & { lsu_wdata_i_t0[23:0], lsu_wdata_i_t0[31:24] };
assign _180_ = { _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_ } & _266_;
assign _034_ = data_rvalid_i & data_bus_err_i_t0;
assign _036_ = data_rvalid_i & data_pmp_err_i_t0;
assign _044_ = _285_ & data_gnt_i_t0;
assign _021_ = _285_ & _290_;
assign _023_ = _285_ & data_pmp_err_i_t0;
assign _007_ = lsu_req_i & lsu_we_i_t0;
assign _010_ = lsu_req_i & data_pmp_err_i_t0;
assign perf_load_o_t0 = _281_ & _007_;
assign _194_ = { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q } & { data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31:24] };
assign _196_ = { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q } & { data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23:16] };
assign _198_ = { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q } & { data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15:8] };
assign _200_ = { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q } & { data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7:0] };
assign _202_ = { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q } & { data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7:0], rdata_q_t0[31:24] };
assign _204_ = { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q } & { data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31:16] };
assign _206_ = { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q } & { data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23:8] };
assign _208_ = { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q } & { data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15:0] };
assign _210_ = { addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o } & { adder_result_ex_i_t0[31:2], 2'h0 };
assign lsu_err_d_t0 = _147_ | _148_;
assign _239_ = _149_ | _150_;
assign pmp_err_d_t0 = _151_ | _152_;
assign _252_ = _153_ | _154_;
assign lsu_rdata_o_t0 = _155_ | _156_;
assign _254_ = _157_ | _158_;
assign _256_ = _159_ | _160_;
assign rdata_b_ext_t0 = _161_ | _162_;
assign _258_ = _163_ | _164_;
assign _260_ = _165_ | _166_;
assign rdata_h_ext_t0 = _167_ | _168_;
assign _262_ = _169_ | _170_;
assign _264_ = _171_ | _172_;
assign rdata_w_ext_t0 = _173_ | _174_;
assign _266_ = _175_ | _176_;
assign _268_ = _177_ | _178_;
assign data_wdata_t0 = _179_ | _180_;
assign _047_ = _193_ | _194_;
assign _038_ = _195_ | _196_;
assign _025_ = _197_ | _198_;
assign _012_ = _199_ | _200_;
assign _049_ = _201_ | _202_;
assign _040_ = _203_ | _204_;
assign _027_ = _205_ | _206_;
assign _014_ = _207_ | _208_;
assign addr_last_d_t0 = _209_ | _210_;
assign _101_ = { _281_, lsu_req_i, data_gnt_i } != 3'h6;
assign _102_ = { _302_, _285_, data_gnt_i } != 3'h4;
assign _103_ = { _281_, lsu_req_i } != 2'h2;
assign _104_ = { _303_, _284_ } != 2'h2;
assign _105_ = { _301_, _284_ } != 2'h2;
assign _106_ = | { _302_, _301_, _281_, _303_ };
assign _107_ = { _300_, data_rvalid_i } != 2'h2;
assign _108_ = { _302_, _285_ } != 2'h2;
assign _109_ = | { _302_, _300_, _281_ };
assign _110_ = & { _101_, _103_, _104_, _106_, _105_, _102_ };
assign _111_ = & { _107_, _109_, _108_ };
assign _112_ = & { _103_, _107_, _109_, _108_ };
assign _113_ = | { _303_, _302_, _301_ };
assign _114_ = | { _303_, _301_ };
assign _094_ = ~ data_bus_err_i;
assign _095_ = ~ lsu_err_q;
assign _096_ = ~ _296_;
assign _097_ = ~ pmp_err_q;
assign _098_ = ~ busy_o;
assign _181_ = data_bus_err_i_t0 & _097_;
assign _295_ = lsu_req_i_t0 & _098_;
assign _184_ = lsu_err_q_t0 & _094_;
assign _187_ = _297_ & _097_;
assign _190_ = data_rvalid_i_t0 & _097_;
assign _182_ = pmp_err_q_t0 & _094_;
assign _185_ = data_bus_err_i_t0 & _095_;
assign _188_ = pmp_err_q_t0 & _096_;
assign _191_ = pmp_err_q_t0 & _090_;
assign _183_ = data_bus_err_i_t0 & pmp_err_q_t0;
assign _186_ = lsu_err_q_t0 & data_bus_err_i_t0;
assign _189_ = _297_ & pmp_err_q_t0;
assign _192_ = data_rvalid_i_t0 & pmp_err_q_t0;
assign _228_ = _181_ | _182_;
assign _229_ = _184_ | _185_;
assign _230_ = _187_ | _188_;
assign _231_ = _190_ | _191_;
assign _290_ = _228_ | _183_;
assign _297_ = _229_ | _186_;
assign data_or_pmp_err_t0 = _230_ | _189_;
assign _299_ = _231_ | _192_;
assign _099_ = | { _302_, _300_ };
assign _100_ = | { _302_, _301_, _300_ };
assign _211_ = _302_ | _301_;
assign _212_ = _308_ | _307_;
assign _213_ = _310_ | _279_;
assign _232_ = _301_ ? _057_ : _045_;
assign _233_ = _300_ ? _058_ : _232_;
assign _234_ = _281_ ? _004_ : 3'h0;
assign _235_ = _303_ ? _032_ : _234_;
assign ls_fsm_ns = _100_ ? _233_ : _235_;
assign _236_ = _302_ ? _020_ : _005_;
assign lsu_err_d = _300_ ? _033_ : _236_;
assign _238_ = _302_ ? _022_ : _009_;
assign pmp_err_d = _300_ ? _035_ : _238_;
assign _240_ = _301_ ? _056_ : _043_;
assign _242_ = _303_ ? _031_ : _003_;
assign handle_misaligned_d = _211_ ? _240_ : _242_;
assign ctrl_update = _114_ ? _029_ : _243_;
assign _244_ = _301_ ? _050_ : _041_;
assign _245_ = _300_ ? _054_ : _244_;
assign _243_ = _281_ ? _000_ : 1'h0;
assign _246_ = _303_ ? _029_ : _243_;
assign addr_update = _100_ ? _245_ : _246_;
assign _247_ = _281_ ? _002_ : 1'h0;
assign data_req_o = _113_ ? 1'h1 : _247_;
assign _248_ = _302_ ? _015_ : 1'h0;
assign rdata_update = _300_ ? _028_ : _248_;
assign _249_ = _301_ ? handle_misaligned_q : 1'h0;
assign addr_incr_req_o = _099_ ? 1'h1 : _249_;
assign _251_ = _306_ ? rdata_h_ext : rdata_w_ext;
assign lsu_rdata_o = _305_ ? rdata_b_ext : _251_;
assign _253_ = _307_ ? _046_ : _037_;
assign _255_ = _309_ ? _024_ : _011_;
assign rdata_b_ext = _212_ ? _253_ : _255_;
assign _257_ = _307_ ? _048_ : _039_;
assign _259_ = _309_ ? _026_ : _013_;
assign rdata_h_ext = _212_ ? _257_ : _259_;
assign _261_ = _307_ ? { data_rdata_i[23:0], rdata_q[31:24] } : { data_rdata_i[15:0], rdata_q[31:16] };
assign _263_ = _309_ ? { data_rdata_i[7:0], rdata_q } : data_rdata_i[31:0];
assign rdata_w_ext = _212_ ? _261_ : _263_;
assign _265_ = _279_ ? { lsu_wdata_i[7:0], lsu_wdata_i[31:8] } : { lsu_wdata_i[15:0], lsu_wdata_i[31:16] };
assign _267_ = _311_ ? { lsu_wdata_i[23:0], lsu_wdata_i[31:24] } : lsu_wdata_i;
assign data_wdata = _213_ ? _265_ : _267_;
assign _269_ = _279_ ? 4'h8 : 4'h4;
assign _270_ = _311_ ? 4'h2 : 4'h1;
assign _055_ = _213_ ? _269_ : _270_;
assign _272_ = _311_ ? 4'h6 : 4'h3;
assign _051_ = _213_ ? _271_ : _272_;
assign _273_ = _279_ ? 4'h7 : 4'h3;
assign _274_ = _311_ ? 4'h1 : 4'h0;
assign _030_ = _213_ ? _273_ : _274_;
assign _271_ = _279_ ? 4'h8 : 4'hc;
assign _275_ = _311_ ? 4'he : 4'hf;
assign _017_ = _213_ ? _271_ : _275_;
assign _276_ = _278_ ? _042_ : _001_;
assign data_be_o = _313_ ? _055_ : _276_;
assign _280_ = ! /* src = "generated/sv2v_out.v:18671.63-18671.80" */ ls_fsm_ns;
assign _282_ = _277_ && /* src = "generated/sv2v_out.v:18591.36-18591.83" */ _286_;
assign _283_ = _278_ && /* src = "generated/sv2v_out.v:18591.89-18591.136" */ _279_;
assign split_misaligned_access = _282_ || /* src = "generated/sv2v_out.v:18591.35-18591.137" */ _283_;
assign _285_ = data_rvalid_i || /* src = "generated/sv2v_out.v:18635.9-18635.35" */ pmp_err_q;
assign _284_ = data_gnt_i || /* src = "generated/sv2v_out.v:18651.9-18651.32" */ pmp_err_q;
assign _286_ = | /* src = "generated/sv2v_out.v:18591.62-18591.82" */ adder_result_ex_i[1:0];
assign busy_o = | /* src = "generated/sv2v_out.v:18709.18-18709.35" */ ls_fsm_cs;
assign _287_ = ~ /* src = "generated/sv2v_out.v:18611.20-18611.29" */ lsu_we_i;
assign _289_ = ~ /* src = "generated/sv2v_out.v:18640.33-18640.62" */ _293_;
assign _291_ = ~ /* src = "generated/sv2v_out.v:18687.71-18687.87" */ data_or_pmp_err;
assign _292_ = ~ /* src = "generated/sv2v_out.v:18687.105-18687.119" */ data_intg_err;
assign _288_ = ~ /* src = "generated/sv2v_out.v:18707.66-18707.76" */ data_we_q;
assign _293_ = data_bus_err_i | /* src = "generated/sv2v_out.v:18640.35-18640.61" */ pmp_err_q;
assign _294_ = lsu_req_i | /* src = "generated/sv2v_out.v:18671.27-18671.58" */ busy_o;
assign _296_ = lsu_err_q | /* src = "generated/sv2v_out.v:18685.28-18685.54" */ data_bus_err_i;
assign data_or_pmp_err = _296_ | /* src = "generated/sv2v_out.v:18685.27-18685.67" */ pmp_err_q;
assign _298_ = data_rvalid_i | /* src = "generated/sv2v_out.v:18686.29-18686.54" */ pmp_err_q;
/* src = "generated/sv2v_out.v:18672.2-18684.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME ls_fsm_cs */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) ls_fsm_cs <= 3'h0;
else ls_fsm_cs <= ls_fsm_ns;
assign _058_ = data_rvalid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18660.9-18660.22|generated/sv2v_out.v:18660.5-18666.8" */ 3'h0 : ls_fsm_cs;
assign _028_ = data_rvalid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18660.9-18660.22|generated/sv2v_out.v:18660.5-18666.8" */ _288_ : 1'h0;
assign _054_ = data_rvalid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18660.9-18660.22|generated/sv2v_out.v:18660.5-18666.8" */ _094_ : 1'h0;
assign _033_ = data_rvalid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18660.9-18660.22|generated/sv2v_out.v:18660.5-18666.8" */ data_bus_err_i : 1'hx;
assign _035_ = data_rvalid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18660.9-18660.22|generated/sv2v_out.v:18660.5-18666.8" */ data_pmp_err_i : 1'hx;
assign _056_ = _284_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18651.9-18651.32|generated/sv2v_out.v:18651.5-18656.8" */ 1'h0 : 1'hx;
assign _057_ = _284_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18651.9-18651.32|generated/sv2v_out.v:18651.5-18656.8" */ 3'h0 : ls_fsm_cs;
assign _050_ = _284_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18651.9-18651.32|generated/sv2v_out.v:18651.5-18656.8" */ _095_ : 1'h0;
assign _052_ = data_gnt_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18643.14-18643.24|generated/sv2v_out.v:18643.10-18646.8" */ 1'h0 : 1'hx;
assign _053_ = data_gnt_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18643.14-18643.24|generated/sv2v_out.v:18643.10-18646.8" */ 3'h4 : ls_fsm_cs;
assign _043_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18635.9-18635.35|generated/sv2v_out.v:18635.5-18646.8" */ _091_ : _052_;
assign _041_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18635.9-18635.35|generated/sv2v_out.v:18635.5-18646.8" */ _059_ : 1'h0;
assign _045_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18635.9-18635.35|generated/sv2v_out.v:18635.5-18646.8" */ _316_ : _053_;
assign _015_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18635.9-18635.35|generated/sv2v_out.v:18635.5-18646.8" */ _288_ : 1'h0;
assign _020_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18635.9-18635.35|generated/sv2v_out.v:18635.5-18646.8" */ _293_ : 1'hx;
assign _022_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18635.9-18635.35|generated/sv2v_out.v:18635.5-18646.8" */ data_pmp_err_i : 1'hx;
assign _032_ = _284_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18625.9-18625.32|generated/sv2v_out.v:18625.5-18630.8" */ 3'h2 : ls_fsm_cs;
assign _031_ = _284_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18625.9-18625.32|generated/sv2v_out.v:18625.5-18630.8" */ 1'h1 : 1'hx;
assign _029_ = _284_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18625.9-18625.32|generated/sv2v_out.v:18625.5-18630.8" */ 1'h1 : 1'h0;
assign _019_ = data_gnt_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18613.10-18613.20|generated/sv2v_out.v:18613.6-18620.59" */ _314_ : _315_;
assign _018_ = data_gnt_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18613.10-18613.20|generated/sv2v_out.v:18613.6-18620.59" */ split_misaligned_access : 1'hx;
assign _016_ = data_gnt_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18613.10-18613.20|generated/sv2v_out.v:18613.6-18620.59" */ 1'h1 : 1'h0;
assign _004_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18607.9-18607.18|generated/sv2v_out.v:18607.5-18621.8" */ _019_ : ls_fsm_cs;
assign _003_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18607.9-18607.18|generated/sv2v_out.v:18607.5-18621.8" */ _018_ : 1'hx;
assign _000_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18607.9-18607.18|generated/sv2v_out.v:18607.5-18621.8" */ _016_ : 1'h0;
assign _008_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18607.9-18607.18|generated/sv2v_out.v:18607.5-18621.8" */ lsu_we_i : 1'h0;
assign _006_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18607.9-18607.18|generated/sv2v_out.v:18607.5-18621.8" */ _287_ : 1'h0;
assign _005_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18607.9-18607.18|generated/sv2v_out.v:18607.5-18621.8" */ 1'h0 : 1'hx;
assign _009_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18607.9-18607.18|generated/sv2v_out.v:18607.5-18621.8" */ data_pmp_err_i : 1'h0;
assign _002_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18607.9-18607.18|generated/sv2v_out.v:18607.5-18621.8" */ 1'h1 : 1'h0;
assign perf_store_o = _281_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18604.3-18669.10" */ _008_ : 1'h0;
assign perf_load_o = _281_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18604.3-18669.10" */ _006_ : 1'h0;
assign _303_ = ls_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18604.3-18669.10" */ 3'h1;
assign _281_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18604.3-18669.10" */ ls_fsm_cs;
assign _300_ = ls_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18604.3-18669.10" */ 3'h4;
assign _301_ = ls_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18604.3-18669.10" */ 3'h3;
assign _302_ = ls_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18604.3-18669.10" */ 3'h2;
assign _305_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18567.3-18572.10" */ _304_;
assign _304_[0] = data_type_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18567.3-18572.10" */ 2'h2;
assign _304_[1] = data_type_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18567.3-18572.10" */ 2'h3;
assign _306_ = data_type_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18567.3-18572.10" */ 2'h1;
assign _046_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18560.9-18560.25|generated/sv2v_out.v:18560.5-18563.67" */ { data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31:24] } : { 24'h000000, data_rdata_i[31:24] };
assign _037_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18555.9-18555.25|generated/sv2v_out.v:18555.5-18558.67" */ { data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23:16] } : { 24'h000000, data_rdata_i[23:16] };
assign _024_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18550.9-18550.25|generated/sv2v_out.v:18550.5-18553.66" */ { data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15:8] } : { 24'h000000, data_rdata_i[15:8] };
assign _011_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18545.9-18545.25|generated/sv2v_out.v:18545.5-18548.64" */ { data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7:0] } : { 24'h000000, data_rdata_i[7:0] };
assign _048_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18536.9-18536.25|generated/sv2v_out.v:18536.5-18539.80" */ { data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7:0], rdata_q[31:24] } : { 16'h0000, data_rdata_i[7:0], rdata_q[31:24] };
assign _039_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18531.9-18531.25|generated/sv2v_out.v:18531.5-18534.67" */ { data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31:16] } : { 16'h0000, data_rdata_i[31:16] };
assign _026_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18526.9-18526.25|generated/sv2v_out.v:18526.5-18529.66" */ { data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23:8] } : { 16'h0000, data_rdata_i[23:8] };
assign _013_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18521.9-18521.25|generated/sv2v_out.v:18521.5-18524.66" */ { data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15:0] } : { 16'h0000, data_rdata_i[15:0] };
assign _307_ = rdata_offset_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18511.3-18517.10" */ 2'h3;
assign _308_ = rdata_offset_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18511.3-18517.10" */ 2'h2;
assign _309_ = rdata_offset_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18511.3-18517.10" */ 2'h1;
assign _313_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18439.3-18477.10" */ _312_;
assign _042_ = handle_misaligned_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18458.9-18458.29|generated/sv2v_out.v:18458.5-18467.24" */ 4'h1 : _051_;
assign _279_ = adder_result_ex_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18442.6-18448.13" */ 2'h3;
assign _310_ = adder_result_ex_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18442.6-18448.13" */ 2'h2;
assign _311_ = adder_result_ex_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18442.6-18448.13" */ 2'h1;
assign _001_ = handle_misaligned_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18441.9-18441.29|generated/sv2v_out.v:18441.5-18456.13" */ _030_ : _017_;
assign _312_[0] = lsu_type_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18439.3-18477.10" */ 2'h2;
assign _312_[1] = lsu_type_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18439.3-18477.10" */ 2'h3;
assign _278_ = lsu_type_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18439.3-18477.10" */ 2'h1;
assign _277_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18439.3-18477.10" */ lsu_type_i;
assign data_intg_err = | /* src = "generated/sv2v_out.v:18585.27-18585.35" */ \g_mem_rdata_ecc.ecc_err ;
assign addr_last_d = addr_incr_req_o ? /* src = "generated/sv2v_out.v:18504.24-18504.73" */ { adder_result_ex_i[31:2], 2'h0 } : adder_result_ex_i;
assign _314_ = split_misaligned_access ? /* src = "generated/sv2v_out.v:18617.20-18617.57" */ 3'h2 : 3'h0;
assign _315_ = split_misaligned_access ? /* src = "generated/sv2v_out.v:18620.20-18620.57" */ 3'h1 : 3'h3;
assign _316_ = data_gnt_i ? /* src = "generated/sv2v_out.v:18639.19-18639.43" */ 3'h0 : 3'h3;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18581.30-18584.5" */
prim_secded_inv_39_32_dec \g_mem_rdata_ecc.u_data_intg_dec  (
.data_i(\g_mem_rdata_ecc.data_rdata_buf ),
.data_i_t0(\g_mem_rdata_ecc.data_rdata_buf_t0 ),
.err_o(\g_mem_rdata_ecc.ecc_err ),
.err_o_t0(\g_mem_rdata_ecc.ecc_err_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18577.37-18580.5" */
\$paramod\prim_buf\Width=32'00000000000000000000000000100111  \g_mem_rdata_ecc.u_prim_buf_instr_rdata  (
.in_i(data_rdata_i),
.in_i_t0(data_rdata_i_t0),
.out_o(\g_mem_rdata_ecc.data_rdata_buf ),
.out_o_t0(\g_mem_rdata_ecc.data_rdata_buf_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18695.30-18698.5" */
prim_secded_inv_39_32_enc \g_mem_wdata_ecc.u_data_gen  (
.data_i(data_wdata),
.data_i_t0(data_wdata_t0),
.data_o(data_wdata_o),
.data_o_t0(data_wdata_o_t0)
);
assign busy_o_t0 = 1'h0;
assign data_addr_o = { adder_result_ex_i[31:2], 2'h0 };
assign data_addr_o_t0 = { adder_result_ex_i_t0[31:2], 2'h0 };
assign data_be_o_t0 = 4'h0;
assign data_req_o_t0 = 1'h0;
assign data_we_o = lsu_we_i;
assign data_we_o_t0 = lsu_we_i_t0;
assign perf_store_o_t0 = perf_load_o_t0;
endmodule

module \$paramod\ibex_prefetch_buffer\ResetAll=1'1 (clk_i, rst_ni, req_i, branch_i, addr_i, ready_i, valid_o, rdata_o, addr_o, err_o, err_plus2_o, instr_req_o, instr_gnt_i, instr_addr_o, instr_rdata_i, instr_err_i, instr_rvalid_i, busy_o, valid_o_t0, req_i_t0, ready_i_t0
, rdata_o_t0, instr_rvalid_i_t0, instr_req_o_t0, instr_rdata_i_t0, instr_gnt_i_t0, instr_err_i_t0, instr_addr_o_t0, err_plus2_o_t0, branch_i_t0, addr_o_t0, addr_i_t0, busy_o_t0, err_o_t0);
/* src = "generated/sv2v_out.v:19990.26-19990.57" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19990.26-19990.57" */
wire _001_;
/* src = "generated/sv2v_out.v:19994.27-19994.55" */
wire _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19994.27-19994.55" */
wire _003_;
/* src = "generated/sv2v_out.v:20031.38-20031.61" */
wire _004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20031.38-20031.61" */
wire _005_;
/* src = "generated/sv2v_out.v:20032.36-20032.77" */
wire _006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20032.36-20032.77" */
wire _007_;
/* src = "generated/sv2v_out.v:20032.82-20032.115" */
wire _008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20032.82-20032.115" */
wire _009_;
/* src = "generated/sv2v_out.v:20035.38-20035.92" */
wire _010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20035.38-20035.92" */
wire _011_;
/* src = "generated/sv2v_out.v:20036.36-20036.108" */
wire _012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20036.36-20036.108" */
wire _013_;
/* src = "generated/sv2v_out.v:20036.113-20036.146" */
wire _014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20036.113-20036.146" */
wire _015_;
wire [31:0] _016_;
wire [31:0] _017_;
wire _018_;
wire _019_;
wire _020_;
wire [31:0] _021_;
wire [31:0] _022_;
wire [1:0] _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire [31:0] _043_;
wire [31:0] _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire [31:0] _079_;
wire [31:0] _080_;
wire [1:0] _081_;
wire [1:0] _082_;
wire [29:0] _083_;
wire [29:0] _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire [31:0] _106_;
wire [31:0] _107_;
wire [31:0] _108_;
wire [31:0] _109_;
wire [31:0] _110_;
wire [1:0] _111_;
wire [1:0] _112_;
wire [1:0] _113_;
wire [1:0] _114_;
wire [31:0] _115_;
wire [31:0] _116_;
wire [31:0] _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire [31:0] _130_;
wire [1:0] _131_;
wire [29:0] _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire [31:0] _141_;
wire [31:0] _142_;
wire [31:0] _143_;
/* src = "generated/sv2v_out.v:19992.35-19992.47" */
wire _144_;
/* src = "generated/sv2v_out.v:19970.25-19970.58" */
wire [1:0] _145_;
/* src = "generated/sv2v_out.v:19990.35-19990.56" */
wire _146_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19990.35-19990.56" */
wire _147_;
/* src = "generated/sv2v_out.v:19993.40-19993.64" */
wire _148_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19993.40-19993.64" */
wire _149_;
/* src = "generated/sv2v_out.v:20032.35-20032.116" */
wire _150_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20032.35-20032.116" */
wire _151_;
/* src = "generated/sv2v_out.v:20036.35-20036.147" */
wire _152_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20036.35-20036.147" */
wire _153_;
/* src = "generated/sv2v_out.v:19962.18-19962.38" */
wire _154_;
/* src = "generated/sv2v_out.v:20011.25-20011.72" */
wire [31:0] _155_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20011.25-20011.72" */
wire [31:0] _156_;
/* src = "generated/sv2v_out.v:20026.54-20026.86" */
wire [31:0] _157_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20026.54-20026.86" */
wire [31:0] _158_;
/* src = "generated/sv2v_out.v:19921.20-19921.26" */
input [31:0] addr_i;
wire [31:0] addr_i;
/* cellift = 32'd1 */
input [31:0] addr_i_t0;
wire [31:0] addr_i_t0;
/* src = "generated/sv2v_out.v:19925.21-19925.27" */
output [31:0] addr_o;
wire [31:0] addr_o;
/* cellift = 32'd1 */
output [31:0] addr_o_t0;
wire [31:0] addr_o_t0;
/* src = "generated/sv2v_out.v:19945.13-19945.29" */
wire [1:0] branch_discard_n;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19945.13-19945.29" */
wire [1:0] branch_discard_n_t0;
/* src = "generated/sv2v_out.v:19947.12-19947.28" */
reg [1:0] branch_discard_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19947.12-19947.28" */
reg [1:0] branch_discard_q_t0;
/* src = "generated/sv2v_out.v:19946.13-19946.29" */
wire [1:0] branch_discard_s;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19946.13-19946.29" */
wire [1:0] branch_discard_s_t0;
/* src = "generated/sv2v_out.v:19920.13-19920.21" */
input branch_i;
wire branch_i;
/* cellift = 32'd1 */
input branch_i_t0;
wire branch_i_t0;
/* src = "generated/sv2v_out.v:19934.14-19934.20" */
output busy_o;
wire busy_o;
/* cellift = 32'd1 */
output busy_o_t0;
wire busy_o_t0;
/* src = "generated/sv2v_out.v:19917.13-19917.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:19940.7-19940.20" */
wire discard_req_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19940.7-19940.20" */
wire discard_req_d_t0;
/* src = "generated/sv2v_out.v:19941.6-19941.19" */
reg discard_req_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19941.6-19941.19" */
reg discard_req_q_t0;
/* src = "generated/sv2v_out.v:19926.14-19926.19" */
output err_o;
wire err_o;
/* cellift = 32'd1 */
output err_o_t0;
wire err_o_t0;
/* src = "generated/sv2v_out.v:19927.14-19927.25" */
output err_plus2_o;
wire err_plus2_o;
/* cellift = 32'd1 */
output err_plus2_o_t0;
wire err_plus2_o_t0;
/* src = "generated/sv2v_out.v:19952.14-19952.26" */
wire [31:0] fetch_addr_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19952.14-19952.26" */
wire [31:0] fetch_addr_d_t0;
/* src = "generated/sv2v_out.v:19954.7-19954.20" */
wire fetch_addr_en;
/* src = "generated/sv2v_out.v:19953.13-19953.25" */
reg [31:0] fetch_addr_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19953.13-19953.25" */
reg [31:0] fetch_addr_q_t0;
/* src = "generated/sv2v_out.v:19961.13-19961.22" */
wire [1:0] fifo_busy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19961.13-19961.22" */
/* unused_bits = "0 1" */
wire [1:0] fifo_busy_t0;
/* src = "generated/sv2v_out.v:19959.7-19959.17" */
wire fifo_ready;
/* src = "generated/sv2v_out.v:19957.7-19957.17" */
wire fifo_valid;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19957.7-19957.17" */
wire fifo_valid_t0;
/* src = "generated/sv2v_out.v:19955.14-19955.24" */
/* unused_bits = "0 1" */
wire [31:0] instr_addr;
/* src = "generated/sv2v_out.v:19930.21-19930.33" */
output [31:0] instr_addr_o;
wire [31:0] instr_addr_o;
/* cellift = 32'd1 */
output [31:0] instr_addr_o_t0;
wire [31:0] instr_addr_o_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19955.14-19955.24" */
/* unused_bits = "0 1" */
wire [31:0] instr_addr_t0;
/* src = "generated/sv2v_out.v:19932.13-19932.24" */
input instr_err_i;
wire instr_err_i;
/* cellift = 32'd1 */
input instr_err_i_t0;
wire instr_err_i_t0;
/* src = "generated/sv2v_out.v:19929.13-19929.24" */
input instr_gnt_i;
wire instr_gnt_i;
/* cellift = 32'd1 */
input instr_gnt_i_t0;
wire instr_gnt_i_t0;
/* src = "generated/sv2v_out.v:19931.20-19931.33" */
input [31:0] instr_rdata_i;
wire [31:0] instr_rdata_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_i_t0;
wire [31:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:19928.14-19928.25" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:19933.13-19933.27" */
input instr_rvalid_i;
wire instr_rvalid_i;
/* cellift = 32'd1 */
input instr_rvalid_i_t0;
wire instr_rvalid_i_t0;
/* src = "generated/sv2v_out.v:19924.21-19924.28" */
output [31:0] rdata_o;
wire [31:0] rdata_o;
/* cellift = 32'd1 */
output [31:0] rdata_o_t0;
wire [31:0] rdata_o_t0;
/* src = "generated/sv2v_out.v:19942.13-19942.32" */
wire [1:0] rdata_outstanding_n;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19942.13-19942.32" */
wire [1:0] rdata_outstanding_n_t0;
/* src = "generated/sv2v_out.v:19944.12-19944.31" */
reg [1:0] rdata_outstanding_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19944.12-19944.31" */
reg [1:0] rdata_outstanding_q_t0;
/* src = "generated/sv2v_out.v:19943.13-19943.32" */
wire [1:0] rdata_outstanding_s;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19943.13-19943.32" */
wire [1:0] rdata_outstanding_s_t0;
/* src = "generated/sv2v_out.v:19922.13-19922.20" */
input ready_i;
wire ready_i;
/* cellift = 32'd1 */
input ready_i_t0;
wire ready_i_t0;
/* src = "generated/sv2v_out.v:19919.13-19919.18" */
input req_i;
wire req_i;
/* cellift = 32'd1 */
input req_i_t0;
wire req_i_t0;
/* src = "generated/sv2v_out.v:19918.13-19918.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:19951.7-19951.21" */
wire stored_addr_en;
/* src = "generated/sv2v_out.v:19950.13-19950.26" */
reg [31:0] stored_addr_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19950.13-19950.26" */
reg [31:0] stored_addr_q_t0;
/* src = "generated/sv2v_out.v:19936.7-19936.20" */
wire valid_new_req;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19936.7-19936.20" */
wire valid_new_req_t0;
/* src = "generated/sv2v_out.v:19923.14-19923.21" */
output valid_o;
wire valid_o;
/* cellift = 32'd1 */
output valid_o_t0;
wire valid_o_t0;
/* src = "generated/sv2v_out.v:19938.7-19938.18" */
wire valid_req_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19938.7-19938.18" */
wire valid_req_d_t0;
/* src = "generated/sv2v_out.v:19939.6-19939.17" */
reg valid_req_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19939.6-19939.17" */
reg valid_req_q_t0;
assign fetch_addr_d = _155_ + /* src = "generated/sv2v_out.v:20011.24-20011.126" */ { 29'h00000000, _002_, 2'h0 };
assign _000_ = req_i & /* src = "generated/sv2v_out.v:19990.26-19990.57" */ _146_;
assign valid_new_req = _000_ & /* src = "generated/sv2v_out.v:19990.25-19990.84" */ _039_;
assign valid_req_d = instr_req_o & /* src = "generated/sv2v_out.v:19992.23-19992.47" */ _144_;
assign discard_req_d = valid_req_q & /* src = "generated/sv2v_out.v:19993.25-19993.65" */ _148_;
assign stored_addr_en = _002_ & /* src = "generated/sv2v_out.v:19994.26-19994.71" */ _144_;
assign _002_ = valid_new_req & /* src = "generated/sv2v_out.v:20011.90-20011.118" */ _024_;
assign _008_ = branch_i & /* src = "generated/sv2v_out.v:20032.82-20032.115" */ rdata_outstanding_q[0];
assign _010_ = _004_ & /* src = "generated/sv2v_out.v:20035.38-20035.92" */ rdata_outstanding_q[0];
assign _004_ = instr_req_o & /* src = "generated/sv2v_out.v:20036.38-20036.61" */ instr_gnt_i;
assign _006_ = _004_ & /* src = "generated/sv2v_out.v:20036.37-20036.78" */ discard_req_d;
assign _012_ = _006_ & /* src = "generated/sv2v_out.v:20036.36-20036.108" */ rdata_outstanding_q[0];
assign _014_ = branch_i & /* src = "generated/sv2v_out.v:20036.113-20036.146" */ rdata_outstanding_q[1];
assign fifo_valid = instr_rvalid_i & /* src = "generated/sv2v_out.v:20042.22-20042.59" */ _038_;
assign _016_ = ~ _156_;
assign _017_ = ~ { 29'h00000000, _003_, 2'h0 };
assign _043_ = _155_ & _016_;
assign _044_ = { 29'h00000000, _002_, 2'h0 } & _017_;
assign _142_ = _043_ + _044_;
assign _115_ = _155_ | _156_;
assign _116_ = { 29'h00000000, _002_, 2'h0 } | { 29'h00000000, _003_, 2'h0 };
assign _143_ = _115_ + _116_;
assign _141_ = _142_ ^ _143_;
assign _117_ = _141_ | _156_;
assign fetch_addr_d_t0 = _117_ | { 29'h00000000, _003_, 2'h0 };
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME valid_req_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) valid_req_q_t0 <= 1'h0;
else valid_req_q_t0 <= valid_req_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME discard_req_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) discard_req_q_t0 <= 1'h0;
else discard_req_q_t0 <= discard_req_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_outstanding_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_outstanding_q_t0 <= 2'h0;
else rdata_outstanding_q_t0 <= rdata_outstanding_s_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME branch_discard_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_discard_q_t0 <= 2'h0;
else branch_discard_q_t0 <= branch_discard_s_t0;
assign _018_ = ~ fetch_addr_en;
assign _019_ = ~ _042_;
assign _020_ = ~ stored_addr_en;
assign _079_ = { fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en } & fetch_addr_d_t0;
assign _081_ = { _042_, _042_ } & _158_[1:0];
assign _083_ = { stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en } & instr_addr_t0[31:2];
assign _080_ = { _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_ } & fetch_addr_q_t0;
assign _082_ = { _019_, _019_ } & stored_addr_q_t0[1:0];
assign _084_ = { _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_ } & stored_addr_q_t0[31:2];
assign _130_ = _079_ | _080_;
assign _131_ = _081_ | _082_;
assign _132_ = _083_ | _084_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME fetch_addr_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) fetch_addr_q_t0 <= 32'd0;
else fetch_addr_q_t0 <= _130_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME stored_addr_q_t0[1:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) stored_addr_q_t0[1:0] <= 2'h0;
else stored_addr_q_t0[1:0] <= _131_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME stored_addr_q_t0[31:2] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) stored_addr_q_t0[31:2] <= 30'h00000000;
else stored_addr_q_t0[31:2] <= _132_;
assign _045_ = req_i_t0 & _146_;
assign _048_ = _001_ & _039_;
assign _051_ = instr_req_o_t0 & _144_;
assign _054_ = valid_req_q_t0 & _148_;
assign _057_ = valid_new_req_t0 & _024_;
assign _060_ = branch_i_t0 & rdata_outstanding_q[0];
assign _063_ = _005_ & rdata_outstanding_q[0];
assign _066_ = instr_req_o_t0 & instr_gnt_i;
assign _067_ = _005_ & discard_req_d;
assign _070_ = _007_ & rdata_outstanding_q[0];
assign _073_ = branch_i_t0 & rdata_outstanding_q[1];
assign _076_ = instr_rvalid_i_t0 & _038_;
assign _046_ = _147_ & req_i;
assign _049_ = rdata_outstanding_q_t0[1] & _000_;
assign _052_ = instr_gnt_i_t0 & instr_req_o;
assign _055_ = _149_ & valid_req_q;
assign _058_ = valid_req_q_t0 & valid_new_req;
assign _061_ = rdata_outstanding_q_t0[0] & branch_i;
assign _064_ = rdata_outstanding_q_t0[0] & _004_;
assign _068_ = discard_req_d_t0 & _004_;
assign _071_ = rdata_outstanding_q_t0[0] & _006_;
assign _074_ = rdata_outstanding_q_t0[1] & branch_i;
assign _077_ = branch_discard_q_t0[0] & instr_rvalid_i;
assign _047_ = req_i_t0 & _147_;
assign _050_ = _001_ & rdata_outstanding_q_t0[1];
assign _053_ = instr_req_o_t0 & instr_gnt_i_t0;
assign _056_ = valid_req_q_t0 & _149_;
assign _059_ = valid_new_req_t0 & valid_req_q_t0;
assign _062_ = branch_i_t0 & rdata_outstanding_q_t0[0];
assign _065_ = _005_ & rdata_outstanding_q_t0[0];
assign _069_ = _005_ & discard_req_d_t0;
assign _072_ = _007_ & rdata_outstanding_q_t0[0];
assign _075_ = branch_i_t0 & rdata_outstanding_q_t0[1];
assign _078_ = instr_rvalid_i_t0 & branch_discard_q_t0[0];
assign _118_ = _045_ | _046_;
assign _119_ = _048_ | _049_;
assign _120_ = _051_ | _052_;
assign _121_ = _054_ | _055_;
assign _122_ = _057_ | _058_;
assign _123_ = _060_ | _061_;
assign _124_ = _063_ | _064_;
assign _125_ = _066_ | _052_;
assign _126_ = _067_ | _068_;
assign _127_ = _070_ | _071_;
assign _128_ = _073_ | _074_;
assign _129_ = _076_ | _077_;
assign _001_ = _118_ | _047_;
assign valid_new_req_t0 = _119_ | _050_;
assign valid_req_d_t0 = _120_ | _053_;
assign discard_req_d_t0 = _121_ | _056_;
assign _003_ = _122_ | _059_;
assign _009_ = _123_ | _062_;
assign _011_ = _124_ | _065_;
assign _005_ = _125_ | _053_;
assign _007_ = _126_ | _069_;
assign _013_ = _127_ | _072_;
assign _015_ = _128_ | _075_;
assign fifo_valid_t0 = _129_ | _078_;
/* src = "generated/sv2v_out.v:20014.4-20018.35" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME fetch_addr_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) fetch_addr_q <= 32'd0;
else if (fetch_addr_en) fetch_addr_q <= fetch_addr_d;
/* src = "generated/sv2v_out.v:19998.4-20002.37" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME stored_addr_q[1:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) stored_addr_q[1:0] <= 2'h0;
else if (_042_) stored_addr_q[1:0] <= _157_[1:0];
/* src = "generated/sv2v_out.v:19998.4-20002.37" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME stored_addr_q[31:2] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) stored_addr_q[31:2] <= 30'h00000000;
else if (stored_addr_en) stored_addr_q[31:2] <= instr_addr[31:2];
assign _021_ = ~ { branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i };
assign _022_ = ~ { valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q };
assign _023_ = ~ { instr_rvalid_i, instr_rvalid_i };
assign _106_ = _021_ & { fetch_addr_q_t0[31:2], 2'h0 };
assign _108_ = _021_ & fetch_addr_q_t0;
assign _109_ = _022_ & _158_;
assign _111_ = _023_ & rdata_outstanding_n_t0;
assign _113_ = _023_ & branch_discard_n_t0;
assign _107_ = { branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i } & addr_i_t0;
assign _110_ = { valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q } & stored_addr_q_t0;
assign _112_ = { instr_rvalid_i, instr_rvalid_i } & { 1'h0, rdata_outstanding_n_t0[1] };
assign _114_ = { instr_rvalid_i, instr_rvalid_i } & { 1'h0, branch_discard_n_t0[1] };
assign _156_ = _106_ | _107_;
assign _158_ = _108_ | _107_;
assign instr_addr_t0 = _109_ | _110_;
assign rdata_outstanding_s_t0 = _111_ | _112_;
assign branch_discard_s_t0 = _113_ | _114_;
assign _024_ = ~ valid_req_q;
assign _042_ = & { _024_, stored_addr_en };
assign _025_ = ~ _154_;
assign _027_ = ~ branch_i;
assign _028_ = ~ _004_;
assign _029_ = ~ _006_;
assign _030_ = ~ _150_;
assign _031_ = ~ _010_;
assign _032_ = ~ _012_;
assign _033_ = ~ _152_;
assign _034_ = ~ valid_new_req;
assign _035_ = ~ discard_req_q;
assign _036_ = ~ rdata_outstanding_q[0];
assign _037_ = ~ _008_;
assign _038_ = ~ branch_discard_q[0];
assign _039_ = ~ rdata_outstanding_q[1];
assign _040_ = ~ _014_;
assign _041_ = ~ branch_discard_q[1];
assign _085_ = valid_req_q_t0 & _034_;
assign _086_ = branch_i_t0 & _035_;
assign _089_ = _005_ & _036_;
assign _091_ = _007_ & _037_;
assign _094_ = _151_ & _038_;
assign _097_ = _011_ & _039_;
assign _100_ = _013_ & _040_;
assign _103_ = _153_ & _041_;
assign busy_o_t0 = instr_req_o_t0 & _025_;
assign _147_ = branch_i_t0 & _026_;
assign _087_ = discard_req_q_t0 & _027_;
assign _090_ = rdata_outstanding_q_t0[0] & _028_;
assign _092_ = _009_ & _029_;
assign _095_ = branch_discard_q_t0[0] & _030_;
assign _098_ = rdata_outstanding_q_t0[1] & _031_;
assign _101_ = _015_ & _032_;
assign _104_ = branch_discard_q_t0[1] & _033_;
assign _088_ = branch_i_t0 & discard_req_q_t0;
assign _093_ = _007_ & _009_;
assign _096_ = _151_ & branch_discard_q_t0[0];
assign _099_ = _011_ & rdata_outstanding_q_t0[1];
assign _102_ = _013_ & _015_;
assign _105_ = _153_ & branch_discard_q_t0[1];
assign _133_ = _085_ | _057_;
assign _134_ = _086_ | _087_;
assign _135_ = _089_ | _090_;
assign _136_ = _091_ | _092_;
assign _137_ = _094_ | _095_;
assign _138_ = _097_ | _098_;
assign _139_ = _100_ | _101_;
assign _140_ = _103_ | _104_;
assign instr_req_o_t0 = _133_ | _059_;
assign _149_ = _134_ | _088_;
assign rdata_outstanding_n_t0[0] = _135_ | _065_;
assign _151_ = _136_ | _093_;
assign branch_discard_n_t0[0] = _137_ | _096_;
assign rdata_outstanding_n_t0[1] = _138_ | _099_;
assign _153_ = _139_ | _102_;
assign branch_discard_n_t0[1] = _140_ | _105_;
assign fifo_ready = ! /* src = "generated/sv2v_out.v:0.0-0.0" */ _026_;
assign _144_ = ~ /* src = "generated/sv2v_out.v:19994.59-19994.71" */ instr_gnt_i;
assign busy_o = _154_ | /* src = "generated/sv2v_out.v:19962.18-19962.52" */ instr_req_o;
assign _145_ = fifo_busy | /* src = "generated/sv2v_out.v:19970.25-19970.58" */ { rdata_outstanding_q[0], rdata_outstanding_q[1] };
assign _146_ = fifo_ready | /* src = "generated/sv2v_out.v:19990.35-19990.56" */ branch_i;
assign instr_req_o = valid_req_q | /* src = "generated/sv2v_out.v:19991.21-19991.48" */ valid_new_req;
assign _148_ = branch_i | /* src = "generated/sv2v_out.v:19993.40-19993.64" */ discard_req_q;
assign fetch_addr_en = branch_i | /* src = "generated/sv2v_out.v:20010.25-20010.66" */ _002_;
assign rdata_outstanding_n[0] = _004_ | /* src = "generated/sv2v_out.v:20031.37-20031.87" */ rdata_outstanding_q[0];
assign _150_ = _006_ | /* src = "generated/sv2v_out.v:20032.35-20032.116" */ _008_;
assign branch_discard_n[0] = _150_ | /* src = "generated/sv2v_out.v:20032.34-20032.139" */ branch_discard_q[0];
assign rdata_outstanding_n[1] = _010_ | /* src = "generated/sv2v_out.v:20035.37-20035.118" */ rdata_outstanding_q[1];
assign _152_ = _012_ | /* src = "generated/sv2v_out.v:20036.35-20036.147" */ _014_;
assign branch_discard_n[1] = _152_ | /* src = "generated/sv2v_out.v:20036.34-20036.170" */ branch_discard_q[1];
/* src = "generated/sv2v_out.v:20044.2-20056.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME valid_req_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) valid_req_q <= 1'h0;
else valid_req_q <= valid_req_d;
/* src = "generated/sv2v_out.v:20044.2-20056.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME discard_req_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) discard_req_q <= 1'h0;
else discard_req_q <= discard_req_d;
/* src = "generated/sv2v_out.v:20044.2-20056.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_outstanding_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_outstanding_q <= 2'h0;
else rdata_outstanding_q <= rdata_outstanding_s;
/* src = "generated/sv2v_out.v:20044.2-20056.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME branch_discard_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_discard_q <= 2'h0;
else branch_discard_q <= branch_discard_s;
assign _026_ = & /* src = "generated/sv2v_out.v:19970.22-19970.59" */ _145_;
assign _154_ = | /* src = "generated/sv2v_out.v:19962.18-19962.38" */ rdata_outstanding_q;
assign _155_ = branch_i ? /* src = "generated/sv2v_out.v:20011.25-20011.72" */ addr_i : { fetch_addr_q[31:2], 2'h0 };
assign _157_ = branch_i ? /* src = "generated/sv2v_out.v:20026.54-20026.86" */ addr_i : fetch_addr_q;
assign instr_addr = valid_req_q ? /* src = "generated/sv2v_out.v:20026.23-20026.87" */ stored_addr_q : _157_;
assign rdata_outstanding_s = instr_rvalid_i ? /* src = "generated/sv2v_out.v:20040.32-20040.103" */ { 1'h0, rdata_outstanding_n[1] } : rdata_outstanding_n;
assign branch_discard_s = instr_rvalid_i ? /* src = "generated/sv2v_out.v:20041.29-20041.94" */ { 1'h0, branch_discard_n[1] } : branch_discard_n;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:19974.4-19989.3" */
\$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  fifo_i (
.busy_o(fifo_busy),
.busy_o_t0(fifo_busy_t0),
.clear_i(branch_i),
.clear_i_t0(branch_i_t0),
.clk_i(clk_i),
.in_addr_i(addr_i),
.in_addr_i_t0(addr_i_t0),
.in_err_i(instr_err_i),
.in_err_i_t0(instr_err_i_t0),
.in_rdata_i(instr_rdata_i),
.in_rdata_i_t0(instr_rdata_i_t0),
.in_valid_i(fifo_valid),
.in_valid_i_t0(fifo_valid_t0),
.out_addr_o(addr_o),
.out_addr_o_t0(addr_o_t0),
.out_err_o(err_o),
.out_err_o_t0(err_o_t0),
.out_err_plus2_o(err_plus2_o),
.out_err_plus2_o_t0(err_plus2_o_t0),
.out_rdata_o(rdata_o),
.out_rdata_o_t0(rdata_o_t0),
.out_ready_i(ready_i),
.out_ready_i_t0(ready_i_t0),
.out_valid_o(valid_o),
.out_valid_o_t0(valid_o_t0),
.rst_ni(rst_ni)
);
assign instr_addr_o = { instr_addr[31:2], 2'h0 };
assign instr_addr_o_t0 = { instr_addr_t0[31:2], 2'h0 };
endmodule

module \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'0\DummyInstructions=1'1 (clk_i, rst_ni, en_wb_i, instr_type_wb_i, pc_id_i, instr_is_compressed_id_i, instr_perf_count_id_i, ready_wb_o, rf_write_wb_o, outstanding_load_wb_o, outstanding_store_wb_o, pc_wb_o, perf_instr_ret_wb_o, perf_instr_ret_compressed_wb_o, perf_instr_ret_wb_spec_o, perf_instr_ret_compressed_wb_spec_o, rf_waddr_id_i, rf_wdata_id_i, rf_we_id_i, dummy_instr_id_i, rf_wdata_lsu_i
, rf_we_lsu_i, rf_wdata_fwd_wb_o, rf_waddr_wb_o, rf_wdata_wb_o, rf_we_wb_o, dummy_instr_wb_o, lsu_resp_valid_i, lsu_resp_err_i, instr_done_wb_o, pc_id_i_t0, lsu_resp_valid_i_t0, dummy_instr_id_i_t0, dummy_instr_wb_o_t0, en_wb_i_t0, instr_done_wb_o_t0, instr_is_compressed_id_i_t0, instr_perf_count_id_i_t0, instr_type_wb_i_t0, lsu_resp_err_i_t0, outstanding_load_wb_o_t0, outstanding_store_wb_o_t0
, pc_wb_o_t0, perf_instr_ret_compressed_wb_o_t0, perf_instr_ret_compressed_wb_spec_o_t0, perf_instr_ret_wb_o_t0, perf_instr_ret_wb_spec_o_t0, ready_wb_o_t0, rf_waddr_id_i_t0, rf_waddr_wb_o_t0, rf_wdata_fwd_wb_o_t0, rf_wdata_id_i_t0, rf_wdata_lsu_i_t0, rf_wdata_wb_o_t0, rf_we_id_i_t0, rf_we_lsu_i_t0, rf_we_wb_o_t0, rf_write_wb_o_t0);
/* src = "generated/sv2v_out.v:21076.34-21076.65" */
wire _00_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21076.34-21076.65" */
wire _01_;
/* src = "generated/sv2v_out.v:21076.71-21076.104" */
wire _02_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21076.71-21076.104" */
wire _03_;
/* src = "generated/sv2v_out.v:21098.26-21098.75" */
wire [31:0] _04_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21098.26-21098.75" */
wire [31:0] _05_;
/* src = "generated/sv2v_out.v:21098.80-21098.129" */
wire [31:0] _06_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21098.80-21098.129" */
wire [31:0] _07_;
wire [31:0] _08_;
wire [31:0] _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire [31:0] _22_;
wire [31:0] _23_;
wire [31:0] _24_;
wire [31:0] _25_;
wire [31:0] _26_;
wire [31:0] _27_;
wire [31:0] _28_;
wire [31:0] _29_;
wire [31:0] _30_;
wire _31_;
wire _32_;
wire _33_;
wire _34_;
wire [31:0] _35_;
wire [31:0] _36_;
wire [31:0] _37_;
/* src = "generated/sv2v_out.v:21076.69-21076.105" */
wire _38_;
/* src = "generated/sv2v_out.v:20947.13-20947.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:20966.13-20966.29" */
input dummy_instr_id_i;
wire dummy_instr_id_i;
/* cellift = 32'd1 */
input dummy_instr_id_i_t0;
wire dummy_instr_id_i_t0;
/* src = "generated/sv2v_out.v:20973.14-20973.30" */
output dummy_instr_wb_o;
wire dummy_instr_wb_o;
/* cellift = 32'd1 */
output dummy_instr_wb_o_t0;
wire dummy_instr_wb_o_t0;
/* src = "generated/sv2v_out.v:20949.13-20949.20" */
input en_wb_i;
wire en_wb_i;
/* cellift = 32'd1 */
input en_wb_i_t0;
wire en_wb_i_t0;
/* src = "generated/sv2v_out.v:20976.14-20976.29" */
output instr_done_wb_o;
wire instr_done_wb_o;
/* cellift = 32'd1 */
output instr_done_wb_o_t0;
wire instr_done_wb_o_t0;
/* src = "generated/sv2v_out.v:20952.13-20952.37" */
input instr_is_compressed_id_i;
wire instr_is_compressed_id_i;
/* cellift = 32'd1 */
input instr_is_compressed_id_i_t0;
wire instr_is_compressed_id_i_t0;
/* src = "generated/sv2v_out.v:20953.13-20953.34" */
input instr_perf_count_id_i;
wire instr_perf_count_id_i;
/* cellift = 32'd1 */
input instr_perf_count_id_i_t0;
wire instr_perf_count_id_i_t0;
/* src = "generated/sv2v_out.v:20950.19-20950.34" */
input [1:0] instr_type_wb_i;
wire [1:0] instr_type_wb_i;
/* cellift = 32'd1 */
input [1:0] instr_type_wb_i_t0;
wire [1:0] instr_type_wb_i_t0;
/* src = "generated/sv2v_out.v:20975.13-20975.27" */
input lsu_resp_err_i;
wire lsu_resp_err_i;
/* cellift = 32'd1 */
input lsu_resp_err_i_t0;
wire lsu_resp_err_i_t0;
/* src = "generated/sv2v_out.v:20974.13-20974.29" */
input lsu_resp_valid_i;
wire lsu_resp_valid_i;
/* cellift = 32'd1 */
input lsu_resp_valid_i_t0;
wire lsu_resp_valid_i_t0;
/* src = "generated/sv2v_out.v:20956.14-20956.35" */
output outstanding_load_wb_o;
wire outstanding_load_wb_o;
/* cellift = 32'd1 */
output outstanding_load_wb_o_t0;
wire outstanding_load_wb_o_t0;
/* src = "generated/sv2v_out.v:20957.14-20957.36" */
output outstanding_store_wb_o;
wire outstanding_store_wb_o;
/* cellift = 32'd1 */
output outstanding_store_wb_o_t0;
wire outstanding_store_wb_o_t0;
/* src = "generated/sv2v_out.v:20951.20-20951.27" */
input [31:0] pc_id_i;
wire [31:0] pc_id_i;
/* cellift = 32'd1 */
input [31:0] pc_id_i_t0;
wire [31:0] pc_id_i_t0;
/* src = "generated/sv2v_out.v:20958.21-20958.28" */
output [31:0] pc_wb_o;
wire [31:0] pc_wb_o;
/* cellift = 32'd1 */
output [31:0] pc_wb_o_t0;
wire [31:0] pc_wb_o_t0;
/* src = "generated/sv2v_out.v:20960.14-20960.44" */
output perf_instr_ret_compressed_wb_o;
wire perf_instr_ret_compressed_wb_o;
/* cellift = 32'd1 */
output perf_instr_ret_compressed_wb_o_t0;
wire perf_instr_ret_compressed_wb_o_t0;
/* src = "generated/sv2v_out.v:20962.14-20962.49" */
output perf_instr_ret_compressed_wb_spec_o;
wire perf_instr_ret_compressed_wb_spec_o;
/* cellift = 32'd1 */
output perf_instr_ret_compressed_wb_spec_o_t0;
wire perf_instr_ret_compressed_wb_spec_o_t0;
/* src = "generated/sv2v_out.v:20959.14-20959.33" */
output perf_instr_ret_wb_o;
wire perf_instr_ret_wb_o;
/* cellift = 32'd1 */
output perf_instr_ret_wb_o_t0;
wire perf_instr_ret_wb_o_t0;
/* src = "generated/sv2v_out.v:20961.14-20961.38" */
output perf_instr_ret_wb_spec_o;
wire perf_instr_ret_wb_spec_o;
/* cellift = 32'd1 */
output perf_instr_ret_wb_spec_o_t0;
wire perf_instr_ret_wb_spec_o_t0;
/* src = "generated/sv2v_out.v:20954.14-20954.24" */
output ready_wb_o;
wire ready_wb_o;
/* cellift = 32'd1 */
output ready_wb_o_t0;
wire ready_wb_o_t0;
/* src = "generated/sv2v_out.v:20963.19-20963.32" */
input [4:0] rf_waddr_id_i;
wire [4:0] rf_waddr_id_i;
/* cellift = 32'd1 */
input [4:0] rf_waddr_id_i_t0;
wire [4:0] rf_waddr_id_i_t0;
/* src = "generated/sv2v_out.v:20970.20-20970.33" */
output [4:0] rf_waddr_wb_o;
wire [4:0] rf_waddr_wb_o;
/* cellift = 32'd1 */
output [4:0] rf_waddr_wb_o_t0;
wire [4:0] rf_waddr_wb_o_t0;
/* src = "generated/sv2v_out.v:20969.21-20969.38" */
output [31:0] rf_wdata_fwd_wb_o;
wire [31:0] rf_wdata_fwd_wb_o;
/* cellift = 32'd1 */
output [31:0] rf_wdata_fwd_wb_o_t0;
wire [31:0] rf_wdata_fwd_wb_o_t0;
/* src = "generated/sv2v_out.v:20964.20-20964.33" */
input [31:0] rf_wdata_id_i;
wire [31:0] rf_wdata_id_i;
/* cellift = 32'd1 */
input [31:0] rf_wdata_id_i_t0;
wire [31:0] rf_wdata_id_i_t0;
/* src = "generated/sv2v_out.v:20967.20-20967.34" */
input [31:0] rf_wdata_lsu_i;
wire [31:0] rf_wdata_lsu_i;
/* cellift = 32'd1 */
input [31:0] rf_wdata_lsu_i_t0;
wire [31:0] rf_wdata_lsu_i_t0;
/* src = "generated/sv2v_out.v:20971.21-20971.34" */
output [31:0] rf_wdata_wb_o;
wire [31:0] rf_wdata_wb_o;
/* cellift = 32'd1 */
output [31:0] rf_wdata_wb_o_t0;
wire [31:0] rf_wdata_wb_o_t0;
/* src = "generated/sv2v_out.v:20965.13-20965.23" */
input rf_we_id_i;
wire rf_we_id_i;
/* cellift = 32'd1 */
input rf_we_id_i_t0;
wire rf_we_id_i_t0;
/* src = "generated/sv2v_out.v:20968.13-20968.24" */
input rf_we_lsu_i;
wire rf_we_lsu_i;
/* cellift = 32'd1 */
input rf_we_lsu_i_t0;
wire rf_we_lsu_i_t0;
/* src = "generated/sv2v_out.v:20972.14-20972.24" */
output rf_we_wb_o;
wire rf_we_wb_o;
/* cellift = 32'd1 */
output rf_we_wb_o_t0;
wire rf_we_wb_o_t0;
/* src = "generated/sv2v_out.v:20955.14-20955.27" */
output rf_write_wb_o;
wire rf_write_wb_o;
/* cellift = 32'd1 */
output rf_write_wb_o_t0;
wire rf_write_wb_o_t0;
/* src = "generated/sv2v_out.v:20948.13-20948.19" */
input rst_ni;
wire rst_ni;
assign _00_ = instr_perf_count_id_i & /* src = "generated/sv2v_out.v:21076.34-21076.65" */ en_wb_i;
assign _02_ = lsu_resp_valid_i & /* src = "generated/sv2v_out.v:21076.71-21076.104" */ lsu_resp_err_i;
assign perf_instr_ret_wb_o = _00_ & /* src = "generated/sv2v_out.v:21076.33-21076.105" */ _38_;
assign perf_instr_ret_compressed_wb_o = perf_instr_ret_wb_o & /* src = "generated/sv2v_out.v:21077.44-21077.90" */ instr_is_compressed_id_i;
assign _04_ = { rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i } & /* src = "generated/sv2v_out.v:21098.26-21098.75" */ rf_wdata_id_i;
assign _06_ = { rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i } & /* src = "generated/sv2v_out.v:21098.80-21098.129" */ rf_wdata_lsu_i;
assign _10_ = instr_perf_count_id_i_t0 & en_wb_i;
assign _13_ = lsu_resp_valid_i_t0 & lsu_resp_err_i;
assign _16_ = _01_ & _38_;
assign _19_ = perf_instr_ret_wb_o_t0 & instr_is_compressed_id_i;
assign _22_ = { rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0 } & rf_wdata_id_i;
assign _25_ = { rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0 } & rf_wdata_lsu_i;
assign _11_ = en_wb_i_t0 & instr_perf_count_id_i;
assign _14_ = lsu_resp_err_i_t0 & lsu_resp_valid_i;
assign _17_ = _03_ & _00_;
assign _20_ = instr_is_compressed_id_i_t0 & perf_instr_ret_wb_o;
assign _23_ = rf_wdata_id_i_t0 & { rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i };
assign _26_ = rf_wdata_lsu_i_t0 & { rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i };
assign _12_ = instr_perf_count_id_i_t0 & en_wb_i_t0;
assign _15_ = lsu_resp_valid_i_t0 & lsu_resp_err_i_t0;
assign _18_ = _01_ & _03_;
assign _21_ = perf_instr_ret_wb_o_t0 & instr_is_compressed_id_i_t0;
assign _24_ = { rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0 } & rf_wdata_id_i_t0;
assign _27_ = { rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0 } & rf_wdata_lsu_i_t0;
assign _31_ = _10_ | _11_;
assign _32_ = _13_ | _14_;
assign _33_ = _16_ | _17_;
assign _34_ = _19_ | _20_;
assign _35_ = _22_ | _23_;
assign _36_ = _25_ | _26_;
assign _01_ = _31_ | _12_;
assign _03_ = _32_ | _15_;
assign perf_instr_ret_wb_o_t0 = _33_ | _18_;
assign perf_instr_ret_compressed_wb_o_t0 = _34_ | _21_;
assign _05_ = _35_ | _24_;
assign _07_ = _36_ | _27_;
assign _08_ = ~ _04_;
assign _09_ = ~ _06_;
assign _28_ = _05_ & _09_;
assign _29_ = _07_ & _08_;
assign _30_ = _05_ & _07_;
assign _37_ = _28_ | _29_;
assign rf_wdata_wb_o_t0 = _37_ | _30_;
assign _38_ = ~ /* src = "generated/sv2v_out.v:21076.69-21076.105" */ _02_;
assign rf_wdata_wb_o = _04_ | /* src = "generated/sv2v_out.v:21098.25-21098.130" */ _06_;
assign rf_we_wb_o = | /* src = "generated/sv2v_out.v:21099.22-21099.41" */ { rf_we_lsu_i, rf_we_id_i };
assign dummy_instr_wb_o = dummy_instr_id_i;
assign dummy_instr_wb_o_t0 = dummy_instr_id_i_t0;
assign instr_done_wb_o = 1'h0;
assign instr_done_wb_o_t0 = 1'h0;
assign outstanding_load_wb_o = 1'h0;
assign outstanding_load_wb_o_t0 = 1'h0;
assign outstanding_store_wb_o = 1'h0;
assign outstanding_store_wb_o_t0 = 1'h0;
assign pc_wb_o = 32'd0;
assign pc_wb_o_t0 = 32'd0;
assign perf_instr_ret_compressed_wb_spec_o = 1'h0;
assign perf_instr_ret_compressed_wb_spec_o_t0 = 1'h0;
assign perf_instr_ret_wb_spec_o = 1'h0;
assign perf_instr_ret_wb_spec_o_t0 = 1'h0;
assign ready_wb_o = 1'h1;
assign ready_wb_o_t0 = 1'h0;
assign rf_waddr_wb_o = rf_waddr_id_i;
assign rf_waddr_wb_o_t0 = rf_waddr_id_i_t0;
assign rf_wdata_fwd_wb_o = 32'd0;
assign rf_wdata_fwd_wb_o_t0 = 32'd0;
assign rf_we_wb_o_t0 = 1'h0;
assign rf_write_wb_o = 1'h0;
assign rf_write_wb_o_t0 = 1'h0;
endmodule

module \$paramod\prim_buf\Width=32'00000000000000000000000000001100 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23046.22-23046.26" */
input [11:0] in_i;
wire [11:0] in_i;
/* cellift = 32'd1 */
input [11:0] in_i_t0;
wire [11:0] in_i_t0;
/* src = "generated/sv2v_out.v:23047.28-23047.33" */
output [11:0] out_o;
wire [11:0] out_o;
/* cellift = 32'd1 */
output [11:0] out_o_t0;
wire [11:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23057.38-23060.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000001100  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_buf\Width=32'00000000000000000000000000100000 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23046.22-23046.26" */
input [31:0] in_i;
wire [31:0] in_i;
/* cellift = 32'd1 */
input [31:0] in_i_t0;
wire [31:0] in_i_t0;
/* src = "generated/sv2v_out.v:23047.28-23047.33" */
output [31:0] out_o;
wire [31:0] out_o;
/* cellift = 32'd1 */
output [31:0] out_o_t0;
wire [31:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23057.38-23060.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000100000  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_buf\Width=32'00000000000000000000000000100111 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23046.22-23046.26" */
input [38:0] in_i;
wire [38:0] in_i;
/* cellift = 32'd1 */
input [38:0] in_i_t0;
wire [38:0] in_i_t0;
/* src = "generated/sv2v_out.v:23047.28-23047.33" */
output [38:0] out_o;
wire [38:0] out_o;
/* cellift = 32'd1 */
output [38:0] out_o_t0;
wire [38:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23057.38-23060.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000100111  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_buf\Width=s32'00000000000000000000000000000100 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23046.22-23046.26" */
input [3:0] in_i;
wire [3:0] in_i;
/* cellift = 32'd1 */
input [3:0] in_i_t0;
wire [3:0] in_i_t0;
/* src = "generated/sv2v_out.v:23047.28-23047.33" */
output [3:0] out_o;
wire [3:0] out_o;
/* cellift = 32'd1 */
output [3:0] out_o_t0;
wire [3:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23057.38-23060.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000000100  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_buf\Width=s32'00000000000000000000000000000111 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23046.22-23046.26" */
input [6:0] in_i;
wire [6:0] in_i;
/* cellift = 32'd1 */
input [6:0] in_i_t0;
wire [6:0] in_i_t0;
/* src = "generated/sv2v_out.v:23047.28-23047.33" */
output [6:0] out_o;
wire [6:0] out_o;
/* cellift = 32'd1 */
output [6:0] out_o_t0;
wire [6:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23057.38-23060.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000000111  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_buf\Width=s32'00000000000000000000000000100000 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23046.22-23046.26" */
input [31:0] in_i;
wire [31:0] in_i;
/* cellift = 32'd1 */
input [31:0] in_i_t0;
wire [31:0] in_i_t0;
/* src = "generated/sv2v_out.v:23047.28-23047.33" */
output [31:0] out_o;
wire [31:0] out_o;
/* cellift = 32'd1 */
output [31:0] out_o_t0;
wire [31:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23057.38-23060.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000100000  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_generic_buf\Width=s32'00000000000000000000000000000100 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:24893.22-24893.26" */
input [3:0] in_i;
wire [3:0] in_i;
/* cellift = 32'd1 */
input [3:0] in_i_t0;
wire [3:0] in_i_t0;
/* src = "generated/sv2v_out.v:24895.21-24895.24" */
wire [3:0] inv;
/* src = "generated/sv2v_out.v:24894.28-24894.33" */
output [3:0] out_o;
wire [3:0] out_o;
/* cellift = 32'd1 */
output [3:0] out_o_t0;
wire [3:0] out_o_t0;
assign inv = ~ /* src = "generated/sv2v_out.v:24896.15-24896.20" */ in_i;
assign out_o = ~ /* src = "generated/sv2v_out.v:24897.17-24897.21" */ inv;
assign out_o_t0 = in_i_t0;
endmodule

module \$paramod\prim_generic_buf\Width=s32'00000000000000000000000000000111 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:24893.22-24893.26" */
input [6:0] in_i;
wire [6:0] in_i;
/* cellift = 32'd1 */
input [6:0] in_i_t0;
wire [6:0] in_i_t0;
/* src = "generated/sv2v_out.v:24895.21-24895.24" */
wire [6:0] inv;
/* src = "generated/sv2v_out.v:24894.28-24894.33" */
output [6:0] out_o;
wire [6:0] out_o;
/* cellift = 32'd1 */
output [6:0] out_o_t0;
wire [6:0] out_o_t0;
assign inv = ~ /* src = "generated/sv2v_out.v:24896.15-24896.20" */ in_i;
assign out_o = ~ /* src = "generated/sv2v_out.v:24897.17-24897.21" */ inv;
assign out_o_t0 = in_i_t0;
endmodule

module \$paramod\prim_generic_buf\Width=s32'00000000000000000000000000001100 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:24893.22-24893.26" */
input [11:0] in_i;
wire [11:0] in_i;
/* cellift = 32'd1 */
input [11:0] in_i_t0;
wire [11:0] in_i_t0;
/* src = "generated/sv2v_out.v:24895.21-24895.24" */
wire [11:0] inv;
/* src = "generated/sv2v_out.v:24894.28-24894.33" */
output [11:0] out_o;
wire [11:0] out_o;
/* cellift = 32'd1 */
output [11:0] out_o_t0;
wire [11:0] out_o_t0;
assign inv = ~ /* src = "generated/sv2v_out.v:24896.15-24896.20" */ in_i;
assign out_o = ~ /* src = "generated/sv2v_out.v:24897.17-24897.21" */ inv;
assign out_o_t0 = in_i_t0;
endmodule

module \$paramod\prim_generic_buf\Width=s32'00000000000000000000000000100000 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:24893.22-24893.26" */
input [31:0] in_i;
wire [31:0] in_i;
/* cellift = 32'd1 */
input [31:0] in_i_t0;
wire [31:0] in_i_t0;
/* src = "generated/sv2v_out.v:24895.21-24895.24" */
wire [31:0] inv;
/* src = "generated/sv2v_out.v:24894.28-24894.33" */
output [31:0] out_o;
wire [31:0] out_o;
/* cellift = 32'd1 */
output [31:0] out_o_t0;
wire [31:0] out_o_t0;
assign inv = ~ /* src = "generated/sv2v_out.v:24896.15-24896.20" */ in_i;
assign out_o = ~ /* src = "generated/sv2v_out.v:24897.17-24897.21" */ inv;
assign out_o_t0 = in_i_t0;
endmodule

module \$paramod\prim_generic_buf\Width=s32'00000000000000000000000000100111 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:24893.22-24893.26" */
input [38:0] in_i;
wire [38:0] in_i;
/* cellift = 32'd1 */
input [38:0] in_i_t0;
wire [38:0] in_i_t0;
/* src = "generated/sv2v_out.v:24895.21-24895.24" */
wire [38:0] inv;
/* src = "generated/sv2v_out.v:24894.28-24894.33" */
output [38:0] out_o;
wire [38:0] out_o;
/* cellift = 32'd1 */
output [38:0] out_o_t0;
wire [38:0] out_o_t0;
assign inv = ~ /* src = "generated/sv2v_out.v:24896.15-24896.20" */ in_i;
assign out_o = ~ /* src = "generated/sv2v_out.v:24897.17-24897.21" */ inv;
assign out_o_t0 = in_i_t0;
endmodule

module ibex_compressed_decoder(clk_i, rst_ni, valid_i, instr_i, instr_o, is_compressed_o, illegal_instr_o, instr_o_t0, instr_i_t0, illegal_instr_o_t0, is_compressed_o_t0, valid_i_t0);
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _000_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _001_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _002_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _003_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _005_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _006_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _007_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _008_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _009_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _010_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _011_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _013_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _014_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _015_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _016_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _017_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _018_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _019_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _020_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _021_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _022_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _023_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _024_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _025_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _026_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _027_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _028_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _029_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _030_;
wire [31:0] _031_;
wire [31:0] _032_;
wire [31:0] _033_;
wire [31:0] _034_;
wire [31:0] _035_;
wire [31:0] _036_;
wire [31:0] _037_;
wire [31:0] _038_;
wire [31:0] _039_;
wire [31:0] _040_;
wire [31:0] _041_;
wire [31:0] _042_;
wire [31:0] _043_;
wire [31:0] _044_;
wire [31:0] _045_;
wire [31:0] _046_;
wire [31:0] _047_;
wire [31:0] _048_;
wire [31:0] _049_;
wire [31:0] _050_;
wire [31:0] _051_;
wire [31:0] _052_;
wire _053_;
wire _054_;
wire _055_;
wire [31:0] _056_;
wire [31:0] _057_;
wire [31:0] _058_;
wire [31:0] _059_;
wire [31:0] _060_;
wire [31:0] _061_;
wire [31:0] _062_;
wire [31:0] _063_;
wire [31:0] _064_;
wire [31:0] _065_;
wire [31:0] _066_;
wire [31:0] _067_;
wire [31:0] _068_;
wire [31:0] _069_;
wire [31:0] _070_;
wire [31:0] _071_;
wire [31:0] _072_;
wire [31:0] _073_;
wire [31:0] _074_;
wire [31:0] _075_;
wire [31:0] _076_;
wire [31:0] _077_;
wire [31:0] _078_;
wire [31:0] _079_;
wire [31:0] _080_;
wire [31:0] _081_;
wire [31:0] _082_;
wire [31:0] _083_;
wire [31:0] _084_;
wire [31:0] _085_;
wire [31:0] _086_;
wire [31:0] _087_;
wire [31:0] _088_;
wire [31:0] _089_;
wire [31:0] _090_;
wire [31:0] _091_;
wire [31:0] _092_;
wire [31:0] _093_;
wire [31:0] _094_;
wire [31:0] _095_;
wire [31:0] _096_;
wire [31:0] _097_;
wire [31:0] _098_;
wire [31:0] _099_;
wire [31:0] _100_;
wire [31:0] _101_;
wire [31:0] _102_;
wire [31:0] _103_;
wire [31:0] _104_;
wire [31:0] _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire [31:0] _113_;
/* cellift = 32'd1 */
wire [31:0] _114_;
wire [31:0] _115_;
/* cellift = 32'd1 */
wire [31:0] _116_;
wire [31:0] _117_;
/* cellift = 32'd1 */
wire [31:0] _118_;
wire [31:0] _119_;
/* cellift = 32'd1 */
wire [31:0] _120_;
wire [31:0] _121_;
/* cellift = 32'd1 */
wire [31:0] _122_;
wire [31:0] _123_;
/* cellift = 32'd1 */
wire [31:0] _124_;
wire _125_;
wire [31:0] _126_;
/* cellift = 32'd1 */
wire [31:0] _127_;
wire [31:0] _128_;
/* cellift = 32'd1 */
wire [31:0] _129_;
wire [31:0] _130_;
/* cellift = 32'd1 */
wire [31:0] _131_;
wire [31:0] _132_;
/* cellift = 32'd1 */
wire [31:0] _133_;
wire [31:0] _134_;
/* cellift = 32'd1 */
wire [31:0] _135_;
wire _136_;
wire _137_;
wire [31:0] _138_;
/* cellift = 32'd1 */
wire [31:0] _139_;
wire [31:0] _140_;
/* cellift = 32'd1 */
wire [31:0] _141_;
wire _142_;
wire _143_;
wire [31:0] _144_;
/* cellift = 32'd1 */
wire [31:0] _145_;
wire [31:0] _146_;
/* cellift = 32'd1 */
wire [31:0] _147_;
/* src = "generated/sv2v_out.v:12058.11-12058.39" */
wire _148_;
/* src = "generated/sv2v_out.v:12073.11-12073.33" */
wire _149_;
/* src = "generated/sv2v_out.v:12075.11-12075.51" */
wire _150_;
/* src = "generated/sv2v_out.v:12109.11-12109.36" */
wire _151_;
/* src = "generated/sv2v_out.v:12114.12-12114.36" */
wire _152_;
/* src = "generated/sv2v_out.v:12069.164-12069.176" */
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire [3:0] _158_;
wire _159_;
wire _160_;
wire [3:0] _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
/* src = "generated/sv2v_out.v:12041.13-12041.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:12047.13-12047.28" */
output illegal_instr_o;
wire illegal_instr_o;
/* cellift = 32'd1 */
output illegal_instr_o_t0;
wire illegal_instr_o_t0;
/* src = "generated/sv2v_out.v:12044.20-12044.27" */
input [31:0] instr_i;
wire [31:0] instr_i;
/* cellift = 32'd1 */
input [31:0] instr_i_t0;
wire [31:0] instr_i_t0;
/* src = "generated/sv2v_out.v:12045.20-12045.27" */
output [31:0] instr_o;
wire [31:0] instr_o;
/* cellift = 32'd1 */
output [31:0] instr_o_t0;
wire [31:0] instr_o_t0;
/* src = "generated/sv2v_out.v:12046.14-12046.29" */
output is_compressed_o;
wire is_compressed_o;
/* cellift = 32'd1 */
output is_compressed_o_t0;
wire is_compressed_o_t0;
/* src = "generated/sv2v_out.v:12042.13-12042.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:12043.13-12043.20" */
input valid_i;
wire valid_i;
/* cellift = 32'd1 */
input valid_i_t0;
wire valid_i_t0;
assign _031_ = ~ { _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_ };
assign _032_ = ~ { _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_ };
assign _033_ = ~ { _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_ };
assign _034_ = ~ { _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_ };
assign _035_ = ~ { _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_ };
assign _036_ = ~ { _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_ };
assign _037_ = ~ { _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_ };
assign _038_ = ~ { _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_ };
assign _039_ = ~ { _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_ };
assign _040_ = ~ { _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_ };
assign _041_ = ~ { _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_ };
assign _042_ = ~ { _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_ };
assign _043_ = ~ { _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_ };
assign _044_ = ~ { _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_ };
assign _045_ = ~ { _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_ };
assign _046_ = ~ { _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_ };
assign _047_ = ~ { _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_ };
assign _048_ = ~ { _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_ };
assign _049_ = ~ { _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_ };
assign _050_ = ~ { _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_ };
assign _051_ = ~ { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12] };
assign _052_ = ~ { _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_ };
assign _056_ = _031_ & { 4'h0, instr_i_t0[8:7], instr_i_t0[12], instr_i_t0[6:2], 8'h00, instr_i_t0[11:9], 9'h000 };
assign _058_ = _032_ & { 7'h00, instr_i_t0[6:2], instr_i_t0[11:7], 3'h0, instr_i_t0[11:7], 7'h00 };
assign _060_ = _033_ & _116_;
assign _062_ = _034_ & _118_;
assign _064_ = _035_ & { 9'h000, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 };
assign _066_ = _036_ & { 9'h000, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 };
assign _068_ = _037_ & _122_;
assign _070_ = _038_ & _124_;
assign _072_ = _039_ & { 1'h0, instr_i_t0[10], 5'h00, instr_i_t0[6:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 };
assign _074_ = _040_ & _127_;
assign _076_ = _033_ & _016_;
assign _078_ = _041_ & _129_;
assign _080_ = _042_ & { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:2], instr_i_t0[11:7], 3'h0, instr_i_t0[11:7], 7'h00 };
assign _082_ = _032_ & _133_;
assign _084_ = _043_ & _135_;
assign _086_ = _044_ & { 5'h00, instr_i_t0[5], instr_i_t0[12], 2'h0, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 3'h0, instr_i_t0[11:10], instr_i_t0[6], 9'h000 };
assign _088_ = _032_ & { 2'h0, instr_i_t0[10:7], instr_i_t0[12:11], instr_i_t0[5], instr_i_t0[6], 12'h000, instr_i_t0[4:2], 7'h00 };
assign _090_ = _045_ & _141_;
assign _092_ = _046_ & _024_;
assign _094_ = _047_ & _010_;
assign _096_ = _048_ & _147_;
assign _005_ = _049_ & { 12'h000, instr_i_t0[11:7], 15'h0000 };
assign _098_ = _050_ & _005_;
assign _100_ = _050_ & { 12'h000, instr_i_t0[11:7], 15'h0000 };
assign _102_ = _051_ & _030_;
assign _104_ = _052_ & { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:2], instr_i_t0[11:7], 7'h00 };
assign _057_ = { _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_ } & instr_i_t0;
assign _059_ = { _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_ } & { 4'h0, instr_i_t0[3:2], instr_i_t0[12], instr_i_t0[6:4], 10'h000, instr_i_t0[11:7], 7'h00 };
assign _061_ = { _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_ } & _027_;
assign _063_ = { _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_ } & _114_;
assign _065_ = { _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_ } & instr_i_t0;
assign _067_ = { _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_ } & { 9'h000, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 };
assign _069_ = { _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_ } & { 9'h000, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 };
assign _071_ = { _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_ } & _120_;
assign _073_ = { _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_ } & { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 };
assign _075_ = { _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_ } & _022_;
assign _077_ = { _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_ } & _019_;
assign _079_ = { _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_ } & { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:5], instr_i_t0[2], 7'h00, instr_i_t0[9:7], 2'h0, instr_i_t0[13], instr_i_t0[11:10], instr_i_t0[4:3], instr_i_t0[12], 7'h00 };
assign _081_ = { _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_ } & { instr_i_t0[12], instr_i_t0[8], instr_i_t0[10:9], instr_i_t0[6], instr_i_t0[7], instr_i_t0[2], instr_i_t0[11], instr_i_t0[5:3], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], 4'h0, instr_i_t0[15], 7'h00 };
assign _083_ = { _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_ } & { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:2], 8'h00, instr_i_t0[11:7], 7'h00 };
assign _085_ = { _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_ } & _131_;
assign _087_ = { _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_ } & instr_i_t0;
assign _089_ = { _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_ } & { 5'h00, instr_i_t0[5], instr_i_t0[12:10], instr_i_t0[6], 4'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[4:2], 7'h00 };
assign _091_ = { _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_ } & _139_;
assign _093_ = { _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_ } & instr_i_t0;
assign _095_ = { _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_ } & _013_;
assign _097_ = { _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_ } & _145_;
assign _099_ = { _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_ } & { 7'h00, instr_i_t0[6:2], instr_i_t0[11:7], 3'h0, instr_i_t0[11:7], 7'h00 };
assign _101_ = { _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_ } & { 7'h00, instr_i_t0[6:2], 8'h00, instr_i_t0[11:7], 7'h00 };
assign _103_ = { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12] } & _002_;
assign _105_ = { _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_ } & { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[4:3], instr_i_t0[5], instr_i_t0[2], instr_i_t0[6], 24'h000000 };
assign _114_ = _056_ | _057_;
assign _116_ = _058_ | _059_;
assign _118_ = _060_ | _061_;
assign _024_ = _062_ | _063_;
assign _120_ = _064_ | _065_;
assign _122_ = _066_ | _067_;
assign _124_ = _068_ | _069_;
assign _022_ = _070_ | _071_;
assign _127_ = _072_ | _073_;
assign _019_ = _074_ | _075_;
assign _129_ = _076_ | _077_;
assign _131_ = _078_ | _079_;
assign _133_ = _080_ | _081_;
assign _135_ = _082_ | _083_;
assign _013_ = _084_ | _085_;
assign _139_ = _086_ | _087_;
assign _141_ = _088_ | _089_;
assign _010_ = _090_ | _091_;
assign _145_ = _092_ | _093_;
assign _147_ = _094_ | _095_;
assign instr_o_t0 = _096_ | _097_;
assign _002_ = _098_ | _099_;
assign _030_ = _100_ | _101_;
assign _027_ = _102_ | _103_;
assign _016_ = _104_ | _105_;
assign _054_ = | { _160_, _156_ };
assign _055_ = | { _160_, _158_[3:2], _158_[0], _157_, _156_ };
assign _106_ = _160_ | _159_;
assign _107_ = _163_ | _162_;
assign _108_ = _160_ | _171_;
assign _109_ = _155_ | _172_;
assign _053_ = | { _160_, _158_[3], _158_[1], _154_ };
assign _110_ = _159_ ? 1'h1 : 1'h0;
assign _111_ = _156_ ? _003_ : _000_;
assign _112_ = _154_ ? _006_ : _111_;
assign _028_ = _106_ ? _110_ : _112_;
assign _113_ = _159_ ? instr_i : { 4'h0, instr_i[8:7], instr_i[12], instr_i[6:2], 8'h12, instr_i[11:9], 9'h023 };
assign _115_ = _156_ ? { 4'h0, instr_i[3:2], instr_i[12], instr_i[6:4], 10'h012, instr_i[11:7], 7'h03 } : { 7'h00, instr_i[6:2], instr_i[11:7], 3'h1, instr_i[11:7], 7'h13 };
assign _117_ = _154_ ? _026_ : _115_;
assign _023_ = _106_ ? _113_ : _117_;
assign _119_ = _162_ ? instr_i : { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h1d, instr_i[9:7], 7'h33 };
assign _121_ = _165_ ? { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h11, instr_i[9:7], 7'h33 } : { 9'h081, instr_i[4:2], 2'h1, instr_i[9:7], 5'h01, instr_i[9:7], 7'h33 };
assign _123_ = _164_ ? { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h19, instr_i[9:7], 7'h33 } : _121_;
assign _021_ = _107_ ? _119_ : _123_;
assign _025_ = _162_ ? 1'h1 : 1'h0;
assign _125_ = _168_ ? 1'h0 : _000_;
assign _020_ = _166_ ? _025_ : _125_;
assign _126_ = _168_ ? { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], 2'h1, instr_i[9:7], 5'h1d, instr_i[9:7], 7'h13 } : { 1'h0, instr_i[10], 5'h00, instr_i[6:2], 2'h1, instr_i[9:7], 5'h15, instr_i[9:7], 7'h13 };
assign _018_ = _166_ ? _021_ : _126_;
assign _128_ = _154_ ? _018_ : _015_;
assign _130_ = _169_ ? { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:5], instr_i[2], 7'h01, instr_i[9:7], 2'h0, instr_i[13], instr_i[11:10], instr_i[4:3], instr_i[12], 7'h63 } : _128_;
assign _132_ = _170_ ? { instr_i[12], instr_i[8], instr_i[10:9], instr_i[6], instr_i[7], instr_i[2], instr_i[11], instr_i[5:3], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], 4'h0, _153_, 7'h6f } : { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], instr_i[11:7], 3'h0, instr_i[11:7], 7'h13 };
assign _134_ = _156_ ? { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], 8'h00, instr_i[11:7], 7'h13 } : _132_;
assign _012_ = _053_ ? _130_ : _134_;
assign _136_ = _154_ ? _020_ : _017_;
assign _014_ = _055_ ? 1'h0 : _136_;
assign _137_ = _054_ ? 1'h0 : _011_;
assign _008_ = _171_ ? 1'h1 : _137_;
assign _138_ = _171_ ? instr_i : { 5'h00, instr_i[5], instr_i[12], 2'h1, instr_i[4:2], 2'h1, instr_i[9:7], 3'h2, instr_i[11:10], instr_i[6], 9'h023 };
assign _140_ = _156_ ? { 5'h00, instr_i[5], instr_i[12:10], instr_i[6], 4'h1, instr_i[9:7], 5'h09, instr_i[4:2], 7'h03 } : { 2'h0, instr_i[10:7], instr_i[12:11], instr_i[5], instr_i[6], 12'h041, instr_i[4:2], 7'h13 };
assign _009_ = _108_ ? _138_ : _140_;
assign _142_ = _172_ ? 1'h0 : _028_;
assign _143_ = _167_ ? _014_ : _008_;
assign illegal_instr_o = _109_ ? _142_ : _143_;
assign _144_ = _172_ ? instr_i : _023_;
assign _146_ = _167_ ? _012_ : _009_;
assign instr_o = _109_ ? _144_ : _146_;
assign _148_ = ! /* src = "generated/sv2v_out.v:12058.11-12058.39" */ instr_i[12:5];
assign _149_ = instr_i[11:7] == /* src = "generated/sv2v_out.v:12073.11-12073.33" */ 5'h02;
assign _150_ = ! /* src = "generated/sv2v_out.v:12075.11-12075.51" */ { instr_i[12], instr_i[6:2] };
assign _151_ = ! /* src = "generated/sv2v_out.v:12124.16-12124.41" */ instr_i[11:7];
assign _152_ = | /* src = "generated/sv2v_out.v:12122.16-12122.40" */ instr_i[6:2];
assign is_compressed_o = instr_i[1:0] != /* src = "generated/sv2v_out.v:12137.27-12137.48" */ 2'h3;
assign _153_ = ~ /* src = "generated/sv2v_out.v:12069.164-12069.176" */ instr_i[15];
assign _004_ = _151_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12124.16-12124.41|generated/sv2v_out.v:12124.12-12127.77" */ 32'd1048691 : { 12'h000, instr_i[11:7], 15'h00e7 };
assign _001_ = _152_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12122.16-12122.40|generated/sv2v_out.v:12122.12-12127.77" */ { 7'h00, instr_i[6:2], instr_i[11:7], 3'h0, instr_i[11:7], 7'h33 } : _004_;
assign _029_ = _152_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12114.12-12114.36|generated/sv2v_out.v:12114.8-12120.11" */ { 7'h00, instr_i[6:2], 8'h00, instr_i[11:7], 7'h33 } : { 12'h000, instr_i[11:7], 15'h0067 };
assign _007_ = _152_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12114.12-12114.36|generated/sv2v_out.v:12114.8-12120.11" */ 1'h0 : _003_;
assign _006_ = instr_i[12] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12113.11-12113.30|generated/sv2v_out.v:12113.7-12127.77" */ 1'h0 : _007_;
assign _026_ = instr_i[12] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12113.11-12113.30|generated/sv2v_out.v:12113.7-12127.77" */ _001_ : _029_;
assign _003_ = _151_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12109.11-12109.36|generated/sv2v_out.v:12109.7-12110.31" */ 1'h1 : 1'h0;
assign _000_ = instr_i[12] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12104.11-12104.30|generated/sv2v_out.v:12104.7-12105.31" */ 1'h1 : 1'h0;
assign _159_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12101.5-12131.12" */ _158_;
assign _162_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12087.9-12094.16" */ _161_;
assign _161_[0] = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12087.9-12094.16" */ 3'h4;
assign _161_[1] = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12087.9-12094.16" */ 3'h5;
assign _161_[2] = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12087.9-12094.16" */ 3'h6;
assign _161_[3] = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12087.9-12094.16" */ 3'h7;
assign _163_ = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12087.9-12094.16" */ 3'h3;
assign _164_ = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12087.9-12094.16" */ 3'h2;
assign _165_ = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12087.9-12094.16" */ 3'h1;
assign _166_ = instr_i[11:10] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12079.7-12096.14" */ 2'h3;
assign _168_ = instr_i[11:10] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12079.7-12096.14" */ 2'h2;
assign _017_ = _150_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12075.11-12075.51|generated/sv2v_out.v:12075.7-12076.31" */ 1'h1 : 1'h0;
assign _015_ = _149_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12073.11-12073.33|generated/sv2v_out.v:12073.7-12074.126" */ { instr_i[12], instr_i[12], instr_i[12], instr_i[4:3], instr_i[5], instr_i[2], instr_i[6], 24'h010113 } : { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], instr_i[11:7], 7'h37 };
assign _169_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12067.5-12099.12" */ { _160_, _158_[3] };
assign _170_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12067.5-12099.12" */ { _158_[2], _158_[0] };
assign _011_ = _148_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12058.11-12058.39|generated/sv2v_out.v:12058.7-12059.31" */ 1'h1 : 1'h0;
assign _171_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ { _158_, _154_ };
assign _158_[0] = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ 3'h1;
assign _158_[1] = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ 3'h3;
assign _154_ = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ 3'h4;
assign _158_[2] = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ 3'h5;
assign _158_[3] = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ 3'h7;
assign _160_ = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ 3'h6;
assign _156_ = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ 3'h2;
assign _157_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ instr_i[15:13];
assign _167_ = instr_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12053.3-12135.10" */ 2'h1;
assign _172_ = instr_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12053.3-12135.10" */ 2'h3;
assign _155_ = instr_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12053.3-12135.10" */ 2'h2;
assign illegal_instr_o_t0 = 1'h0;
assign is_compressed_o_t0 = 1'h0;
endmodule

module ibex_multdiv_slow(clk_i, rst_ni, mult_en_i, div_en_i, mult_sel_i, div_sel_i, operator_i, signed_mode_i, op_a_i, op_b_i, alu_adder_ext_i, alu_adder_i, equal_to_zero_i, data_ind_timing_i, alu_operand_a_o, alu_operand_b_o, imd_val_q_i, imd_val_d_o, imd_val_we_o, multdiv_ready_id_i, multdiv_result_o
, valid_o, valid_o_t0, alu_adder_ext_i_t0, alu_adder_i_t0, alu_operand_a_o_t0, alu_operand_b_o_t0, div_en_i_t0, div_sel_i_t0, equal_to_zero_i_t0, imd_val_d_o_t0, imd_val_q_i_t0, imd_val_we_o_t0, mult_en_i_t0, mult_sel_i_t0, multdiv_ready_id_i_t0, multdiv_result_o_t0, op_a_i_t0, op_b_i_t0, operator_i_t0, signed_mode_i_t0, data_ind_timing_i_t0
);
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _001_;
/* src = "generated/sv2v_out.v:19573.2-19606.5" */
wire [32:0] _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19573.2-19606.5" */
wire [32:0] _003_;
/* src = "generated/sv2v_out.v:19573.2-19606.5" */
wire [32:0] _004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19573.2-19606.5" */
wire [32:0] _005_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [2:0] _006_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [4:0] _007_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire _008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire _009_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _011_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _013_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [31:0] _014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [31:0] _015_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _016_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _017_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire _018_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [2:0] _019_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire _020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire _021_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _022_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _023_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _024_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _025_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _026_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _027_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [2:0] _028_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _029_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _030_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _031_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _032_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _033_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _034_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [2:0] _035_;
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _036_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19620.2-19732.5" */
wire [32:0] _037_;
/* src = "generated/sv2v_out.v:19635.55-19635.88" */
wire [31:0] _038_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19635.55-19635.88" */
wire [31:0] _039_;
/* src = "generated/sv2v_out.v:19635.28-19635.52" */
wire _040_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19635.28-19635.52" */
wire _041_;
/* src = "generated/sv2v_out.v:19641.61-19641.94" */
wire [30:0] _042_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19641.61-19641.94" */
wire [30:0] _043_;
/* src = "generated/sv2v_out.v:19749.43-19749.111" */
wire _044_;
wire _045_;
wire _046_;
wire [32:0] _047_;
wire [32:0] _048_;
wire _049_;
wire [32:0] _050_;
wire [32:0] _051_;
wire [32:0] _052_;
wire [32:0] _053_;
wire [32:0] _054_;
wire [32:0] _055_;
wire [32:0] _056_;
wire [32:0] _057_;
wire [32:0] _058_;
wire [32:0] _059_;
wire _060_;
wire [32:0] _061_;
wire [31:0] _062_;
wire [31:0] _063_;
wire [32:0] _064_;
wire [32:0] _065_;
wire [31:0] _066_;
wire [32:0] _067_;
wire [31:0] _068_;
wire [32:0] _069_;
wire [32:0] _070_;
wire [32:0] _071_;
wire [31:0] _072_;
wire [32:0] _073_;
wire _074_;
wire [32:0] _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire [31:0] _096_;
wire [31:0] _097_;
wire [31:0] _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire [31:0] _108_;
wire [31:0] _109_;
wire [31:0] _110_;
wire [30:0] _111_;
wire [30:0] _112_;
wire [30:0] _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire [32:0] _120_;
wire [32:0] _121_;
wire [32:0] _122_;
wire [32:0] _123_;
wire [32:0] _124_;
wire [32:0] _125_;
wire [32:0] _126_;
wire [32:0] _127_;
wire [32:0] _128_;
wire [32:0] _129_;
wire [32:0] _130_;
wire [32:0] _131_;
wire [32:0] _132_;
wire [32:0] _133_;
wire [32:0] _134_;
wire [32:0] _135_;
wire [32:0] _136_;
wire [32:0] _137_;
wire [32:0] _138_;
wire [32:0] _139_;
wire [32:0] _140_;
wire [32:0] _141_;
wire [32:0] _142_;
wire [32:0] _143_;
wire [32:0] _144_;
wire [32:0] _145_;
wire [32:0] _146_;
wire [32:0] _147_;
wire [32:0] _148_;
wire [32:0] _149_;
wire [32:0] _150_;
wire [32:0] _151_;
wire [32:0] _152_;
wire [32:0] _153_;
wire [32:0] _154_;
wire [32:0] _155_;
wire [32:0] _156_;
wire [32:0] _157_;
wire [32:0] _158_;
wire [32:0] _159_;
wire _160_;
wire _161_;
wire [32:0] _162_;
wire [32:0] _163_;
wire [32:0] _164_;
wire [32:0] _165_;
wire [32:0] _166_;
wire [32:0] _167_;
wire [32:0] _168_;
wire [32:0] _169_;
wire [32:0] _170_;
wire [32:0] _171_;
wire [32:0] _172_;
wire [32:0] _173_;
wire [32:0] _174_;
wire [32:0] _175_;
wire [32:0] _176_;
wire _177_;
wire _178_;
wire _179_;
wire [31:0] _180_;
wire [31:0] _181_;
wire [31:0] _182_;
wire [31:0] _183_;
wire [32:0] _184_;
wire [32:0] _185_;
wire [32:0] _186_;
wire [32:0] _187_;
wire [31:0] _188_;
wire [31:0] _189_;
wire [32:0] _190_;
wire [32:0] _191_;
wire [31:0] _192_;
wire [31:0] _193_;
wire [32:0] _194_;
wire [32:0] _195_;
wire [32:0] _196_;
wire [32:0] _197_;
wire [32:0] _198_;
wire [32:0] _199_;
wire [31:0] _200_;
wire [31:0] _201_;
wire _202_;
wire _203_;
wire _204_;
wire [31:0] _205_;
wire _206_;
wire _207_;
wire _208_;
wire [31:0] _209_;
wire [30:0] _210_;
wire _211_;
wire _212_;
wire [32:0] _213_;
wire [32:0] _214_;
wire [32:0] _215_;
wire _216_;
wire [32:0] _217_;
/* cellift = 32'd1 */
wire [32:0] _218_;
wire [32:0] _219_;
/* cellift = 32'd1 */
wire [32:0] _220_;
wire [32:0] _221_;
/* cellift = 32'd1 */
wire [32:0] _222_;
wire [2:0] _223_;
wire [32:0] _224_;
/* cellift = 32'd1 */
wire [32:0] _225_;
wire [32:0] _226_;
/* cellift = 32'd1 */
wire [32:0] _227_;
wire [32:0] _228_;
/* cellift = 32'd1 */
wire [32:0] _229_;
wire [32:0] _230_;
/* cellift = 32'd1 */
wire [32:0] _231_;
wire [32:0] _232_;
/* cellift = 32'd1 */
wire [32:0] _233_;
wire [32:0] _234_;
/* cellift = 32'd1 */
wire [32:0] _235_;
wire [32:0] _236_;
/* cellift = 32'd1 */
wire [32:0] _237_;
wire [32:0] _238_;
/* cellift = 32'd1 */
wire [32:0] _239_;
wire [2:0] _240_;
wire [2:0] _241_;
wire [2:0] _242_;
wire [2:0] _243_;
wire [2:0] _244_;
wire _245_;
/* cellift = 32'd1 */
wire _246_;
wire [32:0] _247_;
/* cellift = 32'd1 */
wire [32:0] _248_;
wire [32:0] _249_;
/* cellift = 32'd1 */
wire [32:0] _250_;
wire [32:0] _251_;
/* cellift = 32'd1 */
wire [32:0] _252_;
/* src = "generated/sv2v_out.v:19577.29-19577.47" */
wire _253_;
/* src = "generated/sv2v_out.v:19614.29-19614.67" */
wire _254_;
/* src = "generated/sv2v_out.v:19637.45-19637.65" */
wire _255_;
/* src = "generated/sv2v_out.v:19676.46-19676.63" */
wire _256_;
/* src = "generated/sv2v_out.v:19676.70-19676.93" */
wire _257_;
/* src = "generated/sv2v_out.v:19749.20-19749.38" */
wire _258_;
/* src = "generated/sv2v_out.v:19749.68-19749.86" */
wire _259_;
/* src = "generated/sv2v_out.v:19749.91-19749.109" */
wire _260_;
/* src = "generated/sv2v_out.v:19637.22-19637.66" */
wire _261_;
/* src = "generated/sv2v_out.v:19647.22-19647.59" */
wire _262_;
/* src = "generated/sv2v_out.v:19676.23-19676.64" */
wire _263_;
/* src = "generated/sv2v_out.v:19637.22-19637.40" */
wire _264_;
/* src = "generated/sv2v_out.v:19629.7-19629.30" */
wire _265_;
/* src = "generated/sv2v_out.v:19676.22-19676.94" */
wire _266_;
/* src = "generated/sv2v_out.v:19582.26-19582.33" */
wire [31:0] _267_;
/* src = "generated/sv2v_out.v:19586.26-19586.33" */
wire [31:0] _268_;
/* src = "generated/sv2v_out.v:19594.26-19594.47" */
wire [31:0] _269_;
/* src = "generated/sv2v_out.v:19598.26-19598.45" */
wire [31:0] _270_;
/* src = "generated/sv2v_out.v:19614.70-19614.86" */
wire _271_;
/* src = "generated/sv2v_out.v:19618.47-19618.61" */
wire _272_;
/* src = "generated/sv2v_out.v:19635.26-19635.53" */
wire _273_;
/* src = "generated/sv2v_out.v:19698.23-19698.42" */
wire _274_;
/* src = "generated/sv2v_out.v:19617.45-19617.69" */
wire [32:0] _275_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19617.45-19617.69" */
wire [32:0] _276_;
/* src = "generated/sv2v_out.v:19733.23-19733.43" */
wire _277_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19733.23-19733.43" */
wire _278_;
/* src = "generated/sv2v_out.v:19749.67-19749.110" */
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
/* src = "generated/sv2v_out.v:0.0-0.0" */
wire _287_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:0.0-0.0" */
wire _288_;
/* src = "generated/sv2v_out.v:19670.24-19670.47" */
wire [4:0] _289_;
/* src = "generated/sv2v_out.v:19577.29-19577.78" */
wire [32:0] _290_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19577.29-19577.78" */
wire [32:0] _291_;
/* src = "generated/sv2v_out.v:19637.22-19637.80" */
wire [2:0] _292_;
/* src = "generated/sv2v_out.v:19647.22-19647.73" */
wire [2:0] _293_;
/* src = "generated/sv2v_out.v:19661.24-19661.53" */
wire [31:0] _294_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19661.24-19661.53" */
wire [31:0] _295_;
/* src = "generated/sv2v_out.v:19666.22-19666.67" */
wire [32:0] _296_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19666.22-19666.67" */
wire [32:0] _297_;
/* src = "generated/sv2v_out.v:19676.22-19676.108" */
wire [2:0] _298_;
/* src = "generated/sv2v_out.v:19682.22-19682.59" */
wire [2:0] _299_;
/* src = "generated/sv2v_out.v:19720.31-19720.85" */
wire [32:0] _300_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19720.31-19720.85" */
wire [32:0] _301_;
/* src = "generated/sv2v_out.v:19721.31-19721.85" */
wire [32:0] _302_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19721.31-19721.85" */
wire [32:0] _303_;
/* src = "generated/sv2v_out.v:19618.28-19618.43" */
wire _304_;
/* src = "generated/sv2v_out.v:19533.13-19533.27" */
wire [32:0] accum_window_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19533.13-19533.27" */
wire [32:0] accum_window_d_t0;
/* src = "generated/sv2v_out.v:19518.20-19518.35" */
input [33:0] alu_adder_ext_i;
wire [33:0] alu_adder_ext_i;
/* cellift = 32'd1 */
input [33:0] alu_adder_ext_i_t0;
wire [33:0] alu_adder_ext_i_t0;
/* src = "generated/sv2v_out.v:19519.20-19519.31" */
input [31:0] alu_adder_i;
wire [31:0] alu_adder_i;
/* cellift = 32'd1 */
input [31:0] alu_adder_i_t0;
wire [31:0] alu_adder_i_t0;
/* src = "generated/sv2v_out.v:19522.20-19522.35" */
output [32:0] alu_operand_a_o;
wire [32:0] alu_operand_a_o;
/* cellift = 32'd1 */
output [32:0] alu_operand_a_o_t0;
wire [32:0] alu_operand_a_o_t0;
/* src = "generated/sv2v_out.v:19523.20-19523.35" */
output [32:0] alu_operand_b_o;
wire [32:0] alu_operand_b_o;
/* cellift = 32'd1 */
output [32:0] alu_operand_b_o_t0;
wire [32:0] alu_operand_b_o_t0;
/* src = "generated/sv2v_out.v:19508.13-19508.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:19521.13-19521.30" */
input data_ind_timing_i;
wire data_ind_timing_i;
/* cellift = 32'd1 */
input data_ind_timing_i_t0;
wire data_ind_timing_i_t0;
/* src = "generated/sv2v_out.v:19560.6-19560.19" */
reg div_by_zero_q;
/* src = "generated/sv2v_out.v:19557.7-19557.22" */
wire div_change_sign;
/* src = "generated/sv2v_out.v:19511.13-19511.21" */
input div_en_i;
wire div_en_i;
/* cellift = 32'd1 */
input div_en_i_t0;
wire div_en_i_t0;
/* src = "generated/sv2v_out.v:19513.13-19513.22" */
input div_sel_i;
wire div_sel_i;
/* cellift = 32'd1 */
input div_sel_i_t0;
wire div_sel_i_t0;
/* src = "generated/sv2v_out.v:19520.13-19520.28" */
input equal_to_zero_i;
wire equal_to_zero_i;
/* cellift = 32'd1 */
input equal_to_zero_i_t0;
wire equal_to_zero_i_t0;
/* src = "generated/sv2v_out.v:19525.21-19525.32" */
output [67:0] imd_val_d_o;
wire [67:0] imd_val_d_o;
/* cellift = 32'd1 */
output [67:0] imd_val_d_o_t0;
wire [67:0] imd_val_d_o_t0;
/* src = "generated/sv2v_out.v:19524.20-19524.31" */
input [67:0] imd_val_q_i;
wire [67:0] imd_val_q_i;
/* cellift = 32'd1 */
input [67:0] imd_val_q_i_t0;
wire [67:0] imd_val_q_i_t0;
/* src = "generated/sv2v_out.v:19526.20-19526.32" */
output [1:0] imd_val_we_o;
wire [1:0] imd_val_we_o;
/* cellift = 32'd1 */
output [1:0] imd_val_we_o_t0;
wire [1:0] imd_val_we_o_t0;
/* src = "generated/sv2v_out.v:19556.7-19556.23" */
wire is_greater_equal;
/* src = "generated/sv2v_out.v:19530.12-19530.22" */
reg [2:0] md_state_q;
/* src = "generated/sv2v_out.v:19510.13-19510.22" */
input mult_en_i;
wire mult_en_i;
/* cellift = 32'd1 */
input mult_en_i_t0;
wire mult_en_i_t0;
/* src = "generated/sv2v_out.v:19512.13-19512.23" */
input mult_sel_i;
wire mult_sel_i;
/* cellift = 32'd1 */
input mult_sel_i_t0;
wire mult_sel_i_t0;
/* src = "generated/sv2v_out.v:19538.12-19538.27" */
reg [4:0] multdiv_count_q;
/* src = "generated/sv2v_out.v:19562.7-19562.17" */
wire multdiv_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19562.7-19562.17" */
wire multdiv_en_t0;
/* src = "generated/sv2v_out.v:19561.6-19561.18" */
wire multdiv_hold;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19561.6-19561.18" */
wire multdiv_hold_t0;
/* src = "generated/sv2v_out.v:19527.13-19527.31" */
input multdiv_ready_id_i;
wire multdiv_ready_id_i;
/* cellift = 32'd1 */
input multdiv_ready_id_i_t0;
wire multdiv_ready_id_i_t0;
/* src = "generated/sv2v_out.v:19528.21-19528.37" */
output [31:0] multdiv_result_o;
wire [31:0] multdiv_result_o;
/* cellift = 32'd1 */
output [31:0] multdiv_result_o_t0;
wire [31:0] multdiv_result_o_t0;
/* src = "generated/sv2v_out.v:19552.14-19552.27" */
wire [32:0] next_quotient;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19552.14-19552.27" */
wire [32:0] next_quotient_t0;
/* src = "generated/sv2v_out.v:19553.14-19553.28" */
wire [31:0] next_remainder;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19553.14-19553.28" */
wire [31:0] next_remainder_t0;
/* src = "generated/sv2v_out.v:19546.14-19546.23" */
wire [32:0] one_shift;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19546.14-19546.23" */
wire [32:0] one_shift_t0;
/* src = "generated/sv2v_out.v:19548.14-19548.29" */
wire [32:0] op_a_bw_last_pp;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19548.14-19548.29" */
wire [32:0] op_a_bw_last_pp_t0;
/* src = "generated/sv2v_out.v:19547.14-19547.24" */
wire [32:0] op_a_bw_pp;
/* src = "generated/sv2v_out.v:19516.20-19516.26" */
input [31:0] op_a_i;
wire [31:0] op_a_i;
/* cellift = 32'd1 */
input [31:0] op_a_i_t0;
wire [31:0] op_a_i_t0;
/* src = "generated/sv2v_out.v:19542.13-19542.25" */
reg [32:0] op_a_shift_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19542.13-19542.25" */
reg [32:0] op_a_shift_q_t0;
/* src = "generated/sv2v_out.v:19517.20-19517.26" */
input [31:0] op_b_i;
wire [31:0] op_b_i;
/* cellift = 32'd1 */
input [31:0] op_b_i_t0;
wire [31:0] op_b_i_t0;
/* src = "generated/sv2v_out.v:19540.13-19540.25" */
reg [32:0] op_b_shift_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19540.13-19540.25" */
reg [32:0] op_b_shift_q_t0;
/* src = "generated/sv2v_out.v:19555.13-19555.27" */
wire [31:0] op_numerator_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19555.13-19555.27" */
wire [31:0] op_numerator_d_t0;
/* src = "generated/sv2v_out.v:19514.19-19514.29" */
input [1:0] operator_i;
wire [1:0] operator_i;
/* cellift = 32'd1 */
input [1:0] operator_i_t0;
wire [1:0] operator_i_t0;
/* src = "generated/sv2v_out.v:19558.7-19558.22" */
wire rem_change_sign;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19558.7-19558.22" */
wire rem_change_sign_t0;
/* src = "generated/sv2v_out.v:19509.13-19509.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:19551.7-19551.13" */
wire sign_b;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19551.7-19551.13" */
wire sign_b_t0;
/* src = "generated/sv2v_out.v:19515.19-19515.32" */
input [1:0] signed_mode_i;
wire [1:0] signed_mode_i;
/* cellift = 32'd1 */
input [1:0] signed_mode_i_t0;
wire [1:0] signed_mode_i_t0;
/* src = "generated/sv2v_out.v:19529.14-19529.21" */
output valid_o;
wire valid_o;
/* cellift = 32'd1 */
output valid_o_t0;
wire valid_o_t0;
assign op_a_bw_pp[31:0] = op_a_shift_q[31:0] & /* src = "generated/sv2v_out.v:19609.66-19609.90" */ { op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0] };
assign op_a_bw_last_pp[32] = op_a_shift_q[32] & /* src = "generated/sv2v_out.v:19609.28-19609.62" */ op_b_shift_q[0];
assign rem_change_sign = op_a_i[31] & /* src = "generated/sv2v_out.v:19610.18-19610.47" */ signed_mode_i[0];
assign sign_b = op_b_i[31] & /* src = "generated/sv2v_out.v:19611.18-19611.47" */ signed_mode_i[1];
assign div_change_sign = _304_ & /* src = "generated/sv2v_out.v:19618.27-19618.61" */ _272_;
assign _038_ = op_a_i & /* src = "generated/sv2v_out.v:19635.55-19635.88" */ { op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0] };
assign _042_ = op_a_i[31:1] & /* src = "generated/sv2v_out.v:19641.61-19641.94" */ { op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0] };
assign _040_ = rem_change_sign & /* src = "generated/sv2v_out.v:19641.34-19641.58" */ op_b_i[0];
assign multdiv_en = _277_ & /* src = "generated/sv2v_out.v:19733.22-19733.60" */ imd_val_we_o[0];
assign _044_ = _253_ & /* src = "generated/sv2v_out.v:19749.43-19749.111" */ _279_;
assign _045_ = ~ _089_;
assign _046_ = ~ _090_;
assign _120_ = { _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_ } & _013_;
assign _122_ = { _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_ } & _011_;
assign _121_ = { _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_ } & op_b_shift_q_t0;
assign _123_ = { _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_ } & op_a_shift_q_t0;
assign _213_ = _120_ | _121_;
assign _214_ = _122_ | _123_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME op_b_shift_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) op_b_shift_q_t0 <= 33'h000000000;
else op_b_shift_q_t0 <= _213_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME op_a_shift_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) op_a_shift_q_t0 <= 33'h000000000;
else op_a_shift_q_t0 <= _214_;
assign _096_ = op_a_shift_q_t0[31:0] & { op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0] };
assign _099_ = op_a_shift_q_t0[32] & op_b_shift_q[0];
assign _102_ = op_a_i_t0[31] & signed_mode_i[0];
assign _105_ = op_b_i_t0[31] & signed_mode_i[1];
assign _108_ = op_a_i_t0 & { op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0] };
assign _111_ = op_a_i_t0[31:1] & { op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0] };
assign _114_ = rem_change_sign_t0 & op_b_i[0];
assign _117_ = _278_ & imd_val_we_o[0];
assign _097_ = { op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0] } & op_a_shift_q[31:0];
assign _100_ = op_b_shift_q_t0[0] & op_a_shift_q[32];
assign _103_ = signed_mode_i_t0[0] & op_a_i[31];
assign _106_ = signed_mode_i_t0[1] & op_b_i[31];
assign _109_ = { op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0] } & op_a_i;
assign _112_ = { op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0] } & op_a_i[31:1];
assign _115_ = op_b_i_t0[0] & rem_change_sign;
assign _118_ = multdiv_hold_t0 & _277_;
assign _098_ = op_a_shift_q_t0[31:0] & { op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0] };
assign _101_ = op_a_shift_q_t0[32] & op_b_shift_q_t0[0];
assign _104_ = op_a_i_t0[31] & signed_mode_i_t0[0];
assign _107_ = op_b_i_t0[31] & signed_mode_i_t0[1];
assign _110_ = op_a_i_t0 & { op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0] };
assign _113_ = op_a_i_t0[31:1] & { op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0] };
assign _116_ = rem_change_sign_t0 & op_b_i_t0[0];
assign _119_ = _278_ & multdiv_hold_t0;
assign _205_ = _096_ | _097_;
assign _206_ = _099_ | _100_;
assign _207_ = _102_ | _103_;
assign _208_ = _105_ | _106_;
assign _209_ = _108_ | _109_;
assign _210_ = _111_ | _112_;
assign _211_ = _114_ | _115_;
assign _212_ = _117_ | _118_;
assign op_a_bw_last_pp_t0[31:0] = _205_ | _098_;
assign op_a_bw_last_pp_t0[32] = _206_ | _101_;
assign rem_change_sign_t0 = _207_ | _104_;
assign sign_b_t0 = _208_ | _107_;
assign _039_ = _209_ | _110_;
assign _043_ = _210_ | _113_;
assign _041_ = _211_ | _116_;
assign multdiv_en_t0 = _212_ | _119_;
/* src = "generated/sv2v_out.v:19734.2-19748.6" */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME md_state_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) md_state_q <= 3'h0;
else if (_087_) md_state_q <= _006_;
/* src = "generated/sv2v_out.v:19734.2-19748.6" */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME multdiv_count_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) multdiv_count_q <= 5'h00;
else if (_088_) multdiv_count_q <= _007_;
/* src = "generated/sv2v_out.v:19734.2-19748.6" */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME op_b_shift_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) op_b_shift_q <= 33'h000000000;
else if (_089_) op_b_shift_q <= _012_;
/* src = "generated/sv2v_out.v:19734.2-19748.6" */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME op_a_shift_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) op_a_shift_q <= 33'h000000000;
else if (_090_) op_a_shift_q <= _010_;
/* src = "generated/sv2v_out.v:19734.2-19748.6" */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME div_by_zero_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) div_by_zero_q <= 1'h0;
else if (_091_) div_by_zero_q <= _018_;
assign _047_ = ~ { _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_ };
assign _048_ = ~ { _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_ };
assign _049_ = ~ _077_;
assign _050_ = ~ { _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_ };
assign _051_ = ~ { _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_ };
assign _052_ = ~ { _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_ };
assign _053_ = ~ { _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_ };
assign _054_ = ~ { _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_ };
assign _055_ = ~ { _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_ };
assign _056_ = ~ { _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_ };
assign _057_ = ~ { _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_ };
assign _058_ = ~ { _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_ };
assign _059_ = ~ { _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_ };
assign _060_ = ~ _258_;
assign _061_ = ~ { _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_ };
assign _062_ = ~ { _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_ };
assign _063_ = ~ { _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_ };
assign _064_ = ~ { _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_ };
assign _065_ = ~ { _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_ };
assign _066_ = ~ { is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal };
assign _067_ = ~ { is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal };
assign _068_ = ~ { rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign };
assign _069_ = ~ { sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b };
assign _070_ = ~ { div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign };
assign _071_ = ~ { rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign };
assign _072_ = ~ { div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i };
assign _124_ = _047_ & imd_val_q_i_t0[66:34];
assign _126_ = _048_ & _218_;
assign _021_ = _049_ & multdiv_ready_id_i_t0;
assign _128_ = _047_ & alu_adder_ext_i_t0[32:0];
assign _130_ = _048_ & _220_;
assign _132_ = _050_ & { op_a_shift_q_t0[31:0], 1'h0 };
assign _134_ = _051_ & alu_adder_ext_i_t0[32:0];
assign _136_ = _050_ & _222_;
assign _138_ = _051_ & { _041_, _039_ };
assign _140_ = _052_ & _227_;
assign _142_ = _051_ & { op_a_i_t0, 1'h0 };
assign _229_ = _053_ & _023_;
assign _144_ = _054_ & _229_;
assign _146_ = _055_ & _025_;
assign _148_ = _054_ & _231_;
assign _150_ = _056_ & _027_;
assign _152_ = _057_ & _233_;
assign _154_ = _058_ & imd_val_q_i_t0[66:34];
assign _156_ = _055_ & _237_;
assign _158_ = _059_ & _239_;
assign _160_ = _060_ & _246_;
assign _162_ = _057_ & { op_b_i_t0, 1'h0 };
assign _164_ = _053_ & { op_b_shift_q_t0[31:0], 1'h0 };
assign _166_ = _061_ & _250_;
assign _168_ = _051_ & op_a_bw_last_pp_t0;
assign _170_ = _050_ & _252_;
assign _172_ = _050_ & imd_val_q_i_t0[66:34];
assign _180_ = _062_ & imd_val_q_i_t0[31:0];
assign _182_ = _063_ & imd_val_q_i_t0[31:0];
assign _184_ = _064_ & imd_val_q_i_t0[66:34];
assign _003_ = _065_ & { imd_val_q_i_t0[65:34], 1'h0 };
assign _186_ = _056_ & op_a_bw_last_pp_t0;
assign _188_ = _066_ & imd_val_q_i_t0[65:34];
assign _190_ = _067_ & op_a_shift_q_t0;
assign _192_ = _068_ & op_a_i_t0;
assign _194_ = _069_ & { 1'h0, op_b_i_t0 };
assign _196_ = _070_ & imd_val_q_i_t0[66:34];
assign _198_ = _071_ & imd_val_q_i_t0[66:34];
assign _200_ = _072_ & alu_adder_ext_i_t0[31:0];
assign _125_ = { _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_ } & _301_;
assign _127_ = { _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_ } & _303_;
assign _129_ = { _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_ } & next_quotient_t0;
assign _131_ = { _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_ } & { 1'h0, next_remainder_t0 };
assign _133_ = { _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_ } & next_quotient_t0;
assign _135_ = { _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_ } & alu_adder_ext_i_t0[33:1];
assign _137_ = { _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_ } & { next_remainder_t0, _288_ };
assign _225_ = { _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_ } & { rem_change_sign_t0, op_a_i_t0 };
assign _139_ = { _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_ } & { 1'h0, _041_, _043_ };
assign _141_ = { _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_ } & _225_;
assign _143_ = { _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_ } & { rem_change_sign_t0, op_a_i_t0 };
assign _145_ = { _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_ } & _030_;
assign _147_ = { _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_ } & _297_;
assign _149_ = { _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_ } & _032_;
assign _151_ = { _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_ } & _034_;
assign _153_ = { _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_ } & _037_;
assign _155_ = { _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_ } & _017_;
assign _157_ = { _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_ } & { 32'h00000000, imd_val_q_i_t0[31] };
assign _159_ = { _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_ } & _235_;
assign _246_ = _253_ & _021_;
assign _161_ = _258_ & multdiv_ready_id_i_t0;
assign _163_ = { _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_ } & { imd_val_q_i_t0[65:34], 1'h0 };
assign _165_ = { _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_ } & { op_a_i_t0, 1'h0 };
assign _167_ = { _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_ } & _248_;
assign _169_ = { _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_ } & _291_;
assign _171_ = { _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_ } & _005_;
assign _173_ = { _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_ } & _003_;
assign _032_ = { _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_ } & { 1'h0, op_b_shift_q_t0[32:1] };
assign _025_ = { _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_ } & { 1'h0, sign_b_t0, op_b_i_t0[31:1] };
assign _181_ = { _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_ } & _295_;
assign multdiv_hold_t0 = _265_ & _009_;
assign _183_ = { _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_ } & _015_;
assign _185_ = { _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_ } & _001_;
assign _187_ = { _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_ } & op_a_bw_last_pp_t0;
assign _189_ = { is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal } & alu_adder_ext_i_t0[32:1];
assign _191_ = { is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal } & _276_;
assign _193_ = { rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign } & alu_adder_i_t0;
assign _195_ = { sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b } & { 1'h0, alu_adder_i_t0 };
assign _197_ = { div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign } & { 1'h0, alu_adder_i_t0 };
assign _199_ = { rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign } & { 1'h0, alu_adder_i_t0 };
assign _201_ = { div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i } & imd_val_q_i_t0[65:34];
assign _218_ = _124_ | _125_;
assign _037_ = _126_ | _127_;
assign _220_ = _128_ | _129_;
assign _034_ = _130_ | _131_;
assign _030_ = _132_ | _133_;
assign _222_ = _134_ | _135_;
assign _027_ = _136_ | _137_;
assign _227_ = _138_ | _139_;
assign _017_ = _140_ | _141_;
assign _023_ = _142_ | _143_;
assign _011_ = _144_ | _145_;
assign _231_ = _146_ | _147_;
assign _013_ = _148_ | _149_;
assign _233_ = _150_ | _151_;
assign _235_ = _152_ | _153_;
assign _237_ = _154_ | _155_;
assign _239_ = _156_ | _157_;
assign _001_ = _158_ | _159_;
assign _009_ = _160_ | _161_;
assign _248_ = _162_ | _163_;
assign _250_ = _164_ | _165_;
assign _005_ = _166_ | _167_;
assign _252_ = _168_ | _169_;
assign alu_operand_b_o_t0 = _170_ | _171_;
assign alu_operand_a_o_t0 = _172_ | _173_;
assign _015_ = _180_ | _181_;
assign op_numerator_d_t0 = _182_ | _183_;
assign accum_window_d_t0 = _184_ | _185_;
assign _291_ = _186_ | _187_;
assign next_remainder_t0 = _188_ | _189_;
assign next_quotient_t0 = _190_ | _191_;
assign _295_ = _192_ | _193_;
assign _297_ = _194_ | _195_;
assign _301_ = _196_ | _197_;
assign _303_ = _198_ | _199_;
assign multdiv_result_o_t0 = _200_ | _201_;
assign _080_ = | { _284_, _283_ };
assign _081_ = { _283_, _077_ } != 2'h3;
assign _082_ = { _284_, _077_ } != 2'h3;
assign _083_ = | { _286_, _284_, _283_ };
assign _084_ = { _283_, _260_ } != 2'h3;
assign _085_ = | { _285_, _284_, _283_ };
assign _086_ = ~ _092_;
assign _087_ = & { _265_, multdiv_en };
assign _088_ = & { _080_, _265_, multdiv_en };
assign _089_ = & { _265_, multdiv_en, _081_, _082_, _083_ };
assign _090_ = & { _265_, multdiv_en, _082_, _084_, _085_ };
assign _091_ = & { _284_, _265_, multdiv_en, _086_ };
assign _092_ = | { _280_, _260_, _259_ };
assign _094_ = | { _286_, _284_ };
assign _093_ = | { _260_, _259_ };
assign _095_ = | { _281_, _280_, _260_ };
assign _073_ = ~ op_a_shift_q;
assign _074_ = ~ mult_en_i;
assign _075_ = ~ one_shift;
assign _076_ = ~ div_en_i;
assign _174_ = op_a_shift_q_t0 & _075_;
assign _177_ = mult_en_i_t0 & _076_;
assign _175_ = one_shift_t0 & _073_;
assign _178_ = div_en_i_t0 & _074_;
assign _176_ = op_a_shift_q_t0 & one_shift_t0;
assign _179_ = mult_en_i_t0 & div_en_i_t0;
assign _215_ = _174_ | _175_;
assign _216_ = _177_ | _178_;
assign _276_ = _215_ | _176_;
assign _278_ = _216_ | _179_;
assign _077_ = | { _281_, _280_ };
assign _078_ = | { _286_, _285_, _284_, _282_ };
assign _202_ = _281_ | _280_;
assign _203_ = _285_ | _286_;
assign _204_ = _094_ | _282_;
assign _079_ = | { _283_, _282_, _253_ };
assign _217_ = _281_ ? _300_ : imd_val_q_i[66:34];
assign _036_ = _280_ ? _302_ : _217_;
assign _020_ = _077_ ? 1'h0 : _274_;
assign _035_ = _077_ ? 3'h5 : 3'h0;
assign _219_ = _281_ ? next_quotient : alu_adder_ext_i[32:0];
assign _033_ = _280_ ? { 1'h0, next_remainder } : _219_;
assign _028_ = _095_ ? _299_ : _298_;
assign _029_ = _077_ ? next_quotient : { op_a_shift_q[31:0], 1'h0 };
assign _221_ = _260_ ? alu_adder_ext_i[33:1] : alu_adder_ext_i[32:0];
assign _026_ = _077_ ? { next_remainder, _287_ } : _221_;
assign _223_ = _260_ ? 3'h3 : _292_;
assign _019_ = _077_ ? _293_ : _223_;
assign _224_ = _280_ ? { rem_change_sign, op_a_i } : 33'h1ffffffff;
assign _226_ = _260_ ? { 1'h1, _273_, _042_ } : { _273_, _038_ };
assign _016_ = _202_ ? _224_ : _226_;
assign _022_ = _260_ ? { rem_change_sign, op_a_i } : { op_a_i, 1'h0 };
assign _007_ = _283_ ? _289_ : 5'h1f;
assign _228_ = _285_ ? 33'h000000000 : _022_;
assign _010_ = _283_ ? _029_ : _228_;
assign _230_ = _286_ ? _296_ : _024_;
assign _012_ = _283_ ? _031_ : _230_;
assign _232_ = _253_ ? _033_ : _026_;
assign _234_ = _282_ ? _036_ : _232_;
assign _236_ = _284_ ? _016_ : imd_val_q_i[66:34];
assign _238_ = _286_ ? { 32'h00000000, imd_val_q_i[31] } : _236_;
assign _000_ = _079_ ? _234_ : _238_;
assign _240_ = _253_ ? _035_ : _028_;
assign _241_ = _282_ ? 3'h6 : _240_;
assign _242_ = _286_ ? 3'h3 : 3'h2;
assign _243_ = _284_ ? _019_ : 3'h0;
assign _244_ = _203_ ? _242_ : _243_;
assign _006_ = _079_ ? _241_ : _244_;
assign _245_ = _253_ ? _020_ : 1'h0;
assign _008_ = _258_ ? _274_ : _245_;
assign _247_ = _282_ ? { _269_, 1'h1 } : { _267_, 1'h1 };
assign _249_ = _285_ ? { _268_, 1'h1 } : { _270_, 1'h1 };
assign _004_ = _204_ ? _247_ : _249_;
assign _251_ = _260_ ? _290_ : op_a_bw_pp;
assign alu_operand_b_o = _077_ ? _004_ : _251_;
assign alu_operand_a_o = _077_ ? _002_ : imd_val_q_i[66:34];
assign _288_ = imd_val_q_i_t0[31:0] >> _289_;
assign one_shift_t0 = 33'h000000000 << multdiv_count_q;
assign _254_ = imd_val_q_i[65] == /* src = "generated/sv2v_out.v:19614.29-19614.67" */ op_b_shift_q[31];
assign _255_ = ! /* src = "generated/sv2v_out.v:19637.45-19637.65" */ { 1'h0, sign_b, op_b_i[31:1] };
assign _256_ = ! /* src = "generated/sv2v_out.v:19676.46-19676.63" */ { 1'h0, op_b_shift_q[32:1] };
assign _257_ = multdiv_count_q == /* src = "generated/sv2v_out.v:19687.22-19687.45" */ 5'h01;
assign _261_ = _264_ && /* src = "generated/sv2v_out.v:19637.22-19637.66" */ _255_;
assign _262_ = _264_ && /* src = "generated/sv2v_out.v:19652.22-19652.59" */ equal_to_zero_i;
assign _263_ = _264_ && /* src = "generated/sv2v_out.v:19676.23-19676.64" */ _256_;
assign _264_ = ! /* src = "generated/sv2v_out.v:19676.23-19676.41" */ data_ind_timing_i;
assign _265_ = mult_sel_i || /* src = "generated/sv2v_out.v:19629.7-19629.30" */ div_sel_i;
assign _266_ = _263_ || /* src = "generated/sv2v_out.v:19676.22-19676.94" */ _257_;
assign _268_ = ~ /* src = "generated/sv2v_out.v:19586.26-19586.33" */ op_a_i;
assign _267_ = ~ /* src = "generated/sv2v_out.v:19590.26-19590.33" */ op_b_i;
assign _269_ = ~ /* src = "generated/sv2v_out.v:19594.26-19594.47" */ imd_val_q_i[65:34];
assign _270_ = ~ /* src = "generated/sv2v_out.v:19603.24-19603.43" */ op_b_shift_q[31:0];
assign op_a_bw_pp[32] = ~ /* src = "generated/sv2v_out.v:19608.23-19608.60" */ op_a_bw_last_pp[32];
assign op_a_bw_last_pp[31:0] = ~ /* src = "generated/sv2v_out.v:19609.64-19609.91" */ op_a_bw_pp[31:0];
assign _271_ = ~ /* src = "generated/sv2v_out.v:19614.70-19614.86" */ alu_adder_ext_i[32];
assign _272_ = ~ /* src = "generated/sv2v_out.v:19618.47-19618.61" */ div_by_zero_q;
assign _273_ = ~ /* src = "generated/sv2v_out.v:19641.32-19641.59" */ _040_;
assign _274_ = ~ /* src = "generated/sv2v_out.v:19728.21-19728.40" */ multdiv_ready_id_i;
assign imd_val_we_o[0] = ~ /* src = "generated/sv2v_out.v:19733.47-19733.60" */ multdiv_hold;
assign _275_ = op_a_shift_q | /* src = "generated/sv2v_out.v:19617.45-19617.69" */ one_shift;
assign _277_ = mult_en_i | /* src = "generated/sv2v_out.v:19733.23-19733.43" */ div_en_i;
assign _279_ = _259_ | /* src = "generated/sv2v_out.v:19749.67-19749.110" */ _260_;
assign valid_o = _258_ | /* src = "generated/sv2v_out.v:19749.19-19749.112" */ _044_;
assign _031_ = _093_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19671.6-19691.13" */ { 1'h0, op_b_shift_q[32:1] } : 33'hxxxxxxxxx;
assign _024_ = _093_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19632.6-19656.13" */ { 1'h0, sign_b, op_b_i[31:1] } : 33'hxxxxxxxxx;
assign _018_ = _281_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19632.6-19656.13" */ equal_to_zero_i : 1'hx;
assign _283_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19630.4-19731.11" */ 3'h3;
assign _258_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19630.4-19731.11" */ 3'h6;
assign _253_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19630.4-19731.11" */ 3'h4;
assign _014_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19630.4-19731.11" */ _294_ : imd_val_q_i[31:0];
assign multdiv_hold = _265_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:19629.7-19629.30|generated/sv2v_out.v:19629.3-19731.11" */ _008_ : 1'h0;
assign op_numerator_d = _265_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:19629.7-19629.30|generated/sv2v_out.v:19629.3-19731.11" */ _014_ : imd_val_q_i[31:0];
assign accum_window_d = _265_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:19629.7-19629.30|generated/sv2v_out.v:19629.3-19731.11" */ _000_ : imd_val_q_i[66:34];
assign _002_ = _078_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19579.5-19600.12" */ 33'h000000001 : { imd_val_q_i[65:34], 1'h1 };
assign _282_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19579.5-19600.12" */ 3'h5;
assign _286_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19579.5-19600.12" */ 3'h2;
assign _285_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19579.5-19600.12" */ 3'h1;
assign _284_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19579.5-19600.12" */ md_state_q;
assign _260_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19575.3-19605.10" */ 2'h1;
assign _259_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19575.3-19605.10" */ operator_i;
assign _281_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19575.3-19605.10" */ 2'h2;
assign _280_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19575.3-19605.10" */ 2'h3;
wire [31:0] _651_ = imd_val_q_i[31:0];
assign _287_ = _651_[_289_ +: 1];
assign one_shift = 33'h000000001 << /* src = "generated/sv2v_out.v:19615.21-19615.77" */ multdiv_count_q;
assign _289_ = multdiv_count_q - /* src = "generated/sv2v_out.v:19670.24-19670.47" */ 5'h01;
assign _290_ = _253_ ? /* src = "generated/sv2v_out.v:19577.29-19577.78" */ op_a_bw_last_pp : op_a_bw_pp;
assign is_greater_equal = _254_ ? /* src = "generated/sv2v_out.v:19614.29-19614.107" */ _271_ : imd_val_q_i[65];
assign next_remainder = is_greater_equal ? /* src = "generated/sv2v_out.v:19616.27-19616.86" */ alu_adder_ext_i[32:1] : imd_val_q_i[65:34];
assign next_quotient = is_greater_equal ? /* src = "generated/sv2v_out.v:19617.26-19617.84" */ _275_ : op_a_shift_q;
assign _292_ = _261_ ? /* src = "generated/sv2v_out.v:19637.22-19637.80" */ 3'h4 : 3'h3;
assign _293_ = _262_ ? /* src = "generated/sv2v_out.v:19652.22-19652.73" */ 3'h6 : 3'h1;
assign _294_ = rem_change_sign ? /* src = "generated/sv2v_out.v:19661.24-19661.53" */ alu_adder_i : op_a_i;
assign _296_ = sign_b ? /* src = "generated/sv2v_out.v:19666.22-19666.67" */ { 1'h0, alu_adder_i } : { 1'h0, op_b_i };
assign _298_ = _266_ ? /* src = "generated/sv2v_out.v:19676.22-19676.108" */ 3'h4 : 3'h3;
assign _299_ = _257_ ? /* src = "generated/sv2v_out.v:19687.22-19687.59" */ 3'h4 : 3'h3;
assign _300_ = div_change_sign ? /* src = "generated/sv2v_out.v:19720.31-19720.85" */ { 1'h0, alu_adder_i } : imd_val_q_i[66:34];
assign _302_ = rem_change_sign ? /* src = "generated/sv2v_out.v:19721.31-19721.85" */ { 1'h0, alu_adder_i } : imd_val_q_i[66:34];
assign multdiv_result_o = div_en_i ? /* src = "generated/sv2v_out.v:19750.29-19750.80" */ imd_val_q_i[65:34] : alu_adder_ext_i[31:0];
assign _304_ = rem_change_sign ^ /* src = "generated/sv2v_out.v:19618.28-19618.43" */ sign_b;
assign imd_val_d_o = { 1'h0, accum_window_d, 2'h0, op_numerator_d };
assign imd_val_d_o_t0 = { 1'h0, accum_window_d_t0, 2'h0, op_numerator_d_t0 };
assign imd_val_we_o[1] = multdiv_en;
assign imd_val_we_o_t0 = { multdiv_en_t0, multdiv_hold_t0 };
assign valid_o_t0 = 1'h0;
endmodule

module ibex_top(clk_i, rst_ni, test_en_i, ram_cfg_i, hart_id_i, boot_addr_i, instr_req_o, instr_gnt_i, instr_rvalid_i, instr_addr_o, instr_rdata_i, instr_rdata_intg_i, instr_err_i, data_req_o, data_gnt_i, data_rvalid_i, data_we_o, data_be_o, data_addr_o, data_wdata_o, data_wdata_intg_o
, data_rdata_i, data_rdata_intg_i, data_err_i, irq_software_i, irq_timer_i, irq_external_i, irq_fast_i, irq_nm_i, scramble_key_valid_i, scramble_key_i, scramble_nonce_i, scramble_req_o, debug_req_i, crash_dump_o, double_fault_seen_o, fetch_enable_i, alert_minor_o, alert_major_internal_o, alert_major_bus_o, core_sleep_o, scan_rst_ni
, instr_rvalid_i_t0, instr_req_o_t0, instr_rdata_i_t0, instr_gnt_i_t0, instr_err_i_t0, instr_addr_o_t0, data_we_o_t0, data_req_o_t0, debug_req_i_t0, data_rdata_i_t0, data_gnt_i_t0, data_be_o_t0, data_addr_o_t0, data_rvalid_i_t0, data_wdata_o_t0, irq_nm_i_t0, boot_addr_i_t0, test_en_i_t0, double_fault_seen_o_t0, hart_id_i_t0, irq_external_i_t0
, irq_fast_i_t0, irq_software_i_t0, irq_timer_i_t0, alert_major_bus_o_t0, alert_major_internal_o_t0, alert_minor_o_t0, crash_dump_o_t0, data_err_i_t0, fetch_enable_i_t0, core_sleep_o_t0, data_rdata_intg_i_t0, data_wdata_intg_o_t0, instr_rdata_intg_i_t0, ram_cfg_i_t0, scan_rst_ni_t0, scramble_key_i_t0, scramble_key_valid_i_t0, scramble_nonce_i_t0, scramble_req_o_t0);
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
/* src = "generated/sv2v_out.v:20366.25-20366.60" */
wire _19_;
/* src = "generated/sv2v_out.v:20366.24-20366.75" */
wire _20_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20366.24-20366.75" */
wire _21_;
/* src = "generated/sv2v_out.v:20366.23-20366.90" */
wire _22_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20366.23-20366.90" */
wire _23_;
/* src = "generated/sv2v_out.v:20281.14-20281.31" */
output alert_major_bus_o;
wire alert_major_bus_o;
/* cellift = 32'd1 */
output alert_major_bus_o_t0;
wire alert_major_bus_o_t0;
/* src = "generated/sv2v_out.v:20280.14-20280.36" */
output alert_major_internal_o;
wire alert_major_internal_o;
/* cellift = 32'd1 */
output alert_major_internal_o_t0;
wire alert_major_internal_o_t0;
/* src = "generated/sv2v_out.v:20279.14-20279.27" */
output alert_minor_o;
wire alert_minor_o;
/* cellift = 32'd1 */
output alert_minor_o_t0;
wire alert_minor_o_t0;
/* src = "generated/sv2v_out.v:20247.20-20247.31" */
input [31:0] boot_addr_i;
wire [31:0] boot_addr_i;
/* cellift = 32'd1 */
input [31:0] boot_addr_i_t0;
wire [31:0] boot_addr_i_t0;
/* src = "generated/sv2v_out.v:20309.7-20309.10" */
wire clk;
/* src = "generated/sv2v_out.v:20242.13-20242.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:20312.7-20312.15" */
wire clock_en;
/* src = "generated/sv2v_out.v:20339.7-20339.32" */
wire core_alert_major_internal;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20339.7-20339.32" */
wire core_alert_major_internal_t0;
/* src = "generated/sv2v_out.v:20310.13-20310.24" */
wire [3:0] core_busy_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20310.13-20310.24" */
wire [3:0] core_busy_d_t0;
/* src = "generated/sv2v_out.v:20311.12-20311.23" */
wire [3:0] core_busy_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20311.12-20311.23" */
/* unused_bits = "0 1 2 3" */
wire [3:0] core_busy_q_t0;
/* src = "generated/sv2v_out.v:20282.14-20282.26" */
output core_sleep_o;
wire core_sleep_o;
/* cellift = 32'd1 */
output core_sleep_o_t0;
wire core_sleep_o_t0;
/* src = "generated/sv2v_out.v:20276.22-20276.34" */
output [159:0] crash_dump_o;
wire [159:0] crash_dump_o;
/* cellift = 32'd1 */
output [159:0] crash_dump_o_t0;
wire [159:0] crash_dump_o_t0;
/* src = "generated/sv2v_out.v:20260.21-20260.32" */
output [31:0] data_addr_o;
wire [31:0] data_addr_o;
/* cellift = 32'd1 */
output [31:0] data_addr_o_t0;
wire [31:0] data_addr_o_t0;
/* src = "generated/sv2v_out.v:20259.20-20259.29" */
output [3:0] data_be_o;
wire [3:0] data_be_o;
/* cellift = 32'd1 */
output [3:0] data_be_o_t0;
wire [3:0] data_be_o_t0;
/* src = "generated/sv2v_out.v:20265.13-20265.23" */
input data_err_i;
wire data_err_i;
/* cellift = 32'd1 */
input data_err_i_t0;
wire data_err_i_t0;
/* src = "generated/sv2v_out.v:20256.13-20256.23" */
input data_gnt_i;
wire data_gnt_i;
/* cellift = 32'd1 */
input data_gnt_i_t0;
wire data_gnt_i_t0;
/* src = "generated/sv2v_out.v:20263.20-20263.32" */
input [31:0] data_rdata_i;
wire [31:0] data_rdata_i;
/* cellift = 32'd1 */
input [31:0] data_rdata_i_t0;
wire [31:0] data_rdata_i_t0;
/* src = "generated/sv2v_out.v:20264.19-20264.36" */
input [6:0] data_rdata_intg_i;
wire [6:0] data_rdata_intg_i;
/* cellift = 32'd1 */
input [6:0] data_rdata_intg_i_t0;
wire [6:0] data_rdata_intg_i_t0;
/* src = "generated/sv2v_out.v:20255.14-20255.24" */
output data_req_o;
wire data_req_o;
/* cellift = 32'd1 */
output data_req_o_t0;
wire data_req_o_t0;
/* src = "generated/sv2v_out.v:20257.13-20257.26" */
input data_rvalid_i;
wire data_rvalid_i;
/* cellift = 32'd1 */
input data_rvalid_i_t0;
wire data_rvalid_i_t0;
/* src = "generated/sv2v_out.v:20325.28-20325.43" */
wire [38:0] data_wdata_core;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20325.28-20325.43" */
wire [38:0] data_wdata_core_t0;
/* src = "generated/sv2v_out.v:20262.20-20262.37" */
output [6:0] data_wdata_intg_o;
wire [6:0] data_wdata_intg_o;
/* cellift = 32'd1 */
output [6:0] data_wdata_intg_o_t0;
wire [6:0] data_wdata_intg_o_t0;
/* src = "generated/sv2v_out.v:20261.21-20261.33" */
output [31:0] data_wdata_o;
wire [31:0] data_wdata_o;
/* cellift = 32'd1 */
output [31:0] data_wdata_o_t0;
wire [31:0] data_wdata_o_t0;
/* src = "generated/sv2v_out.v:20258.14-20258.23" */
output data_we_o;
wire data_we_o;
/* cellift = 32'd1 */
output data_we_o_t0;
wire data_we_o_t0;
/* src = "generated/sv2v_out.v:20275.13-20275.24" */
input debug_req_i;
wire debug_req_i;
/* cellift = 32'd1 */
input debug_req_i_t0;
wire debug_req_i_t0;
/* src = "generated/sv2v_out.v:20277.14-20277.33" */
output double_fault_seen_o;
wire double_fault_seen_o;
/* cellift = 32'd1 */
output double_fault_seen_o_t0;
wire double_fault_seen_o_t0;
/* src = "generated/sv2v_out.v:20314.7-20314.21" */
wire dummy_instr_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20314.7-20314.21" */
wire dummy_instr_id_t0;
/* src = "generated/sv2v_out.v:20315.7-20315.21" */
wire dummy_instr_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20315.7-20315.21" */
wire dummy_instr_wb_t0;
/* src = "generated/sv2v_out.v:20351.13-20351.29" */
wire [3:0] fetch_enable_buf;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20351.13-20351.29" */
wire [3:0] fetch_enable_buf_t0;
/* src = "generated/sv2v_out.v:20278.19-20278.33" */
input [3:0] fetch_enable_i;
wire [3:0] fetch_enable_i;
/* cellift = 32'd1 */
input [3:0] fetch_enable_i_t0;
wire [3:0] fetch_enable_i_t0;
/* src = "generated/sv2v_out.v:20246.20-20246.29" */
input [31:0] hart_id_i;
wire [31:0] hart_id_i;
/* cellift = 32'd1 */
input [31:0] hart_id_i_t0;
wire [31:0] hart_id_i_t0;
/* src = "generated/sv2v_out.v:20335.35-20335.47" */
/* unused_bits = "0 1 2 3 4 5 6 7" */
wire [7:0] ic_data_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20335.35-20335.47" */
/* unused_bits = "0 1 2 3 4 5 6 7" */
wire [7:0] ic_data_addr_t0;
/* src = "generated/sv2v_out.v:20333.13-20333.24" */
/* unused_bits = "0 1" */
wire [1:0] ic_data_req;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20333.13-20333.24" */
/* unused_bits = "0 1" */
wire [1:0] ic_data_req_t0;
/* src = "generated/sv2v_out.v:20336.27-20336.40" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63" */
wire [63:0] ic_data_wdata;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20336.27-20336.40" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63" */
wire [63:0] ic_data_wdata_t0;
/* src = "generated/sv2v_out.v:20334.7-20334.20" */
/* unused_bits = "0" */
wire ic_data_write;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20334.7-20334.20" */
/* unused_bits = "0" */
wire ic_data_write_t0;
/* src = "generated/sv2v_out.v:20338.7-20338.21" */
/* unused_bits = "0" */
wire ic_scr_key_req;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20338.7-20338.21" */
/* unused_bits = "0" */
wire ic_scr_key_req_t0;
/* src = "generated/sv2v_out.v:20330.35-20330.46" */
/* unused_bits = "0 1 2 3 4 5 6 7" */
wire [7:0] ic_tag_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20330.35-20330.46" */
/* unused_bits = "0 1 2 3 4 5 6 7" */
wire [7:0] ic_tag_addr_t0;
/* src = "generated/sv2v_out.v:20328.13-20328.23" */
/* unused_bits = "0 1" */
wire [1:0] ic_tag_req;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20328.13-20328.23" */
/* unused_bits = "0 1" */
wire [1:0] ic_tag_req_t0;
/* src = "generated/sv2v_out.v:20331.26-20331.38" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21" */
wire [21:0] ic_tag_wdata;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20331.26-20331.38" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21" */
wire [21:0] ic_tag_wdata_t0;
/* src = "generated/sv2v_out.v:20329.7-20329.19" */
/* unused_bits = "0" */
wire ic_tag_write;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20329.7-20329.19" */
/* unused_bits = "0" */
wire ic_tag_write_t0;
/* src = "generated/sv2v_out.v:20251.21-20251.33" */
output [31:0] instr_addr_o;
wire [31:0] instr_addr_o;
/* cellift = 32'd1 */
output [31:0] instr_addr_o_t0;
wire [31:0] instr_addr_o_t0;
/* src = "generated/sv2v_out.v:20254.13-20254.24" */
input instr_err_i;
wire instr_err_i;
/* cellift = 32'd1 */
input instr_err_i_t0;
wire instr_err_i_t0;
/* src = "generated/sv2v_out.v:20249.13-20249.24" */
input instr_gnt_i;
wire instr_gnt_i;
/* cellift = 32'd1 */
input instr_gnt_i_t0;
wire instr_gnt_i_t0;
/* src = "generated/sv2v_out.v:20252.20-20252.33" */
input [31:0] instr_rdata_i;
wire [31:0] instr_rdata_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_i_t0;
wire [31:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:20253.19-20253.37" */
input [6:0] instr_rdata_intg_i;
wire [6:0] instr_rdata_intg_i;
/* cellift = 32'd1 */
input [6:0] instr_rdata_intg_i_t0;
wire [6:0] instr_rdata_intg_i_t0;
/* src = "generated/sv2v_out.v:20248.14-20248.25" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:20250.13-20250.27" */
input instr_rvalid_i;
wire instr_rvalid_i;
/* cellift = 32'd1 */
input instr_rvalid_i_t0;
wire instr_rvalid_i_t0;
/* src = "generated/sv2v_out.v:20268.13-20268.27" */
input irq_external_i;
wire irq_external_i;
/* cellift = 32'd1 */
input irq_external_i_t0;
wire irq_external_i_t0;
/* src = "generated/sv2v_out.v:20269.20-20269.30" */
input [14:0] irq_fast_i;
wire [14:0] irq_fast_i;
/* cellift = 32'd1 */
input [14:0] irq_fast_i_t0;
wire [14:0] irq_fast_i_t0;
/* src = "generated/sv2v_out.v:20270.13-20270.21" */
input irq_nm_i;
wire irq_nm_i;
/* cellift = 32'd1 */
input irq_nm_i_t0;
wire irq_nm_i_t0;
/* src = "generated/sv2v_out.v:20313.7-20313.18" */
wire irq_pending;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20313.7-20313.18" */
wire irq_pending_t0;
/* src = "generated/sv2v_out.v:20266.13-20266.27" */
input irq_software_i;
wire irq_software_i;
/* cellift = 32'd1 */
input irq_software_i_t0;
wire irq_software_i_t0;
/* src = "generated/sv2v_out.v:20267.13-20267.24" */
input irq_timer_i;
wire irq_timer_i;
/* cellift = 32'd1 */
input irq_timer_i_t0;
wire irq_timer_i_t0;
/* src = "generated/sv2v_out.v:20245.19-20245.28" */
input [9:0] ram_cfg_i;
wire [9:0] ram_cfg_i;
/* cellift = 32'd1 */
input [9:0] ram_cfg_i_t0;
wire [9:0] ram_cfg_i_t0;
/* src = "generated/sv2v_out.v:20496.7-20496.30" */
wire rf_alert_major_internal;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20496.7-20496.30" */
wire rf_alert_major_internal_t0;
/* src = "generated/sv2v_out.v:20316.13-20316.23" */
wire [4:0] rf_raddr_a;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20316.13-20316.23" */
wire [4:0] rf_raddr_a_t0;
/* src = "generated/sv2v_out.v:20317.13-20317.23" */
wire [4:0] rf_raddr_b;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20317.13-20317.23" */
wire [4:0] rf_raddr_b_t0;
/* src = "generated/sv2v_out.v:20321.32-20321.46" */
wire [38:0] rf_rdata_a_ecc;
/* src = "generated/sv2v_out.v:20322.32-20322.50" */
wire [38:0] rf_rdata_a_ecc_buf;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20322.32-20322.50" */
wire [38:0] rf_rdata_a_ecc_buf_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20321.32-20321.46" */
wire [38:0] rf_rdata_a_ecc_t0;
/* src = "generated/sv2v_out.v:20323.32-20323.46" */
wire [38:0] rf_rdata_b_ecc;
/* src = "generated/sv2v_out.v:20324.32-20324.50" */
wire [38:0] rf_rdata_b_ecc_buf;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20324.32-20324.50" */
wire [38:0] rf_rdata_b_ecc_buf_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20323.32-20323.46" */
wire [38:0] rf_rdata_b_ecc_t0;
/* src = "generated/sv2v_out.v:20318.13-20318.24" */
wire [4:0] rf_waddr_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20318.13-20318.24" */
wire [4:0] rf_waddr_wb_t0;
/* src = "generated/sv2v_out.v:20320.32-20320.47" */
wire [38:0] rf_wdata_wb_ecc;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20320.32-20320.47" */
wire [38:0] rf_wdata_wb_ecc_t0;
/* src = "generated/sv2v_out.v:20319.7-20319.15" */
wire rf_we_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20319.7-20319.15" */
wire rf_we_wb_t0;
/* src = "generated/sv2v_out.v:20243.13-20243.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:20283.13-20283.24" */
input scan_rst_ni;
wire scan_rst_ni;
/* cellift = 32'd1 */
input scan_rst_ni_t0;
wire scan_rst_ni_t0;
/* src = "generated/sv2v_out.v:20272.21-20272.35" */
input [127:0] scramble_key_i;
wire [127:0] scramble_key_i;
/* cellift = 32'd1 */
input [127:0] scramble_key_i_t0;
wire [127:0] scramble_key_i_t0;
/* src = "generated/sv2v_out.v:20271.13-20271.33" */
input scramble_key_valid_i;
wire scramble_key_valid_i;
/* cellift = 32'd1 */
input scramble_key_valid_i_t0;
wire scramble_key_valid_i_t0;
/* src = "generated/sv2v_out.v:20273.20-20273.36" */
input [63:0] scramble_nonce_i;
wire [63:0] scramble_nonce_i;
/* cellift = 32'd1 */
input [63:0] scramble_nonce_i_t0;
wire [63:0] scramble_nonce_i_t0;
/* src = "generated/sv2v_out.v:20274.14-20274.28" */
output scramble_req_o;
wire scramble_req_o;
/* cellift = 32'd1 */
output scramble_req_o_t0;
wire scramble_req_o_t0;
/* src = "generated/sv2v_out.v:20244.13-20244.22" */
input test_en_i;
wire test_en_i;
/* cellift = 32'd1 */
input test_en_i_t0;
wire test_en_i_t0;
assign _00_ = ~ _19_;
assign _01_ = ~ _20_;
assign _02_ = ~ _22_;
assign _03_ = ~ core_alert_major_internal;
assign _04_ = ~ irq_pending;
assign _05_ = ~ irq_nm_i;
assign _06_ = ~ rf_alert_major_internal;
assign _07_ = _21_ & _04_;
assign _10_ = _23_ & _05_;
assign _13_ = core_alert_major_internal_t0 & _06_;
assign _21_ = debug_req_i_t0 & _00_;
assign _08_ = irq_pending_t0 & _01_;
assign _11_ = irq_nm_i_t0 & _02_;
assign _14_ = rf_alert_major_internal_t0 & _03_;
assign _09_ = _21_ & irq_pending_t0;
assign _12_ = _23_ & irq_nm_i_t0;
assign _15_ = core_alert_major_internal_t0 & rf_alert_major_internal_t0;
assign _16_ = _07_ | _08_;
assign _17_ = _10_ | _11_;
assign _18_ = _13_ | _14_;
assign _23_ = _16_ | _09_;
assign core_sleep_o_t0 = _17_ | _12_;
assign alert_major_internal_o_t0 = _18_ | _15_;
assign _19_ = core_busy_q != /* src = "generated/sv2v_out.v:20366.25-20366.60" */ 4'ha;
assign core_sleep_o = ~ /* src = "generated/sv2v_out.v:20379.24-20379.33" */ clock_en;
assign _20_ = _19_ | /* src = "generated/sv2v_out.v:20366.24-20366.75" */ debug_req_i;
assign _22_ = _20_ | /* src = "generated/sv2v_out.v:20366.23-20366.90" */ irq_pending;
assign clock_en = _22_ | /* src = "generated/sv2v_out.v:20366.22-20366.102" */ irq_nm_i;
assign alert_major_internal_o = core_alert_major_internal | /* src = "generated/sv2v_out.v:20908.34-20908.119" */ rf_alert_major_internal;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20380.20-20385.3" */
prim_clock_gating core_clock_gate_i (
.clk_i(clk_i),
.clk_o(clk),
.en_i(clock_en),
.en_i_t0(core_sleep_o_t0),
.test_en_i(test_en_i),
.test_en_i_t0(test_en_i_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20360.6-20365.5" */
\$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_flop  \g_clock_en_secure.u_prim_core_busy_flop  (
.clk_i(clk_i),
.d_i(core_busy_d),
.d_i_t0(core_busy_d_t0),
.q_o(core_busy_q),
.q_o_t0(core_busy_q_t0),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20719.26-20722.5" */
\$paramod\prim_buf\Width=s32'00000000000000000000000000000111  \gen_mem_wdata_ecc.u_prim_buf_data_wdata_intg  (
.in_i(data_wdata_core[38:32]),
.in_i_t0(data_wdata_core_t0[38:32]),
.out_o(data_wdata_intg_o),
.out_o_t0(data_wdata_intg_o_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20510.6-20524.5" */
\$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  \gen_regfile_ff.register_file_i  (
.clk_i(clk),
.dummy_instr_id_i(dummy_instr_id),
.dummy_instr_id_i_t0(dummy_instr_id_t0),
.dummy_instr_wb_i(dummy_instr_wb),
.dummy_instr_wb_i_t0(dummy_instr_wb_t0),
.err_o(rf_alert_major_internal),
.err_o_t0(rf_alert_major_internal_t0),
.raddr_a_i(rf_raddr_a),
.raddr_a_i_t0(rf_raddr_a_t0),
.raddr_b_i(rf_raddr_b),
.raddr_b_i_t0(rf_raddr_b_t0),
.rdata_a_o(rf_rdata_a_ecc),
.rdata_a_o_t0(rf_rdata_a_ecc_t0),
.rdata_b_o(rf_rdata_b_ecc),
.rdata_b_o_t0(rf_rdata_b_ecc_t0),
.rst_ni(rst_ni),
.test_en_i(test_en_i),
.test_en_i_t0(test_en_i_t0),
.waddr_a_i(rf_waddr_wb),
.waddr_a_i_t0(rf_waddr_wb_t0),
.wdata_a_i(rf_wdata_wb_ecc),
.wdata_a_i_t0(rf_wdata_wb_ecc_t0),
.we_a_i(rf_we_wb),
.we_a_i_t0(rf_we_wb_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20386.24-20389.3" */
\$paramod\prim_buf\Width=s32'00000000000000000000000000000100  u_fetch_enable_buf (
.in_i(fetch_enable_i),
.in_i_t0(fetch_enable_i_t0),
.out_o(fetch_enable_buf),
.out_o_t0(fetch_enable_buf_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20440.4-20495.3" */
\$paramod$5c0dc9f9e0551018f7d8916b4fcabdef94a17390\ibex_core  u_ibex_core (
.alert_major_bus_o(alert_major_bus_o),
.alert_major_bus_o_t0(alert_major_bus_o_t0),
.alert_major_internal_o(core_alert_major_internal),
.alert_major_internal_o_t0(core_alert_major_internal_t0),
.alert_minor_o(alert_minor_o),
.alert_minor_o_t0(alert_minor_o_t0),
.boot_addr_i(boot_addr_i),
.boot_addr_i_t0(boot_addr_i_t0),
.clk_i(clk),
.core_busy_o(core_busy_d),
.core_busy_o_t0(core_busy_d_t0),
.crash_dump_o(crash_dump_o),
.crash_dump_o_t0(crash_dump_o_t0),
.data_addr_o(data_addr_o),
.data_addr_o_t0(data_addr_o_t0),
.data_be_o(data_be_o),
.data_be_o_t0(data_be_o_t0),
.data_err_i(data_err_i),
.data_err_i_t0(data_err_i_t0),
.data_gnt_i(data_gnt_i),
.data_gnt_i_t0(data_gnt_i_t0),
.data_rdata_i({ data_rdata_intg_i, data_rdata_i }),
.data_rdata_i_t0({ data_rdata_intg_i_t0, data_rdata_i_t0 }),
.data_req_o(data_req_o),
.data_req_o_t0(data_req_o_t0),
.data_rvalid_i(data_rvalid_i),
.data_rvalid_i_t0(data_rvalid_i_t0),
.data_wdata_o(data_wdata_core),
.data_wdata_o_t0(data_wdata_core_t0),
.data_we_o(data_we_o),
.data_we_o_t0(data_we_o_t0),
.debug_req_i(debug_req_i),
.debug_req_i_t0(debug_req_i_t0),
.double_fault_seen_o(double_fault_seen_o),
.double_fault_seen_o_t0(double_fault_seen_o_t0),
.dummy_instr_id_o(dummy_instr_id),
.dummy_instr_id_o_t0(dummy_instr_id_t0),
.dummy_instr_wb_o(dummy_instr_wb),
.dummy_instr_wb_o_t0(dummy_instr_wb_t0),
.fetch_enable_i(fetch_enable_buf),
.fetch_enable_i_t0(fetch_enable_buf_t0),
.hart_id_i(hart_id_i),
.hart_id_i_t0(hart_id_i_t0),
.ic_data_addr_o(ic_data_addr),
.ic_data_addr_o_t0(ic_data_addr_t0),
.ic_data_rdata_i(128'h00000000000000000000000000000000),
.ic_data_rdata_i_t0(128'h00000000000000000000000000000000),
.ic_data_req_o(ic_data_req),
.ic_data_req_o_t0(ic_data_req_t0),
.ic_data_wdata_o(ic_data_wdata),
.ic_data_wdata_o_t0(ic_data_wdata_t0),
.ic_data_write_o(ic_data_write),
.ic_data_write_o_t0(ic_data_write_t0),
.ic_scr_key_req_o(ic_scr_key_req),
.ic_scr_key_req_o_t0(ic_scr_key_req_t0),
.ic_scr_key_valid_i(1'h1),
.ic_scr_key_valid_i_t0(1'h0),
.ic_tag_addr_o(ic_tag_addr),
.ic_tag_addr_o_t0(ic_tag_addr_t0),
.ic_tag_rdata_i(44'h00000000000),
.ic_tag_rdata_i_t0(44'h00000000000),
.ic_tag_req_o(ic_tag_req),
.ic_tag_req_o_t0(ic_tag_req_t0),
.ic_tag_wdata_o(ic_tag_wdata),
.ic_tag_wdata_o_t0(ic_tag_wdata_t0),
.ic_tag_write_o(ic_tag_write),
.ic_tag_write_o_t0(ic_tag_write_t0),
.instr_addr_o(instr_addr_o),
.instr_addr_o_t0(instr_addr_o_t0),
.instr_err_i(instr_err_i),
.instr_err_i_t0(instr_err_i_t0),
.instr_gnt_i(instr_gnt_i),
.instr_gnt_i_t0(instr_gnt_i_t0),
.instr_rdata_i({ instr_rdata_intg_i, instr_rdata_i }),
.instr_rdata_i_t0({ instr_rdata_intg_i_t0, instr_rdata_i_t0 }),
.instr_req_o(instr_req_o),
.instr_req_o_t0(instr_req_o_t0),
.instr_rvalid_i(instr_rvalid_i),
.instr_rvalid_i_t0(instr_rvalid_i_t0),
.irq_external_i(irq_external_i),
.irq_external_i_t0(irq_external_i_t0),
.irq_fast_i(irq_fast_i),
.irq_fast_i_t0(irq_fast_i_t0),
.irq_nm_i(irq_nm_i),
.irq_nm_i_t0(irq_nm_i_t0),
.irq_pending_o(irq_pending),
.irq_pending_o_t0(irq_pending_t0),
.irq_software_i(irq_software_i),
.irq_software_i_t0(irq_software_i_t0),
.irq_timer_i(irq_timer_i),
.irq_timer_i_t0(irq_timer_i_t0),
.rf_raddr_a_o(rf_raddr_a),
.rf_raddr_a_o_t0(rf_raddr_a_t0),
.rf_raddr_b_o(rf_raddr_b),
.rf_raddr_b_o_t0(rf_raddr_b_t0),
.rf_rdata_a_ecc_i(rf_rdata_a_ecc_buf),
.rf_rdata_a_ecc_i_t0(rf_rdata_a_ecc_buf_t0),
.rf_rdata_b_ecc_i(rf_rdata_b_ecc_buf),
.rf_rdata_b_ecc_i_t0(rf_rdata_b_ecc_buf_t0),
.rf_waddr_wb_o(rf_waddr_wb),
.rf_waddr_wb_o_t0(rf_waddr_wb_t0),
.rf_wdata_wb_ecc_o(rf_wdata_wb_ecc),
.rf_wdata_wb_ecc_o_t0(rf_wdata_wb_ecc_t0),
.rf_we_wb_o(rf_we_wb),
.rf_we_wb_o_t0(rf_we_wb_t0),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20390.39-20393.3" */
\$paramod\prim_buf\Width=32'00000000000000000000000000100111  u_rf_rdata_a_ecc_buf (
.in_i(rf_rdata_a_ecc),
.in_i_t0(rf_rdata_a_ecc_t0),
.out_o(rf_rdata_a_ecc_buf),
.out_o_t0(rf_rdata_a_ecc_buf_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20394.39-20397.3" */
\$paramod\prim_buf\Width=32'00000000000000000000000000100111  u_rf_rdata_b_ecc_buf (
.in_i(rf_rdata_b_ecc),
.in_i_t0(rf_rdata_b_ecc_t0),
.out_o(rf_rdata_b_ecc_buf),
.out_o_t0(rf_rdata_b_ecc_buf_t0)
);
assign data_wdata_o = data_wdata_core[31:0];
assign data_wdata_o_t0 = data_wdata_core_t0[31:0];
assign scramble_req_o = 1'h0;
assign scramble_req_o_t0 = 1'h0;
endmodule

module prim_clock_gating(clk_i, en_i, test_en_i, clk_o, clk_o_t0, en_i_t0, test_en_i_t0);
/* src = "generated/sv2v_out.v:23091.2-23093.32" */
wire _00_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:23091.2-23093.32" */
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
/* src = "generated/sv2v_out.v:23086.8-23086.13" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:23089.14-23089.19" */
output clk_o;
wire clk_o;
/* cellift = 32'd1 */
output clk_o_t0;
wire clk_o_t0;
/* src = "generated/sv2v_out.v:23087.8-23087.12" */
input en_i;
wire en_i;
/* cellift = 32'd1 */
input en_i_t0;
wire en_i_t0;
/* src = "generated/sv2v_out.v:23090.6-23090.14" */
reg en_latch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:23090.6-23090.14" */
reg en_latch_t0;
/* src = "generated/sv2v_out.v:23088.8-23088.17" */
input test_en_i;
wire test_en_i;
/* cellift = 32'd1 */
input test_en_i_t0;
wire test_en_i_t0;
assign clk_o = en_latch & /* src = "generated/sv2v_out.v:23094.17-23094.33" */ clk_i;
assign clk_o_t0 = en_latch_t0 & clk_i;
/* taint_latch = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME prim_clock_gating */
/* PC_TAINT_INFO STATE_NAME en_latch_t0 */
always_latch
if (!clk_i) en_latch_t0 = _01_;
assign _02_ = ~ en_i;
assign _03_ = ~ test_en_i;
assign _04_ = en_i_t0 & _03_;
assign _05_ = test_en_i_t0 & _02_;
assign _06_ = en_i_t0 & test_en_i_t0;
assign _07_ = _04_ | _05_;
assign _01_ = _07_ | _06_;
/* src = "generated/sv2v_out.v:23091.2-23093.32" */
/* PC_TAINT_INFO MODULE_NAME prim_clock_gating */
/* PC_TAINT_INFO STATE_NAME en_latch */
always_latch
if (!clk_i) en_latch = _00_;
assign _00_ = en_i | /* src = "generated/sv2v_out.v:23093.15-23093.31" */ test_en_i;
endmodule

module prim_secded_inv_39_32_dec(data_i, data_o, syndrome_o, err_o, syndrome_o_t0, err_o_t0, data_o_t0, data_i_t0);
/* src = "generated/sv2v_out.v:29304.21-29304.63" */
wire [38:0] _000_;
/* src = "generated/sv2v_out.v:29306.21-29306.63" */
wire [38:0] _001_;
/* src = "generated/sv2v_out.v:29308.21-29308.63" */
wire [38:0] _002_;
/* src = "generated/sv2v_out.v:29310.16-29310.35" */
wire _003_;
/* src = "generated/sv2v_out.v:29311.16-29311.35" */
wire _004_;
/* src = "generated/sv2v_out.v:29312.16-29312.35" */
wire _005_;
/* src = "generated/sv2v_out.v:29313.16-29313.35" */
wire _006_;
/* src = "generated/sv2v_out.v:29314.16-29314.35" */
wire _007_;
/* src = "generated/sv2v_out.v:29315.16-29315.35" */
wire _008_;
/* src = "generated/sv2v_out.v:29316.16-29316.35" */
wire _009_;
/* src = "generated/sv2v_out.v:29317.16-29317.35" */
wire _010_;
/* src = "generated/sv2v_out.v:29318.16-29318.35" */
wire _011_;
/* src = "generated/sv2v_out.v:29319.16-29319.35" */
wire _012_;
/* src = "generated/sv2v_out.v:29320.17-29320.36" */
wire _013_;
/* src = "generated/sv2v_out.v:29321.17-29321.36" */
wire _014_;
/* src = "generated/sv2v_out.v:29322.17-29322.36" */
wire _015_;
/* src = "generated/sv2v_out.v:29323.17-29323.36" */
wire _016_;
/* src = "generated/sv2v_out.v:29324.17-29324.36" */
wire _017_;
/* src = "generated/sv2v_out.v:29325.17-29325.36" */
wire _018_;
/* src = "generated/sv2v_out.v:29326.17-29326.36" */
wire _019_;
/* src = "generated/sv2v_out.v:29327.17-29327.36" */
wire _020_;
/* src = "generated/sv2v_out.v:29328.17-29328.36" */
wire _021_;
/* src = "generated/sv2v_out.v:29329.17-29329.36" */
wire _022_;
/* src = "generated/sv2v_out.v:29330.17-29330.36" */
wire _023_;
/* src = "generated/sv2v_out.v:29331.17-29331.36" */
wire _024_;
/* src = "generated/sv2v_out.v:29332.17-29332.36" */
wire _025_;
/* src = "generated/sv2v_out.v:29333.17-29333.36" */
wire _026_;
/* src = "generated/sv2v_out.v:29334.17-29334.36" */
wire _027_;
/* src = "generated/sv2v_out.v:29335.17-29335.36" */
wire _028_;
/* src = "generated/sv2v_out.v:29336.17-29336.36" */
wire _029_;
/* src = "generated/sv2v_out.v:29337.17-29337.36" */
wire _030_;
/* src = "generated/sv2v_out.v:29338.17-29338.36" */
wire _031_;
/* src = "generated/sv2v_out.v:29339.17-29339.36" */
wire _032_;
/* src = "generated/sv2v_out.v:29340.17-29340.36" */
wire _033_;
/* src = "generated/sv2v_out.v:29341.17-29341.36" */
wire _034_;
/* src = "generated/sv2v_out.v:29343.14-29343.23" */
wire _035_;
/* src = "generated/sv2v_out.v:29343.26-29343.37" */
wire _036_;
/* src = "generated/sv2v_out.v:29298.15-29298.21" */
input [38:0] data_i;
wire [38:0] data_i;
/* cellift = 32'd1 */
input [38:0] data_i_t0;
wire [38:0] data_i_t0;
/* src = "generated/sv2v_out.v:29299.20-29299.26" */
output [31:0] data_o;
wire [31:0] data_o;
/* cellift = 32'd1 */
output [31:0] data_o_t0;
wire [31:0] data_o_t0;
/* src = "generated/sv2v_out.v:29301.19-29301.24" */
output [1:0] err_o;
wire [1:0] err_o;
/* cellift = 32'd1 */
output [1:0] err_o_t0;
wire [1:0] err_o_t0;
/* src = "generated/sv2v_out.v:29300.19-29300.29" */
output [6:0] syndrome_o;
wire [6:0] syndrome_o;
/* cellift = 32'd1 */
output [6:0] syndrome_o_t0;
wire [6:0] syndrome_o_t0;
assign err_o[1] = _035_ & /* src = "generated/sv2v_out.v:29343.14-29343.37" */ _036_;
assign { _002_[37], _001_[35], _000_[33] } = ~ { data_i[37], data_i[35], data_i[33] };
assign _003_ = syndrome_o == /* src = "generated/sv2v_out.v:29310.16-29310.35" */ 7'h19;
assign _004_ = syndrome_o == /* src = "generated/sv2v_out.v:29311.16-29311.35" */ 7'h54;
assign _005_ = syndrome_o == /* src = "generated/sv2v_out.v:29312.16-29312.35" */ 7'h61;
assign _006_ = syndrome_o == /* src = "generated/sv2v_out.v:29313.16-29313.35" */ 7'h34;
assign _007_ = syndrome_o == /* src = "generated/sv2v_out.v:29314.16-29314.35" */ 7'h1a;
assign _008_ = syndrome_o == /* src = "generated/sv2v_out.v:29315.16-29315.35" */ 7'h15;
assign _009_ = syndrome_o == /* src = "generated/sv2v_out.v:29316.16-29316.35" */ 7'h2a;
assign _010_ = syndrome_o == /* src = "generated/sv2v_out.v:29317.16-29317.35" */ 7'h4c;
assign _011_ = syndrome_o == /* src = "generated/sv2v_out.v:29318.16-29318.35" */ 7'h45;
assign _012_ = syndrome_o == /* src = "generated/sv2v_out.v:29319.16-29319.35" */ 7'h38;
assign _013_ = syndrome_o == /* src = "generated/sv2v_out.v:29320.17-29320.36" */ 7'h49;
assign _014_ = syndrome_o == /* src = "generated/sv2v_out.v:29321.17-29321.36" */ 7'h0d;
assign _015_ = syndrome_o == /* src = "generated/sv2v_out.v:29322.17-29322.36" */ 7'h51;
assign _016_ = syndrome_o == /* src = "generated/sv2v_out.v:29323.17-29323.36" */ 7'h31;
assign _017_ = syndrome_o == /* src = "generated/sv2v_out.v:29324.17-29324.36" */ 7'h68;
assign _018_ = syndrome_o == /* src = "generated/sv2v_out.v:29325.17-29325.36" */ 7'h07;
assign _019_ = syndrome_o == /* src = "generated/sv2v_out.v:29326.17-29326.36" */ 7'h1c;
assign _020_ = syndrome_o == /* src = "generated/sv2v_out.v:29327.17-29327.36" */ 7'h0b;
assign _021_ = syndrome_o == /* src = "generated/sv2v_out.v:29328.17-29328.36" */ 7'h25;
assign _022_ = syndrome_o == /* src = "generated/sv2v_out.v:29329.17-29329.36" */ 7'h26;
assign _023_ = syndrome_o == /* src = "generated/sv2v_out.v:29330.17-29330.36" */ 7'h46;
assign _024_ = syndrome_o == /* src = "generated/sv2v_out.v:29331.17-29331.36" */ 7'h0e;
assign _025_ = syndrome_o == /* src = "generated/sv2v_out.v:29332.17-29332.36" */ 7'h70;
assign _026_ = syndrome_o == /* src = "generated/sv2v_out.v:29333.17-29333.36" */ 7'h32;
assign _027_ = syndrome_o == /* src = "generated/sv2v_out.v:29334.17-29334.36" */ 7'h2c;
assign _028_ = syndrome_o == /* src = "generated/sv2v_out.v:29335.17-29335.36" */ 7'h13;
assign _029_ = syndrome_o == /* src = "generated/sv2v_out.v:29336.17-29336.36" */ 7'h23;
assign _030_ = syndrome_o == /* src = "generated/sv2v_out.v:29337.17-29337.36" */ 7'h62;
assign _031_ = syndrome_o == /* src = "generated/sv2v_out.v:29338.17-29338.36" */ 7'h4a;
assign _032_ = syndrome_o == /* src = "generated/sv2v_out.v:29339.17-29339.36" */ 7'h29;
assign _033_ = syndrome_o == /* src = "generated/sv2v_out.v:29340.17-29340.36" */ 7'h16;
assign _034_ = syndrome_o == /* src = "generated/sv2v_out.v:29341.17-29341.36" */ 7'h52;
assign _035_ = ~ /* src = "generated/sv2v_out.v:29343.14-29343.23" */ err_o[0];
assign _036_ = | /* src = "generated/sv2v_out.v:29343.26-29343.37" */ syndrome_o;
assign syndrome_o[0] = ^ /* src = "generated/sv2v_out.v:29303.19-29303.64" */ { 6'h00, data_i[32], 2'h0, data_i[29], 2'h0, data_i[26:25], 6'h00, data_i[18:17], 1'h0, data_i[15], 1'h0, data_i[13:10], 1'h0, data_i[8], 2'h0, data_i[5], 2'h0, data_i[2], 1'h0, data_i[0] };
assign syndrome_o[1] = ^ /* src = "generated/sv2v_out.v:29304.19-29304.64" */ { 5'h00, _000_[33], 1'h0, data_i[31:30], 1'h0, data_i[28:25], 1'h0, data_i[23], 1'h0, data_i[21:19], 1'h0, data_i[17], 1'h0, data_i[15], 8'h00, data_i[6], 1'h0, data_i[4], 4'h0 };
assign syndrome_o[2] = ^ /* src = "generated/sv2v_out.v:29305.19-29305.64" */ { 4'h0, data_i[34], 3'h0, data_i[30], 5'h00, data_i[24], 2'h0, data_i[21:18], 1'h0, data_i[16:15], 3'h0, data_i[11], 2'h0, data_i[8:7], 1'h0, data_i[5], 1'h0, data_i[3], 1'h0, data_i[1], 1'h0 };
assign syndrome_o[3] = ^ /* src = "generated/sv2v_out.v:29306.19-29306.64" */ { 3'h0, _001_[35], 5'h00, data_i[29:28], 3'h0, data_i[24], 2'h0, data_i[21], 3'h0, data_i[17:16], 1'h0, data_i[14], 2'h0, data_i[11:9], 1'h0, data_i[7:6], 1'h0, data_i[4], 3'h0, data_i[0] };
assign syndrome_o[4] = ^ /* src = "generated/sv2v_out.v:29307.19-29307.64" */ { 2'h0, data_i[36], 4'h0, data_i[31:30], 4'h0, data_i[25], 1'h0, data_i[23:22], 5'h00, data_i[16], 2'h0, data_i[13:12], 2'h0, data_i[9], 3'h0, data_i[5:3], 1'h0, data_i[1:0] };
assign syndrome_o[5] = ^ /* src = "generated/sv2v_out.v:29308.19-29308.64" */ { 1'h0, _002_[37], 7'h00, data_i[29], 1'h0, data_i[27:26], 1'h0, data_i[24:22], 2'h0, data_i[19:18], 3'h0, data_i[14:13], 3'h0, data_i[9], 2'h0, data_i[6], 2'h0, data_i[3:2], 2'h0 };
assign syndrome_o[6] = ^ /* src = "generated/sv2v_out.v:29309.19-29309.64" */ { data_i[38], 6'h00, data_i[31], 2'h0, data_i[28:27], 4'h0, data_i[22], 1'h0, data_i[20], 5'h00, data_i[14], 1'h0, data_i[12], 1'h0, data_i[10], 1'h0, data_i[8:7], 4'h0, data_i[2:1], 1'h0 };
assign err_o[0] = ^ /* src = "generated/sv2v_out.v:29342.14-29342.25" */ syndrome_o;
assign data_o[0] = _003_ ^ /* src = "generated/sv2v_out.v:29310.15-29310.48" */ data_i[0];
assign data_o[1] = _004_ ^ /* src = "generated/sv2v_out.v:29311.15-29311.48" */ data_i[1];
assign data_o[2] = _005_ ^ /* src = "generated/sv2v_out.v:29312.15-29312.48" */ data_i[2];
assign data_o[3] = _006_ ^ /* src = "generated/sv2v_out.v:29313.15-29313.48" */ data_i[3];
assign data_o[4] = _007_ ^ /* src = "generated/sv2v_out.v:29314.15-29314.48" */ data_i[4];
assign data_o[5] = _008_ ^ /* src = "generated/sv2v_out.v:29315.15-29315.48" */ data_i[5];
assign data_o[6] = _009_ ^ /* src = "generated/sv2v_out.v:29316.15-29316.48" */ data_i[6];
assign data_o[7] = _010_ ^ /* src = "generated/sv2v_out.v:29317.15-29317.48" */ data_i[7];
assign data_o[8] = _011_ ^ /* src = "generated/sv2v_out.v:29318.15-29318.48" */ data_i[8];
assign data_o[9] = _012_ ^ /* src = "generated/sv2v_out.v:29319.15-29319.48" */ data_i[9];
assign data_o[10] = _013_ ^ /* src = "generated/sv2v_out.v:29320.16-29320.50" */ data_i[10];
assign data_o[11] = _014_ ^ /* src = "generated/sv2v_out.v:29321.16-29321.50" */ data_i[11];
assign data_o[12] = _015_ ^ /* src = "generated/sv2v_out.v:29322.16-29322.50" */ data_i[12];
assign data_o[13] = _016_ ^ /* src = "generated/sv2v_out.v:29323.16-29323.50" */ data_i[13];
assign data_o[14] = _017_ ^ /* src = "generated/sv2v_out.v:29324.16-29324.50" */ data_i[14];
assign data_o[15] = _018_ ^ /* src = "generated/sv2v_out.v:29325.16-29325.50" */ data_i[15];
assign data_o[16] = _019_ ^ /* src = "generated/sv2v_out.v:29326.16-29326.50" */ data_i[16];
assign data_o[17] = _020_ ^ /* src = "generated/sv2v_out.v:29327.16-29327.50" */ data_i[17];
assign data_o[18] = _021_ ^ /* src = "generated/sv2v_out.v:29328.16-29328.50" */ data_i[18];
assign data_o[19] = _022_ ^ /* src = "generated/sv2v_out.v:29329.16-29329.50" */ data_i[19];
assign data_o[20] = _023_ ^ /* src = "generated/sv2v_out.v:29330.16-29330.50" */ data_i[20];
assign data_o[21] = _024_ ^ /* src = "generated/sv2v_out.v:29331.16-29331.50" */ data_i[21];
assign data_o[22] = _025_ ^ /* src = "generated/sv2v_out.v:29332.16-29332.50" */ data_i[22];
assign data_o[23] = _026_ ^ /* src = "generated/sv2v_out.v:29333.16-29333.50" */ data_i[23];
assign data_o[24] = _027_ ^ /* src = "generated/sv2v_out.v:29334.16-29334.50" */ data_i[24];
assign data_o[25] = _028_ ^ /* src = "generated/sv2v_out.v:29335.16-29335.50" */ data_i[25];
assign data_o[26] = _029_ ^ /* src = "generated/sv2v_out.v:29336.16-29336.50" */ data_i[26];
assign data_o[27] = _030_ ^ /* src = "generated/sv2v_out.v:29337.16-29337.50" */ data_i[27];
assign data_o[28] = _031_ ^ /* src = "generated/sv2v_out.v:29338.16-29338.50" */ data_i[28];
assign data_o[29] = _032_ ^ /* src = "generated/sv2v_out.v:29339.16-29339.50" */ data_i[29];
assign data_o[30] = _033_ ^ /* src = "generated/sv2v_out.v:29340.16-29340.50" */ data_i[30];
assign data_o[31] = _034_ ^ /* src = "generated/sv2v_out.v:29341.16-29341.50" */ data_i[31];
assign { _000_[38:34], _000_[32:0] } = { 6'h00, data_i[31:30], 1'h0, data_i[28:25], 1'h0, data_i[23], 1'h0, data_i[21:19], 1'h0, data_i[17], 1'h0, data_i[15], 8'h00, data_i[6], 1'h0, data_i[4], 4'h0 };
assign { _001_[38:36], _001_[34:0] } = { 8'h00, data_i[29:28], 3'h0, data_i[24], 2'h0, data_i[21], 3'h0, data_i[17:16], 1'h0, data_i[14], 2'h0, data_i[11:9], 1'h0, data_i[7:6], 1'h0, data_i[4], 3'h0, data_i[0] };
assign { _002_[38], _002_[36:0] } = { 8'h00, data_i[29], 1'h0, data_i[27:26], 1'h0, data_i[24:22], 2'h0, data_i[19:18], 3'h0, data_i[14:13], 3'h0, data_i[9], 2'h0, data_i[6], 2'h0, data_i[3:2], 2'h0 };
assign data_o_t0 = data_i_t0[31:0];
assign err_o_t0 = 2'h0;
assign syndrome_o_t0 = 7'h00;
endmodule

module prim_secded_inv_39_32_enc(data_i, data_o, data_o_t0, data_i_t0);
/* src = "generated/sv2v_out.v:29359.16-29359.42" */
wire _00_;
/* src = "generated/sv2v_out.v:29361.16-29361.42" */
wire _01_;
/* src = "generated/sv2v_out.v:29363.16-29363.42" */
wire _02_;
/* src = "generated/sv2v_out.v:29350.15-29350.21" */
input [31:0] data_i;
wire [31:0] data_i;
/* cellift = 32'd1 */
input [31:0] data_i_t0;
wire [31:0] data_i_t0;
/* src = "generated/sv2v_out.v:29351.20-29351.26" */
output [38:0] data_o;
wire [38:0] data_o;
/* cellift = 32'd1 */
output [38:0] data_o_t0;
wire [38:0] data_o_t0;
assign { data_o[37], data_o[35], data_o[33] } = ~ { _02_, _01_, _00_ };
assign data_o[32] = ^ /* src = "generated/sv2v_out.v:29358.16-29358.42" */ { 9'h000, data_i[29], 2'h0, data_i[26:25], 6'h00, data_i[18:17], 1'h0, data_i[15], 1'h0, data_i[13:10], 1'h0, data_i[8], 2'h0, data_i[5], 2'h0, data_i[2], 1'h0, data_i[0] };
assign _00_ = ^ /* src = "generated/sv2v_out.v:29359.16-29359.42" */ { 7'h00, data_i[31:30], 1'h0, data_i[28:25], 1'h0, data_i[23], 1'h0, data_i[21:19], 1'h0, data_i[17], 1'h0, data_i[15], 8'h00, data_i[6], 1'h0, data_i[4], 4'h0 };
assign data_o[34] = ^ /* src = "generated/sv2v_out.v:29360.16-29360.42" */ { 8'h00, data_i[30], 5'h00, data_i[24], 2'h0, data_i[21:18], 1'h0, data_i[16:15], 3'h0, data_i[11], 2'h0, data_i[8:7], 1'h0, data_i[5], 1'h0, data_i[3], 1'h0, data_i[1], 1'h0 };
assign _01_ = ^ /* src = "generated/sv2v_out.v:29361.16-29361.42" */ { 9'h000, data_i[29:28], 3'h0, data_i[24], 2'h0, data_i[21], 3'h0, data_i[17:16], 1'h0, data_i[14], 2'h0, data_i[11:9], 1'h0, data_i[7:6], 1'h0, data_i[4], 3'h0, data_i[0] };
assign data_o[36] = ^ /* src = "generated/sv2v_out.v:29362.16-29362.42" */ { 7'h00, data_i[31:30], 4'h0, data_i[25], 1'h0, data_i[23:22], 5'h00, data_i[16], 2'h0, data_i[13:12], 2'h0, data_i[9], 3'h0, data_i[5:3], 1'h0, data_i[1:0] };
assign _02_ = ^ /* src = "generated/sv2v_out.v:29363.16-29363.42" */ { 9'h000, data_i[29], 1'h0, data_i[27:26], 1'h0, data_i[24:22], 2'h0, data_i[19:18], 3'h0, data_i[14:13], 3'h0, data_i[9], 2'h0, data_i[6], 2'h0, data_i[3:2], 2'h0 };
assign data_o[38] = ^ /* src = "generated/sv2v_out.v:29364.16-29364.42" */ { 7'h00, data_i[31], 2'h0, data_i[28:27], 4'h0, data_i[22], 1'h0, data_i[20], 5'h00, data_i[14], 1'h0, data_i[12], 1'h0, data_i[10], 1'h0, data_i[8:7], 4'h0, data_i[2:1], 1'h0 };
assign data_o[31:0] = data_i;
assign data_o_t0 = { 7'h00, data_i_t0 };
endmodule