`include "formal/assumptions/cellift_data_flow_picorv32_di_asm.sv"
`include "formal/assumptions/cellift_data_flow_picorv32_ti_asm.sv"
