asm_declass_cpuregs_wrdata_t0: assume property(!cpuregs_wrdata_t0);
