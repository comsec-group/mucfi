asm_declass_u_ibex_core__rf_wdata_wb_ecc_o_t0: assume property(!u_ibex_core__rf_wdata_wb_ecc_o_t0);
asm_declass_u_ibex_core__wb_stage_i__rf_wdata_fwd_wb_o_t0: assume property(!u_ibex_core__wb_stage_i__rf_wdata_fwd_wb_o_t0);
