bit gen_uc_rs1;
assign gen_uc_rs1 = ((((| { (| { (| { ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1e) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1f)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1d), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1c) }), ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1a) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1b)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h19), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h18) }), (| { ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h16) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h17)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h15), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h14) }), ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h12) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h13)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h11), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h10) }) & (((| { (| { ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1e) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1f)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1d), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1c) }), ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1a) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1b)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h19), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h18) }) & (((| { ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1e) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1f)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1d), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1c) }) & ((((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1e) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1f)) & (((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1f)) | ((~ (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1f))))) | ((~ ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1e) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1f))) & (((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1d)) | ((~ (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1d))))))) | ((~ (| { ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1e) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1f)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1d), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1c) })) & ((((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1a) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1b)) & (((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1b)) | ((~ (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1b))))) | ((~ ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1a) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1b))) & (((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h19)) | ((~ (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h19))))))))) | ((~ (| { (| { ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1e) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1f)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1d), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1c) }), ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1a) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1b)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h19), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h18) })) & (((| { ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h16) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h17)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h15), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h14) }) & ((((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h16) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h17)) & (((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h17)) | ((~ (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h17))))) | ((~ ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h16) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h17))) & (((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h15)) | ((~ (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h15))))))) | ((~ (| { ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h16) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h17)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h15), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h14) })) & ((((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h12) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h13)) & (((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h13)) | ((~ (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h13))))) | ((~ ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h12) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h13))) & (((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h11)) | ((~ (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h11))))))))))) | ((~ (| { (| { (| { ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1e) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1f)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1d), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1c) }), ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1a) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h1b)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h19), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h18) }), (| { ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h16) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h17)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h15), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h14) }), ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h12) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h13)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h11), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h10) })) & (((| { (| { ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0e) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0f)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0d), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0c) }), ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0a) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0b)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h09), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h08) }) & (((| { ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0e) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0f)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0d), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0c) }) & ((((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0e) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0f)) & (((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0f)) | ((~ (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0f))))) | ((~ ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0e) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0f))) & (((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0d)) | ((~ (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0d))))))) | ((~ (| { ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0e) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0f)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0d), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0c) })) & ((((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0a) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0b)) & (((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0b)) | ((~ (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0b))))) | ((~ ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0a) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0b))) & (((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h09)) | ((~ (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h09))))))))) | ((~ (| { (| { ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0e) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0f)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0d), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0c) }), ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0a) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h0b)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h09), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h08) })) & (((| { ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h06) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h07)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h05), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h04) }) & ((((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h06) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h07)) & (((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h07)) | ((~ (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h07))))) | ((~ ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h06) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h07))) & (((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h05)) | ((~ (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h05))))))) | ((~ (| { ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h06) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h07)), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h05), (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h04) })) & ((((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h02) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h03)) & (((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h03)) | ((~ (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h03))))) | ((~ ((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h02) | (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h03))) & (((gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h01)) | ((~ (gen_regfile_ff__register_file_i__raddr_a_i  ==  5'h01)) & ((gen_regfile_ff__register_file_i__dummy_instr_id_i ) | ((~ gen_regfile_ff__register_file_i__dummy_instr_id_i ))))))))))))));
