// kceesay@ee-tik-cn105:/data/kceesay/workspace/cellift-designs/cellift-picorv32/cellift/generated$ git log -1
// commit eb41d95179d5064eb1a8f435df46879702022c92 (HEAD -> master, origin/master, origin/HEAD)
// Author: Flavien Solt <flsolt@ethz.ch>
// Date:   Thu Nov 16 10:41:00 2023 +0100

//     Accelerate mem bandwidth by using the lookahead interface
// kceesay@ee-tik-cn105:/data/kceesay/workspace/cellift-designs/cellift-picorv32/cellift/generated$ git branch
// * master

// update condition Yosys

/* Generated by Yosys 0.29+11 (git sha1 eb3eaeb79, gcc 11.4.0-1ubuntu1~22.04 -Og -fPIC) */
// cellift-picorv32 git commit eb41d95179d5064eb1a8f435df46879702022c92

/* cellift =  1  */
/* dynports =  1  */
/* hdlname = "\\picorv32" */
/* src = "generated/out/vanilla.sv:1.1-1811.10" */
module cellift_data_flow_picorv32 (clk, resetn, trap, mem_valid, mem_instr, mem_ready, mem_addr, mem_wdata, mem_wstrb, mem_rdata, mem_la_read, mem_la_write, mem_la_addr, mem_la_wdata, mem_la_wstrb, pcpi_valid, pcpi_insn, pcpi_rs1, pcpi_rs2, pcpi_wr, pcpi_rd
, pcpi_wait, pcpi_ready, irq, eoi, rvfi_valid, rvfi_order, rvfi_insn, rvfi_trap, rvfi_halt, rvfi_intr, rvfi_mode, rvfi_ixl, rvfi_rs1_addr, rvfi_rs2_addr, rvfi_rs1_rdata, rvfi_rs2_rdata, rvfi_rd_addr, rvfi_rd_wdata, rvfi_pc_rdata, rvfi_pc_wdata, rvfi_mem_addr
, rvfi_mem_rmask, rvfi_mem_wmask, rvfi_mem_rdata, rvfi_mem_wdata, rvfi_csr_mcycle_rmask, rvfi_csr_mcycle_wmask, rvfi_csr_mcycle_rdata, rvfi_csr_mcycle_wdata, rvfi_csr_minstret_rmask, rvfi_csr_minstret_wmask, rvfi_csr_minstret_rdata, rvfi_csr_minstret_wdata, trace_valid, trace_data, trap_t0, trace_valid_t0, trace_data_t0, rvfi_valid_t0, rvfi_trap_t0, rvfi_rs2_rdata_t0, rvfi_rs2_addr_t0
, rvfi_rs1_rdata_t0, rvfi_rs1_addr_t0, rvfi_rd_wdata_t0, rvfi_rd_addr_t0, rvfi_pc_wdata_t0, rvfi_pc_rdata_t0, rvfi_order_t0, rvfi_mode_t0, rvfi_mem_wmask_t0, rvfi_mem_wdata_t0, rvfi_mem_rmask_t0, rvfi_mem_rdata_t0, rvfi_mem_addr_t0, rvfi_ixl_t0, rvfi_intr_t0, rvfi_insn_t0, rvfi_halt_t0, rvfi_csr_minstret_wmask_t0, rvfi_csr_minstret_wdata_t0, rvfi_csr_minstret_rmask_t0, rvfi_csr_minstret_rdata_t0
, rvfi_csr_mcycle_wmask_t0, rvfi_csr_mcycle_wdata_t0, rvfi_csr_mcycle_rmask_t0, rvfi_csr_mcycle_rdata_t0, mem_wstrb_t0, mem_wdata_t0, mem_valid_t0, mem_ready_t0, mem_rdata_t0, mem_la_wstrb_t0, mem_la_write_t0, mem_la_wdata_t0, mem_la_read_t0, mem_la_addr_t0, mem_instr_t0, mem_addr_t0, irq_t0, eoi_t0, pcpi_insn_t0, pcpi_rd_t0, pcpi_ready_t0
, pcpi_rs1_t0, pcpi_rs2_t0, pcpi_valid_t0, pcpi_wait_t0, pcpi_wr_t0);
  /* src = "generated/out/vanilla.sv:1180.2-1182.42" */
  wire [4:0] _0000_;
  /* src = "generated/out/vanilla.sv:1180.2-1182.42" */
  wire [31:0] _0001_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1180.2-1182.42" */
  wire [31:0] _0002_;
  /* src = "generated/out/vanilla.sv:1180.2-1182.42" */
  wire [31:0] _0003_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [31:0] _0004_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [31:0] _0005_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _0006_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [31:0] _0007_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [31:0] _0008_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _0009_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _0010_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
  wire _0011_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
  wire _0012_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
  wire _0013_;
  /* src = "generated/out/vanilla.sv:339.2-446.5" */
  /* unused_bits = "0 1 2 3 4 5 6" */
  wire [31:0] _0014_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:339.2-446.5" */
  /* unused_bits = "0 1 2 3 4 5 6" */
  wire [31:0] _0015_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
  wire [1:0] _0016_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
  wire _0017_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [31:0] _0018_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [31:0] _0019_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [4:0] _0020_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
  wire _0021_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _0022_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _0023_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _0024_;
  /* src = "generated/out/vanilla.sv:1144.2-1150.5" */
  wire _0025_;
  /* src = "generated/out/vanilla.sv:1156.2-1179.5" */
  wire [31:0] _0026_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1156.2-1179.5" */
  wire [31:0] _0027_;
  /* src = "generated/out/vanilla.sv:1156.2-1179.5" */
  wire _0028_;
  /* src = "generated/out/vanilla.sv:761.2-788.5" */
  wire [31:0] _0029_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:761.2-788.5" */
  wire [31:0] _0030_;
  /* src = "generated/out/vanilla.sv:761.2-788.5" */
  wire [4:0] _0031_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:761.2-788.5" */
  wire [4:0] _0032_;
  /* src = "generated/out/vanilla.sv:761.2-788.5" */
  wire [4:0] _0033_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:761.2-788.5" */
  wire [4:0] _0034_;
  /* src = "generated/out/vanilla.sv:312.2-338.10" */
  wire [31:0] _0035_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:312.2-338.10" */
  wire [31:0] _0036_;
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _0037_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _0038_;
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _0039_;
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _0040_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _0041_;
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _0042_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _0043_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _0044_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _0045_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [31:0] _0046_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire [31:0] _0047_;
  /* src = "generated/out/vanilla.sv:761.2-788.5" */
  wire [31:0] _0048_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:761.2-788.5" */
  wire [31:0] _0049_;
  /* src = "generated/out/vanilla.sv:312.2-338.10" */
  wire [31:0] _0050_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:312.2-338.10" */
  wire [31:0] _0051_;
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _0052_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _0053_;
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _0054_;
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _0055_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _0056_;
  /* src = "generated/out/vanilla.sv:1782.2-1810.5" */
  wire [63:0] _0057_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _0058_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _0059_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _0060_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _0061_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _0062_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
  wire _0063_;
  reg [4:0] _0064_;
  reg [4:0] _0065_;
  /* src = "generated/out/vanilla.sv:1110.52-1110.69" */
  wire [31:0] _0066_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1110.52-1110.69" */
  wire [31:0] _0067_;
  /* src = "generated/out/vanilla.sv:1163.23-1163.55" */
  wire [31:0] _0068_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1163.23-1163.55" */
  wire [31:0] _0069_;
  /* src = "generated/out/vanilla.sv:1223.29-1223.44" */
  wire [63:0] _0070_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1223.29-1223.44" */
  wire [63:0] _0071_;
  /* src = "generated/out/vanilla.sv:1323.23-1323.62" */
  wire [31:0] _0072_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1323.23-1323.62" */
  wire [31:0] _0073_;
  /* src = "generated/out/vanilla.sv:1335.23-1335.38" */
  wire [63:0] _0074_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1335.23-1335.38" */
  wire [63:0] _0075_;
  /* src = "generated/out/vanilla.sv:1341.23-1341.49" */
  wire [31:0] _0076_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1341.23-1341.49" */
  wire [31:0] _0077_;
  /* src = "generated/out/vanilla.sv:1554.17-1554.37" */
  wire [31:0] _0078_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1554.17-1554.37" */
  wire [31:0] _0079_;
  /* src = "generated/out/vanilla.sv:1618.19-1618.40" */
  wire [31:0] _0080_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1618.19-1618.40" */
  wire [31:0] _0081_;
  /* src = "generated/out/vanilla.sv:1716.27-1716.50" */
  wire [63:0] _0082_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1716.27-1716.50" */
  wire [63:0] _0083_;
  /* src = "generated/out/vanilla.sv:299.59-299.96" */
  wire [29:0] _0084_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:299.59-299.96" */
  wire [29:0] _0085_;
  /* src = "generated/out/vanilla.sv:829.23-829.49" */
  /* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _0086_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:829.23-829.49" */
  /* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _0087_;
  /* src = "generated/out/vanilla.sv:833.24-833.50" */
  /* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _0088_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:833.24-833.50" */
  /* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _0089_;
  /* src = "generated/out/vanilla.sv:1137.39-1137.56" */
  wire [31:0] _0090_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1137.39-1137.56" */
  wire [31:0] _0091_;
  /* src = "generated/out/vanilla.sv:1280.53-1280.95" */
  wire [31:0] _0092_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1280.53-1280.95" */
  wire [31:0] _0093_;
  /* src = "generated/out/vanilla.sv:472.18-472.51" */
  wire [3:0] _0094_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:472.18-472.51" */
  wire [3:0] _0095_;
  wire [31:0] _0096_;
  wire [31:0] _0097_;
  wire [63:0] _0098_;
  wire [31:0] _0099_;
  wire [63:0] _0100_;
  wire [63:0] _0101_;
  wire [29:0] _0102_;
  wire [31:0] _0103_;
  wire [31:0] _0104_;
  wire [31:0] _0105_;
  wire [31:0] _0106_;
  wire [31:0] _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire [31:0] _0155_;
  wire [31:0] _0156_;
  wire [31:0] _0157_;
  wire [31:0] _0158_;
  wire [31:0] _0159_;
  wire [31:0] _0160_;
  wire [31:0] _0161_;
  wire [31:0] _0162_;
  wire [31:0] _0163_;
  wire [31:0] _0164_;
  wire [4:0] _0165_;
  wire [31:0] _0166_;
  wire [31:0] _0167_;
  wire [31:0] _0168_;
  wire [31:0] _0169_;
  wire [31:0] _0170_;
  wire [31:0] _0171_;
  wire [31:0] _0172_;
  wire [31:0] _0173_;
  wire [31:0] _0174_;
  wire [31:0] _0175_;
  wire [31:0] _0176_;
  wire [31:0] _0177_;
  wire [31:0] _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire [3:0] _0186_;
  wire [3:0] _0187_;
  wire [3:0] _0188_;
  wire [3:0] _0189_;
  wire [3:0] _0190_;
  wire [3:0] _0191_;
  wire [3:0] _0192_;
  wire [3:0] _0193_;
  wire [3:0] _0194_;
  wire _0195_;
  wire [31:0] _0196_;
  wire [31:0] _0197_;
  wire [31:0] _0198_;
  wire [31:0] _0199_;
  wire [31:0] _0200_;
  wire [4:0] _0201_;
  wire [4:0] _0202_;
  wire [4:0] _0203_;
  wire [4:0] _0204_;
  wire [4:0] _0205_;
  wire [4:0] _0206_;
  wire [4:0] _0207_;
  wire [4:0] _0208_;
  wire [4:0] _0209_;
  wire [4:0] _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire [4:0] _0214_;
  wire [2:0] _0215_;
  wire [2:0] _0216_;
  wire [2:0] _0217_;
  wire [2:0] _0218_;
  wire [2:0] _0219_;
  wire [2:0] _0220_;
  wire [2:0] _0221_;
  wire [2:0] _0222_;
  wire [2:0] _0223_;
  wire [5:0] _0224_;
  wire [5:0] _0225_;
  wire [5:0] _0226_;
  wire [5:0] _0227_;
  wire [5:0] _0228_;
  wire [5:0] _0229_;
  wire [5:0] _0230_;
  wire [5:0] _0231_;
  wire [5:0] _0232_;
  wire [5:0] _0233_;
  wire [5:0] _0234_;
  wire [5:0] _0235_;
  wire [31:0] _0236_;
  wire [31:0] _0237_;
  wire [31:0] _0238_;
  wire [31:0] _0239_;
  wire [31:0] _0240_;
  wire [31:0] _0241_;
  wire [31:0] _0242_;
  wire [31:0] _0243_;
  wire [31:0] _0244_;
  wire [31:0] _0245_;
  wire [31:0] _0246_;
  wire [31:0] _0247_;
  wire [31:0] _0248_;
  wire [31:0] _0249_;
  wire [31:0] _0250_;
  wire [31:0] _0251_;
  wire [31:0] _0252_;
  wire _0253_;
  wire [31:0] _0254_;
  wire [31:0] _0255_;
  wire _0256_;
  wire [31:0] _0257_;
  wire _0258_;
  wire [31:0] _0259_;
  wire [31:0] _0260_;
  wire [31:0] _0261_;
  wire [31:0] _0262_;
  wire [31:0] _0263_;
  wire [31:0] _0264_;
  wire [31:0] _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire [2:0] _0274_;
  wire [1:0] _0275_;
  wire [11:0] _0276_;
  wire [3:0] _0277_;
  wire [3:0] _0278_;
  wire [3:0] _0279_;
  wire [3:0] _0280_;
  wire [3:0] _0281_;
  wire [3:0] _0282_;
  wire [3:0] _0283_;
  wire _0284_;
  wire [4:0] _0285_;
  wire [4:0] _0286_;
  wire [4:0] _0287_;
  wire [4:0] _0288_;
  wire [7:0] _0289_;
  wire [4:0] _0290_;
  wire [4:0] _0291_;
  wire [4:0] _0292_;
  wire [31:0] _0293_;
  wire [4:0] _0294_;
  wire [31:0] _0295_;
  wire [31:0] _0296_;
  wire [15:0] _0297_;
  wire [15:0] _0298_;
  wire [15:0] _0299_;
  wire _0300_;
  wire [3:0] _0301_;
  wire [3:0] _0302_;
  wire [3:0] _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire [4:0] _0308_;
  wire [4:0] _0309_;
  wire [4:0] _0310_;
  wire [4:0] _0311_;
  wire [4:0] _0312_;
  wire [4:0] _0313_;
  wire [2:0] _0314_;
  wire [2:0] _0315_;
  wire [2:0] _0316_;
  wire [2:0] _0317_;
  wire [2:0] _0318_;
  wire [2:0] _0319_;
  wire [2:0] _0320_;
  wire [2:0] _0321_;
  wire [2:0] _0322_;
  wire [2:0] _0323_;
  wire [2:0] _0324_;
  wire [2:0] _0325_;
  wire [2:0] _0326_;
  wire [2:0] _0327_;
  wire [2:0] _0328_;
  wire [3:0] _0329_;
  wire [3:0] _0330_;
  wire [5:0] _0331_;
  wire [5:0] _0332_;
  wire [5:0] _0333_;
  wire [5:0] _0334_;
  wire [5:0] _0335_;
  wire [5:0] _0336_;
  wire [5:0] _0337_;
  wire [5:0] _0338_;
  wire [5:0] _0339_;
  wire [5:0] _0340_;
  wire [5:0] _0341_;
  wire [63:0] _0342_;
  wire [63:0] _0343_;
  wire [31:0] _0344_;
  wire [31:0] _0345_;
  wire [31:0] _0346_;
  wire [31:0] _0347_;
  wire [31:0] _0348_;
  wire [31:0] _0349_;
  wire [31:0] _0350_;
  wire [31:0] _0351_;
  wire [31:0] _0352_;
  wire [31:0] _0353_;
  wire _0354_;
  wire [31:0] _0355_;
  wire [31:0] _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire [31:0] _0454_;
  wire [31:0] _0455_;
  wire [31:0] _0456_;
  wire [31:0] _0457_;
  wire [31:0] _0458_;
  wire [31:0] _0459_;
  wire [31:0] _0460_;
  wire [31:0] _0461_;
  wire [31:0] _0462_;
  wire [31:0] _0463_;
  wire [31:0] _0464_;
  wire [31:0] _0465_;
  wire [31:0] _0466_;
  wire [31:0] _0467_;
  wire [31:0] _0468_;
  wire [31:0] _0469_;
  wire [31:0] _0470_;
  wire [31:0] _0471_;
  wire [31:0] _0472_;
  wire [31:0] _0473_;
  wire [31:0] _0474_;
  wire [31:0] _0475_;
  wire [31:0] _0476_;
  wire [31:0] _0477_;
  wire [31:0] _0478_;
  wire [31:0] _0479_;
  wire [31:0] _0480_;
  wire [31:0] _0481_;
  wire [4:0] _0482_;
  wire [31:0] _0483_;
  wire [31:0] _0484_;
  wire [31:0] _0485_;
  wire [31:0] _0486_;
  wire [31:0] _0487_;
  wire [31:0] _0488_;
  wire [31:0] _0489_;
  wire [31:0] _0490_;
  wire [31:0] _0491_;
  wire [31:0] _0492_;
  wire [31:0] _0493_;
  wire [31:0] _0494_;
  wire [31:0] _0495_;
  wire [31:0] _0496_;
  wire [31:0] _0497_;
  wire [31:0] _0498_;
  wire [31:0] _0499_;
  wire [31:0] _0500_;
  wire [31:0] _0501_;
  wire [31:0] _0502_;
  wire [31:0] _0503_;
  wire [31:0] _0504_;
  wire [31:0] _0505_;
  wire [31:0] _0506_;
  wire [31:0] _0507_;
  wire [31:0] _0508_;
  wire [31:0] _0509_;
  wire [31:0] _0510_;
  wire [31:0] _0511_;
  wire [31:0] _0512_;
  wire [31:0] _0513_;
  wire [31:0] _0514_;
  wire [31:0] _0515_;
  wire [31:0] _0516_;
  wire [31:0] _0517_;
  wire [31:0] _0518_;
  wire [31:0] _0519_;
  wire [31:0] _0520_;
  wire [31:0] _0521_;
  wire [31:0] _0522_;
  wire [31:0] _0523_;
  wire [31:0] _0524_;
  wire [31:0] _0525_;
  wire [31:0] _0526_;
  wire [31:0] _0527_;
  wire [31:0] _0528_;
  wire [31:0] _0529_;
  wire [31:0] _0530_;
  wire [31:0] _0531_;
  wire [31:0] _0532_;
  wire [31:0] _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire [3:0] _0546_;
  wire [3:0] _0547_;
  wire [3:0] _0548_;
  wire [3:0] _0549_;
  wire [3:0] _0550_;
  wire [3:0] _0551_;
  wire [3:0] _0552_;
  wire [3:0] _0553_;
  wire [3:0] _0554_;
  wire [3:0] _0555_;
  wire [3:0] _0556_;
  wire [3:0] _0557_;
  wire [31:0] _0558_;
  wire [31:0] _0559_;
  wire [31:0] _0560_;
  wire [31:0] _0561_;
  wire [31:0] _0562_;
  wire [31:0] _0563_;
  wire [31:0] _0564_;
  wire [31:0] _0565_;
  wire [4:0] _0566_;
  wire [4:0] _0567_;
  wire [4:0] _0568_;
  wire [4:0] _0569_;
  wire [4:0] _0570_;
  wire [4:0] _0571_;
  wire [4:0] _0572_;
  wire [4:0] _0573_;
  wire [4:0] _0574_;
  wire [4:0] _0575_;
  wire [4:0] _0576_;
  wire [4:0] _0577_;
  wire [4:0] _0578_;
  wire [4:0] _0579_;
  wire [4:0] _0580_;
  wire [4:0] _0581_;
  wire [4:0] _0582_;
  wire [4:0] _0583_;
  wire [4:0] _0584_;
  wire [4:0] _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire [4:0] _0601_;
  wire [4:0] _0602_;
  wire [4:0] _0603_;
  wire [4:0] _0604_;
  wire [4:0] _0605_;
  wire [4:0] _0606_;
  wire [4:0] _0607_;
  wire [4:0] _0608_;
  wire [4:0] _0609_;
  wire [4:0] _0610_;
  wire [4:0] _0611_;
  wire [4:0] _0612_;
  wire [4:0] _0613_;
  wire [4:0] _0614_;
  wire [4:0] _0615_;
  wire [4:0] _0616_;
  wire [4:0] _0617_;
  wire [4:0] _0618_;
  wire [4:0] _0619_;
  wire [4:0] _0620_;
  wire [2:0] _0621_;
  wire [2:0] _0622_;
  wire [2:0] _0623_;
  wire [2:0] _0624_;
  wire [2:0] _0625_;
  wire [2:0] _0626_;
  wire [2:0] _0627_;
  wire [2:0] _0628_;
  wire [2:0] _0629_;
  wire [2:0] _0630_;
  wire [2:0] _0631_;
  wire [2:0] _0632_;
  wire [3:0] _0633_;
  wire [3:0] _0634_;
  wire [3:0] _0635_;
  wire [3:0] _0636_;
  wire [3:0] _0637_;
  wire [3:0] _0638_;
  wire [5:0] _0639_;
  wire [5:0] _0640_;
  wire [5:0] _0641_;
  wire [5:0] _0642_;
  wire [5:0] _0643_;
  wire [5:0] _0644_;
  wire [5:0] _0645_;
  wire [5:0] _0646_;
  wire [5:0] _0647_;
  wire [5:0] _0648_;
  wire [5:0] _0649_;
  wire [5:0] _0650_;
  wire [5:0] _0651_;
  wire [5:0] _0652_;
  wire [5:0] _0653_;
  wire [5:0] _0654_;
  wire [5:0] _0655_;
  wire [5:0] _0656_;
  wire [5:0] _0657_;
  wire [5:0] _0658_;
  wire [5:0] _0659_;
  wire [5:0] _0660_;
  wire [5:0] _0661_;
  wire [31:0] _0662_;
  wire [31:0] _0663_;
  wire [31:0] _0664_;
  wire [31:0] _0665_;
  wire [31:0] _0666_;
  wire [31:0] _0667_;
  wire [31:0] _0668_;
  wire [31:0] _0669_;
  wire [31:0] _0670_;
  wire [31:0] _0671_;
  wire [31:0] _0672_;
  wire [31:0] _0673_;
  wire [31:0] _0674_;
  wire [31:0] _0675_;
  wire [31:0] _0676_;
  wire [31:0] _0677_;
  wire [31:0] _0678_;
  wire [31:0] _0679_;
  wire [31:0] _0680_;
  wire [31:0] _0681_;
  wire [31:0] _0682_;
  wire [31:0] _0683_;
  wire [31:0] _0684_;
  wire [31:0] _0685_;
  wire [31:0] _0686_;
  wire [31:0] _0687_;
  wire [31:0] _0688_;
  wire [31:0] _0689_;
  wire [31:0] _0690_;
  wire [31:0] _0691_;
  wire [31:0] _0692_;
  wire [31:0] _0693_;
  wire [31:0] _0694_;
  wire [31:0] _0695_;
  wire [31:0] _0696_;
  wire [31:0] _0697_;
  wire [31:0] _0698_;
  wire [31:0] _0699_;
  wire [31:0] _0700_;
  wire [31:0] _0701_;
  wire [31:0] _0702_;
  wire [31:0] _0703_;
  wire [31:0] _0704_;
  wire [31:0] _0705_;
  wire [31:0] _0706_;
  wire [31:0] _0707_;
  wire [31:0] _0708_;
  wire [31:0] _0709_;
  wire [31:0] _0710_;
  wire [31:0] _0711_;
  wire [31:0] _0712_;
  wire [31:0] _0713_;
  wire [31:0] _0714_;
  wire [31:0] _0715_;
  wire [31:0] _0716_;
  wire [31:0] _0717_;
  wire [31:0] _0718_;
  wire [31:0] _0719_;
  wire [31:0] _0720_;
  wire [31:0] _0721_;
  wire [31:0] _0722_;
  wire [31:0] _0723_;
  wire [31:0] _0724_;
  wire [31:0] _0725_;
  wire [31:0] _0726_;
  wire [31:0] _0727_;
  wire [31:0] _0728_;
  wire [31:0] _0729_;
  wire [31:0] _0730_;
  wire [31:0] _0731_;
  wire [31:0] _0732_;
  wire [31:0] _0733_;
  wire [31:0] _0734_;
  wire [31:0] _0735_;
  wire [31:0] _0736_;
  wire [31:0] _0737_;
  wire [31:0] _0738_;
  wire [31:0] _0739_;
  wire [31:0] _0740_;
  wire [31:0] _0741_;
  wire [31:0] _0742_;
  wire [31:0] _0743_;
  wire [31:0] _0744_;
  wire [31:0] _0745_;
  wire [31:0] _0746_;
  wire [31:0] _0747_;
  wire [31:0] _0748_;
  wire [31:0] _0749_;
  wire [31:0] _0750_;
  wire [31:0] _0751_;
  wire [31:0] _0752_;
  wire [31:0] _0753_;
  wire [31:0] _0754_;
  wire [31:0] _0755_;
  wire [31:0] _0756_;
  wire [31:0] _0757_;
  wire [31:0] _0758_;
  wire [31:0] _0759_;
  wire [31:0] _0760_;
  wire [31:0] _0761_;
  wire [31:0] _0762_;
  wire [31:0] _0763_;
  wire [31:0] _0764_;
  wire [31:0] _0765_;
  wire [31:0] _0766_;
  wire [31:0] _0767_;
  wire [31:0] _0768_;
  wire [31:0] _0769_;
  wire [31:0] _0770_;
  wire [31:0] _0771_;
  wire [31:0] _0772_;
  wire [31:0] _0773_;
  wire [31:0] _0774_;
  wire [31:0] _0775_;
  wire [31:0] _0776_;
  wire [31:0] _0777_;
  wire [31:0] _0778_;
  wire [31:0] _0779_;
  wire [31:0] _0780_;
  wire [31:0] _0781_;
  wire [31:0] _0782_;
  wire [31:0] _0783_;
  wire [31:0] _0784_;
  wire [31:0] _0785_;
  wire [31:0] _0786_;
  wire [31:0] _0787_;
  wire [31:0] _0788_;
  wire [31:0] _0789_;
  wire [31:0] _0790_;
  wire [31:0] _0791_;
  wire [31:0] _0792_;
  wire [31:0] _0793_;
  wire [31:0] _0794_;
  wire [31:0] _0795_;
  wire [31:0] _0796_;
  wire [31:0] _0797_;
  wire [31:0] _0798_;
  wire [31:0] _0799_;
  wire [31:0] _0800_;
  wire [31:0] _0801_;
  wire [31:0] _0802_;
  wire [31:0] _0803_;
  wire [31:0] _0804_;
  wire [31:0] _0805_;
  wire [31:0] _0806_;
  wire [31:0] _0807_;
  wire [31:0] _0808_;
  wire [31:0] _0809_;
  wire [31:0] _0810_;
  wire [31:0] _0811_;
  wire [31:0] _0812_;
  wire [31:0] _0813_;
  wire [31:0] _0814_;
  wire [31:0] _0815_;
  wire [31:0] _0816_;
  wire [31:0] _0817_;
  wire [31:0] _0818_;
  wire [31:0] _0819_;
  wire [31:0] _0820_;
  wire [31:0] _0821_;
  wire [31:0] _0822_;
  wire [31:0] _0823_;
  wire [31:0] _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire [2:0] _0841_;
  wire [2:0] _0842_;
  wire _0843_;
  wire _0844_;
  wire [1:0] _0845_;
  wire [1:0] _0846_;
  wire [11:0] _0847_;
  wire [11:0] _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire [3:0] _0853_;
  wire [3:0] _0854_;
  wire [3:0] _0855_;
  wire [3:0] _0856_;
  wire [3:0] _0857_;
  wire [3:0] _0858_;
  wire [3:0] _0859_;
  wire [3:0] _0860_;
  wire [3:0] _0861_;
  wire [3:0] _0862_;
  wire [4:0] _0863_;
  wire [4:0] _0864_;
  wire [4:0] _0865_;
  wire [4:0] _0866_;
  wire [4:0] _0867_;
  wire [4:0] _0868_;
  wire [7:0] _0869_;
  wire [7:0] _0870_;
  wire [4:0] _0871_;
  wire [4:0] _0872_;
  wire [4:0] _0873_;
  wire [4:0] _0874_;
  wire [4:0] _0875_;
  wire [4:0] _0876_;
  wire [4:0] _0877_;
  wire [4:0] _0878_;
  wire [4:0] _0879_;
  wire [4:0] _0880_;
  wire [4:0] _0881_;
  wire [4:0] _0882_;
  wire [31:0] _0883_;
  wire [31:0] _0884_;
  wire [4:0] _0885_;
  wire [4:0] _0886_;
  wire [4:0] _0887_;
  wire [4:0] _0888_;
  wire [31:0] _0889_;
  wire [31:0] _0890_;
  wire [31:0] _0891_;
  wire [31:0] _0892_;
  wire [15:0] _0893_;
  wire [15:0] _0894_;
  wire [3:0] _0895_;
  wire [3:0] _0896_;
  wire [3:0] _0897_;
  wire [3:0] _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire [4:0] _0911_;
  wire [4:0] _0912_;
  wire [4:0] _0913_;
  wire [4:0] _0914_;
  wire [4:0] _0915_;
  wire [4:0] _0916_;
  wire [4:0] _0917_;
  wire [4:0] _0918_;
  wire [4:0] _0919_;
  wire [4:0] _0920_;
  wire [4:0] _0921_;
  wire [4:0] _0922_;
  wire [4:0] _0923_;
  wire [4:0] _0924_;
  wire [4:0] _0925_;
  wire [4:0] _0926_;
  wire [4:0] _0927_;
  wire [4:0] _0928_;
  wire [2:0] _0929_;
  wire [2:0] _0930_;
  wire [2:0] _0931_;
  wire [2:0] _0932_;
  wire [2:0] _0933_;
  wire [2:0] _0934_;
  wire [3:0] _0935_;
  wire [3:0] _0936_;
  wire [3:0] _0937_;
  wire [3:0] _0938_;
  wire [3:0] _0939_;
  wire [3:0] _0940_;
  wire [3:0] _0941_;
  wire [3:0] _0942_;
  wire [3:0] _0943_;
  wire [5:0] _0944_;
  wire [5:0] _0945_;
  wire [5:0] _0946_;
  wire [5:0] _0947_;
  wire [5:0] _0948_;
  wire [5:0] _0949_;
  wire [5:0] _0950_;
  wire [5:0] _0951_;
  wire [63:0] _0952_;
  wire [63:0] _0953_;
  wire [63:0] _0954_;
  wire [63:0] _0955_;
  wire [31:0] _0956_;
  wire [31:0] _0957_;
  wire [31:0] _0958_;
  wire [31:0] _0959_;
  wire [31:0] _0960_;
  wire [31:0] _0961_;
  wire [31:0] _0962_;
  wire [31:0] _0963_;
  wire [31:0] _0964_;
  wire [31:0] _0965_;
  wire [31:0] _0966_;
  wire [31:0] _0967_;
  wire [31:0] _0968_;
  wire [31:0] _0969_;
  wire [31:0] _0970_;
  wire [31:0] _0971_;
  wire [31:0] _0972_;
  wire [31:0] _0973_;
  wire [31:0] _0974_;
  wire [31:0] _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire [31:0] _1024_;
  wire [31:0] _1025_;
  wire [63:0] _1026_;
  wire [31:0] _1027_;
  wire [31:0] _1028_;
  wire [63:0] _1029_;
  wire [31:0] _1030_;
  wire [31:0] _1031_;
  wire [63:0] _1032_;
  wire [29:0] _1033_;
  wire [31:0] _1034_;
  wire [31:0] _1035_;
  wire [31:0] _1036_;
  wire [31:0] _1037_;
  wire [6:0] _1038_;
  wire [6:0] _1039_;
  wire [31:0] _1040_;
  wire [31:0] _1041_;
  wire [15:0] _1042_;
  wire [15:0] _1043_;
  wire [3:0] _1044_;
  wire [3:0] _1045_;
  wire _1046_;
  wire [31:0] _1047_;
  wire [31:0] _1048_;
  wire [31:0] _1049_;
  wire [31:0] _1050_;
  wire _1051_;
  wire [4:0] _1052_;
  wire [4:0] _1053_;
  wire [4:0] _1054_;
  wire [4:0] _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire [2:0] _1062_;
  wire [2:0] _1063_;
  wire _1064_;
  wire _1065_;
  wire [1:0] _1066_;
  wire [1:0] _1067_;
  wire [11:0] _1068_;
  wire [11:0] _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire [7:0] _1074_;
  wire [7:0] _1075_;
  wire [31:0] _1076_;
  wire [31:0] _1077_;
  wire [4:0] _1078_;
  wire [31:0] _1079_;
  wire [31:0] _1080_;
  wire [31:0] _1081_;
  wire [31:0] _1082_;
  wire _1083_;
  wire _1084_;
  wire [3:0] _1085_;
  wire [3:0] _1086_;
  wire [4:0] _1087_;
  wire [4:0] _1088_;
  wire [31:0] _1089_;
  wire [31:0] _1090_;
  wire [4:0] _1091_;
  wire [4:0] _1092_;
  wire [31:0] _1093_;
  wire [31:0] _1094_;
  wire [31:0] _1095_;
  wire [31:0] _1096_;
  wire [3:0] _1097_;
  wire [3:0] _1098_;
  wire [3:0] _1099_;
  wire [31:0] _1100_;
  wire [31:0] _1101_;
  wire _1102_;
  wire _1103_;
  wire [30:0] _1104_;
  wire [30:0] _1105_;
  wire [31:0] _1106_;
  wire [31:0] _1107_;
  wire [31:0] _1108_;
  wire [31:0] _1109_;
  wire [31:0] _1110_;
  wire [31:0] _1111_;
  wire [4:0] _1112_;
  wire [4:0] _1113_;
  wire [7:0] _1114_;
  wire [7:0] _1115_;
  wire [63:0] _1116_;
  wire [63:0] _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire [30:0] _1121_;
  wire [30:0] _1122_;
  wire [31:0] _1123_;
  wire [31:0] _1124_;
  wire [31:0] _1125_;
  wire [31:0] _1126_;
  wire [31:0] _1127_;
  wire [31:0] _1128_;
  wire [31:0] _1129_;
  wire [31:0] _1130_;
  wire [31:0] _1131_;
  wire [31:0] _1132_;
  wire [31:0] _1133_;
  wire [31:0] _1134_;
  wire [31:0] _1135_;
  wire [31:0] _1136_;
  wire [31:0] _1137_;
  wire [31:0] _1138_;
  wire [31:0] _1139_;
  wire [31:0] _1140_;
  wire [31:0] _1141_;
  wire [31:0] _1142_;
  wire [31:0] _1143_;
  wire [31:0] _1144_;
  wire [31:0] _1145_;
  wire [31:0] _1146_;
  wire [31:0] _1147_;
  wire [31:0] _1148_;
  wire [31:0] _1149_;
  wire [31:0] _1150_;
  wire [31:0] _1151_;
  wire [31:0] _1152_;
  wire [31:0] _1153_;
  wire [31:0] _1154_;
  wire [31:0] _1155_;
  wire [31:0] _1156_;
  wire [31:0] _1157_;
  wire [31:0] _1158_;
  wire [31:0] _1159_;
  wire [31:0] _1160_;
  wire [31:0] _1161_;
  wire [31:0] _1162_;
  wire [31:0] _1163_;
  wire [31:0] _1164_;
  wire [31:0] _1165_;
  wire [31:0] _1166_;
  wire [31:0] _1167_;
  wire [31:0] _1168_;
  wire [31:0] _1169_;
  wire [31:0] _1170_;
  wire [31:0] _1171_;
  wire [31:0] _1172_;
  wire [31:0] _1173_;
  wire [31:0] _1174_;
  wire [31:0] _1175_;
  wire [31:0] _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire [31:0] _1195_;
  wire [31:0] _1196_;
  wire [63:0] _1197_;
  wire [31:0] _1198_;
  wire [63:0] _1199_;
  wire [31:0] _1200_;
  wire [31:0] _1201_;
  wire [31:0] _1202_;
  wire [31:0] _1203_;
  wire [31:0] _1204_;
  wire [63:0] _1205_;
  wire [29:0] _1206_;
  wire [31:0] _1207_;
  wire [31:0] _1208_;
  wire [31:0] _1209_;
  wire [31:0] _1210_;
  wire [31:0] _1211_;
  wire [6:0] _1212_;
  wire [31:0] _1213_;
  wire [15:0] _1214_;
  wire [3:0] _1215_;
  wire [31:0] _1216_;
  wire [31:0] _1217_;
  wire [4:0] _1218_;
  wire [4:0] _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire [2:0] _1223_;
  wire _1224_;
  wire [1:0] _1225_;
  wire [11:0] _1226_;
  wire _1227_;
  wire _1228_;
  wire [7:0] _1229_;
  wire [31:0] _1230_;
  wire [4:0] _1231_;
  wire [31:0] _1232_;
  wire [31:0] _1233_;
  wire _1234_;
  wire [3:0] _1235_;
  wire [4:0] _1236_;
  wire [31:0] _1237_;
  wire [4:0] _1238_;
  wire [31:0] _1239_;
  wire [31:0] _1240_;
  wire [3:0] _1241_;
  wire [31:0] _1242_;
  wire _1243_;
  wire [30:0] _1244_;
  wire [31:0] _1245_;
  wire [31:0] _1246_;
  wire [31:0] _1247_;
  wire [4:0] _1248_;
  wire [7:0] _1249_;
  wire [63:0] _1250_;
  wire _1251_;
  wire [30:0] _1252_;
  wire [31:0] _1253_;
  wire [31:0] _1254_;
  wire [31:0] _1255_;
  wire [31:0] _1256_;
  wire [31:0] _1257_;
  wire [31:0] _1258_;
  wire [31:0] _1259_;
  wire [31:0] _1260_;
  wire [31:0] _1261_;
  wire [31:0] _1262_;
  wire [31:0] _1263_;
  wire [31:0] _1264_;
  wire [31:0] _1265_;
  wire [31:0] _1266_;
  wire [31:0] _1267_;
  wire [31:0] _1268_;
  wire [31:0] _1269_;
  wire [31:0] _1270_;
  wire [31:0] _1271_;
  wire [31:0] _1272_;
  wire [31:0] _1273_;
  wire [63:0] _1274_;
  wire [31:0] _1275_;
  wire [63:0] _1276_;
  wire [31:0] _1277_;
  wire [31:0] _1278_;
  wire [31:0] _1279_;
  wire [63:0] _1280_;
  wire [29:0] _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire [31:0] _1287_;
  wire [31:0] _1288_;
  wire [31:0] _1289_;
  wire [31:0] _1290_;
  wire [63:0] _1291_;
  wire [63:0] _1292_;
  wire [31:0] _1293_;
  wire [31:0] _1294_;
  wire [63:0] _1295_;
  wire [63:0] _1296_;
  wire [31:0] _1297_;
  wire [31:0] _1298_;
  wire [31:0] _1299_;
  wire [31:0] _1300_;
  wire [31:0] _1301_;
  wire [31:0] _1302_;
  wire [63:0] _1303_;
  wire [63:0] _1304_;
  wire [29:0] _1305_;
  wire [29:0] _1306_;
  wire [31:0] _1307_;
  wire [31:0] _1308_;
  wire [31:0] _1309_;
  wire [31:0] _1310_;
  wire [31:0] _1311_;
  wire [31:0] _1312_;
  wire [4:0] _1313_;
  wire [4:0] _1314_;
  wire _1315_;
  wire _1316_;
  wire [31:0] _1317_;
  /* cellift = 32'd1 */
  wire [31:0] _1318_;
  wire [31:0] _1319_;
  /* cellift = 32'd1 */
  wire [31:0] _1320_;
  wire [31:0] _1321_;
  /* cellift = 32'd1 */
  wire [31:0] _1322_;
  wire [31:0] _1323_;
  /* cellift = 32'd1 */
  wire [31:0] _1324_;
  wire [31:0] _1325_;
  /* cellift = 32'd1 */
  wire [31:0] _1326_;
  wire [31:0] _1327_;
  /* cellift = 32'd1 */
  wire [31:0] _1328_;
  wire [31:0] _1329_;
  /* cellift = 32'd1 */
  wire [31:0] _1330_;
  wire [31:0] _1331_;
  /* cellift = 32'd1 */
  wire [31:0] _1332_;
  wire [31:0] _1333_;
  /* cellift = 32'd1 */
  wire [31:0] _1334_;
  wire [31:0] _1335_;
  /* cellift = 32'd1 */
  wire [31:0] _1336_;
  wire [4:0] _1337_;
  wire [4:0] _1338_;
  wire [4:0] _1339_;
  wire [4:0] _1340_;
  wire [4:0] _1341_;
  /* cellift = 32'd1 */
  wire [4:0] _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire [7:0] _1352_;
  wire [7:0] _1353_;
  wire [7:0] _1354_;
  wire [7:0] _1355_;
  wire [7:0] _1356_;
  wire [7:0] _1357_;
  wire [7:0] _1358_;
  wire [7:0] _1359_;
  wire [7:0] _1360_;
  wire [7:0] _1361_;
  wire [7:0] _1362_;
  wire [7:0] _1363_;
  wire [7:0] _1364_;
  wire [7:0] _1365_;
  wire [7:0] _1366_;
  wire [7:0] _1367_;
  wire _1368_;
  wire _1369_;
  wire [31:0] _1370_;
  /* cellift = 32'd1 */
  wire [31:0] _1371_;
  wire [31:0] _1372_;
  /* cellift = 32'd1 */
  wire [31:0] _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire [1:0] _1386_;
  wire [1:0] _1387_;
  wire [1:0] _1388_;
  wire [1:0] _1389_;
  wire [1:0] _1390_;
  wire [1:0] _1391_;
  wire [31:0] _1392_;
  /* cellift = 32'd1 */
  wire [31:0] _1393_;
  wire [31:0] _1394_;
  /* cellift = 32'd1 */
  wire [31:0] _1395_;
  wire [31:0] _1396_;
  /* cellift = 32'd1 */
  wire [31:0] _1397_;
  wire [31:0] _1398_;
  /* cellift = 32'd1 */
  wire [31:0] _1399_;
  wire [31:0] _1400_;
  /* cellift = 32'd1 */
  wire [31:0] _1401_;
  wire [31:0] _1402_;
  /* cellift = 32'd1 */
  wire [31:0] _1403_;
  wire [31:0] _1404_;
  /* cellift = 32'd1 */
  wire [31:0] _1405_;
  wire [31:0] _1406_;
  /* cellift = 32'd1 */
  wire [31:0] _1407_;
  wire [31:0] _1408_;
  /* cellift = 32'd1 */
  wire [31:0] _1409_;
  wire [31:0] _1410_;
  /* cellift = 32'd1 */
  wire [31:0] _1411_;
  wire [31:0] _1412_;
  /* cellift = 32'd1 */
  wire [31:0] _1413_;
  wire [31:0] _1414_;
  /* cellift = 32'd1 */
  wire [31:0] _1415_;
  wire [31:0] _1416_;
  /* cellift = 32'd1 */
  wire [31:0] _1417_;
  wire [31:0] _1418_;
  /* cellift = 32'd1 */
  wire [31:0] _1419_;
  wire [31:0] _1420_;
  /* cellift = 32'd1 */
  wire [31:0] _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  /* cellift = 32'd1 */
  wire _1427_;
  wire _1428_;
  /* cellift = 32'd1 */
  wire _1429_;
  wire _1430_;
  /* cellift = 32'd1 */
  wire _1431_;
  wire _1432_;
  /* cellift = 32'd1 */
  wire _1433_;
  wire _1434_;
  /* cellift = 32'd1 */
  wire _1435_;
  wire _1436_;
  /* cellift = 32'd1 */
  wire _1437_;
  wire _1438_;
  /* cellift = 32'd1 */
  wire _1439_;
  wire _1440_;
  /* cellift = 32'd1 */
  wire _1441_;
  wire _1442_;
  /* cellift = 32'd1 */
  wire _1443_;
  wire [3:0] _1444_;
  /* cellift = 32'd1 */
  wire [3:0] _1445_;
  wire [3:0] _1446_;
  /* cellift = 32'd1 */
  wire [3:0] _1447_;
  wire [3:0] _1448_;
  /* cellift = 32'd1 */
  wire [3:0] _1449_;
  wire [3:0] _1450_;
  /* cellift = 32'd1 */
  wire [3:0] _1451_;
  wire [3:0] _1452_;
  /* cellift = 32'd1 */
  wire [3:0] _1453_;
  wire [3:0] _1454_;
  /* cellift = 32'd1 */
  wire [3:0] _1455_;
  wire [3:0] _1456_;
  /* cellift = 32'd1 */
  wire [3:0] _1457_;
  wire [3:0] _1458_;
  /* cellift = 32'd1 */
  wire [3:0] _1459_;
  wire [3:0] _1460_;
  /* cellift = 32'd1 */
  wire [3:0] _1461_;
  wire [3:0] _1462_;
  /* cellift = 32'd1 */
  wire [3:0] _1463_;
  wire [3:0] _1464_;
  /* cellift = 32'd1 */
  wire [3:0] _1465_;
  wire [3:0] _1466_;
  wire [3:0] _1467_;
  /* cellift = 32'd1 */
  wire [3:0] _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire [31:0] _1479_;
  /* cellift = 32'd1 */
  wire [31:0] _1480_;
  wire [31:0] _1481_;
  /* cellift = 32'd1 */
  wire [31:0] _1482_;
  wire [31:0] _1483_;
  /* cellift = 32'd1 */
  wire [31:0] _1484_;
  wire [31:0] _1485_;
  /* cellift = 32'd1 */
  wire [31:0] _1486_;
  wire [31:0] _1487_;
  /* cellift = 32'd1 */
  wire [31:0] _1488_;
  wire [4:0] _1489_;
  /* cellift = 32'd1 */
  wire [4:0] _1490_;
  wire [4:0] _1491_;
  /* cellift = 32'd1 */
  wire [4:0] _1492_;
  wire [4:0] _1493_;
  /* cellift = 32'd1 */
  wire [4:0] _1494_;
  wire [4:0] _1495_;
  /* cellift = 32'd1 */
  wire [4:0] _1496_;
  wire [4:0] _1497_;
  /* cellift = 32'd1 */
  wire [4:0] _1498_;
  wire [4:0] _1499_;
  /* cellift = 32'd1 */
  wire [4:0] _1500_;
  wire [4:0] _1501_;
  /* cellift = 32'd1 */
  wire [4:0] _1502_;
  wire [4:0] _1503_;
  /* cellift = 32'd1 */
  wire [4:0] _1504_;
  wire [4:0] _1505_;
  /* cellift = 32'd1 */
  wire [4:0] _1506_;
  wire [4:0] _1507_;
  /* cellift = 32'd1 */
  wire [4:0] _1508_;
  wire [4:0] _1509_;
  /* cellift = 32'd1 */
  wire [4:0] _1510_;
  wire [4:0] _1511_;
  /* cellift = 32'd1 */
  wire [4:0] _1512_;
  wire [4:0] _1513_;
  /* cellift = 32'd1 */
  wire [4:0] _1514_;
  wire [4:0] _1515_;
  wire [4:0] _1516_;
  /* cellift = 32'd1 */
  wire [4:0] _1517_;
  wire [4:0] _1518_;
  /* cellift = 32'd1 */
  wire [4:0] _1519_;
  wire [1:0] _1520_;
  wire [1:0] _1521_;
  wire [1:0] _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  /* cellift = 32'd1 */
  wire _1526_;
  wire _1527_;
  /* cellift = 32'd1 */
  wire _1528_;
  wire _1529_;
  /* cellift = 32'd1 */
  wire _1530_;
  wire _1531_;
  /* cellift = 32'd1 */
  wire _1532_;
  wire _1533_;
  /* cellift = 32'd1 */
  wire _1534_;
  wire _1535_;
  /* cellift = 32'd1 */
  wire _1536_;
  wire _1537_;
  /* cellift = 32'd1 */
  wire _1538_;
  wire _1539_;
  /* cellift = 32'd1 */
  wire _1540_;
  wire _1541_;
  /* cellift = 32'd1 */
  wire _1542_;
  wire [4:0] _1543_;
  /* cellift = 32'd1 */
  wire [4:0] _1544_;
  wire [4:0] _1545_;
  /* cellift = 32'd1 */
  wire [4:0] _1546_;
  wire [4:0] _1547_;
  /* cellift = 32'd1 */
  wire [4:0] _1548_;
  wire [4:0] _1549_;
  /* cellift = 32'd1 */
  wire [4:0] _1550_;
  wire [4:0] _1551_;
  /* cellift = 32'd1 */
  wire [4:0] _1552_;
  wire [4:0] _1553_;
  /* cellift = 32'd1 */
  wire [4:0] _1554_;
  wire [4:0] _1555_;
  /* cellift = 32'd1 */
  wire [4:0] _1556_;
  wire [4:0] _1557_;
  /* cellift = 32'd1 */
  wire [4:0] _1558_;
  wire [4:0] _1559_;
  /* cellift = 32'd1 */
  wire [4:0] _1560_;
  wire [4:0] _1561_;
  /* cellift = 32'd1 */
  wire [4:0] _1562_;
  wire [2:0] _1563_;
  /* cellift = 32'd1 */
  wire [2:0] _1564_;
  wire [2:0] _1565_;
  /* cellift = 32'd1 */
  wire [2:0] _1566_;
  wire [2:0] _1567_;
  /* cellift = 32'd1 */
  wire [2:0] _1568_;
  wire [2:0] _1569_;
  /* cellift = 32'd1 */
  wire [2:0] _1570_;
  wire [2:0] _1571_;
  /* cellift = 32'd1 */
  wire [2:0] _1572_;
  wire [2:0] _1573_;
  /* cellift = 32'd1 */
  wire [2:0] _1574_;
  wire [2:0] _1575_;
  wire [2:0] _1576_;
  /* cellift = 32'd1 */
  wire [2:0] _1577_;
  wire [2:0] _1578_;
  /* cellift = 32'd1 */
  wire [2:0] _1579_;
  wire [2:0] _1580_;
  /* cellift = 32'd1 */
  wire [2:0] _1581_;
  wire [2:0] _1582_;
  wire [2:0] _1583_;
  /* cellift = 32'd1 */
  wire [2:0] _1584_;
  wire [3:0] _1585_;
  /* cellift = 32'd1 */
  wire [3:0] _1586_;
  wire [3:0] _1587_;
  /* cellift = 32'd1 */
  wire [3:0] _1588_;
  wire [3:0] _1589_;
  /* cellift = 32'd1 */
  wire [3:0] _1590_;
  wire [5:0] _1591_;
  /* cellift = 32'd1 */
  wire [5:0] _1592_;
  wire [5:0] _1593_;
  /* cellift = 32'd1 */
  wire [5:0] _1594_;
  wire [5:0] _1595_;
  /* cellift = 32'd1 */
  wire [5:0] _1596_;
  wire [5:0] _1597_;
  /* cellift = 32'd1 */
  wire [5:0] _1598_;
  wire [5:0] _1599_;
  /* cellift = 32'd1 */
  wire [5:0] _1600_;
  wire [5:0] _1601_;
  /* cellift = 32'd1 */
  wire [5:0] _1602_;
  wire [5:0] _1603_;
  /* cellift = 32'd1 */
  wire [5:0] _1604_;
  wire [5:0] _1605_;
  /* cellift = 32'd1 */
  wire [5:0] _1606_;
  wire [5:0] _1607_;
  /* cellift = 32'd1 */
  wire [5:0] _1608_;
  wire [5:0] _1609_;
  /* cellift = 32'd1 */
  wire [5:0] _1610_;
  wire [5:0] _1611_;
  /* cellift = 32'd1 */
  wire [5:0] _1612_;
  wire [5:0] _1613_;
  /* cellift = 32'd1 */
  wire [5:0] _1614_;
  wire [5:0] _1615_;
  /* cellift = 32'd1 */
  wire [5:0] _1616_;
  wire [31:0] _1617_;
  /* cellift = 32'd1 */
  wire [31:0] _1618_;
  wire [31:0] _1619_;
  /* cellift = 32'd1 */
  wire [31:0] _1620_;
  wire [31:0] _1621_;
  /* cellift = 32'd1 */
  wire [31:0] _1622_;
  wire [3:0] _1623_;
  wire [31:0] _1624_;
  /* cellift = 32'd1 */
  wire [31:0] _1625_;
  wire _1626_;
  /* src = "generated/out/vanilla.sv:1050.7-1050.34" */
  wire _1627_;
  /* src = "generated/out/vanilla.sv:1052.7-1052.35" */
  wire _1628_;
  /* src = "generated/out/vanilla.sv:1054.7-1054.36" */
  wire _1629_;
  /* src = "generated/out/vanilla.sv:1056.7-1056.36" */
  wire _1630_;
  /* src = "generated/out/vanilla.sv:1058.7-1058.34" */
  wire _1631_;
  /* src = "generated/out/vanilla.sv:1060.7-1060.35" */
  wire _1632_;
  /* src = "generated/out/vanilla.sv:1062.7-1062.35" */
  wire _1633_;
  /* src = "generated/out/vanilla.sv:1064.7-1064.35" */
  wire _1634_;
  /* src = "generated/out/vanilla.sv:1579.10-1579.21" */
  wire _1635_;
  /* src = "generated/out/vanilla.sv:1669.9-1669.26" */
  wire _1636_;
  /* src = "generated/out/vanilla.sv:1674.9-1674.26" */
  wire _1637_;
  /* src = "generated/out/vanilla.sv:1792.23-1792.51" */
  wire _1638_;
  /* src = "generated/out/vanilla.sv:1792.58-1792.84" */
  wire _1639_;
  /* src = "generated/out/vanilla.sv:1793.8-1793.35" */
  wire _1640_;
  /* src = "generated/out/vanilla.sv:1797.8-1797.35" */
  wire _1641_;
  /* src = "generated/out/vanilla.sv:1801.8-1801.35" */
  wire _1642_;
  /* src = "generated/out/vanilla.sv:1805.8-1805.35" */
  wire _1643_;
  /* src = "generated/out/vanilla.sv:372.12-372.40" */
  wire _1644_;
  /* src = "generated/out/vanilla.sv:379.12-379.45" */
  wire _1645_;
  /* src = "generated/out/vanilla.sv:383.12-383.45" */
  wire _1646_;
  /* src = "generated/out/vanilla.sv:387.12-387.45" */
  wire _1647_;
  /* src = "generated/out/vanilla.sv:391.12-391.46" */
  wire _1648_;
  /* src = "generated/out/vanilla.sv:392.13-392.44" */
  wire _1649_;
  /* src = "generated/out/vanilla.sv:394.13-394.44" */
  wire _1650_;
  /* src = "generated/out/vanilla.sv:396.13-396.44" */
  wire _1651_;
  /* src = "generated/out/vanilla.sv:398.13-398.44" */
  wire _1652_;
  /* src = "generated/out/vanilla.sv:423.45-423.72" */
  wire _1653_;
  /* src = "generated/out/vanilla.sv:457.9-457.23" */
  wire _1654_;
  /* src = "generated/out/vanilla.sv:457.29-457.43" */
  wire _1655_;
  /* src = "generated/out/vanilla.sv:797.17-797.53" */
  wire _1656_;
  /* src = "generated/out/vanilla.sv:798.19-798.55" */
  wire _1657_;
  /* src = "generated/out/vanilla.sv:799.17-799.53" */
  wire _1658_;
  /* src = "generated/out/vanilla.sv:800.19-800.55" */
  wire _1659_;
  /* src = "generated/out/vanilla.sv:800.61-800.95" */
  wire _1660_;
  /* src = "generated/out/vanilla.sv:803.36-803.72" */
  wire _1661_;
  /* src = "generated/out/vanilla.sv:804.27-804.63" */
  wire _1662_;
  /* src = "generated/out/vanilla.sv:805.19-805.55" */
  wire _1663_;
  /* src = "generated/out/vanilla.sv:806.22-806.58" */
  wire _1664_;
  /* src = "generated/out/vanilla.sv:807.22-807.58" */
  wire _1665_;
  /* src = "generated/out/vanilla.sv:951.50-951.78" */
  wire _1666_;
  /* src = "generated/out/vanilla.sv:952.50-952.78" */
  wire _1667_;
  /* src = "generated/out/vanilla.sv:953.50-953.78" */
  wire _1668_;
  /* src = "generated/out/vanilla.sv:954.50-954.78" */
  wire _1669_;
  /* src = "generated/out/vanilla.sv:955.51-955.79" */
  wire _1670_;
  /* src = "generated/out/vanilla.sv:956.51-956.79" */
  wire _1671_;
  /* src = "generated/out/vanilla.sv:959.40-959.68" */
  wire _1672_;
  /* src = "generated/out/vanilla.sv:967.38-967.66" */
  wire _1673_;
  /* src = "generated/out/vanilla.sv:971.73-971.105" */
  wire _1674_;
  /* src = "generated/out/vanilla.sv:973.73-973.105" */
  wire _1675_;
  /* src = "generated/out/vanilla.sv:984.25-984.55" */
  wire _1676_;
  /* src = "generated/out/vanilla.sv:984.61-984.97" */
  wire _1677_;
  /* src = "generated/out/vanilla.sv:984.174-984.210" */
  wire _1678_;
  /* src = "generated/out/vanilla.sv:985.63-985.99" */
  wire _1679_;
  /* src = "generated/out/vanilla.sv:985.176-985.212" */
  wire _1680_;
  /* src = "generated/out/vanilla.sv:986.60-986.96" */
  wire _1681_;
  /* src = "generated/out/vanilla.sv:987.62-987.98" */
  wire _1682_;
  /* src = "generated/out/vanilla.sv:988.131-988.160" */
  wire _1683_;
  /* src = "generated/out/vanilla.sv:989.20-989.50" */
  wire _1684_;
  /* src = "generated/out/vanilla.sv:1584.35-1584.46" */
  wire _1685_;
  /* src = "generated/out/vanilla.sv:1080.20-1080.51" */
  wire _1686_;
  /* src = "generated/out/vanilla.sv:1166.5-1166.37" */
  wire _1687_;
  /* src = "generated/out/vanilla.sv:1181.8-1181.31" */
  wire _1688_;
  /* src = "generated/out/vanilla.sv:1181.7-1181.46" */
  wire _1689_;
  /* src = "generated/out/vanilla.sv:1214.9-1214.29" */
  wire _1690_;
  /* src = "generated/out/vanilla.sv:1214.8-1214.48" */
  wire _1691_;
  /* src = "generated/out/vanilla.sv:1234.22-1234.46" */
  wire _1692_;
  /* src = "generated/out/vanilla.sv:1275.22-1275.53" */
  wire _1693_;
  /* src = "generated/out/vanilla.sv:1346.27-1346.55" */
  wire _1694_;
  /* src = "generated/out/vanilla.sv:1374.19-1374.72" */
  wire _1695_;
  /* src = "generated/out/vanilla.sv:1454.7-1454.41" */
  wire _1696_;
  /* src = "generated/out/vanilla.sv:1621.11-1621.39" */
  wire _1697_;
  /* src = "generated/out/vanilla.sv:1668.7-1668.67" */
  wire _1698_;
  /* src = "generated/out/vanilla.sv:1669.8-1669.50" */
  wire _1699_;
  /* src = "generated/out/vanilla.sv:1674.8-1674.48" */
  wire _1700_;
  /* src = "generated/out/vanilla.sv:1680.8-1680.50" */
  wire _1701_;
  /* src = "generated/out/vanilla.sv:1680.7-1680.98" */
  wire _1702_;
  /* src = "generated/out/vanilla.sv:1715.18-1715.54" */
  wire _1703_;
  /* src = "generated/out/vanilla.sv:1774.13-1774.43" */
  wire _1704_;
  /* src = "generated/out/vanilla.sv:1792.8-1792.52" */
  wire _1705_;
  /* src = "generated/out/vanilla.sv:1792.7-1792.85" */
  wire _1706_;
  /* src = "generated/out/vanilla.sv:286.28-286.79" */
  wire _1707_;
  /* src = "generated/out/vanilla.sv:286.27-286.94" */
  wire _1708_;
  /* src = "generated/out/vanilla.sv:293.42-293.102" */
  wire _1709_;
  /* src = "generated/out/vanilla.sv:294.49-294.96" */
  wire _1710_;
  /* src = "generated/out/vanilla.sv:296.32-296.54" */
  wire _1711_;
  /* src = "generated/out/vanilla.sv:296.31-296.107" */
  wire _1712_;
  /* src = "generated/out/vanilla.sv:296.113-296.139" */
  wire _1713_;
  /* src = "generated/out/vanilla.sv:296.19-296.141" */
  wire _1714_;
  /* src = "generated/out/vanilla.sv:296.169-296.205" */
  wire _1715_;
  /* src = "generated/out/vanilla.sv:297.25-297.45" */
  wire _1716_;
  /* src = "generated/out/vanilla.sv:298.36-298.82" */
  wire _1717_;
  /* src = "generated/out/vanilla.sv:298.35-298.138" */
  wire _1718_;
  /* src = "generated/out/vanilla.sv:298.145-298.260" */
  wire _1719_;
  /* src = "generated/out/vanilla.sv:298.144-298.288" */
  wire _1720_;
  /* src = "generated/out/vanilla.sv:310.22-310.45" */
  wire _1721_;
  /* src = "generated/out/vanilla.sv:344.7-344.72" */
  wire _1722_;
  /* src = "generated/out/vanilla.sv:423.12-423.73" */
  wire _1723_;
  /* src = "generated/out/vanilla.sv:427.12-427.73" */
  wire _1724_;
  /* src = "generated/out/vanilla.sv:431.13-431.75" */
  wire _1725_;
  /* src = "generated/out/vanilla.sv:431.12-431.109" */
  wire _1726_;
  /* src = "generated/out/vanilla.sv:435.12-435.73" */
  wire _1727_;
  /* src = "generated/out/vanilla.sv:800.18-800.96" */
  wire _1728_;
  /* src = "generated/out/vanilla.sv:817.8-817.59" */
  wire _1729_;
  /* src = "generated/out/vanilla.sv:871.13-871.61" */
  wire _1730_;
  /* src = "generated/out/vanilla.sv:917.14-917.76" */
  wire _1731_;
  /* src = "generated/out/vanilla.sv:917.13-917.110" */
  wire _1732_;
  /* src = "generated/out/vanilla.sv:949.7-949.49" */
  wire _1733_;
  /* src = "generated/out/vanilla.sv:951.17-951.79" */
  wire _1734_;
  /* src = "generated/out/vanilla.sv:952.17-952.79" */
  wire _1735_;
  /* src = "generated/out/vanilla.sv:953.17-953.79" */
  wire _1736_;
  /* src = "generated/out/vanilla.sv:954.17-954.79" */
  wire _1737_;
  /* src = "generated/out/vanilla.sv:955.18-955.80" */
  wire _1738_;
  /* src = "generated/out/vanilla.sv:956.18-956.80" */
  wire _1739_;
  /* src = "generated/out/vanilla.sv:957.16-957.69" */
  wire _1740_;
  /* src = "generated/out/vanilla.sv:958.16-958.69" */
  wire _1741_;
  /* src = "generated/out/vanilla.sv:959.16-959.69" */
  wire _1742_;
  /* src = "generated/out/vanilla.sv:960.17-960.70" */
  wire _1743_;
  /* src = "generated/out/vanilla.sv:961.17-961.70" */
  wire _1744_;
  /* src = "generated/out/vanilla.sv:962.16-962.61" */
  wire _1745_;
  /* src = "generated/out/vanilla.sv:963.16-963.61" */
  wire _1746_;
  /* src = "generated/out/vanilla.sv:964.16-964.61" */
  wire _1747_;
  /* src = "generated/out/vanilla.sv:965.18-965.66" */
  wire _1748_;
  /* src = "generated/out/vanilla.sv:966.18-966.66" */
  wire _1749_;
  /* src = "generated/out/vanilla.sv:967.19-967.67" */
  wire _1750_;
  /* src = "generated/out/vanilla.sv:968.18-968.66" */
  wire _1751_;
  /* src = "generated/out/vanilla.sv:969.17-969.65" */
  wire _1752_;
  /* src = "generated/out/vanilla.sv:970.18-970.66" */
  wire _1753_;
  /* src = "generated/out/vanilla.sv:971.19-971.67" */
  wire _1754_;
  /* src = "generated/out/vanilla.sv:971.18-971.106" */
  wire _1755_;
  /* src = "generated/out/vanilla.sv:972.19-972.67" */
  wire _1756_;
  /* src = "generated/out/vanilla.sv:972.18-972.106" */
  wire _1757_;
  /* src = "generated/out/vanilla.sv:973.18-973.106" */
  wire _1758_;
  /* src = "generated/out/vanilla.sv:974.18-974.66" */
  wire _1759_;
  /* src = "generated/out/vanilla.sv:974.17-974.105" */
  wire _1760_;
  /* src = "generated/out/vanilla.sv:975.17-975.105" */
  wire _1761_;
  /* src = "generated/out/vanilla.sv:976.18-976.66" */
  wire _1762_;
  /* src = "generated/out/vanilla.sv:976.17-976.105" */
  wire _1763_;
  /* src = "generated/out/vanilla.sv:977.18-977.66" */
  wire _1764_;
  /* src = "generated/out/vanilla.sv:977.17-977.105" */
  wire _1765_;
  /* src = "generated/out/vanilla.sv:978.19-978.67" */
  wire _1766_;
  /* src = "generated/out/vanilla.sv:978.18-978.106" */
  wire _1767_;
  /* src = "generated/out/vanilla.sv:979.18-979.66" */
  wire _1768_;
  /* src = "generated/out/vanilla.sv:979.17-979.105" */
  wire _1769_;
  /* src = "generated/out/vanilla.sv:980.18-980.66" */
  wire _1770_;
  /* src = "generated/out/vanilla.sv:980.17-980.105" */
  wire _1771_;
  /* src = "generated/out/vanilla.sv:981.17-981.105" */
  wire _1772_;
  /* src = "generated/out/vanilla.sv:982.17-982.65" */
  wire _1773_;
  /* src = "generated/out/vanilla.sv:982.16-982.104" */
  wire _1774_;
  /* src = "generated/out/vanilla.sv:983.18-983.66" */
  wire _1775_;
  /* src = "generated/out/vanilla.sv:983.17-983.105" */
  wire _1776_;
  /* src = "generated/out/vanilla.sv:984.24-984.98" */
  wire _1777_;
  /* src = "generated/out/vanilla.sv:984.23-984.130" */
  wire _1778_;
  /* src = "generated/out/vanilla.sv:984.137-984.211" */
  wire _1779_;
  /* src = "generated/out/vanilla.sv:984.136-984.243" */
  wire _1780_;
  /* src = "generated/out/vanilla.sv:984.21-984.264" */
  wire _1781_;
  /* src = "generated/out/vanilla.sv:985.26-985.100" */
  wire _1782_;
  /* src = "generated/out/vanilla.sv:985.25-985.132" */
  wire _1783_;
  /* src = "generated/out/vanilla.sv:985.139-985.213" */
  wire _1784_;
  /* src = "generated/out/vanilla.sv:985.138-985.245" */
  wire _1785_;
  /* src = "generated/out/vanilla.sv:985.23-985.266" */
  wire _1786_;
  /* src = "generated/out/vanilla.sv:986.23-986.97" */
  wire _1787_;
  /* src = "generated/out/vanilla.sv:986.22-986.129" */
  wire _1788_;
  /* src = "generated/out/vanilla.sv:987.25-987.99" */
  wire _1789_;
  /* src = "generated/out/vanilla.sv:987.24-987.131" */
  wire _1790_;
  /* src = "generated/out/vanilla.sv:988.28-988.83" */
  wire _1791_;
  /* src = "generated/out/vanilla.sv:988.27-988.106" */
  wire _1792_;
  /* src = "generated/out/vanilla.sv:989.19-989.74" */
  wire _1793_;
  /* src = "generated/out/vanilla.sv:994.185-994.253" */
  wire _1794_;
  /* src = "generated/out/vanilla.sv:994.115-994.183" */
  wire _1795_;
  /* src = "generated/out/vanilla.sv:994.45-994.113" */
  wire _1796_;
  /* src = "generated/out/vanilla.sv:994.25-994.254" */
  wire _1797_;
  /* src = "generated/out/vanilla.sv:995.60-995.259" */
  wire _1798_;
  /* src = "generated/out/vanilla.sv:996.22-996.251" */
  wire _1799_;
  /* src = "generated/out/vanilla.sv:0.0-0.0" */
  wire _1800_;
  /* src = "generated/out/vanilla.sv:0.0-0.0" */
  wire _1801_;
  /* src = "generated/out/vanilla.sv:1009.7-1009.14" */
  wire _1802_;
  /* src = "generated/out/vanilla.sv:1124.27-1124.34" */
  wire _1803_;
  /* src = "generated/out/vanilla.sv:1125.27-1125.35" */
  wire _1804_;
  /* src = "generated/out/vanilla.sv:1126.28-1126.36" */
  wire _1805_;
  /* src = "generated/out/vanilla.sv:1166.22-1166.37" */
  wire _1806_;
  /* src = "generated/out/vanilla.sv:1214.34-1214.48" */
  wire _1807_;
  /* src = "generated/out/vanilla.sv:1220.20-1220.41" */
  wire _1808_;
  /* src = "generated/out/vanilla.sv:1454.30-1454.41" */
  wire _1809_;
  /* src = "generated/out/vanilla.sv:1606.10-1606.26" */
  wire _1810_;
  /* src = "generated/out/vanilla.sv:286.99-286.117" */
  wire _1811_;
  /* src = "generated/out/vanilla.sv:293.107-293.134" */
  wire _1812_;
  /* src = "generated/out/vanilla.sv:296.147-296.164" */
  wire _1813_;
  /* src = "generated/out/vanilla.sv:297.35-297.45" */
  wire _1814_;
  /* src = "generated/out/vanilla.sv:298.36-298.68" */
  wire _1815_;
  /* src = "generated/out/vanilla.sv:310.35-310.45" */
  wire _1816_;
  /* src = "generated/out/vanilla.sv:871.13-871.35" */
  wire _1817_;
  /* src = "generated/out/vanilla.sv:871.39-871.61" */
  wire _1818_;
  /* src = "generated/out/vanilla.sv:949.26-949.49" */
  wire _1819_;
  /* src = "generated/out/vanilla.sv:988.64-988.83" */
  wire _1820_;
  /* src = "generated/out/vanilla.sv:988.88-988.106" */
  wire _1821_;
  /* src = "generated/out/vanilla.sv:989.55-989.74" */
  wire _1822_;
  /* src = "generated/out/vanilla.sv:1115.25-1115.48" */
  wire _1823_;
  /* src = "generated/out/vanilla.sv:1135.4-1135.27" */
  wire _1824_;
  /* src = "generated/out/vanilla.sv:1136.4-1136.25" */
  wire _1825_;
  /* src = "generated/out/vanilla.sv:1137.4-1137.27" */
  wire _1826_;
  /* src = "generated/out/vanilla.sv:1138.23-1138.46" */
  wire _1827_;
  /* src = "generated/out/vanilla.sv:1139.25-1139.48" */
  wire _1828_;
  /* src = "generated/out/vanilla.sv:1148.8-1148.35" */
  wire _1829_;
  /* src = "generated/out/vanilla.sv:1148.7-1148.47" */
  wire _1830_;
  /* src = "generated/out/vanilla.sv:1606.10-1606.38" */
  wire _1831_;
  /* src = "generated/out/vanilla.sv:1634.9-1634.30" */
  wire _1832_;
  /* src = "generated/out/vanilla.sv:1635.9-1635.30" */
  wire _1833_;
  /* src = "generated/out/vanilla.sv:1668.38-1668.66" */
  wire _1834_;
  /* src = "generated/out/vanilla.sv:1687.7-1687.26" */
  wire _1835_;
  /* src = "generated/out/vanilla.sv:1715.29-1715.53" */
  wire _1836_;
  /* src = "generated/out/vanilla.sv:296.61-296.89" */
  wire _1837_;
  /* src = "generated/out/vanilla.sv:296.60-296.106" */
  wire _1838_;
  /* src = "generated/out/vanilla.sv:296.30-296.140" */
  wire _1839_;
  /* src = "generated/out/vanilla.sv:296.147-296.206" */
  wire _1840_;
  /* src = "generated/out/vanilla.sv:298.88-298.137" */
  wire _1841_;
  /* src = "generated/out/vanilla.sv:298.34-298.289" */
  wire _1842_;
  /* src = "generated/out/vanilla.sv:461.7-461.22" */
  wire _1843_;
  /* src = "generated/out/vanilla.sv:464.8-464.28" */
  wire _1844_;
  /* src = "generated/out/vanilla.sv:470.8-470.35" */
  wire _1845_;
  /* src = "generated/out/vanilla.sv:506.13-506.50" */
  wire _1846_;
  /* src = "generated/out/vanilla.sv:859.13-859.60" */
  wire _1847_;
  /* src = "generated/out/vanilla.sv:988.26-988.162" */
  wire _1848_;
  /* src = "generated/out/vanilla.sv:995.45-995.260" */
  wire _1849_;
  wire [31:0] _1850_;
  /* cellift = 32'd1 */
  wire [31:0] _1851_;
  wire [31:0] _1852_;
  /* cellift = 32'd1 */
  wire [31:0] _1853_;
  wire [31:0] _1854_;
  /* cellift = 32'd1 */
  wire [31:0] _1855_;
  wire [31:0] _1856_;
  /* cellift = 32'd1 */
  wire [31:0] _1857_;
  wire [31:0] _1858_;
  /* cellift = 32'd1 */
  wire [31:0] _1859_;
  wire [31:0] _1860_;
  /* cellift = 32'd1 */
  wire [31:0] _1861_;
  wire [31:0] _1862_;
  /* cellift = 32'd1 */
  wire [31:0] _1863_;
  wire [31:0] _1864_;
  /* cellift = 32'd1 */
  wire [31:0] _1865_;
  wire [31:0] _1866_;
  /* cellift = 32'd1 */
  wire [31:0] _1867_;
  wire [31:0] _1868_;
  /* cellift = 32'd1 */
  wire [31:0] _1869_;
  wire [31:0] _1870_;
  /* cellift = 32'd1 */
  wire [31:0] _1871_;
  wire [31:0] _1872_;
  /* cellift = 32'd1 */
  wire [31:0] _1873_;
  wire [31:0] _1874_;
  /* cellift = 32'd1 */
  wire [31:0] _1875_;
  wire [31:0] _1876_;
  /* cellift = 32'd1 */
  wire [31:0] _1877_;
  wire [31:0] _1878_;
  /* cellift = 32'd1 */
  wire [31:0] _1879_;
  wire [31:0] _1880_;
  /* cellift = 32'd1 */
  wire [31:0] _1881_;
  wire [31:0] _1882_;
  /* cellift = 32'd1 */
  wire [31:0] _1883_;
  wire [31:0] _1884_;
  /* cellift = 32'd1 */
  wire [31:0] _1885_;
  wire [31:0] _1886_;
  /* cellift = 32'd1 */
  wire [31:0] _1887_;
  wire [31:0] _1888_;
  /* cellift = 32'd1 */
  wire [31:0] _1889_;
  wire [31:0] _1890_;
  /* cellift = 32'd1 */
  wire [31:0] _1891_;
  wire [31:0] _1892_;
  /* cellift = 32'd1 */
  wire [31:0] _1893_;
  wire [31:0] _1894_;
  /* cellift = 32'd1 */
  wire [31:0] _1895_;
  wire [31:0] _1896_;
  /* cellift = 32'd1 */
  wire [31:0] _1897_;
  wire [31:0] _1898_;
  /* cellift = 32'd1 */
  wire [31:0] _1899_;
  wire [31:0] _1900_;
  /* cellift = 32'd1 */
  wire [31:0] _1901_;
  wire [31:0] _1902_;
  /* cellift = 32'd1 */
  wire [31:0] _1903_;
  wire [31:0] _1904_;
  /* cellift = 32'd1 */
  wire [31:0] _1905_;
  wire [31:0] _1906_;
  /* cellift = 32'd1 */
  wire [31:0] _1907_;
  wire [31:0] _1908_;
  /* cellift = 32'd1 */
  wire [31:0] _1909_;
  wire [31:0] _1910_;
  /* cellift = 32'd1 */
  wire [31:0] _1911_;
  wire [31:0] _1912_;
  /* cellift = 32'd1 */
  wire [31:0] _1913_;
  wire [31:0] _1914_;
  /* cellift = 32'd1 */
  wire [31:0] _1915_;
  wire [31:0] _1916_;
  /* cellift = 32'd1 */
  wire [31:0] _1917_;
  wire [31:0] _1918_;
  /* cellift = 32'd1 */
  wire [31:0] _1919_;
  wire [31:0] _1920_;
  /* cellift = 32'd1 */
  wire [31:0] _1921_;
  wire [31:0] _1922_;
  /* cellift = 32'd1 */
  wire [31:0] _1923_;
  wire [31:0] _1924_;
  /* cellift = 32'd1 */
  wire [31:0] _1925_;
  wire [31:0] _1926_;
  /* cellift = 32'd1 */
  wire [31:0] _1927_;
  wire [31:0] _1928_;
  /* cellift = 32'd1 */
  wire [31:0] _1929_;
  wire [31:0] _1930_;
  /* cellift = 32'd1 */
  wire [31:0] _1931_;
  wire [31:0] _1932_;
  /* cellift = 32'd1 */
  wire [31:0] _1933_;
  wire [31:0] _1934_;
  /* cellift = 32'd1 */
  wire [31:0] _1935_;
  wire [31:0] _1936_;
  /* cellift = 32'd1 */
  wire [31:0] _1937_;
  wire [31:0] _1938_;
  /* cellift = 32'd1 */
  wire [31:0] _1939_;
  wire [31:0] _1940_;
  /* cellift = 32'd1 */
  wire [31:0] _1941_;
  wire [31:0] _1942_;
  /* cellift = 32'd1 */
  wire [31:0] _1943_;
  wire [31:0] _1944_;
  /* cellift = 32'd1 */
  wire [31:0] _1945_;
  wire [31:0] _1946_;
  /* cellift = 32'd1 */
  wire [31:0] _1947_;
  wire [31:0] _1948_;
  /* cellift = 32'd1 */
  wire [31:0] _1949_;
  wire [31:0] _1950_;
  /* cellift = 32'd1 */
  wire [31:0] _1951_;
  wire [31:0] _1952_;
  /* cellift = 32'd1 */
  wire [31:0] _1953_;
  wire [31:0] _1954_;
  /* cellift = 32'd1 */
  wire [31:0] _1955_;
  wire [31:0] _1956_;
  /* cellift = 32'd1 */
  wire [31:0] _1957_;
  wire [31:0] _1958_;
  /* cellift = 32'd1 */
  wire [31:0] _1959_;
  wire [31:0] _1960_;
  /* cellift = 32'd1 */
  wire [31:0] _1961_;
  wire [31:0] _1962_;
  /* cellift = 32'd1 */
  wire [31:0] _1963_;
  wire [31:0] _1964_;
  /* cellift = 32'd1 */
  wire [31:0] _1965_;
  wire [31:0] _1966_;
  /* cellift = 32'd1 */
  wire [31:0] _1967_;
  wire [31:0] _1968_;
  /* cellift = 32'd1 */
  wire [31:0] _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  /* src = "generated/out/vanilla.sv:1186.33-1186.40" */
  wire [31:0] _2002_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1186.33-1186.40" */
  wire [31:0] _2003_;
  /* src = "generated/out/vanilla.sv:1187.33-1187.40" */
  wire [31:0] _2004_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1187.33-1187.40" */
  wire [31:0] _2005_;
  /* src = "generated/out/vanilla.sv:1669.32-1669.49" */
  wire _2006_;
  /* src = "generated/out/vanilla.sv:427.45-427.72" */
  wire _2007_;
  /* src = "generated/out/vanilla.sv:431.46-431.74" */
  wire _2008_;
  /* src = "generated/out/vanilla.sv:984.104-984.129" */
  wire _2009_;
  /* src = "generated/out/vanilla.sv:1136.37-1136.54" */
  wire [31:0] _2010_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1136.37-1136.54" */
  wire [31:0] _2011_;
  wire _2012_;
  wire _2013_;
  wire [31:0] _2014_;
  /* cellift = 32'd1 */
  wire [31:0] _2015_;
  wire [31:0] _2016_;
  /* cellift = 32'd1 */
  wire [31:0] _2017_;
  wire [3:0] _2018_;
  /* cellift = 32'd1 */
  wire [3:0] _2019_;
  wire [3:0] _2020_;
  wire [31:0] _2021_;
  /* cellift = 32'd1 */
  wire [31:0] _2022_;
  wire [31:0] _2023_;
  wire [31:0] _2024_;
  /* cellift = 32'd1 */
  wire [31:0] _2025_;
  wire _2026_;
  wire [4:0] _2027_;
  wire [4:0] _2028_;
  /* cellift = 32'd1 */
  wire [4:0] _2029_;
  wire [31:0] _2030_;
  /* cellift = 32'd1 */
  wire [31:0] _2031_;
  wire [31:0] _2032_;
  /* cellift = 32'd1 */
  wire [31:0] _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire [31:0] _2039_;
  /* cellift = 32'd1 */
  wire [31:0] _2040_;
  wire [31:0] _2041_;
  /* cellift = 32'd1 */
  wire [31:0] _2042_;
  wire [31:0] _2043_;
  /* cellift = 32'd1 */
  wire [31:0] _2044_;
  wire [31:0] _2045_;
  /* cellift = 32'd1 */
  wire [31:0] _2046_;
  wire [31:0] _2047_;
  /* cellift = 32'd1 */
  wire [31:0] _2048_;
  wire [4:0] _2049_;
  wire [4:0] _2050_;
  wire _2051_;
  wire _2052_;
  wire [4:0] _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire [7:0] _2065_;
  wire [7:0] _2066_;
  wire [7:0] _2067_;
  wire [7:0] _2068_;
  wire [7:0] _2069_;
  wire [7:0] _2070_;
  wire [7:0] _2071_;
  wire [7:0] _2072_;
  wire [7:0] _2073_;
  wire [7:0] _2074_;
  wire [7:0] _2075_;
  wire [7:0] _2076_;
  wire [7:0] _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire [31:0] _2083_;
  /* cellift = 32'd1 */
  wire [31:0] _2084_;
  wire [31:0] _2085_;
  /* cellift = 32'd1 */
  wire [31:0] _2086_;
  wire [31:0] _2087_;
  /* cellift = 32'd1 */
  wire [31:0] _2088_;
  wire [31:0] _2089_;
  /* cellift = 32'd1 */
  wire [31:0] _2090_;
  wire [31:0] _2091_;
  /* cellift = 32'd1 */
  wire [31:0] _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire [1:0] _2098_;
  wire [1:0] _2099_;
  wire [1:0] _2100_;
  wire [1:0] _2101_;
  wire [31:0] _2102_;
  /* cellift = 32'd1 */
  wire [31:0] _2103_;
  wire [31:0] _2104_;
  /* cellift = 32'd1 */
  wire [31:0] _2105_;
  wire [31:0] _2106_;
  /* cellift = 32'd1 */
  wire [31:0] _2107_;
  wire [31:0] _2108_;
  /* cellift = 32'd1 */
  wire [31:0] _2109_;
  wire [31:0] _2110_;
  /* cellift = 32'd1 */
  wire [31:0] _2111_;
  wire [31:0] _2112_;
  /* cellift = 32'd1 */
  wire [31:0] _2113_;
  wire [31:0] _2114_;
  /* cellift = 32'd1 */
  wire [31:0] _2115_;
  wire [31:0] _2116_;
  /* cellift = 32'd1 */
  wire [31:0] _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  /* cellift = 32'd1 */
  wire _2123_;
  wire _2124_;
  /* cellift = 32'd1 */
  wire _2125_;
  wire _2126_;
  /* cellift = 32'd1 */
  wire _2127_;
  wire _2128_;
  /* cellift = 32'd1 */
  wire _2129_;
  wire _2130_;
  wire _2131_;
  /* cellift = 32'd1 */
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  /* cellift = 32'd1 */
  wire _2138_;
  wire _2139_;
  /* cellift = 32'd1 */
  wire _2140_;
  wire _2141_;
  /* cellift = 32'd1 */
  wire _2142_;
  wire _2143_;
  /* cellift = 32'd1 */
  wire _2144_;
  wire _2145_;
  /* cellift = 32'd1 */
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  /* cellift = 32'd1 */
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  /* cellift = 32'd1 */
  wire _2154_;
  wire _2155_;
  /* cellift = 32'd1 */
  wire _2156_;
  wire _2157_;
  /* cellift = 32'd1 */
  wire _2158_;
  wire _2159_;
  /* cellift = 32'd1 */
  wire _2160_;
  wire [2:0] _2161_;
  /* cellift = 32'd1 */
  wire [2:0] _2162_;
  wire _2163_;
  /* cellift = 32'd1 */
  wire _2164_;
  wire [1:0] _2165_;
  /* cellift = 32'd1 */
  wire [1:0] _2166_;
  wire [11:0] _2167_;
  /* cellift = 32'd1 */
  wire [11:0] _2168_;
  wire _2169_;
  /* cellift = 32'd1 */
  wire _2170_;
  wire _2171_;
  /* cellift = 32'd1 */
  wire _2172_;
  wire [3:0] _2173_;
  /* cellift = 32'd1 */
  wire [3:0] _2174_;
  wire [3:0] _2175_;
  /* cellift = 32'd1 */
  wire [3:0] _2176_;
  wire [3:0] _2177_;
  /* cellift = 32'd1 */
  wire [3:0] _2178_;
  wire [3:0] _2179_;
  /* cellift = 32'd1 */
  wire [3:0] _2180_;
  wire [3:0] _2181_;
  wire [3:0] _2182_;
  /* cellift = 32'd1 */
  wire [3:0] _2183_;
  wire [3:0] _2184_;
  /* cellift = 32'd1 */
  wire [3:0] _2185_;
  wire [3:0] _2186_;
  /* cellift = 32'd1 */
  wire [3:0] _2187_;
  wire [3:0] _2188_;
  /* cellift = 32'd1 */
  wire [3:0] _2189_;
  wire [3:0] _2190_;
  /* cellift = 32'd1 */
  wire [3:0] _2191_;
  wire [3:0] _2192_;
  /* cellift = 32'd1 */
  wire [3:0] _2193_;
  wire [3:0] _2194_;
  /* cellift = 32'd1 */
  wire [3:0] _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  wire _2214_;
  wire _2215_;
  wire _2216_;
  wire _2217_;
  wire _2218_;
  wire _2219_;
  wire _2220_;
  wire _2221_;
  wire [4:0] _2222_;
  /* cellift = 32'd1 */
  wire [4:0] _2223_;
  wire [4:0] _2224_;
  /* cellift = 32'd1 */
  wire [4:0] _2225_;
  wire [4:0] _2226_;
  /* cellift = 32'd1 */
  wire [4:0] _2227_;
  wire [4:0] _2228_;
  /* cellift = 32'd1 */
  wire [4:0] _2229_;
  wire [4:0] _2230_;
  /* cellift = 32'd1 */
  wire [4:0] _2231_;
  wire [4:0] _2232_;
  /* cellift = 32'd1 */
  wire [4:0] _2233_;
  wire [4:0] _2234_;
  /* cellift = 32'd1 */
  wire [4:0] _2235_;
  wire [4:0] _2236_;
  /* cellift = 32'd1 */
  wire [4:0] _2237_;
  wire [7:0] _2238_;
  /* cellift = 32'd1 */
  wire [7:0] _2239_;
  wire [4:0] _2240_;
  /* cellift = 32'd1 */
  wire [4:0] _2241_;
  wire [4:0] _2242_;
  /* cellift = 32'd1 */
  wire [4:0] _2243_;
  wire [4:0] _2244_;
  /* cellift = 32'd1 */
  wire [4:0] _2245_;
  wire [4:0] _2246_;
  /* cellift = 32'd1 */
  wire [4:0] _2247_;
  wire [4:0] _2248_;
  /* cellift = 32'd1 */
  wire [4:0] _2249_;
  wire [4:0] _2250_;
  /* cellift = 32'd1 */
  wire [4:0] _2251_;
  wire [4:0] _2252_;
  /* cellift = 32'd1 */
  wire [4:0] _2253_;
  wire [4:0] _2254_;
  /* cellift = 32'd1 */
  wire [4:0] _2255_;
  wire [4:0] _2256_;
  /* cellift = 32'd1 */
  wire [4:0] _2257_;
  wire _2258_;
  wire [4:0] _2259_;
  /* cellift = 32'd1 */
  wire [4:0] _2260_;
  wire [4:0] _2261_;
  /* cellift = 32'd1 */
  wire [4:0] _2262_;
  wire _2263_;
  wire _2264_;
  wire _2265_;
  wire _2266_;
  wire _2267_;
  wire _2268_;
  wire _2269_;
  wire _2270_;
  wire _2271_;
  wire _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire [15:0] _2278_;
  /* cellift = 32'd1 */
  wire [15:0] _2279_;
  wire [15:0] _2280_;
  /* cellift = 32'd1 */
  wire [15:0] _2281_;
  wire [15:0] _2282_;
  /* cellift = 32'd1 */
  wire [15:0] _2283_;
  wire [15:0] _2284_;
  /* cellift = 32'd1 */
  wire [15:0] _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire [1:0] _2289_;
  wire [1:0] _2290_;
  wire [1:0] _2291_;
  wire [1:0] _2292_;
  wire [1:0] _2293_;
  wire [1:0] _2294_;
  wire [1:0] _2295_;
  wire [3:0] _2296_;
  /* cellift = 32'd1 */
  wire [3:0] _2297_;
  wire [3:0] _2298_;
  /* cellift = 32'd1 */
  wire [3:0] _2299_;
  wire [3:0] _2300_;
  /* cellift = 32'd1 */
  wire [3:0] _2301_;
  wire _2302_;
  wire _2303_;
  wire _2304_;
  wire _2305_;
  wire _2306_;
  wire _2307_;
  wire _2308_;
  /* cellift = 32'd1 */
  wire _2309_;
  wire _2310_;
  /* cellift = 32'd1 */
  wire _2311_;
  wire _2312_;
  /* cellift = 32'd1 */
  wire _2313_;
  wire _2314_;
  /* cellift = 32'd1 */
  wire _2315_;
  wire _2316_;
  /* cellift = 32'd1 */
  wire _2317_;
  wire _2318_;
  /* cellift = 32'd1 */
  wire _2319_;
  wire _2320_;
  /* cellift = 32'd1 */
  wire _2321_;
  wire _2322_;
  /* cellift = 32'd1 */
  wire _2323_;
  wire _2324_;
  /* cellift = 32'd1 */
  wire _2325_;
  wire _2326_;
  /* cellift = 32'd1 */
  wire _2327_;
  wire _2328_;
  /* cellift = 32'd1 */
  wire _2329_;
  wire _2330_;
  /* cellift = 32'd1 */
  wire _2331_;
  wire _2332_;
  /* cellift = 32'd1 */
  wire _2333_;
  wire [4:0] _2334_;
  /* cellift = 32'd1 */
  wire [4:0] _2335_;
  wire [4:0] _2336_;
  /* cellift = 32'd1 */
  wire [4:0] _2337_;
  wire [4:0] _2338_;
  /* cellift = 32'd1 */
  wire [4:0] _2339_;
  wire [4:0] _2340_;
  /* cellift = 32'd1 */
  wire [4:0] _2341_;
  wire [4:0] _2342_;
  /* cellift = 32'd1 */
  wire [4:0] _2343_;
  wire [4:0] _2344_;
  /* cellift = 32'd1 */
  wire [4:0] _2345_;
  wire [4:0] _2346_;
  /* cellift = 32'd1 */
  wire [4:0] _2347_;
  wire [4:0] _2348_;
  /* cellift = 32'd1 */
  wire [4:0] _2349_;
  wire [4:0] _2350_;
  /* cellift = 32'd1 */
  wire [4:0] _2351_;
  wire [2:0] _2352_;
  /* cellift = 32'd1 */
  wire [2:0] _2353_;
  wire [2:0] _2354_;
  /* cellift = 32'd1 */
  wire [2:0] _2355_;
  wire [2:0] _2356_;
  /* cellift = 32'd1 */
  wire [2:0] _2357_;
  wire [2:0] _2358_;
  /* cellift = 32'd1 */
  wire [2:0] _2359_;
  wire [2:0] _2360_;
  /* cellift = 32'd1 */
  wire [2:0] _2361_;
  wire [2:0] _2362_;
  /* cellift = 32'd1 */
  wire [2:0] _2363_;
  wire [2:0] _2364_;
  /* cellift = 32'd1 */
  wire [2:0] _2365_;
  wire [2:0] _2366_;
  /* cellift = 32'd1 */
  wire [2:0] _2367_;
  wire [2:0] _2368_;
  /* cellift = 32'd1 */
  wire [2:0] _2369_;
  wire [2:0] _2370_;
  /* cellift = 32'd1 */
  wire [2:0] _2371_;
  wire [2:0] _2372_;
  /* cellift = 32'd1 */
  wire [2:0] _2373_;
  wire [2:0] _2374_;
  /* cellift = 32'd1 */
  wire [2:0] _2375_;
  wire [2:0] _2376_;
  /* cellift = 32'd1 */
  wire [2:0] _2377_;
  wire [2:0] _2378_;
  /* cellift = 32'd1 */
  wire [2:0] _2379_;
  wire [3:0] _2380_;
  /* cellift = 32'd1 */
  wire [3:0] _2381_;
  wire [3:0] _2382_;
  /* cellift = 32'd1 */
  wire [3:0] _2383_;
  wire [3:0] _2384_;
  /* cellift = 32'd1 */
  wire [3:0] _2385_;
  wire [3:0] _2386_;
  /* cellift = 32'd1 */
  wire [3:0] _2387_;
  wire [5:0] _2388_;
  /* cellift = 32'd1 */
  wire [5:0] _2389_;
  wire [5:0] _2390_;
  /* cellift = 32'd1 */
  wire [5:0] _2391_;
  wire [5:0] _2392_;
  /* cellift = 32'd1 */
  wire [5:0] _2393_;
  wire [5:0] _2394_;
  /* cellift = 32'd1 */
  wire [5:0] _2395_;
  wire [5:0] _2396_;
  /* cellift = 32'd1 */
  wire [5:0] _2397_;
  wire [5:0] _2398_;
  /* cellift = 32'd1 */
  wire [5:0] _2399_;
  wire [5:0] _2400_;
  /* cellift = 32'd1 */
  wire [5:0] _2401_;
  wire [5:0] _2402_;
  /* cellift = 32'd1 */
  wire [5:0] _2403_;
  wire [5:0] _2404_;
  /* cellift = 32'd1 */
  wire [5:0] _2405_;
  wire [5:0] _2406_;
  /* cellift = 32'd1 */
  wire [5:0] _2407_;
  wire _2408_;
  wire _2409_;
  wire _2410_;
  wire _2411_;
  wire _2412_;
  /* src = "generated/out/vanilla.sv:296.113-296.123" */
  wire _2413_;
  /* src = "generated/out/vanilla.sv:296.169-296.193" */
  wire _2414_;
  /* src = "generated/out/vanilla.sv:506.13-506.29" */
  wire _2415_;
  /* src = "generated/out/vanilla.sv:1186.19-1186.57" */
  wire _2416_;
  /* src = "generated/out/vanilla.sv:1187.19-1187.57" */
  wire _2417_;
  /* src = "generated/out/vanilla.sv:1746.22-1746.53" */
  wire _2418_;
  /* src = "generated/out/vanilla.sv:1776.24-1776.46" */
  wire _2419_;
  /* src = "generated/out/vanilla.sv:296.44-296.54" */
  wire _2420_;
  /* src = "generated/out/vanilla.sv:795.17-795.96" */
  wire _2421_;
  /* src = "generated/out/vanilla.sv:827.27-827.51" */
  wire _2422_;
  /* src = "generated/out/vanilla.sv:994.43-994.254" */
  wire _2423_;
  /* src = "generated/out/vanilla.sv:995.78-995.259" */
  wire _2424_;
  /* src = "generated/out/vanilla.sv:330.20-330.43" */
  wire [3:0] _2425_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:330.20-330.43" */
  wire [3:0] _2426_;
  /* src = "generated/out/vanilla.sv:1110.32-1110.49" */
  wire [31:0] _2427_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1110.32-1110.49" */
  wire [31:0] _2428_;
  /* src = "generated/out/vanilla.sv:1216.30-1216.54" */
  /* unused_bits = "4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _2429_;
  /* src = "generated/out/vanilla.sv:1591.17-1591.27" */
  /* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _2430_;
  /* src = "generated/out/vanilla.sv:1600.17-1600.27" */
  /* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _2431_;
  /* src = "generated/out/vanilla.sv:1167.24-1167.59" */
  wire [31:0] _2432_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1167.24-1167.59" */
  wire [31:0] _2433_;
  /* src = "generated/out/vanilla.sv:1280.37-1280.109" */
  wire [31:0] _2434_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1280.37-1280.109" */
  wire [31:0] _2435_;
  /* src = "generated/out/vanilla.sv:1405.20-1405.42" */
  wire [31:0] _2436_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1405.20-1405.42" */
  wire [31:0] _2437_;
  /* src = "generated/out/vanilla.sv:1746.22-1746.53" */
  wire [31:0] _2438_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1746.22-1746.53" */
  wire [31:0] _2439_;
  /* src = "generated/out/vanilla.sv:1776.24-1776.46" */
  /* unused_bits = "4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _2440_;
  /* src = "generated/out/vanilla.sv:301.221-301.346" */
  wire [31:0] _2441_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:301.221-301.346" */
  wire [31:0] _2442_;
  /* src = "generated/out/vanilla.sv:301.126-301.347" */
  wire [31:0] _2443_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:301.126-301.347" */
  wire [31:0] _2444_;
  /* src = "generated/out/vanilla.sv:322.21-322.51" */
  wire [3:0] _2445_;
  /* src = "generated/out/vanilla.sv:400.32-400.89" */
  wire [6:0] _2446_;
  /* src = "generated/out/vanilla.sv:512.22-512.58" */
  /* unused_bits = "2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _2447_;
  /* src = "generated/out/vanilla.sv:1135.39-1135.56" */
  wire [31:0] _2448_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1135.39-1135.56" */
  wire [31:0] _2449_;
  /* src = "generated/out/vanilla.sv:1091.13-1091.24" */
  wire [31:0] alu_add_sub;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1091.13-1091.24" */
  wire [31:0] alu_add_sub_t0;
  /* src = "generated/out/vanilla.sv:1094.6-1094.12" */
  wire alu_eq;
  /* src = "generated/out/vanilla.sv:1096.6-1096.13" */
  wire alu_lts;
  /* src = "generated/out/vanilla.sv:1095.6-1095.13" */
  wire alu_ltu;
  /* src = "generated/out/vanilla.sv:1085.13-1085.20" */
  wire [31:0] alu_out;
  /* src = "generated/out/vanilla.sv:1087.6-1087.15" */
  wire alu_out_0;
  /* src = "generated/out/vanilla.sv:1086.13-1086.22" */
  reg [31:0] alu_out_q;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1086.13-1086.22" */
  reg [31:0] alu_out_q_t0;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1085.13-1085.20" */
  wire [31:0] alu_out_t0;
  /* src = "generated/out/vanilla.sv:731.13-731.31" */
  reg [31:0] cached_insn_opcode;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:731.13-731.31" */
  reg [31:0] cached_insn_opcode_t0;
  /* src = "generated/out/vanilla.sv:732.12-732.27" */
  reg [4:0] cached_insn_rs1;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:732.12-732.27" */
  reg [4:0] cached_insn_rs1_t0;
  /* src = "generated/out/vanilla.sv:733.12-733.27" */
  reg [4:0] cached_insn_rs2;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:733.12-733.27" */
  reg [4:0] cached_insn_rs2_t0;
  /* src = "generated/out/vanilla.sv:289.6-289.32" */
  wire clear_prefetched_high_word;
  /* src = "generated/out/vanilla.sv:1142.6-1142.34" */
  reg clear_prefetched_high_word_q;
  /* src = "generated/out/vanilla.sv:85.8-85.11" */
  input clk;
  wire clk;
  /* src = "generated/out/vanilla.sv:593.6-593.22" */
  reg compressed_instr;
  /* src = "generated/out/vanilla.sv:151.13-151.24" */
  reg [63:0] count_cycle;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:151.13-151.24" */
  reg [63:0] count_cycle_t0;
  /* src = "generated/out/vanilla.sv:152.13-152.24" */
  reg [63:0] count_instr;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:152.13-152.24" */
  reg [63:0] count_instr_t0;
  /* src = "generated/out/vanilla.sv:1045.12-1045.21" */
  reg [7:0] cpu_state;
  reg [31:0] \cpuregs[0] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[0]_t0 ;
  reg [31:0] \cpuregs[10] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[10]_t0 ;
  reg [31:0] \cpuregs[11] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[11]_t0 ;
  reg [31:0] \cpuregs[12] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[12]_t0 ;
  reg [31:0] \cpuregs[13] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[13]_t0 ;
  reg [31:0] \cpuregs[14] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[14]_t0 ;
  reg [31:0] \cpuregs[15] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[15]_t0 ;
  reg [31:0] \cpuregs[16] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[16]_t0 ;
  reg [31:0] \cpuregs[17] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[17]_t0 ;
  reg [31:0] \cpuregs[18] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[18]_t0 ;
  reg [31:0] \cpuregs[19] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[19]_t0 ;
  reg [31:0] \cpuregs[1] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[1]_t0 ;
  reg [31:0] \cpuregs[20] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[20]_t0 ;
  reg [31:0] \cpuregs[21] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[21]_t0 ;
  reg [31:0] \cpuregs[22] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[22]_t0 ;
  reg [31:0] \cpuregs[23] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[23]_t0 ;
  reg [31:0] \cpuregs[24] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[24]_t0 ;
  reg [31:0] \cpuregs[25] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[25]_t0 ;
  reg [31:0] \cpuregs[26] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[26]_t0 ;
  reg [31:0] \cpuregs[27] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[27]_t0 ;
  reg [31:0] \cpuregs[28] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[28]_t0 ;
  reg [31:0] \cpuregs[29] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[29]_t0 ;
  reg [31:0] \cpuregs[2] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[2]_t0 ;
  reg [31:0] \cpuregs[30] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[30]_t0 ;
  reg [31:0] \cpuregs[31] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[31]_t0 ;
  reg [31:0] \cpuregs[3] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[3]_t0 ;
  reg [31:0] \cpuregs[4] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[4]_t0 ;
  reg [31:0] \cpuregs[5] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[5]_t0 ;
  reg [31:0] \cpuregs[6] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[6]_t0 ;
  reg [31:0] \cpuregs[7] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[7]_t0 ;
  reg [31:0] \cpuregs[8] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[8]_t0 ;
  reg [31:0] \cpuregs[9] ;
  /* cellift = 32'd1 */
  reg [31:0] \cpuregs[9]_t0 ;
  /* src = "generated/out/vanilla.sv:1153.13-1153.24" */
  wire [31:0] cpuregs_rs1;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1153.13-1153.24" */
  wire [31:0] cpuregs_rs1_t0;
  /* src = "generated/out/vanilla.sv:1154.13-1154.24" */
  wire [31:0] cpuregs_rs2;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1154.13-1154.24" */
  wire [31:0] cpuregs_rs2_t0;
  /* src = "generated/out/vanilla.sv:1152.13-1152.27" */
  wire [31:0] cpuregs_wrdata;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1152.13-1152.27" */
  wire [31:0] cpuregs_wrdata_t0;
  /* src = "generated/out/vanilla.sv:1151.6-1151.19" */
  wire cpuregs_write;
  /* src = "generated/out/vanilla.sv:160.13-160.28" */
  wire [31:0] dbg_insn_opcode;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:160.13-160.28" */
  wire [31:0] dbg_insn_opcode_t0;
  /* src = "generated/out/vanilla.sv:614.12-614.24" */
  wire [4:0] dbg_insn_rs1;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:614.12-614.24" */
  wire [4:0] dbg_insn_rs1_t0;
  /* src = "generated/out/vanilla.sv:615.12-615.24" */
  wire [4:0] dbg_insn_rs2;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:615.12-615.24" */
  wire [4:0] dbg_insn_rs2_t0;
  /* src = "generated/out/vanilla.sv:726.6-726.14" */
  reg dbg_next;
  /* src = "generated/out/vanilla.sv:617.13-617.23" */
  reg [31:0] dbg_rs1val;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:617.13-617.23" */
  reg [31:0] dbg_rs1val_t0;
  /* src = "generated/out/vanilla.sv:619.6-619.22" */
  reg dbg_rs1val_valid;
  /* src = "generated/out/vanilla.sv:618.13-618.23" */
  reg [31:0] dbg_rs2val;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:618.13-618.23" */
  reg [31:0] dbg_rs2val_t0;
  /* src = "generated/out/vanilla.sv:620.6-620.22" */
  reg dbg_rs2val_valid;
  /* src = "generated/out/vanilla.sv:728.6-728.20" */
  reg dbg_valid_insn;
  /* src = "generated/out/vanilla.sv:587.13-587.24" */
  reg [31:0] decoded_imm;
  /* src = "generated/out/vanilla.sv:588.13-588.26" */
  wire [31:0] decoded_imm_j;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:588.13-588.26" */
  wire [31:0] decoded_imm_j_t0;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:587.13-587.24" */
  reg [31:0] decoded_imm_t0;
  /* src = "generated/out/vanilla.sv:584.28-584.38" */
  reg [4:0] decoded_rd;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:584.28-584.38" */
  reg [4:0] decoded_rd_t0;
  /* src = "generated/out/vanilla.sv:585.28-585.39" */
  reg [4:0] decoded_rs1;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:585.28-585.39" */
  reg [4:0] decoded_rs1_t0;
  /* src = "generated/out/vanilla.sv:586.28-586.39" */
  reg [4:0] decoded_rs2;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:586.28-586.39" */
  reg [4:0] decoded_rs2_t0;
  /* src = "generated/out/vanilla.sv:591.6-591.28" */
  reg decoder_pseudo_trigger;
  /* src = "generated/out/vanilla.sv:592.6-592.30" */
  reg decoder_pseudo_trigger_q;
  /* src = "generated/out/vanilla.sv:589.6-589.21" */
  reg decoder_trigger;
  /* src = "generated/out/vanilla.sv:590.6-590.23" */
  reg decoder_trigger_q;
  /* src = "generated/out/vanilla.sv:109.20-109.23" */
  output [31:0] eoi;
  wire [31:0] eoi;
  /* cellift = 32'd1 */
  output [31:0] eoi_t0;
  wire [31:0] eoi_t0;
  /* src = "generated/out/vanilla.sv:561.6-561.15" */
  reg instr_add;
  /* src = "generated/out/vanilla.sv:552.6-552.16" */
  reg instr_addi;
  /* src = "generated/out/vanilla.sv:570.6-570.15" */
  reg instr_and;
  /* src = "generated/out/vanilla.sv:557.6-557.16" */
  reg instr_andi;
  /* src = "generated/out/vanilla.sv:535.6-535.17" */
  reg instr_auipc;
  /* src = "generated/out/vanilla.sv:538.6-538.15" */
  reg instr_beq;
  /* src = "generated/out/vanilla.sv:541.6-541.15" */
  reg instr_bge;
  /* src = "generated/out/vanilla.sv:543.6-543.16" */
  reg instr_bgeu;
  /* src = "generated/out/vanilla.sv:540.6-540.15" */
  reg instr_blt;
  /* src = "generated/out/vanilla.sv:542.6-542.16" */
  reg instr_bltu;
  /* src = "generated/out/vanilla.sv:539.6-539.15" */
  reg instr_bne;
  /* src = "generated/out/vanilla.sv:575.6-575.24" */
  reg instr_ecall_ebreak;
  /* src = "generated/out/vanilla.sv:576.6-576.17" */
  reg instr_fence;
  /* src = "generated/out/vanilla.sv:536.6-536.15" */
  reg instr_jal;
  /* src = "generated/out/vanilla.sv:537.6-537.16" */
  reg instr_jalr;
  /* src = "generated/out/vanilla.sv:544.6-544.14" */
  reg instr_lb;
  /* src = "generated/out/vanilla.sv:547.6-547.15" */
  reg instr_lbu;
  /* src = "generated/out/vanilla.sv:545.6-545.14" */
  reg instr_lh;
  /* src = "generated/out/vanilla.sv:548.6-548.15" */
  reg instr_lhu;
  /* src = "generated/out/vanilla.sv:534.6-534.15" */
  reg instr_lui;
  /* src = "generated/out/vanilla.sv:546.6-546.14" */
  reg instr_lw;
  /* src = "generated/out/vanilla.sv:569.6-569.14" */
  reg instr_or;
  /* src = "generated/out/vanilla.sv:556.6-556.15" */
  reg instr_ori;
  /* src = "generated/out/vanilla.sv:571.6-571.19" */
  reg instr_rdcycle;
  /* src = "generated/out/vanilla.sv:572.6-572.20" */
  reg instr_rdcycleh;
  /* src = "generated/out/vanilla.sv:573.6-573.19" */
  reg instr_rdinstr;
  /* src = "generated/out/vanilla.sv:574.6-574.20" */
  reg instr_rdinstrh;
  /* src = "generated/out/vanilla.sv:549.6-549.14" */
  reg instr_sb;
  /* src = "generated/out/vanilla.sv:550.6-550.14" */
  reg instr_sh;
  /* src = "generated/out/vanilla.sv:563.6-563.15" */
  reg instr_sll;
  /* src = "generated/out/vanilla.sv:558.6-558.16" */
  reg instr_slli;
  /* src = "generated/out/vanilla.sv:564.6-564.15" */
  reg instr_slt;
  /* src = "generated/out/vanilla.sv:553.6-553.16" */
  reg instr_slti;
  /* src = "generated/out/vanilla.sv:554.6-554.17" */
  reg instr_sltiu;
  /* src = "generated/out/vanilla.sv:565.6-565.16" */
  reg instr_sltu;
  /* src = "generated/out/vanilla.sv:568.6-568.15" */
  reg instr_sra;
  /* src = "generated/out/vanilla.sv:560.6-560.16" */
  reg instr_srai;
  /* src = "generated/out/vanilla.sv:567.6-567.15" */
  reg instr_srl;
  /* src = "generated/out/vanilla.sv:559.6-559.16" */
  reg instr_srli;
  /* src = "generated/out/vanilla.sv:562.6-562.15" */
  reg instr_sub;
  /* src = "generated/out/vanilla.sv:551.6-551.14" */
  reg instr_sw;
  /* src = "generated/out/vanilla.sv:583.7-583.17" */
  wire instr_trap;
  /* src = "generated/out/vanilla.sv:566.6-566.15" */
  reg instr_xor;
  /* src = "generated/out/vanilla.sv:555.6-555.16" */
  reg instr_xori;
  /* src = "generated/out/vanilla.sv:108.15-108.18" */
  input [31:0] irq;
  wire [31:0] irq;
  /* cellift = 32'd1 */
  input [31:0] irq_t0;
  wire [31:0] irq_t0;
  /* src = "generated/out/vanilla.sv:605.6-605.20" */
  reg is_alu_reg_imm;
  /* src = "generated/out/vanilla.sv:606.6-606.20" */
  reg is_alu_reg_reg;
  /* src = "generated/out/vanilla.sv:603.6-603.34" */
  reg is_beq_bne_blt_bge_bltu_bgeu;
  /* src = "generated/out/vanilla.sv:607.6-607.16" */
  reg is_compare;
  /* src = "generated/out/vanilla.sv:597.6-597.43" */
  reg is_jalr_addi_slti_sltiu_xori_ori_andi;
  /* src = "generated/out/vanilla.sv:595.6-595.25" */
  reg is_lb_lh_lw_lbu_lhu;
  /* src = "generated/out/vanilla.sv:594.6-594.22" */
  reg is_lui_auipc_jal;
  /* src = "generated/out/vanilla.sv:609.7-609.43" */
  wire is_rdcycle_rdcycleh_rdinstr_rdinstrh;
  /* src = "generated/out/vanilla.sv:598.6-598.17" */
  reg is_sb_sh_sw;
  /* src = "generated/out/vanilla.sv:599.6-599.20" */
  reg is_sll_srl_sra;
  /* src = "generated/out/vanilla.sv:596.6-596.23" */
  reg is_slli_srli_srai;
  /* src = "generated/out/vanilla.sv:601.6-601.21" */
  reg is_slti_blt_slt;
  /* src = "generated/out/vanilla.sv:602.6-602.24" */
  reg is_sltiu_bltu_sltu;
  /* src = "generated/out/vanilla.sv:285.6-285.20" */
  reg last_mem_valid;
  /* src = "generated/out/vanilla.sv:1072.6-1072.20" */
  reg latched_branch;
  /* src = "generated/out/vanilla.sv:1073.6-1073.19" */
  reg latched_compr;
  /* src = "generated/out/vanilla.sv:1077.6-1077.19" */
  reg latched_is_lb;
  /* src = "generated/out/vanilla.sv:1076.6-1076.19" */
  reg latched_is_lh;
  /* src = "generated/out/vanilla.sv:1078.28-1078.38" */
  reg [4:0] latched_rd;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1078.28-1078.38" */
  reg [4:0] latched_rd_t0;
  /* src = "generated/out/vanilla.sv:1071.6-1071.19" */
  reg latched_stalu;
  /* src = "generated/out/vanilla.sv:1070.6-1070.19" */
  reg latched_store;
  /* src = "generated/out/vanilla.sv:727.7-727.23" */
  wire launch_next_insn;
  /* src = "generated/out/vanilla.sv:290.13-290.29" */
  reg [15:0] mem_16bit_buffer;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:290.13-290.29" */
  reg [15:0] mem_16bit_buffer_t0;
  /* src = "generated/out/vanilla.sv:91.20-91.28" */
  output [31:0] mem_addr;
  reg [31:0] mem_addr;
  /* cellift = 32'd1 */
  output [31:0] mem_addr_t0;
  reg [31:0] mem_addr_t0;
  /* src = "generated/out/vanilla.sv:278.6-278.21" */
  reg mem_do_prefetch;
  /* src = "generated/out/vanilla.sv:280.6-280.18" */
  reg mem_do_rdata;
  /* src = "generated/out/vanilla.sv:279.6-279.18" */
  reg mem_do_rinst;
  /* src = "generated/out/vanilla.sv:281.6-281.18" */
  reg mem_do_wdata;
  /* src = "generated/out/vanilla.sv:296.7-296.15" */
  wire mem_done;
  /* src = "generated/out/vanilla.sv:89.13-89.22" */
  output mem_instr;
  reg mem_instr;
  /* cellift = 32'd1 */
  output mem_instr_t0;
  reg mem_instr_t0;
  /* src = "generated/out/vanilla.sv:97.21-97.32" */
  output [31:0] mem_la_addr;
  wire [31:0] mem_la_addr;
  /* cellift = 32'd1 */
  output [31:0] mem_la_addr_t0;
  wire [31:0] mem_la_addr_t0;
  /* src = "generated/out/vanilla.sv:286.7-286.23" */
  wire mem_la_firstword;
  /* src = "generated/out/vanilla.sv:284.6-284.26" */
  reg mem_la_firstword_reg;
  /* src = "generated/out/vanilla.sv:287.7-287.28" */
  wire mem_la_firstword_xfer;
  /* src = "generated/out/vanilla.sv:95.14-95.25" */
  output mem_la_read;
  wire mem_la_read;
  /* cellift = 32'd1 */
  output mem_la_read_t0;
  wire mem_la_read_t0;
  /* src = "generated/out/vanilla.sv:283.6-283.23" */
  reg mem_la_secondword;
  /* src = "generated/out/vanilla.sv:293.7-293.38" */
  wire mem_la_use_prefetched_high_word;
  /* src = "generated/out/vanilla.sv:98.20-98.32" */
  output [31:0] mem_la_wdata;
  wire [31:0] mem_la_wdata;
  /* cellift = 32'd1 */
  output [31:0] mem_la_wdata_t0;
  wire [31:0] mem_la_wdata_t0;
  /* src = "generated/out/vanilla.sv:96.14-96.26" */
  output mem_la_write;
  wire mem_la_write;
  /* cellift = 32'd1 */
  output mem_la_write_t0;
  wire mem_la_write_t0;
  /* src = "generated/out/vanilla.sv:99.19-99.31" */
  output [3:0] mem_la_wstrb;
  wire [3:0] mem_la_wstrb;
  /* cellift = 32'd1 */
  output [3:0] mem_la_wstrb_t0;
  wire [3:0] mem_la_wstrb_t0;
  /* src = "generated/out/vanilla.sv:94.15-94.24" */
  input [31:0] mem_rdata;
  wire [31:0] mem_rdata;
  /* src = "generated/out/vanilla.sv:292.14-292.31" */
  wire [31:0] mem_rdata_latched;
  /* src = "generated/out/vanilla.sv:291.14-291.41" */
  wire [31:0] mem_rdata_latched_noshuffle;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:291.14-291.41" */
  wire [31:0] mem_rdata_latched_noshuffle_t0;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:292.14-292.31" */
  wire [31:0] mem_rdata_latched_t0;
  /* src = "generated/out/vanilla.sv:277.13-277.24" */
  reg [31:0] mem_rdata_q;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:277.13-277.24" */
  reg [31:0] mem_rdata_q_t0;
  /* cellift = 32'd1 */
  input [31:0] mem_rdata_t0;
  wire [31:0] mem_rdata_t0;
  /* src = "generated/out/vanilla.sv:276.13-276.27" */
  wire [31:0] mem_rdata_word;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:276.13-276.27" */
  wire [31:0] mem_rdata_word_t0;
  /* src = "generated/out/vanilla.sv:90.8-90.17" */
  input mem_ready;
  wire mem_ready;
  /* cellift = 32'd1 */
  input mem_ready_t0;
  wire mem_ready_t0;
  /* src = "generated/out/vanilla.sv:274.12-274.21" */
  reg [1:0] mem_state;
  /* src = "generated/out/vanilla.sv:88.13-88.22" */
  output mem_valid;
  reg mem_valid;
  /* cellift = 32'd1 */
  output mem_valid_t0;
  reg mem_valid_t0;
  /* src = "generated/out/vanilla.sv:92.20-92.29" */
  output [31:0] mem_wdata;
  reg [31:0] mem_wdata;
  /* cellift = 32'd1 */
  output [31:0] mem_wdata_t0;
  reg [31:0] mem_wdata_t0;
  /* src = "generated/out/vanilla.sv:275.12-275.24" */
  reg [1:0] mem_wordsize;
  /* src = "generated/out/vanilla.sv:93.19-93.28" */
  output [3:0] mem_wstrb;
  reg [3:0] mem_wstrb;
  /* cellift = 32'd1 */
  output [3:0] mem_wstrb_t0;
  reg [3:0] mem_wstrb_t0;
  /* src = "generated/out/vanilla.sv:282.7-282.15" */
  wire mem_xfer;
  /* src = "generated/out/vanilla.sv:159.13-159.29" */
  reg [31:0] next_insn_opcode;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:159.13-159.29" */
  reg [31:0] next_insn_opcode_t0;
  /* src = "generated/out/vanilla.sv:171.14-171.21" */
  /* unused_bits = "0" */
  wire [31:0] next_pc /* verilator public */;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:171.14-171.21" */
  /* unused_bits = "0" */
  wire [31:0] next_pc_t0 /* verilator public */;
  /* src = "generated/out/vanilla.sv:190.14-190.25" */
  wire [31:0] pcpi_div_rd;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:190.14-190.25" */
  wire [31:0] pcpi_div_rd_t0;
  /* src = "generated/out/vanilla.sv:192.7-192.21" */
  wire pcpi_div_ready;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:192.7-192.21" */
  /* unused_bits = "0" */
  wire pcpi_div_ready_t0;
  /* src = "generated/out/vanilla.sv:191.7-191.20" */
  wire pcpi_div_wait;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:191.7-191.20" */
  /* unused_bits = "0" */
  wire pcpi_div_wait_t0;
  /* src = "generated/out/vanilla.sv:189.7-189.18" */
  wire pcpi_div_wr;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:189.7-189.18" */
  /* unused_bits = "0" */
  wire pcpi_div_wr_t0;
  /* src = "generated/out/vanilla.sv:101.20-101.29" */
  output [31:0] pcpi_insn;
  reg [31:0] pcpi_insn;
  /* cellift = 32'd1 */
  output [31:0] pcpi_insn_t0;
  reg [31:0] pcpi_insn_t0;
  /* src = "generated/out/vanilla.sv:194.13-194.24" */
  wire [31:0] pcpi_int_rd;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:194.13-194.24" */
  wire [31:0] pcpi_int_rd_t0;
  /* src = "generated/out/vanilla.sv:196.6-196.20" */
  wire pcpi_int_ready;
  /* src = "generated/out/vanilla.sv:195.6-195.19" */
  wire pcpi_int_wait;
  /* src = "generated/out/vanilla.sv:193.6-193.17" */
  wire pcpi_int_wr;
  /* src = "generated/out/vanilla.sv:186.14-186.25" */
  wire [31:0] pcpi_mul_rd;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:186.14-186.25" */
  wire [31:0] pcpi_mul_rd_t0;
  /* src = "generated/out/vanilla.sv:188.7-188.21" */
  wire pcpi_mul_ready;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:188.7-188.21" */
  /* unused_bits = "0" */
  wire pcpi_mul_ready_t0;
  /* src = "generated/out/vanilla.sv:187.7-187.20" */
  wire pcpi_mul_wait;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:187.7-187.20" */
  /* unused_bits = "0" */
  wire pcpi_mul_wait_t0;
  /* src = "generated/out/vanilla.sv:185.7-185.18" */
  wire pcpi_mul_wr;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:185.7-185.18" */
  /* unused_bits = "0" */
  wire pcpi_mul_wr_t0;
  /* src = "generated/out/vanilla.sv:105.15-105.22" */
  input [31:0] pcpi_rd;
  wire [31:0] pcpi_rd;
  /* cellift = 32'd1 */
  input [31:0] pcpi_rd_t0;
  wire [31:0] pcpi_rd_t0;
  /* src = "generated/out/vanilla.sv:107.8-107.18" */
  input pcpi_ready;
  wire pcpi_ready;
  /* cellift = 32'd1 */
  input pcpi_ready_t0;
  wire pcpi_ready_t0;
  /* src = "generated/out/vanilla.sv:102.21-102.29" */
  output [31:0] pcpi_rs1;
  reg [31:0] pcpi_rs1;
  /* cellift = 32'd1 */
  output [31:0] pcpi_rs1_t0;
  reg [31:0] pcpi_rs1_t0;
  /* src = "generated/out/vanilla.sv:103.21-103.29" */
  output [31:0] pcpi_rs2;
  reg [31:0] pcpi_rs2;
  /* cellift = 32'd1 */
  output [31:0] pcpi_rs2_t0;
  reg [31:0] pcpi_rs2_t0;
  /* src = "generated/out/vanilla.sv:1082.6-1082.18" */
  reg pcpi_timeout;
  /* src = "generated/out/vanilla.sv:1081.12-1081.32" */
  reg [3:0] pcpi_timeout_counter;
  /* src = "generated/out/vanilla.sv:100.13-100.23" */
  output pcpi_valid;
  reg pcpi_valid;
  /* cellift = 32'd1 */
  output pcpi_valid_t0;
  reg pcpi_valid_t0;
  /* src = "generated/out/vanilla.sv:106.8-106.17" */
  input pcpi_wait;
  wire pcpi_wait;
  /* cellift = 32'd1 */
  input pcpi_wait_t0;
  wire pcpi_wait_t0;
  /* src = "generated/out/vanilla.sv:104.8-104.15" */
  input pcpi_wr;
  wire pcpi_wr;
  /* cellift = 32'd1 */
  input pcpi_wr_t0;
  wire pcpi_wr_t0;
  /* src = "generated/out/vanilla.sv:288.6-288.26" */
  reg prefetched_high_word;
  /* src = "generated/out/vanilla.sv:723.12-723.22" */
  reg [4:0] q_insn_rs1;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:723.12-723.22" */
  reg [4:0] q_insn_rs1_t0;
  /* src = "generated/out/vanilla.sv:724.12-724.22" */
  reg [4:0] q_insn_rs2;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:724.12-724.22" */
  reg [4:0] q_insn_rs2_t0;
  /* src = "generated/out/vanilla.sv:154.13-154.24" */
  reg [31:0] reg_next_pc;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:154.13-154.24" */
  reg [31:0] reg_next_pc_t0;
  /* src = "generated/out/vanilla.sv:157.13-157.20" */
  reg [31:0] reg_out;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:157.13-157.20" */
  reg [31:0] reg_out_t0;
  /* src = "generated/out/vanilla.sv:153.13-153.19" */
  reg [31:0] reg_pc;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:153.13-153.19" */
  reg [31:0] reg_pc_t0;
  /* src = "generated/out/vanilla.sv:158.12-158.18" */
  reg [4:0] reg_sh;
  /* src = "generated/out/vanilla.sv:86.8-86.14" */
  input resetn;
  wire resetn;
  /* src = "generated/out/vanilla.sv:133.20-133.41" */
  output [63:0] rvfi_csr_mcycle_rdata;
  wire [63:0] rvfi_csr_mcycle_rdata;
  /* cellift = 32'd1 */
  output [63:0] rvfi_csr_mcycle_rdata_t0;
  wire [63:0] rvfi_csr_mcycle_rdata_t0;
  /* src = "generated/out/vanilla.sv:131.20-131.41" */
  output [63:0] rvfi_csr_mcycle_rmask;
  wire [63:0] rvfi_csr_mcycle_rmask;
  /* cellift = 32'd1 */
  output [63:0] rvfi_csr_mcycle_rmask_t0;
  wire [63:0] rvfi_csr_mcycle_rmask_t0;
  /* src = "generated/out/vanilla.sv:134.20-134.41" */
  output [63:0] rvfi_csr_mcycle_wdata;
  wire [63:0] rvfi_csr_mcycle_wdata;
  /* cellift = 32'd1 */
  output [63:0] rvfi_csr_mcycle_wdata_t0;
  wire [63:0] rvfi_csr_mcycle_wdata_t0;
  /* src = "generated/out/vanilla.sv:132.20-132.41" */
  output [63:0] rvfi_csr_mcycle_wmask;
  wire [63:0] rvfi_csr_mcycle_wmask;
  /* cellift = 32'd1 */
  output [63:0] rvfi_csr_mcycle_wmask_t0;
  wire [63:0] rvfi_csr_mcycle_wmask_t0;
  /* src = "generated/out/vanilla.sv:137.20-137.43" */
  output [63:0] rvfi_csr_minstret_rdata;
  wire [63:0] rvfi_csr_minstret_rdata;
  /* cellift = 32'd1 */
  output [63:0] rvfi_csr_minstret_rdata_t0;
  wire [63:0] rvfi_csr_minstret_rdata_t0;
  /* src = "generated/out/vanilla.sv:135.20-135.43" */
  output [63:0] rvfi_csr_minstret_rmask;
  wire [63:0] rvfi_csr_minstret_rmask;
  /* cellift = 32'd1 */
  output [63:0] rvfi_csr_minstret_rmask_t0;
  wire [63:0] rvfi_csr_minstret_rmask_t0;
  /* src = "generated/out/vanilla.sv:138.20-138.43" */
  output [63:0] rvfi_csr_minstret_wdata;
  wire [63:0] rvfi_csr_minstret_wdata;
  /* cellift = 32'd1 */
  output [63:0] rvfi_csr_minstret_wdata_t0;
  wire [63:0] rvfi_csr_minstret_wdata_t0;
  /* src = "generated/out/vanilla.sv:136.20-136.43" */
  output [63:0] rvfi_csr_minstret_wmask;
  wire [63:0] rvfi_csr_minstret_wmask;
  /* cellift = 32'd1 */
  output [63:0] rvfi_csr_minstret_wmask_t0;
  wire [63:0] rvfi_csr_minstret_wmask_t0;
  /* src = "generated/out/vanilla.sv:114.13-114.22" */
  output rvfi_halt;
  reg rvfi_halt;
  /* cellift = 32'd1 */
  output rvfi_halt_t0;
  wire rvfi_halt_t0;
  /* src = "generated/out/vanilla.sv:112.20-112.29" */
  output [31:0] rvfi_insn;
  wire [31:0] rvfi_insn;
  /* cellift = 32'd1 */
  output [31:0] rvfi_insn_t0;
  wire [31:0] rvfi_insn_t0;
  /* src = "generated/out/vanilla.sv:115.13-115.22" */
  output rvfi_intr;
  wire rvfi_intr;
  /* cellift = 32'd1 */
  output rvfi_intr_t0;
  wire rvfi_intr_t0;
  /* src = "generated/out/vanilla.sv:117.19-117.27" */
  output [1:0] rvfi_ixl;
  wire [1:0] rvfi_ixl;
  /* cellift = 32'd1 */
  output [1:0] rvfi_ixl_t0;
  wire [1:0] rvfi_ixl_t0;
  /* src = "generated/out/vanilla.sv:126.20-126.33" */
  output [31:0] rvfi_mem_addr;
  reg [31:0] rvfi_mem_addr;
  /* cellift = 32'd1 */
  output [31:0] rvfi_mem_addr_t0;
  reg [31:0] rvfi_mem_addr_t0;
  /* src = "generated/out/vanilla.sv:129.20-129.34" */
  output [31:0] rvfi_mem_rdata;
  reg [31:0] rvfi_mem_rdata;
  /* cellift = 32'd1 */
  output [31:0] rvfi_mem_rdata_t0;
  reg [31:0] rvfi_mem_rdata_t0;
  /* src = "generated/out/vanilla.sv:127.19-127.33" */
  output [3:0] rvfi_mem_rmask;
  reg [3:0] rvfi_mem_rmask;
  /* cellift = 32'd1 */
  output [3:0] rvfi_mem_rmask_t0;
  reg [3:0] rvfi_mem_rmask_t0;
  /* src = "generated/out/vanilla.sv:130.20-130.34" */
  output [31:0] rvfi_mem_wdata;
  reg [31:0] rvfi_mem_wdata;
  /* cellift = 32'd1 */
  output [31:0] rvfi_mem_wdata_t0;
  reg [31:0] rvfi_mem_wdata_t0;
  /* src = "generated/out/vanilla.sv:128.19-128.33" */
  output [3:0] rvfi_mem_wmask;
  reg [3:0] rvfi_mem_wmask;
  /* cellift = 32'd1 */
  output [3:0] rvfi_mem_wmask_t0;
  reg [3:0] rvfi_mem_wmask_t0;
  /* src = "generated/out/vanilla.sv:116.19-116.28" */
  output [1:0] rvfi_mode;
  wire [1:0] rvfi_mode;
  /* cellift = 32'd1 */
  output [1:0] rvfi_mode_t0;
  wire [1:0] rvfi_mode_t0;
  /* src = "generated/out/vanilla.sv:111.20-111.30" */
  output [63:0] rvfi_order;
  reg [63:0] rvfi_order;
  /* cellift = 32'd1 */
  output [63:0] rvfi_order_t0;
  reg [63:0] rvfi_order_t0;
  /* src = "generated/out/vanilla.sv:124.20-124.33" */
  output [31:0] rvfi_pc_rdata;
  reg [31:0] rvfi_pc_rdata;
  /* cellift = 32'd1 */
  output [31:0] rvfi_pc_rdata_t0;
  reg [31:0] rvfi_pc_rdata_t0;
  /* src = "generated/out/vanilla.sv:125.20-125.33" */
  output [31:0] rvfi_pc_wdata;
  reg [31:0] rvfi_pc_wdata;
  /* cellift = 32'd1 */
  output [31:0] rvfi_pc_wdata_t0;
  reg [31:0] rvfi_pc_wdata_t0;
  /* src = "generated/out/vanilla.sv:122.19-122.31" */
  output [4:0] rvfi_rd_addr;
  reg [4:0] rvfi_rd_addr;
  /* cellift = 32'd1 */
  output [4:0] rvfi_rd_addr_t0;
  reg [4:0] rvfi_rd_addr_t0;
  /* src = "generated/out/vanilla.sv:123.20-123.33" */
  output [31:0] rvfi_rd_wdata;
  reg [31:0] rvfi_rd_wdata;
  /* cellift = 32'd1 */
  output [31:0] rvfi_rd_wdata_t0;
  reg [31:0] rvfi_rd_wdata_t0;
  /* src = "generated/out/vanilla.sv:118.19-118.32" */
  output [4:0] rvfi_rs1_addr;
  reg [4:0] rvfi_rs1_addr;
  /* cellift = 32'd1 */
  output [4:0] rvfi_rs1_addr_t0;
  reg [4:0] rvfi_rs1_addr_t0;
  /* src = "generated/out/vanilla.sv:120.20-120.34" */
  output [31:0] rvfi_rs1_rdata;
  reg [31:0] rvfi_rs1_rdata;
  /* cellift = 32'd1 */
  output [31:0] rvfi_rs1_rdata_t0;
  reg [31:0] rvfi_rs1_rdata_t0;
  /* src = "generated/out/vanilla.sv:119.19-119.32" */
  output [4:0] rvfi_rs2_addr;
  reg [4:0] rvfi_rs2_addr;
  /* cellift = 32'd1 */
  output [4:0] rvfi_rs2_addr_t0;
  reg [4:0] rvfi_rs2_addr_t0;
  /* src = "generated/out/vanilla.sv:121.20-121.34" */
  output [31:0] rvfi_rs2_rdata;
  reg [31:0] rvfi_rs2_rdata;
  /* cellift = 32'd1 */
  output [31:0] rvfi_rs2_rdata_t0;
  reg [31:0] rvfi_rs2_rdata_t0;
  /* src = "generated/out/vanilla.sv:113.13-113.22" */
  output rvfi_trap;
  wire rvfi_trap;
  /* cellift = 32'd1 */
  output rvfi_trap_t0;
  wire rvfi_trap_t0;
  /* src = "generated/out/vanilla.sv:110.13-110.23" */
  output rvfi_valid;
  reg rvfi_valid;
  /* cellift = 32'd1 */
  output rvfi_valid_t0;
  wire rvfi_valid_t0;
  /* src = "generated/out/vanilla.sv:140.20-140.30" */
  output [35:0] trace_data;
  wire [35:0] trace_data;
  /* cellift = 32'd1 */
  output [35:0] trace_data_t0;
  wire [35:0] trace_data_t0;
  /* src = "generated/out/vanilla.sv:139.13-139.24" */
  output trace_valid;
  wire trace_valid;
  /* cellift = 32'd1 */
  output trace_valid_t0;
  wire trace_valid_t0;
  /* src = "generated/out/vanilla.sv:87.13-87.17" */
  output trap;
  reg trap;
  /* cellift = 32'd1 */
  output trap_t0;
  wire trap_t0;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME _0064_ */
  always_ff @(posedge clk)
    _0064_ <= _1313_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME _0065_ */
  always_ff @(posedge clk)
    _0065_ <= _1314_;
  assign _0066_ = pcpi_rs1 + /* src = "generated/out/vanilla.sv:1110.52-1110.69" */ pcpi_rs2;
  assign _0068_ = reg_pc + /* src = "generated/out/vanilla.sv:1163.23-1163.55" */ _1025_;
  assign _0070_ = count_cycle + /* src = "generated/out/vanilla.sv:1223.29-1223.44" */ 32'd1;
  assign _0072_ = _0046_ + /* src = "generated/out/vanilla.sv:1331.22-1331.61" */ _1028_;
  assign _0074_ = count_instr + /* src = "generated/out/vanilla.sv:1335.23-1335.38" */ 32'd1;
  assign _0076_ = _0046_ + /* src = "generated/out/vanilla.sv:1341.23-1341.49" */ { decoded_imm_j[31:1], 1'h0 };
  assign _0078_ = reg_pc + /* src = "generated/out/vanilla.sv:1554.17-1554.37" */ decoded_imm;
  assign _0080_ = pcpi_rs1 + /* src = "generated/out/vanilla.sv:1645.19-1645.40" */ decoded_imm;
  assign _0082_ = rvfi_order + /* src = "generated/out/vanilla.sv:1716.27-1716.50" */ rvfi_valid;
  assign _0084_ = next_pc[31:2] + /* src = "generated/out/vanilla.sv:299.59-299.96" */ mem_la_firstword_xfer;
  assign _0086_ = 32'd8 + /* src = "generated/out/vanilla.sv:886.25-886.51" */ mem_rdata_latched[4:2];
  assign _0088_ = 32'd8 + /* src = "generated/out/vanilla.sv:897.24-897.50" */ mem_rdata_latched[9:7];
  assign _0090_ = pcpi_rs1 & /* src = "generated/out/vanilla.sv:1137.39-1137.56" */ pcpi_rs2;
  assign _0094_ = mem_la_wstrb & /* src = "generated/out/vanilla.sv:472.18-472.51" */ { mem_la_write, mem_la_write, mem_la_write, mem_la_write };
  assign _0096_ = ~ pcpi_rs1_t0;
  assign _0097_ = ~ reg_pc_t0;
  assign _0098_ = ~ count_cycle_t0;
  assign _0099_ = ~ _0047_;
  assign _0100_ = ~ count_instr_t0;
  assign _0101_ = ~ rvfi_order_t0;
  assign _0102_ = ~ next_pc_t0[31:2];
  assign _0103_ = ~ pcpi_rs2_t0;
  assign _0104_ = ~ { decoded_imm_j_t0[31:1], 1'h0 };
  assign _0105_ = ~ decoded_imm_t0;
  assign _0106_ = ~ { 29'h00000000, mem_rdata_latched_t0[4:2] };
  assign _0107_ = ~ { 29'h00000000, mem_rdata_latched_t0[9:7] };
  assign _0956_ = pcpi_rs1 & _0096_;
  assign _1024_ = reg_pc & _0097_;
  assign _1026_ = count_cycle & _0098_;
  assign _1027_ = _0046_ & _0099_;
  assign _1029_ = count_instr & _0100_;
  assign _1032_ = rvfi_order & _0101_;
  assign _1033_ = next_pc[31:2] & _0102_;
  assign _0957_ = pcpi_rs2 & _0103_;
  assign _1030_ = { decoded_imm_j[31:1], 1'h0 } & _0104_;
  assign _1031_ = decoded_imm & _0105_;
  assign _1034_ = { 29'h00000000, mem_rdata_latched[4:2] } & _0106_;
  assign _1035_ = { 29'h00000000, mem_rdata_latched[9:7] } & _0107_;
  assign _1287_ = _0956_ + _0957_;
  assign _1289_ = _1024_ + _1025_;
  assign _1291_ = _1026_ + 64'h0000000000000001;
  assign _1293_ = _1027_ + _1028_;
  assign _1295_ = _1029_ + 64'h0000000000000001;
  assign _1297_ = _1027_ + _1030_;
  assign _1299_ = _1024_ + _1031_;
  assign _1301_ = _0956_ + _1031_;
  assign _1303_ = _1032_ + { 63'h0000000000000000, rvfi_valid };
  assign _1305_ = _1033_ + { 29'h00000000, mem_la_firstword_xfer };
  assign _1307_ = 32'd8 + _1034_;
  assign _1309_ = 32'd8 + _1035_;
  assign _1196_ = reg_pc | reg_pc_t0;
  assign _1197_ = count_cycle | count_cycle_t0;
  assign _1199_ = count_instr | count_instr_t0;
  assign _1198_ = _0046_ | _0047_;
  assign _1174_ = pcpi_rs1 | pcpi_rs1_t0;
  assign _1205_ = rvfi_order | rvfi_order_t0;
  assign _1206_ = next_pc[31:2] | next_pc_t0[31:2];
  assign _1175_ = pcpi_rs2 | pcpi_rs2_t0;
  assign _1200_ = { decoded_imm_j[31:1], 1'h0 } | { decoded_imm_j_t0[31:1], 1'h0 };
  assign _1202_ = decoded_imm | decoded_imm_t0;
  assign _1207_ = { 29'h00000000, mem_rdata_latched[4:2] } | { 29'h00000000, mem_rdata_latched_t0[4:2] };
  assign _1209_ = { 29'h00000000, mem_rdata_latched[9:7] } | { 29'h00000000, mem_rdata_latched_t0[9:7] };
  assign _1288_ = _1174_ + _1175_;
  assign _1290_ = _1196_ + _1025_;
  assign _1292_ = _1197_ + 64'h0000000000000001;
  assign _1294_ = _1198_ + _1028_;
  assign _1296_ = _1199_ + 64'h0000000000000001;
  assign _1298_ = _1198_ + _1200_;
  assign _1300_ = _1196_ + _1202_;
  assign _1302_ = _1174_ + _1202_;
  assign _1304_ = _1205_ + { 63'h0000000000000000, rvfi_valid };
  assign _1306_ = _1206_ + { 29'h00000000, mem_la_firstword_xfer };
  assign _1308_ = 32'd8 + _1207_;
  assign _1310_ = 32'd8 + _1209_;
  assign _1272_ = _1287_ ^ _1288_;
  assign _1273_ = _1289_ ^ _1290_;
  assign _1274_ = _1291_ ^ _1292_;
  assign _1275_ = _1293_ ^ _1294_;
  assign _1276_ = _1295_ ^ _1296_;
  assign _1277_ = _1297_ ^ _1298_;
  assign _1278_ = _1299_ ^ _1300_;
  assign _1279_ = _1301_ ^ _1302_;
  assign _1280_ = _1303_ ^ _1304_;
  assign _1281_ = _1305_ ^ _1306_;
  assign _1208_ = _1307_ ^ _1308_;
  assign _1210_ = _1309_ ^ _1310_;
  assign _1195_ = _1272_ | pcpi_rs1_t0;
  assign _0069_ = _1273_ | reg_pc_t0;
  assign _0071_ = _1274_ | count_cycle_t0;
  assign _0073_ = _1275_ | _0047_;
  assign _0075_ = _1276_ | count_instr_t0;
  assign _1201_ = _1277_ | _0047_;
  assign _1203_ = _1278_ | reg_pc_t0;
  assign _1204_ = _1279_ | pcpi_rs1_t0;
  assign _0083_ = _1280_ | rvfi_order_t0;
  assign _0085_ = _1281_ | next_pc_t0[31:2];
  assign _0067_ = _1195_ | pcpi_rs2_t0;
  assign _0077_ = _1201_ | { decoded_imm_j_t0[31:1], 1'h0 };
  assign _0079_ = _1203_ | decoded_imm_t0;
  assign _0081_ = _1204_ | decoded_imm_t0;
  assign _0087_ = _1208_ | { 29'h00000000, mem_rdata_latched_t0[4:2] };
  assign _0089_ = _1210_ | { 29'h00000000, mem_rdata_latched_t0[9:7] };
  assign _1036_ = pcpi_rs1_t0 & pcpi_rs2;
  assign _0095_ = mem_la_wstrb_t0 & { mem_la_write, mem_la_write, mem_la_write, mem_la_write };
  assign _1037_ = pcpi_rs2_t0 & pcpi_rs1;
  assign _0806_ = pcpi_rs1_t0 & pcpi_rs2_t0;
  assign _1211_ = _1036_ | _1037_;
  assign _0091_ = _1211_ | _0806_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_pc_rdata_t0 */
  always_ff @(posedge clk)
    rvfi_pc_rdata_t0 <= rvfi_pc_wdata_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME reg_out_t0 */
  always_ff @(posedge clk)
    reg_out_t0 <= _0019_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_rs1val_t0 */
  always_ff @(posedge clk)
    dbg_rs1val_t0 <= _0005_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_rs2val_t0 */
  always_ff @(posedge clk)
    dbg_rs2val_t0 <= _0008_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME alu_out_q_t0 */
  always_ff @(posedge clk)
    alu_out_q_t0 <= alu_out_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME q_insn_rs1_t0 */
  always_ff @(posedge clk)
    q_insn_rs1_t0 <= dbg_insn_rs1_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME q_insn_rs2_t0 */
  always_ff @(posedge clk)
    q_insn_rs2_t0 <= dbg_insn_rs2_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_rdata_q_t0[31:7] */
  always_ff @(posedge clk)
    mem_rdata_q_t0[31:7] <= _0015_[31:7];
  reg [23:0] _2568_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME _2568_ */
  always_ff @(posedge clk)
    _2568_ <= { dbg_insn_opcode_t0[31:25], dbg_insn_opcode_t0[19:15], dbg_insn_opcode_t0[11:0] };
  assign { rvfi_insn_t0[31:25], rvfi_insn_t0[19:15], rvfi_insn_t0[11:0] } = _2568_;
  assign _0108_ = ~ _1983_;
  assign _0109_ = ~ _1982_;
  assign _0110_ = ~ _1981_;
  assign _0111_ = ~ _1980_;
  assign _0112_ = ~ _1979_;
  assign _0113_ = ~ _1978_;
  assign _0114_ = ~ _1977_;
  assign _0115_ = ~ _1976_;
  assign _0116_ = ~ _1975_;
  assign _0117_ = ~ _1974_;
  assign _0118_ = ~ _1973_;
  assign _0119_ = ~ _1972_;
  assign _0120_ = ~ _1971_;
  assign _0121_ = ~ _1970_;
  assign _0123_ = ~ _0415_;
  assign _0125_ = ~ _0420_;
  assign _0126_ = ~ decoder_trigger_q;
  assign _0127_ = ~ _0421_;
  assign _0128_ = ~ _1692_;
  assign _0130_ = ~ _0422_;
  assign _0129_ = ~ _1733_;
  assign _0131_ = ~ _0423_;
  assign _0132_ = ~ _0429_;
  assign _0133_ = ~ _0430_;
  assign _0134_ = ~ _0431_;
  assign _0135_ = ~ dbg_next;
  assign _0137_ = ~ _2001_;
  assign _0138_ = ~ _2000_;
  assign _0139_ = ~ _1999_;
  assign _0140_ = ~ _1998_;
  assign _0141_ = ~ _1997_;
  assign _0142_ = ~ _1996_;
  assign _0143_ = ~ _1995_;
  assign _0144_ = ~ _1994_;
  assign _0145_ = ~ _1993_;
  assign _0146_ = ~ _1992_;
  assign _0147_ = ~ _1991_;
  assign _0148_ = ~ _1990_;
  assign _0149_ = ~ _1989_;
  assign _0150_ = ~ _1988_;
  assign _0151_ = ~ _1987_;
  assign _0152_ = ~ _1986_;
  assign _0153_ = ~ _1985_;
  assign _0154_ = ~ _1984_;
  assign _0454_ = { _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_, _1983_ } & _0002_;
  assign _0456_ = { _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_, _1982_ } & _0002_;
  assign _0458_ = { _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_, _1981_ } & _0002_;
  assign _0460_ = { _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_, _1980_ } & _0002_;
  assign _0462_ = { _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_, _1979_ } & _0002_;
  assign _0464_ = { _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_, _1978_ } & _0002_;
  assign _0466_ = { _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_, _1977_ } & _0002_;
  assign _0468_ = { _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_, _1976_ } & _0002_;
  assign _0470_ = { _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_, _1975_ } & _0002_;
  assign _0472_ = { _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_, _1974_ } & _0002_;
  assign _0474_ = { _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_, _1973_ } & _0002_;
  assign _0476_ = { _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_, _1972_ } & _0002_;
  assign _0478_ = { _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_, _1971_ } & _0002_;
  assign _0480_ = { _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_, _1970_ } & _0002_;
  assign _1038_ = { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer } & mem_rdata_latched_t0[6:0];
  assign _1040_ = { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer } & mem_rdata_latched_t0;
  assign _1042_ = { _0415_, _0415_, _0415_, _0415_, _0415_, _0415_, _0415_, _0415_, _0415_, _0415_, _0415_, _0415_, _0415_, _0415_, _0415_, _0415_ } & _2285_;
  assign _1044_ = { _0124_, _0124_, _0124_, _0124_ } & _2301_;
  assign _1047_ = { _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_, _0420_ } & mem_la_addr_t0;
  assign _1049_ = { decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q } & _0049_;
  assign _1052_ = { decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q } & decoded_rs2_t0;
  assign _1054_ = { decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q, decoder_trigger_q } & decoded_rs1_t0;
  assign _1056_ = _1692_ & _2156_;
  assign _1058_ = _1692_ & _2158_;
  assign _1060_ = _1692_ & _2160_;
  assign _1062_ = { _1692_, _1692_, _1692_ } & _2162_;
  assign _1064_ = _1692_ & _2164_;
  assign _1066_ = { _1692_, _1692_ } & _2166_;
  assign _1068_ = { _1692_, _1692_, _1692_, _1692_, _1692_, _1692_, _1692_, _1692_, _1692_, _1692_, _1692_, _1692_ } & _2168_;
  assign _1070_ = _1692_ & _2170_;
  assign _1072_ = _1692_ & _2172_;
  assign _1074_ = { _1692_, _1692_, _1692_, _1692_, _1692_, _1692_, _1692_, _1692_ } & _2239_;
  assign _1076_ = { _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_ } & _1488_;
  assign _1081_ = { _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_ } & mem_la_wdata_t0;
  assign _1083_ = _1692_ & _2154_;
  assign _1085_ = { _1692_, _1692_, _1692_, _1692_ } & _2195_;
  assign _1087_ = { _1692_, _1692_, _1692_, _1692_, _1692_ } & _2262_;
  assign _1089_ = { _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_, _1733_ } & mem_rdata_q_t0;
  assign _1091_ = { _0423_, _0423_, _0423_, _0423_, _0423_ } & _1342_;
  assign _1100_ = { _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_, _0429_ } & _1393_;
  assign _1102_ = _0430_ & _1403_[31];
  assign _1104_ = { _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_ } & _1403_[30:0];
  assign _1114_ = { dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next } & { dbg_insn_opcode_t0[24:20], dbg_insn_opcode_t0[14:12] };
  assign _1121_ = { launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn } & next_pc_t0[31:1];
  assign _1123_ = { _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_, _2001_ } & _0002_;
  assign _1125_ = { _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_, _2000_ } & _0002_;
  assign _1127_ = { _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_, _1999_ } & _0002_;
  assign _1129_ = { _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_, _1998_ } & _0002_;
  assign _1131_ = { _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_, _1997_ } & _0002_;
  assign _1133_ = { _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_, _1996_ } & _0002_;
  assign _1135_ = { _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_, _1995_ } & _0002_;
  assign _1137_ = { _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_, _1994_ } & _0002_;
  assign _1139_ = { _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_, _1993_ } & _0002_;
  assign _1141_ = { _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_, _1992_ } & _0002_;
  assign _1143_ = { _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_, _1991_ } & _0002_;
  assign _1145_ = { _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_, _1990_ } & _0002_;
  assign _1147_ = { _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_, _1989_ } & _0002_;
  assign _1149_ = { _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_, _1988_ } & _0002_;
  assign _1151_ = { _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_, _1987_ } & _0002_;
  assign _1153_ = { _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_, _1986_ } & _0002_;
  assign _1155_ = { _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_, _1985_ } & _0002_;
  assign _1157_ = { _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_, _1984_ } & _0002_;
  assign _0455_ = { _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_, _0108_ } & \cpuregs[21]_t0 ;
  assign _0457_ = { _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_, _0109_ } & \cpuregs[20]_t0 ;
  assign _0459_ = { _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_, _0110_ } & \cpuregs[1]_t0 ;
  assign _0461_ = { _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_, _0111_ } & \cpuregs[19]_t0 ;
  assign _0463_ = { _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_ } & \cpuregs[18]_t0 ;
  assign _0465_ = { _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_, _0113_ } & \cpuregs[17]_t0 ;
  assign _0467_ = { _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_, _0114_ } & \cpuregs[16]_t0 ;
  assign _0469_ = { _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_, _0115_ } & \cpuregs[15]_t0 ;
  assign _0471_ = { _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_, _0116_ } & \cpuregs[14]_t0 ;
  assign _0473_ = { _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_, _0117_ } & \cpuregs[13]_t0 ;
  assign _0475_ = { _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_, _0118_ } & \cpuregs[12]_t0 ;
  assign _0477_ = { _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_, _0119_ } & \cpuregs[11]_t0 ;
  assign _0479_ = { _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_, _0120_ } & \cpuregs[10]_t0 ;
  assign _0481_ = { _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_, _0121_ } & \cpuregs[0]_t0 ;
  assign _1039_ = { _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_ } & mem_rdata_q_t0[6:0];
  assign _1041_ = { _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_, _0122_ } & next_insn_opcode_t0;
  assign _1043_ = { _0123_, _0123_, _0123_, _0123_, _0123_, _0123_, _0123_, _0123_, _0123_, _0123_, _0123_, _0123_, _0123_, _0123_, _0123_, _0123_ } & mem_16bit_buffer_t0;
  assign _1045_ = { _1843_, _1843_, _1843_, _1843_ } & mem_wstrb_t0;
  assign _1048_ = { _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_, _0125_ } & mem_addr_t0;
  assign _1050_ = { _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_, _0126_ } & cached_insn_opcode_t0;
  assign _1051_ = _0127_ & mem_valid_t0;
  assign _1053_ = { _0126_, _0126_, _0126_, _0126_, _0126_ } & cached_insn_rs2_t0;
  assign _1055_ = { _0126_, _0126_, _0126_, _0126_, _0126_ } & cached_insn_rs1_t0;
  assign _1057_ = _0128_ & decoded_imm_j_t0[10];
  assign _1059_ = _0128_ & decoded_imm_j_t0[7];
  assign _1061_ = _0128_ & decoded_imm_j_t0[6];
  assign _1063_ = { _0128_, _0128_, _0128_ } & decoded_imm_j_t0[3:1];
  assign _1065_ = _0128_ & decoded_imm_j_t0[5];
  assign _1067_ = { _0128_, _0128_ } & decoded_imm_j_t0[9:8];
  assign _1069_ = { _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_ } & decoded_imm_j_t0[31:20];
  assign _1071_ = _0128_ & decoded_imm_j_t0[4];
  assign _1073_ = _0128_ & decoded_imm_j_t0[11];
  assign _1075_ = { _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_ } & decoded_imm_j_t0[19:12];
  assign _1077_ = { _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_ } & decoded_imm_t0;
  assign _1078_ = { _0128_, _0128_, _0128_, _0128_, _0128_ } & decoded_rs2_t0;
  assign _1082_ = { _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_, _0130_ } & mem_wdata_t0;
  assign _1084_ = _0128_ & decoded_rs1_t0[4];
  assign _1086_ = { _0128_, _0128_, _0128_, _0128_ } & decoded_rs1_t0[3:0];
  assign _1088_ = { _0128_, _0128_, _0128_, _0128_, _0128_ } & decoded_rd_t0;
  assign _1090_ = { _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_, _0129_ } & pcpi_insn_t0;
  assign _1092_ = { _0131_, _0131_, _0131_, _0131_, _0131_ } & latched_rd_t0;
  assign _1101_ = { _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_, _0132_ } & pcpi_rs2_t0;
  assign _1103_ = _0133_ & pcpi_rs1_t0[31];
  assign _1105_ = { _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_, _0134_ } & pcpi_rs1_t0[30:0];
  assign _1115_ = { _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_, _0135_ } & { rvfi_insn_t0[24:20], rvfi_insn_t0[14:12] };
  assign _1122_ = { _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_, _0136_ } & rvfi_pc_wdata_t0[31:1];
  assign _1124_ = { _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_, _0137_ } & \cpuregs[9]_t0 ;
  assign _1126_ = { _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_, _0138_ } & \cpuregs[8]_t0 ;
  assign _1128_ = { _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_, _0139_ } & \cpuregs[7]_t0 ;
  assign _1130_ = { _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_, _0140_ } & \cpuregs[6]_t0 ;
  assign _1132_ = { _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_, _0141_ } & \cpuregs[5]_t0 ;
  assign _1134_ = { _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_ } & \cpuregs[4]_t0 ;
  assign _1136_ = { _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_, _0143_ } & \cpuregs[3]_t0 ;
  assign _1138_ = { _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_, _0144_ } & \cpuregs[31]_t0 ;
  assign _1140_ = { _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_, _0145_ } & \cpuregs[30]_t0 ;
  assign _1142_ = { _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_, _0146_ } & \cpuregs[2]_t0 ;
  assign _1144_ = { _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_, _0147_ } & \cpuregs[29]_t0 ;
  assign _1146_ = { _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_, _0148_ } & \cpuregs[28]_t0 ;
  assign _1148_ = { _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_, _0149_ } & \cpuregs[27]_t0 ;
  assign _1150_ = { _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_, _0150_ } & \cpuregs[26]_t0 ;
  assign _1152_ = { _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_, _0151_ } & \cpuregs[25]_t0 ;
  assign _1154_ = { _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_ } & \cpuregs[24]_t0 ;
  assign _1156_ = { _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_ } & \cpuregs[23]_t0 ;
  assign _1158_ = { _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_, _0154_ } & \cpuregs[22]_t0 ;
  assign _1159_ = _0454_ | _0455_;
  assign _1160_ = _0456_ | _0457_;
  assign _1161_ = _0458_ | _0459_;
  assign _1162_ = _0460_ | _0461_;
  assign _1163_ = _0462_ | _0463_;
  assign _1164_ = _0464_ | _0465_;
  assign _1165_ = _0466_ | _0467_;
  assign _1166_ = _0468_ | _0469_;
  assign _1167_ = _0470_ | _0471_;
  assign _1168_ = _0472_ | _0473_;
  assign _1169_ = _0474_ | _0475_;
  assign _1170_ = _0476_ | _0477_;
  assign _1171_ = _0478_ | _0479_;
  assign _1172_ = _0480_ | _0481_;
  assign _1212_ = _1038_ | _1039_;
  assign _1213_ = _1040_ | _1041_;
  assign _1214_ = _1042_ | _1043_;
  assign _1215_ = _1044_ | _1045_;
  assign _1216_ = _1047_ | _1048_;
  assign _1217_ = _1049_ | _1050_;
  assign _1218_ = _1052_ | _1053_;
  assign _1219_ = _1054_ | _1055_;
  assign _1220_ = _1056_ | _1057_;
  assign _1221_ = _1058_ | _1059_;
  assign _1222_ = _1060_ | _1061_;
  assign _1223_ = _1062_ | _1063_;
  assign _1224_ = _1064_ | _1065_;
  assign _1225_ = _1066_ | _1067_;
  assign _1226_ = _1068_ | _1069_;
  assign _1227_ = _1070_ | _1071_;
  assign _1228_ = _1072_ | _1073_;
  assign _1229_ = _1074_ | _1075_;
  assign _1230_ = _1076_ | _1077_;
  assign _1231_ = _0482_ | _1078_;
  assign _1233_ = _1081_ | _1082_;
  assign _1234_ = _1083_ | _1084_;
  assign _1235_ = _1085_ | _1086_;
  assign _1236_ = _1087_ | _1088_;
  assign _1237_ = _1089_ | _1090_;
  assign _1238_ = _1091_ | _1092_;
  assign _1242_ = _1100_ | _1101_;
  assign _1243_ = _1102_ | _1103_;
  assign _1244_ = _1104_ | _1105_;
  assign _1249_ = _1114_ | _1115_;
  assign _1252_ = _1121_ | _1122_;
  assign _1253_ = _1123_ | _1124_;
  assign _1254_ = _1125_ | _1126_;
  assign _1255_ = _1127_ | _1128_;
  assign _1256_ = _1129_ | _1130_;
  assign _1257_ = _1131_ | _1132_;
  assign _1258_ = _1133_ | _1134_;
  assign _1259_ = _1135_ | _1136_;
  assign _1260_ = _1137_ | _1138_;
  assign _1261_ = _1139_ | _1140_;
  assign _1262_ = _1141_ | _1142_;
  assign _1263_ = _1143_ | _1144_;
  assign _1264_ = _1145_ | _1146_;
  assign _1265_ = _1147_ | _1148_;
  assign _1266_ = _1149_ | _1150_;
  assign _1267_ = _1151_ | _1152_;
  assign _1268_ = _1153_ | _1154_;
  assign _1269_ = _1155_ | _1156_;
  assign _1270_ = _1157_ | _1158_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[21]_t0  */
  always_ff @(posedge clk)
    \cpuregs[21]_t0  <= _1159_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[20]_t0  */
  always_ff @(posedge clk)
    \cpuregs[20]_t0  <= _1160_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[1]_t0  */
  always_ff @(posedge clk)
    \cpuregs[1]_t0  <= _1161_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[19]_t0  */
  always_ff @(posedge clk)
    \cpuregs[19]_t0  <= _1162_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[18]_t0  */
  always_ff @(posedge clk)
    \cpuregs[18]_t0  <= _1163_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[17]_t0  */
  always_ff @(posedge clk)
    \cpuregs[17]_t0  <= _1164_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[16]_t0  */
  always_ff @(posedge clk)
    \cpuregs[16]_t0  <= _1165_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[15]_t0  */
  always_ff @(posedge clk)
    \cpuregs[15]_t0  <= _1166_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[14]_t0  */
  always_ff @(posedge clk)
    \cpuregs[14]_t0  <= _1167_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[13]_t0  */
  always_ff @(posedge clk)
    \cpuregs[13]_t0  <= _1168_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[12]_t0  */
  always_ff @(posedge clk)
    \cpuregs[12]_t0  <= _1169_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[11]_t0  */
  always_ff @(posedge clk)
    \cpuregs[11]_t0  <= _1170_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[10]_t0  */
  always_ff @(posedge clk)
    \cpuregs[10]_t0  <= _1171_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[0]_t0  */
  always_ff @(posedge clk)
    \cpuregs[0]_t0  <= _1172_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_rdata_q_t0[6:0] */
  always_ff @(posedge clk)
    mem_rdata_q_t0[6:0] <= _1212_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME next_insn_opcode_t0 */
  always_ff @(posedge clk)
    next_insn_opcode_t0 <= _1213_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_16bit_buffer_t0 */
  always_ff @(posedge clk)
    mem_16bit_buffer_t0 <= _1214_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_wstrb_t0 */
  always_ff @(posedge clk)
    mem_wstrb_t0 <= _1215_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_addr_t0 */
  always_ff @(posedge clk)
    mem_addr_t0 <= _1216_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME cached_insn_opcode_t0 */
  always_ff @(posedge clk)
    cached_insn_opcode_t0 <= _1217_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_valid_t0 */
  always_ff @(posedge clk)
    mem_valid_t0 <= _1051_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME cached_insn_rs2_t0 */
  always_ff @(posedge clk)
    cached_insn_rs2_t0 <= _1218_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME cached_insn_rs1_t0 */
  always_ff @(posedge clk)
    cached_insn_rs1_t0 <= _1219_;
  reg \decoded_imm_j_t0_reg[10] ;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_t0_reg[10]  */
  always_ff @(posedge clk)
    \decoded_imm_j_t0_reg[10]  <= _1220_;
  assign decoded_imm_j_t0[10] = \decoded_imm_j_t0_reg[10] ;
  reg \decoded_imm_j_t0_reg[7] ;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_t0_reg[7]  */
  always_ff @(posedge clk)
    \decoded_imm_j_t0_reg[7]  <= _1221_;
  assign decoded_imm_j_t0[7] = \decoded_imm_j_t0_reg[7] ;
  reg \decoded_imm_j_t0_reg[6] ;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_t0_reg[6]  */
  always_ff @(posedge clk)
    \decoded_imm_j_t0_reg[6]  <= _1222_;
  assign decoded_imm_j_t0[6] = \decoded_imm_j_t0_reg[6] ;
  reg [2:0] _2828_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME _2828_ */
  always_ff @(posedge clk)
    _2828_ <= _1223_;
  assign decoded_imm_j_t0[3:1] = _2828_;
  reg \decoded_imm_j_t0_reg[5] ;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_t0_reg[5]  */
  always_ff @(posedge clk)
    \decoded_imm_j_t0_reg[5]  <= _1224_;
  assign decoded_imm_j_t0[5] = \decoded_imm_j_t0_reg[5] ;
  reg [1:0] _2830_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME _2830_ */
  always_ff @(posedge clk)
    _2830_ <= _1225_;
  assign decoded_imm_j_t0[9:8] = _2830_;
  reg [11:0] _2831_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME _2831_ */
  always_ff @(posedge clk)
    _2831_ <= _1226_;
  assign decoded_imm_j_t0[31:20] = _2831_;
  reg \decoded_imm_j_t0_reg[4] ;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_t0_reg[4]  */
  always_ff @(posedge clk)
    \decoded_imm_j_t0_reg[4]  <= _1227_;
  assign decoded_imm_j_t0[4] = \decoded_imm_j_t0_reg[4] ;
  reg \decoded_imm_j_t0_reg[11] ;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_t0_reg[11]  */
  always_ff @(posedge clk)
    \decoded_imm_j_t0_reg[11]  <= _1228_;
  assign decoded_imm_j_t0[11] = \decoded_imm_j_t0_reg[11] ;
  reg [7:0] _2834_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME _2834_ */
  always_ff @(posedge clk)
    _2834_ <= _1229_;
  assign decoded_imm_j_t0[19:12] = _2834_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_imm_t0 */
  always_ff @(posedge clk)
    decoded_imm_t0 <= _1230_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_rs2_t0 */
  always_ff @(posedge clk)
    decoded_rs2_t0 <= _1231_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_wdata_t0 */
  always_ff @(posedge clk)
    mem_wdata_t0 <= _1233_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_rs1_t0[4] */
  always_ff @(posedge clk)
    decoded_rs1_t0[4] <= _1234_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_rs1_t0[3:0] */
  always_ff @(posedge clk)
    decoded_rs1_t0[3:0] <= _1235_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_rd_t0 */
  always_ff @(posedge clk)
    decoded_rd_t0 <= _1236_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_insn_t0 */
  always_ff @(posedge clk)
    pcpi_insn_t0 <= _1237_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_rd_t0 */
  always_ff @(posedge clk)
    latched_rd_t0 <= _1238_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_rs2_t0 */
  always_ff @(posedge clk)
    pcpi_rs2_t0 <= _1242_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_rs1_t0[31] */
  always_ff @(posedge clk)
    pcpi_rs1_t0[31] <= _1243_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_rs1_t0[30:0] */
  always_ff @(posedge clk)
    pcpi_rs1_t0[30:0] <= _1244_;
  reg [7:0] _2846_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME _2846_ */
  always_ff @(posedge clk)
    _2846_ <= _1249_;
  assign { rvfi_insn_t0[24:20], rvfi_insn_t0[14:12] } = _2846_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_pc_wdata_t0[31:1] */
  always_ff @(posedge clk)
    rvfi_pc_wdata_t0[31:1] <= _1252_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[9]_t0  */
  always_ff @(posedge clk)
    \cpuregs[9]_t0  <= _1253_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[8]_t0  */
  always_ff @(posedge clk)
    \cpuregs[8]_t0  <= _1254_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[7]_t0  */
  always_ff @(posedge clk)
    \cpuregs[7]_t0  <= _1255_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[6]_t0  */
  always_ff @(posedge clk)
    \cpuregs[6]_t0  <= _1256_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[5]_t0  */
  always_ff @(posedge clk)
    \cpuregs[5]_t0  <= _1257_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[4]_t0  */
  always_ff @(posedge clk)
    \cpuregs[4]_t0  <= _1258_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[3]_t0  */
  always_ff @(posedge clk)
    \cpuregs[3]_t0  <= _1259_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[31]_t0  */
  always_ff @(posedge clk)
    \cpuregs[31]_t0  <= _1260_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[30]_t0  */
  always_ff @(posedge clk)
    \cpuregs[30]_t0  <= _1261_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[2]_t0  */
  always_ff @(posedge clk)
    \cpuregs[2]_t0  <= _1262_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[29]_t0  */
  always_ff @(posedge clk)
    \cpuregs[29]_t0  <= _1263_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[28]_t0  */
  always_ff @(posedge clk)
    \cpuregs[28]_t0  <= _1264_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[27]_t0  */
  always_ff @(posedge clk)
    \cpuregs[27]_t0  <= _1265_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[26]_t0  */
  always_ff @(posedge clk)
    \cpuregs[26]_t0  <= _1266_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[25]_t0  */
  always_ff @(posedge clk)
    \cpuregs[25]_t0  <= _1267_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[24]_t0  */
  always_ff @(posedge clk)
    \cpuregs[24]_t0  <= _1268_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[23]_t0  */
  always_ff @(posedge clk)
    \cpuregs[23]_t0  <= _1269_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[22]_t0  */
  always_ff @(posedge clk)
    \cpuregs[22]_t0  <= _1270_;
  /* src = "generated/out/vanilla.sv:302.2-311.6" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME last_mem_valid */
  always_ff @(posedge clk)
    if (!resetn) last_mem_valid <= 1'h0;
    else last_mem_valid <= _1721_;
  /* src = "generated/out/vanilla.sv:302.2-311.6" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_la_firstword_reg */
  always_ff @(posedge clk)
    if (!resetn) mem_la_firstword_reg <= 1'h0;
    else mem_la_firstword_reg <= _2412_;
  /* src = "generated/out/vanilla.sv:339.2-446.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_rdata_q[6:0] */
  always_ff @(posedge clk)
    if (mem_xfer) mem_rdata_q[6:0] <= mem_rdata_latched[6:0];
  /* src = "generated/out/vanilla.sv:339.2-446.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_rdata_q[31:7] */
  always_ff @(posedge clk)
    mem_rdata_q[31:7] <= _0014_[31:7];
  /* src = "generated/out/vanilla.sv:339.2-446.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME next_insn_opcode */
  always_ff @(posedge clk)
    if (mem_xfer) next_insn_opcode <= mem_rdata_latched;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_16bit_buffer */
  always_ff @(posedge clk)
    if (_0415_) mem_16bit_buffer <= _2284_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME prefetched_high_word */
  always_ff @(posedge clk)
    if (_0436_) prefetched_high_word <= 1'h0;
    else if (_0416_) prefetched_high_word <= _2287_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_la_secondword */
  always_ff @(posedge clk)
    if (_1843_) mem_la_secondword <= 1'h0;
    else if (_0417_) mem_la_secondword <= _2288_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_state */
  always_ff @(posedge clk)
    if (_0418_) mem_state <= _0016_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_wstrb */
  always_ff @(posedge clk)
    if (!_1843_) mem_wstrb <= _2300_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_instr */
  always_ff @(posedge clk)
    if (_0419_)
      if (mem_do_wdata) mem_instr <= 1'h0;
      else mem_instr <= _2302_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_addr */
  always_ff @(posedge clk)
    if (_0420_) mem_addr <= mem_la_addr;
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME cached_insn_opcode */
  always_ff @(posedge clk)
    if (decoder_trigger_q) cached_insn_opcode <= _0048_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_valid */
  always_ff @(posedge clk)
    if (_0421_) mem_valid <= _0017_;
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME cached_insn_rs2 */
  always_ff @(posedge clk)
    if (decoder_trigger_q) cached_insn_rs2 <= decoded_rs2;
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME cached_insn_rs1 */
  always_ff @(posedge clk)
    if (decoder_trigger_q) cached_insn_rs1 <= decoded_rs1;
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_valid_insn */
  always_ff @(posedge clk)
    if (_1843_) dbg_valid_insn <= 1'h0;
    else if (launch_next_insn) dbg_valid_insn <= 1'h1;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME is_compare */
  always_ff @(posedge clk)
    if (_0437_) is_compare <= 1'h0;
    else is_compare <= _2421_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME is_alu_reg_reg */
  always_ff @(posedge clk)
    if (_1692_) is_alu_reg_reg <= _2201_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME is_alu_reg_imm */
  always_ff @(posedge clk)
    if (_1692_) is_alu_reg_imm <= _2209_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_fence */
  always_ff @(posedge clk)
    if (!resetn) instr_fence <= 1'h0;
    else if (_1733_) instr_fence <= _1793_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_ecall_ebreak */
  always_ff @(posedge clk)
    if (_1733_) instr_ecall_ebreak <= _1848_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME is_beq_bne_blt_bge_bltu_bgeu */
  always_ff @(posedge clk)
    if (!resetn) is_beq_bne_blt_bge_bltu_bgeu <= 1'h0;
    else if (_1692_) is_beq_bne_blt_bge_bltu_bgeu <= _2212_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME is_sll_srl_sra */
  always_ff @(posedge clk)
    if (_1733_) is_sll_srl_sra <= _1799_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME is_sb_sh_sw */
  always_ff @(posedge clk)
    if (_1692_) is_sb_sh_sw <= _2215_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME is_jalr_addi_slti_sltiu_xori_ori_andi */
  always_ff @(posedge clk)
    if (_1733_) is_jalr_addi_slti_sltiu_xori_ori_andi <= _1849_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME is_slli_srli_srai */
  always_ff @(posedge clk)
    if (_1733_) is_slli_srli_srai <= _1797_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME is_lb_lh_lw_lbu_lhu */
  always_ff @(posedge clk)
    if (_1692_) is_lb_lh_lw_lbu_lhu <= _2219_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME compressed_instr */
  always_ff @(posedge clk)
    if (_1692_) compressed_instr <= _2220_;
  reg \decoded_imm_j_reg[10] ;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_reg[10]  */
  always_ff @(posedge clk)
    if (_1692_) \decoded_imm_j_reg[10]  <= _2155_;
  assign decoded_imm_j[10] = \decoded_imm_j_reg[10] ;
  reg \decoded_imm_j_reg[7] ;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_reg[7]  */
  always_ff @(posedge clk)
    if (_1692_) \decoded_imm_j_reg[7]  <= _2157_;
  assign decoded_imm_j[7] = \decoded_imm_j_reg[7] ;
  reg \decoded_imm_j_reg[6] ;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_reg[6]  */
  always_ff @(posedge clk)
    if (_1692_) \decoded_imm_j_reg[6]  <= _2159_;
  assign decoded_imm_j[6] = \decoded_imm_j_reg[6] ;
  reg [2:0] _2898_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME _2898_ */
  always_ff @(posedge clk)
    if (_1692_) _2898_ <= _2161_;
  assign decoded_imm_j[3:1] = _2898_;
  reg \decoded_imm_j_reg[5] ;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_reg[5]  */
  always_ff @(posedge clk)
    if (_1692_) \decoded_imm_j_reg[5]  <= _2163_;
  assign decoded_imm_j[5] = \decoded_imm_j_reg[5] ;
  reg [1:0] _2900_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME _2900_ */
  always_ff @(posedge clk)
    if (_1692_) _2900_ <= _2165_;
  assign decoded_imm_j[9:8] = _2900_;
  reg [11:0] _2901_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME _2901_ */
  always_ff @(posedge clk)
    if (_1692_) _2901_ <= _2167_;
  assign decoded_imm_j[31:20] = _2901_;
  reg \decoded_imm_j_reg[4] ;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_reg[4]  */
  always_ff @(posedge clk)
    if (_1692_) \decoded_imm_j_reg[4]  <= _2169_;
  assign decoded_imm_j[4] = \decoded_imm_j_reg[4] ;
  reg \decoded_imm_j_reg[11] ;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \decoded_imm_j_reg[11]  */
  always_ff @(posedge clk)
    if (_1692_) \decoded_imm_j_reg[11]  <= _2171_;
  assign decoded_imm_j[11] = \decoded_imm_j_reg[11] ;
  reg [7:0] _2904_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME _2904_ */
  always_ff @(posedge clk)
    if (_1692_) _2904_ <= _2238_;
  assign decoded_imm_j[19:12] = _2904_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_imm */
  always_ff @(posedge clk)
    if (_1733_) decoded_imm <= _1487_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_rs2 */
  always_ff @(posedge clk)
    if (_1692_) decoded_rs2 <= _2236_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME trap */
  always_ff @(posedge clk)
    if (!resetn) trap <= 1'h0;
    else trap <= _2051_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_wdata */
  always_ff @(posedge clk)
    if (_0386_)
      if (mem_instr) rvfi_mem_wdata <= 32'd0;
      else rvfi_mem_wdata <= _2014_;
  /* src = "generated/out/vanilla.sv:460.2-533.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_wdata */
  always_ff @(posedge clk)
    if (_0422_) mem_wdata <= mem_la_wdata;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_rs1[4] */
  always_ff @(posedge clk)
    if (_1692_) decoded_rs1[4] <= _2153_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_rs1[3:0] */
  always_ff @(posedge clk)
    if (_1692_) decoded_rs1[3:0] <= _2194_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME decoded_rd */
  always_ff @(posedge clk)
    if (_1692_) decoded_rd <= _2261_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_rdinstrh */
  always_ff @(posedge clk)
    if (_1733_) instr_rdinstrh <= _1790_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_rdinstr */
  always_ff @(posedge clk)
    if (_1733_) instr_rdinstr <= _1788_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_rdcycleh */
  always_ff @(posedge clk)
    if (_1733_) instr_rdcycleh <= _1786_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_rdcycle */
  always_ff @(posedge clk)
    if (_1733_) instr_rdcycle <= _1781_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_and */
  always_ff @(posedge clk)
    if (!resetn) instr_and <= 1'h0;
    else if (_1733_) instr_and <= _1776_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_or */
  always_ff @(posedge clk)
    if (!resetn) instr_or <= 1'h0;
    else if (_1733_) instr_or <= _1774_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sra */
  always_ff @(posedge clk)
    if (!resetn) instr_sra <= 1'h0;
    else if (_1733_) instr_sra <= _1772_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_srl */
  always_ff @(posedge clk)
    if (!resetn) instr_srl <= 1'h0;
    else if (_1733_) instr_srl <= _1771_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_xor */
  always_ff @(posedge clk)
    if (!resetn) instr_xor <= 1'h0;
    else if (_1733_) instr_xor <= _1769_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sltu */
  always_ff @(posedge clk)
    if (!resetn) instr_sltu <= 1'h0;
    else if (_1733_) instr_sltu <= _1767_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_slt */
  always_ff @(posedge clk)
    if (!resetn) instr_slt <= 1'h0;
    else if (_1733_) instr_slt <= _1765_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sub */
  always_ff @(posedge clk)
    if (!resetn) instr_sub <= 1'h0;
    else if (_1733_) instr_sub <= _1761_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_add */
  always_ff @(posedge clk)
    if (!resetn) instr_add <= 1'h0;
    else if (_1733_) instr_add <= _1760_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_srai */
  always_ff @(posedge clk)
    if (_1733_) instr_srai <= _1758_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_srli */
  always_ff @(posedge clk)
    if (_1733_) instr_srli <= _1757_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_slli */
  always_ff @(posedge clk)
    if (_1733_) instr_slli <= _1755_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_andi */
  always_ff @(posedge clk)
    if (!resetn) instr_andi <= 1'h0;
    else if (_1733_) instr_andi <= _1753_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_ori */
  always_ff @(posedge clk)
    if (!resetn) instr_ori <= 1'h0;
    else if (_1733_) instr_ori <= _1752_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_xori */
  always_ff @(posedge clk)
    if (!resetn) instr_xori <= 1'h0;
    else if (_1733_) instr_xori <= _1751_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sltiu */
  always_ff @(posedge clk)
    if (!resetn) instr_sltiu <= 1'h0;
    else if (_1733_) instr_sltiu <= _1750_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_slti */
  always_ff @(posedge clk)
    if (!resetn) instr_slti <= 1'h0;
    else if (_1733_) instr_slti <= _1749_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_addi */
  always_ff @(posedge clk)
    if (!resetn) instr_addi <= 1'h0;
    else if (_1733_) instr_addi <= _1748_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sw */
  always_ff @(posedge clk)
    if (_1733_) instr_sw <= _1747_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sh */
  always_ff @(posedge clk)
    if (_1733_) instr_sh <= _1746_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sb */
  always_ff @(posedge clk)
    if (_1733_) instr_sb <= _1745_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lhu */
  always_ff @(posedge clk)
    if (_1733_) instr_lhu <= _1744_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lbu */
  always_ff @(posedge clk)
    if (_1733_) instr_lbu <= _1743_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lw */
  always_ff @(posedge clk)
    if (_1733_) instr_lw <= _1742_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lh */
  always_ff @(posedge clk)
    if (_1733_) instr_lh <= _1741_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lb */
  always_ff @(posedge clk)
    if (_1733_) instr_lb <= _1740_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_bgeu */
  always_ff @(posedge clk)
    if (!resetn) instr_bgeu <= 1'h0;
    else if (_1733_) instr_bgeu <= _1739_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_bltu */
  always_ff @(posedge clk)
    if (!resetn) instr_bltu <= 1'h0;
    else if (_1733_) instr_bltu <= _1738_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_bge */
  always_ff @(posedge clk)
    if (!resetn) instr_bge <= 1'h0;
    else if (_1733_) instr_bge <= _1737_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_blt */
  always_ff @(posedge clk)
    if (!resetn) instr_blt <= 1'h0;
    else if (_1733_) instr_blt <= _1736_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_bne */
  always_ff @(posedge clk)
    if (!resetn) instr_bne <= 1'h0;
    else if (_1733_) instr_bne <= _1735_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_beq */
  always_ff @(posedge clk)
    if (!resetn) instr_beq <= 1'h0;
    else if (_1733_) instr_beq <= _1734_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_jalr */
  always_ff @(posedge clk)
    if (_1692_) instr_jalr <= _2267_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_jal */
  always_ff @(posedge clk)
    if (_1692_) instr_jal <= _2271_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_auipc */
  always_ff @(posedge clk)
    if (_1692_) instr_auipc <= _1657_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_lui */
  always_ff @(posedge clk)
    if (_1692_) instr_lui <= _2276_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_insn */
  always_ff @(posedge clk)
    if (_1733_) pcpi_insn <= mem_rdata_q;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_timeout */
  always_ff @(posedge clk)
    if (!resetn) pcpi_timeout <= 1'h0;
    else pcpi_timeout <= _1808_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_timeout_counter */
  always_ff @(posedge clk)
    if (!_1691_) pcpi_timeout_counter <= 4'hf;
    else if (_2052_) pcpi_timeout_counter <= _2429_[3:0];
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_rd */
  always_ff @(posedge clk)
    if (_0423_) latched_rd <= _1341_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_is_lb */
  always_ff @(posedge clk)
    if (!resetn) latched_is_lb <= 1'h0;
    else if (_0424_) latched_is_lb <= _1343_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_is_lh */
  always_ff @(posedge clk)
    if (!resetn) latched_is_lh <= 1'h0;
    else if (_0424_) latched_is_lh <= _1344_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_compr */
  always_ff @(posedge clk)
    if (_0425_) latched_compr <= compressed_instr;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_branch */
  always_ff @(posedge clk)
    if (!resetn) latched_branch <= 1'h0;
    else if (_0388_) latched_branch <= _1345_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_stalu */
  always_ff @(posedge clk)
    if (!resetn) latched_stalu <= 1'h0;
    else if (_0426_) latched_stalu <= _1346_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME latched_store */
  always_ff @(posedge clk)
    if (!resetn) latched_store <= 1'h0;
    else if (_0427_) latched_store <= _1350_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME count_cycle */
  always_ff @(posedge clk)
    if (!resetn) count_cycle <= 64'h0000000000000000;
    else count_cycle <= _0070_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME reg_pc */
  always_ff @(posedge clk)
    if (!resetn) reg_pc <= 32'd2147483648;
    else if (_1628_) reg_pc <= _0046_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME reg_next_pc */
  always_ff @(posedge clk)
    if (!resetn) reg_next_pc <= 32'd2147483648;
    else if (_1628_) reg_next_pc <= _2116_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_wmask */
  always_ff @(posedge clk)
    if (_0386_)
      if (mem_instr) rvfi_mem_wmask <= 4'h0;
      else rvfi_mem_wmask <= _2018_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_rmask */
  always_ff @(posedge clk)
    if (_0386_)
      if (mem_instr) rvfi_mem_rmask <= 4'h0;
      else rvfi_mem_rmask <= _2020_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_do_wdata */
  always_ff @(posedge clk)
    if (_0024_) mem_do_wdata <= 1'h1;
    else if (_1835_) mem_do_wdata <= 1'h0;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_do_rdata */
  always_ff @(posedge clk)
    if (_0022_) mem_do_rdata <= 1'h1;
    else if (_1835_) mem_do_rdata <= 1'h0;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_do_rinst */
  always_ff @(posedge clk)
    if (_0023_) mem_do_rinst <= 1'h1;
    else if (_0428_) mem_do_rinst <= _2097_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_rs2 */
  always_ff @(posedge clk)
    if (_0429_) pcpi_rs2 <= _1392_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_rs1[31] */
  always_ff @(posedge clk)
    if (_0430_) pcpi_rs1[31] <= _1402_[31];
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_rs1[30:0] */
  always_ff @(posedge clk)
    if (_0431_) pcpi_rs1[30:0] <= _1402_[30:0];
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_rdata */
  always_ff @(posedge clk)
    if (_0386_)
      if (mem_instr) rvfi_mem_rdata <= 32'd0;
      else rvfi_mem_rdata <= _2016_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_wordsize */
  always_ff @(posedge clk)
    if (_0432_) mem_wordsize <= _1389_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME instr_sll */
  always_ff @(posedge clk)
    if (!resetn) instr_sll <= 1'h0;
    else if (_1733_) instr_sll <= _1763_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_addr */
  always_ff @(posedge clk)
    if (_0386_)
      if (mem_instr) rvfi_mem_addr <= 32'd0;
      else rvfi_mem_addr <= _2021_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rd_wdata */
  always_ff @(posedge clk)
    if (_0438_) rvfi_rd_wdata <= 32'd0;
    else if (_0413_) rvfi_rd_wdata <= _2024_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rd_addr */
  always_ff @(posedge clk)
    if (_0438_) rvfi_rd_addr <= 5'h00;
    else if (_0413_) rvfi_rd_addr <= _2028_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rs2_rdata */
  always_ff @(posedge clk)
    if (!dbg_rs2val_valid) rvfi_rs2_rdata <= 32'd0;
    else rvfi_rs2_rdata <= dbg_rs2val;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rs1_rdata */
  always_ff @(posedge clk)
    if (_0439_) rvfi_rs1_rdata <= 32'd0;
    else rvfi_rs1_rdata <= dbg_rs1val;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rs2_addr */
  always_ff @(posedge clk)
    if (!dbg_rs2val_valid) rvfi_rs2_addr <= 5'h00;
    else rvfi_rs2_addr <= dbg_insn_rs2;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rs1_addr */
  always_ff @(posedge clk)
    if (_0439_) rvfi_rs1_addr <= 5'h00;
    else rvfi_rs1_addr <= dbg_insn_rs1;
  reg [7:0] _2984_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME _2984_ */
  always_ff @(posedge clk)
    if (dbg_next) _2984_ <= { dbg_insn_opcode[24:20], dbg_insn_opcode[14:12] };
  assign { rvfi_insn[24:20], rvfi_insn[14:12] } = _2984_;
  reg [23:0] _2985_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME _2985_ */
  always_ff @(posedge clk)
    _2985_ <= { dbg_insn_opcode[31:25], dbg_insn_opcode[19:15], dbg_insn_opcode[11:0] };
  assign { rvfi_insn[31:25], rvfi_insn[19:15], rvfi_insn[11:0] } = _2985_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_order */
  always_ff @(posedge clk)
    if (!resetn) rvfi_order <= 64'h0000000000000000;
    else rvfi_order <= _0082_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME cpu_state */
  always_ff @(posedge clk)
    if (_1702_) cpu_state <= 8'h80;
    else cpu_state <= _2077_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_do_prefetch */
  always_ff @(posedge clk)
    if (_1835_) mem_do_prefetch <= 1'h0;
    else if (_0433_) mem_do_prefetch <= _1694_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME decoder_pseudo_trigger */
  always_ff @(posedge clk)
    if (!_0440_) decoder_pseudo_trigger <= 1'h0;
    else decoder_pseudo_trigger <= _2034_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME count_instr */
  always_ff @(posedge clk)
    if (!resetn) count_instr <= 64'h0000000000000000;
    else if (_0434_) count_instr <= _0074_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_valid */
  always_ff @(posedge clk)
    if (!resetn) pcpi_valid <= 1'h0;
    else if (_0435_) pcpi_valid <= _2121_;
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_pc_wdata[0] */
  always_ff @(posedge clk)
    if (launch_next_insn)
      if (_1686_) rvfi_pc_wdata[0] <= 1'h0;
      else rvfi_pc_wdata[0] <= reg_next_pc[0];
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_pc_wdata[31:1] */
  always_ff @(posedge clk)
    if (launch_next_insn) rvfi_pc_wdata[31:1] <= next_pc[31:1];
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[9]  */
  always_ff @(posedge clk)
    if (_2001_) \cpuregs[9]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[8]  */
  always_ff @(posedge clk)
    if (_2000_) \cpuregs[8]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[7]  */
  always_ff @(posedge clk)
    if (_1999_) \cpuregs[7]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[6]  */
  always_ff @(posedge clk)
    if (_1998_) \cpuregs[6]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[5]  */
  always_ff @(posedge clk)
    if (_1997_) \cpuregs[5]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[4]  */
  always_ff @(posedge clk)
    if (_1996_) \cpuregs[4]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[3]  */
  always_ff @(posedge clk)
    if (_1995_) \cpuregs[3]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[31]  */
  always_ff @(posedge clk)
    if (_1994_) \cpuregs[31]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[30]  */
  always_ff @(posedge clk)
    if (_1993_) \cpuregs[30]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[2]  */
  always_ff @(posedge clk)
    if (_1992_) \cpuregs[2]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[29]  */
  always_ff @(posedge clk)
    if (_1991_) \cpuregs[29]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[28]  */
  always_ff @(posedge clk)
    if (_1990_) \cpuregs[28]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[27]  */
  always_ff @(posedge clk)
    if (_1989_) \cpuregs[27]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[26]  */
  always_ff @(posedge clk)
    if (_1988_) \cpuregs[26]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[25]  */
  always_ff @(posedge clk)
    if (_1987_) \cpuregs[25]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[24]  */
  always_ff @(posedge clk)
    if (_1986_) \cpuregs[24]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[23]  */
  always_ff @(posedge clk)
    if (_1985_) \cpuregs[23]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[22]  */
  always_ff @(posedge clk)
    if (_1984_) \cpuregs[22]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[21]  */
  always_ff @(posedge clk)
    if (_1983_) \cpuregs[21]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[20]  */
  always_ff @(posedge clk)
    if (_1982_) \cpuregs[20]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[1]  */
  always_ff @(posedge clk)
    if (_1981_) \cpuregs[1]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[19]  */
  always_ff @(posedge clk)
    if (_1980_) \cpuregs[19]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[18]  */
  always_ff @(posedge clk)
    if (_1979_) \cpuregs[18]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[17]  */
  always_ff @(posedge clk)
    if (_1978_) \cpuregs[17]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[16]  */
  always_ff @(posedge clk)
    if (_1977_) \cpuregs[16]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[15]  */
  always_ff @(posedge clk)
    if (_1976_) \cpuregs[15]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[14]  */
  always_ff @(posedge clk)
    if (_1975_) \cpuregs[14]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[13]  */
  always_ff @(posedge clk)
    if (_1974_) \cpuregs[13]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[12]  */
  always_ff @(posedge clk)
    if (_1973_) \cpuregs[12]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[11]  */
  always_ff @(posedge clk)
    if (_1972_) \cpuregs[11]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[10]  */
  always_ff @(posedge clk)
    if (_1971_) \cpuregs[10]  <= _0001_;
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME \cpuregs[0]  */
  always_ff @(posedge clk)
    if (_1970_) \cpuregs[0]  <= _0001_;
  assign _1313_ = _1692_ ? _2236_ : decoded_rs2;
  assign _1314_ = _1692_ ? { _2153_, _2194_ } : decoded_rs1;
  assign _1282_ = ~ _0000_[0];
  assign _1283_ = ~ _0000_[1];
  assign _1284_ = ~ _0000_[2];
  assign _1285_ = ~ _0000_[3];
  assign _1286_ = ~ _0000_[4];
  assign _0976_ = _1282_ & _1283_;
  assign _0977_ = _1285_ & _1286_;
  assign _0978_ = _1284_ & _0977_;
  assign _0979_ = _0976_ & _0978_;
  assign _0980_ = _0000_[0] & _1283_;
  assign _0981_ = _0980_ & _0978_;
  assign _0982_ = _1282_ & _0000_[1];
  assign _0983_ = _0982_ & _0978_;
  assign _0984_ = _0000_[0] & _0000_[1];
  assign _0985_ = _0984_ & _0978_;
  assign _0986_ = _0000_[2] & _0977_;
  assign _0987_ = _0976_ & _0986_;
  assign _0988_ = _0980_ & _0986_;
  assign _0989_ = _0982_ & _0986_;
  assign _0990_ = _0984_ & _0986_;
  assign _0991_ = _0000_[3] & _1286_;
  assign _0992_ = _1284_ & _0991_;
  assign _0993_ = _0976_ & _0992_;
  assign _0994_ = _0980_ & _0992_;
  assign _0995_ = _0982_ & _0992_;
  assign _0996_ = _0984_ & _0992_;
  assign _0997_ = _0000_[2] & _0991_;
  assign _0998_ = _0976_ & _0997_;
  assign _0999_ = _0980_ & _0997_;
  assign _1000_ = _0982_ & _0997_;
  assign _1001_ = _0984_ & _0997_;
  assign _1002_ = _1285_ & _0000_[4];
  assign _1003_ = _1284_ & _1002_;
  assign _1004_ = _0976_ & _1003_;
  assign _1005_ = _0980_ & _1003_;
  assign _1006_ = _0982_ & _1003_;
  assign _1007_ = _0984_ & _1003_;
  assign _1008_ = _0000_[2] & _1002_;
  assign _1009_ = _0976_ & _1008_;
  assign _1010_ = _0980_ & _1008_;
  assign _1011_ = _0982_ & _1008_;
  assign _1012_ = _0984_ & _1008_;
  assign _1013_ = _0000_[3] & _0000_[4];
  assign _1014_ = _1284_ & _1013_;
  assign _1015_ = _0976_ & _1014_;
  assign _1016_ = _0980_ & _1014_;
  assign _1017_ = _0982_ & _1014_;
  assign _1018_ = _0984_ & _1014_;
  assign _1019_ = _0000_[2] & _1013_;
  assign _1020_ = _0976_ & _1019_;
  assign _1021_ = _0980_ & _1019_;
  assign _1022_ = _0982_ & _1019_;
  assign _1023_ = _0984_ & _1019_;
  assign _0155_ = ~ { latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh };
  assign _0156_ = ~ { latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb };
  assign _0157_ = ~ { _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_ };
  assign _0158_ = ~ { _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_ };
  assign _0159_ = ~ { _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_ };
  assign _0160_ = ~ { _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_ };
  assign _0161_ = ~ { is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh };
  assign _0162_ = ~ { instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh };
  assign _0163_ = ~ { instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh };
  assign _0164_ = ~ { _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_ };
  assign _0165_ = ~ { _1631_, _1631_, _1631_, _1631_, _1631_ };
  assign _0166_ = ~ { _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_ };
  assign _0167_ = ~ { _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_, _0452_ };
  assign _0168_ = ~ { _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_ };
  assign _0169_ = ~ { _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_ };
  assign _0170_ = ~ { _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_ };
  assign _0171_ = ~ { _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_ };
  assign _0172_ = ~ { _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_ };
  assign _0173_ = ~ { is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal };
  assign _0174_ = ~ { _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_ };
  assign _0175_ = ~ { _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_ };
  assign _0176_ = ~ { is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare, is_compare };
  assign _0177_ = ~ { _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_ };
  assign _0178_ = ~ { _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_ };
  assign _0179_ = ~ _2130_;
  assign _0180_ = ~ _2134_;
  assign _0181_ = ~ _2152_;
  assign _0182_ = ~ _1186_;
  assign _0183_ = ~ _0442_;
  assign _0184_ = ~ _2147_;
  assign _0185_ = ~ _1187_;
  assign _0186_ = ~ { _2136_, _2136_, _2136_, _2136_ };
  assign _0187_ = ~ { _2151_, _2151_, _2151_, _2151_ };
  assign _0188_ = ~ { _1188_, _1188_, _1188_, _1188_ };
  assign _0189_ = ~ { _2134_, _2134_, _2134_, _2134_ };
  assign _0190_ = ~ { _2152_, _2152_, _2152_, _2152_ };
  assign _0191_ = ~ { _1186_, _1186_, _1186_, _1186_ };
  assign _0192_ = ~ { _0442_, _0442_, _0442_, _0442_ };
  assign _0193_ = ~ { _2147_, _2147_, _2147_, _2147_ };
  assign _0194_ = ~ { _1187_, _1187_, _1187_, _1187_ };
  assign _0195_ = ~ _2148_;
  assign _0196_ = ~ { is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu };
  assign _0197_ = ~ { is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw };
  assign _0198_ = ~ { instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal };
  assign _0199_ = ~ { _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_ };
  assign _0200_ = ~ { _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_ };
  assign _0201_ = ~ { _2136_, _2136_, _2136_, _2136_, _2136_ };
  assign _0202_ = ~ { _2133_, _2133_, _2133_, _2133_, _2133_ };
  assign _0203_ = ~ { _1188_, _1188_, _1188_, _1188_, _1188_ };
  assign _0204_ = ~ { _2134_, _2134_, _2134_, _2134_, _2134_ };
  assign _0205_ = ~ { _2152_, _2152_, _2152_, _2152_, _2152_ };
  assign _0206_ = ~ { _1186_, _1186_, _1186_, _1186_, _1186_ };
  assign _0207_ = ~ { _2130_, _2130_, _2130_, _2130_, _2130_ };
  assign _0208_ = ~ { _1190_, _1190_, _1190_, _1190_, _1190_ };
  assign _0209_ = ~ { _0362_, _0362_, _0362_, _0362_, _0362_ };
  assign _0210_ = ~ { _1189_, _1189_, _1189_, _1189_, _1189_ };
  assign _0211_ = ~ _0360_;
  assign _0212_ = ~ _0449_;
  assign _0213_ = ~ _0361_;
  assign _0214_ = ~ { _2151_, _2151_, _2151_, _2151_, _2151_ };
  assign _0215_ = ~ { _0441_, _0441_, _0441_ };
  assign _0216_ = ~ { _2133_, _2133_, _2133_ };
  assign _0217_ = ~ { _1192_, _1192_, _1192_ };
  assign _0218_ = ~ { _2134_, _2134_, _2134_ };
  assign _0219_ = ~ { _2152_, _2152_, _2152_ };
  assign _0220_ = ~ { _1186_, _1186_, _1186_ };
  assign _0221_ = ~ { _2147_, _2147_, _2147_ };
  assign _0222_ = ~ { _2130_, _2130_, _2130_ };
  assign _0223_ = ~ { _1193_, _1193_, _1193_ };
  assign _0224_ = ~ { _2136_, _2136_, _2136_, _2136_, _2136_, _2136_ };
  assign _0225_ = ~ { _2133_, _2133_, _2133_, _2133_, _2133_, _2133_ };
  assign _0226_ = ~ { _2151_, _2151_, _2151_, _2151_, _2151_, _2151_ };
  assign _0227_ = ~ { _1188_, _1188_, _1188_, _1188_, _1188_, _1188_ };
  assign _0228_ = ~ { _2134_, _2134_, _2134_, _2134_, _2134_, _2134_ };
  assign _0229_ = ~ { _2152_, _2152_, _2152_, _2152_, _2152_, _2152_ };
  assign _0230_ = ~ { _1186_, _1186_, _1186_, _1186_, _1186_, _1186_ };
  assign _0231_ = ~ { _0442_, _0442_, _0442_, _0442_, _0442_, _0442_ };
  assign _0232_ = ~ { _0362_, _0362_, _0362_, _0362_, _0362_, _0362_ };
  assign _0233_ = ~ { _2147_, _2147_, _2147_, _2147_, _2147_, _2147_ };
  assign _0234_ = ~ { _1187_, _1187_, _1187_, _1187_, _1187_, _1187_ };
  assign _0235_ = ~ { _0441_, _0441_, _0441_, _0441_, _0441_, _0441_ };
  assign _0236_ = ~ { _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_ };
  assign _0237_ = ~ { _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_ };
  assign _0238_ = ~ { _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_ };
  assign _0239_ = ~ { pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1] };
  assign _0240_ = ~ { _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_ };
  assign _0241_ = ~ { _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_ };
  assign _0242_ = ~ { pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready };
  assign _0243_ = ~ { _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4] };
  assign _0244_ = ~ { _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3] };
  assign _0245_ = ~ { _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2] };
  assign _0246_ = ~ { _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1] };
  assign _0247_ = ~ { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] };
  assign _0248_ = ~ { _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4] };
  assign _0249_ = ~ { _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3] };
  assign _0250_ = ~ { _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2] };
  assign _0251_ = ~ { _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1] };
  assign _0252_ = ~ { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] };
  assign _0253_ = ~ mem_do_rdata;
  assign _0254_ = ~ { latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch };
  assign _0255_ = ~ { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn };
  assign _0256_ = ~ resetn;
  assign _0257_ = ~ { _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_ };
  assign _0258_ = ~ instr_jal;
  assign _0136_ = ~ launch_next_insn;
  assign _0259_ = ~ { launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn, launch_next_insn };
  assign _0260_ = ~ { _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_ };
  assign _0261_ = ~ { _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_ };
  assign _0262_ = ~ { mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata };
  assign _0263_ = ~ { mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata, mem_do_wdata };
  assign _0264_ = ~ { _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_ };
  assign _0265_ = ~ { decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger };
  assign _0266_ = ~ _1628_;
  assign _0267_ = ~ _1724_;
  assign _0268_ = ~ _1726_;
  assign _0269_ = ~ _1727_;
  assign _0270_ = ~ mem_rdata_latched[12];
  assign _0271_ = ~ _1647_;
  assign _0272_ = ~ _1648_;
  assign _0273_ = ~ _1729_;
  assign _0274_ = ~ { _1729_, _1729_, _1729_ };
  assign _0275_ = ~ { _1729_, _1729_ };
  assign _0276_ = ~ { _1729_, _1729_, _1729_, _1729_, _1729_, _1729_, _1729_, _1729_, _1729_, _1729_, _1729_, _1729_ };
  assign _0277_ = ~ { _1724_, _1724_, _1724_, _1724_ };
  assign _0278_ = ~ { _1726_, _1726_, _1726_, _1726_ };
  assign _0279_ = ~ { _1727_, _1727_, _1727_, _1727_ };
  assign _0280_ = ~ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] };
  assign _0281_ = ~ { _1647_, _1647_, _1647_, _1647_ };
  assign _0282_ = ~ { _1648_, _1648_, _1648_, _1648_ };
  assign _0283_ = ~ { _1729_, _1729_, _1729_, _1729_ };
  assign _0284_ = ~ _2136_;
  assign _0285_ = ~ { _1727_, _1727_, _1727_, _1727_, _1727_ };
  assign _0286_ = ~ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] };
  assign _0287_ = ~ { _1648_, _1648_, _1648_, _1648_, _1648_ };
  assign _0288_ = ~ { _1729_, _1729_, _1729_, _1729_, _1729_ };
  assign _0289_ = ~ { _1729_, _1729_, _1729_, _1729_, _1729_, _1729_, _1729_, _1729_ };
  assign _0290_ = ~ { _1726_, _1726_, _1726_, _1726_, _1726_ };
  assign _0291_ = ~ { _1647_, _1647_, _1647_, _1647_, _1647_ };
  assign _0292_ = ~ { decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q };
  assign _0293_ = ~ { decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q };
  assign _0294_ = ~ { dbg_next, dbg_next, dbg_next, dbg_next, dbg_next };
  assign _0295_ = ~ { dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next };
  assign _0296_ = ~ { _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_ };
  assign _0297_ = ~ { mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata, mem_do_rdata };
  assign _0298_ = ~ { mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word };
  assign _0299_ = ~ { mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read };
  assign _0300_ = ~ mem_la_read;
  assign _0301_ = ~ { _1845_, _1845_, _1845_, _1845_ };
  assign _0302_ = ~ { _1841_, _1841_, _1841_, _1841_ };
  assign _0303_ = ~ { _1814_, _1814_, _1814_, _1814_ };
  assign _0122_ = ~ mem_xfer;
  assign _0124_ = ~ _1843_;
  assign _0304_ = ~ _1723_;
  assign _0305_ = ~ _1645_;
  assign _0306_ = ~ _1646_;
  assign _0307_ = ~ _1722_;
  assign _0308_ = ~ { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer };
  assign _0309_ = ~ { _1723_, _1723_, _1723_, _1723_, _1723_ };
  assign _0310_ = ~ { _1644_, _1644_, _1644_, _1644_, _1644_ };
  assign _0311_ = ~ { _1722_, _1722_, _1722_, _1722_, _1722_ };
  assign _0312_ = ~ { _2147_, _2147_, _2147_, _2147_, _2147_ };
  assign _0313_ = ~ { _2148_, _2148_, _2148_, _2148_, _2148_ };
  assign _0314_ = ~ { mem_xfer, mem_xfer, mem_xfer };
  assign _0315_ = ~ { _1723_, _1723_, _1723_ };
  assign _0316_ = ~ { _1724_, _1724_, _1724_ };
  assign _0317_ = ~ { _1726_, _1726_, _1726_ };
  assign _0318_ = ~ { _1727_, _1727_, _1727_ };
  assign _0319_ = ~ { _1645_, _1645_, _1645_ };
  assign _0320_ = ~ { _1646_, _1646_, _1646_ };
  assign _0321_ = ~ { _1647_, _1647_, _1647_ };
  assign _0322_ = ~ { _1649_, _1649_, _1649_ };
  assign _0323_ = ~ { _1650_, _1650_, _1650_ };
  assign _0324_ = ~ { _1651_, _1651_, _1651_ };
  assign _0325_ = ~ { _1652_, _1652_, _1652_ };
  assign _0326_ = ~ { _1648_, _1648_, _1648_ };
  assign _0327_ = ~ { _1644_, _1644_, _1644_ };
  assign _0328_ = ~ { _1722_, _1722_, _1722_ };
  assign _0329_ = ~ { mem_xfer, mem_xfer, mem_xfer, mem_xfer };
  assign _0330_ = ~ { _1722_, _1722_, _1722_, _1722_ };
  assign _0331_ = ~ { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer };
  assign _0332_ = ~ { _1723_, _1723_, _1723_, _1723_, _1723_, _1723_ };
  assign _0333_ = ~ { _1724_, _1724_, _1724_, _1724_, _1724_, _1724_ };
  assign _0334_ = ~ { _1726_, _1726_, _1726_, _1726_, _1726_, _1726_ };
  assign _0335_ = ~ { _1727_, _1727_, _1727_, _1727_, _1727_, _1727_ };
  assign _0336_ = ~ { _1645_, _1645_, _1645_, _1645_, _1645_, _1645_ };
  assign _0337_ = ~ { _1646_, _1646_, _1646_, _1646_, _1646_, _1646_ };
  assign _0338_ = ~ { _1647_, _1647_, _1647_, _1647_, _1647_, _1647_ };
  assign _0339_ = ~ { _1648_, _1648_, _1648_, _1648_, _1648_, _1648_ };
  assign _0340_ = ~ { _1644_, _1644_, _1644_, _1644_, _1644_, _1644_ };
  assign _0341_ = ~ { _1722_, _1722_, _1722_, _1722_, _1722_, _1722_ };
  assign _0342_ = ~ { _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_ };
  assign _0343_ = ~ { _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_ };
  assign _0344_ = ~ { _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_ };
  assign _0345_ = ~ { instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub };
  assign _0346_ = ~ { latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store };
  assign _0347_ = ~ { latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu };
  assign _0348_ = ~ { instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui, instr_lui };
  assign _0349_ = ~ { _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_ };
  assign _0350_ = ~ { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer };
  assign _0351_ = ~ { mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word };
  assign _0352_ = ~ { mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword };
  assign _0353_ = ~ { mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword };
  assign _0483_ = _0155_ & mem_rdata_word_t0;
  assign _0485_ = _0156_ & _1318_;
  assign _0487_ = _0157_ & _2044_;
  assign _0489_ = _0158_ & _1330_;
  assign _0491_ = _0159_ & _1324_;
  assign _0493_ = _0160_ & _1326_;
  assign _0495_ = _0161_ & _2046_;
  assign _0497_ = _0162_ & count_instr_t0[31:0];
  assign _0499_ = _0163_ & count_cycle_t0[31:0];
  assign _0501_ = _0164_ & _1334_;
  assign _1342_ = _0165_ & decoded_rd_t0;
  assign _0503_ = _0166_ & _2084_;
  assign _0505_ = _0158_ & _1371_;
  assign _0507_ = _0158_ & _1397_;
  assign _1395_ = _0167_ & cpuregs_rs2_t0;
  assign _0508_ = _0168_ & _1395_;
  assign _0510_ = _0157_ & _2109_;
  assign _0512_ = _0169_ & _1415_;
  assign _0514_ = _0170_ & _1401_;
  assign _0516_ = _0171_ & { pcpi_rs1_t0[30:0], 1'h0 };
  assign _0518_ = _0172_ & _1405_;
  assign _0520_ = _0171_ & { pcpi_rs1_t0[27:0], 4'h0 };
  assign _0522_ = _0172_ & _1409_;
  assign _1413_ = _0161_ & cpuregs_rs1_t0;
  assign _0524_ = _0173_ & _1413_;
  assign _0526_ = _0174_ & _0069_;
  assign _0528_ = _0175_ & _2011_;
  assign _1419_ = _0176_ & alu_add_sub_t0;
  assign _0530_ = _0177_ & _1419_;
  assign _0532_ = _0178_ & _1421_;
  assign _0534_ = _0179_ & _1427_;
  assign _0536_ = _0180_ & _1443_;
  assign _0538_ = _0182_ & _1433_;
  assign _0540_ = _0183_ & _2142_;
  assign _0542_ = _0184_ & _1439_;
  assign _0544_ = _0185_ & _1441_;
  assign _1445_ = _0186_ & _2180_;
  assign _1449_ = _0187_ & _1447_;
  assign _0546_ = _0188_ & _1449_;
  assign _0548_ = _0189_ & _1465_;
  assign _0550_ = _0191_ & _1455_;
  assign _0552_ = _0192_ & _2189_;
  assign _0554_ = _0193_ & _1461_;
  assign _0556_ = _0194_ & _1463_;
  assign _0558_ = _0196_ & { mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31:20] };
  assign _0560_ = _0197_ & _1480_;
  assign _0562_ = _0199_ & _1484_;
  assign _0564_ = _0200_ & _1486_;
  assign _0566_ = _0201_ & _2225_;
  assign _0568_ = _0203_ & _1492_;
  assign _0570_ = _0204_ & _2233_;
  assign _0572_ = _0206_ & _1498_;
  assign _0574_ = _0207_ & _2247_;
  assign _0576_ = _0208_ & _1504_;
  assign _0578_ = _0204_ & _1519_;
  assign _0580_ = _0206_ & _1510_;
  assign _0582_ = _0207_ & _2257_;
  assign _0584_ = _0210_ & _1517_;
  assign _0586_ = _0179_ & _2309_;
  assign _1528_ = _0211_ & _1526_;
  assign _0588_ = _0180_ & _1538_;
  assign _0590_ = _0181_ & _2309_;
  assign _0592_ = _0182_ & _1532_;
  assign _0595_ = _0212_ & _1536_;
  assign _0597_ = _0195_ & _2329_;
  assign _0599_ = _0213_ & _1540_;
  assign _0601_ = _0214_ & _2335_;
  assign _0603_ = _0207_ & _1544_;
  assign _0605_ = _0204_ & _1558_;
  assign _0607_ = _0205_ & _2335_;
  assign _0609_ = _0206_ & _1550_;
  assign _0611_ = _0207_ & _2343_;
  assign _0613_ = _0209_ & _2335_;
  assign _0615_ = _0210_ & _1556_;
  assign _0617_ = _0202_ & _2335_;
  assign _0619_ = _0214_ & _1560_;
  assign _1564_ = _0215_ & _2361_;
  assign _1566_ = _0216_ & _2353_;
  assign _0621_ = _0217_ & _1566_;
  assign _0623_ = _0218_ & _1581_;
  assign _0625_ = _0219_ & _2353_;
  assign _0627_ = _0220_ & _1572_;
  assign _0629_ = _0221_ & _2353_;
  assign _0631_ = _0222_ & _1577_;
  assign _1581_ = _0223_ & _1579_;
  assign _1584_ = _0215_ & _1566_;
  assign _0633_ = _0189_ & _2385_;
  assign _0635_ = _0190_ & _2381_;
  assign _0637_ = _0191_ & _1588_;
  assign _0639_ = _0224_ & _2397_;
  assign _1594_ = _0225_ & _2389_;
  assign _0641_ = _0226_ & _1594_;
  assign _0643_ = _0227_ & _1596_;
  assign _0645_ = _0228_ & _1612_;
  assign _0647_ = _0229_ & _2389_;
  assign _0649_ = _0230_ & _1602_;
  assign _0651_ = _0231_ & _2405_;
  assign _0653_ = _0232_ & _2389_;
  assign _0655_ = _0233_ & _1608_;
  assign _0657_ = _0234_ & _1610_;
  assign _0660_ = _0235_ & _1614_;
  assign _0662_ = _0236_ & { 24'h000000, mem_rdata_t0[23:16] };
  assign _0664_ = _0237_ & { 24'h000000, mem_rdata_t0[7:0] };
  assign _0666_ = _0238_ & _1620_;
  assign _0668_ = _0239_ & { 16'h0000, mem_rdata_t0[15:0] };
  assign _0670_ = _0240_ & mem_rdata_t0;
  assign _0672_ = _0241_ & _1622_;
  assign _0674_ = _0240_ & pcpi_rs2_t0;
  assign _0676_ = _0241_ & _1625_;
  assign _0678_ = _0242_ & pcpi_mul_rd_t0;
  assign _0680_ = _0243_ & _1851_;
  assign _0682_ = _0244_ & _1855_;
  assign _0684_ = _0244_ & _1859_;
  assign _0686_ = _0245_ & _1863_;
  assign _0688_ = _0245_ & _1867_;
  assign _0690_ = _0245_ & _1871_;
  assign _0692_ = _0245_ & _1875_;
  assign _0694_ = _0246_ & _1879_;
  assign _0696_ = _0246_ & _1883_;
  assign _0698_ = _0246_ & _1887_;
  assign _0700_ = _0246_ & _1891_;
  assign _0702_ = _0246_ & _1895_;
  assign _0704_ = _0246_ & _1899_;
  assign _0706_ = _0246_ & _1903_;
  assign _0708_ = _0246_ & _1907_;
  assign _0710_ = _0247_ & \cpuregs[0]_t0 ;
  assign _0712_ = _0247_ & \cpuregs[20]_t0 ;
  assign _0714_ = _0247_ & \cpuregs[22]_t0 ;
  assign _0716_ = _0247_ & \cpuregs[24]_t0 ;
  assign _0718_ = _0247_ & \cpuregs[26]_t0 ;
  assign _0720_ = _0247_ & \cpuregs[28]_t0 ;
  assign _0722_ = _0247_ & \cpuregs[30]_t0 ;
  assign _0724_ = _0247_ & \cpuregs[2]_t0 ;
  assign _0726_ = _0247_ & \cpuregs[4]_t0 ;
  assign _0728_ = _0247_ & \cpuregs[6]_t0 ;
  assign _0730_ = _0247_ & \cpuregs[8]_t0 ;
  assign _0732_ = _0247_ & \cpuregs[10]_t0 ;
  assign _0734_ = _0247_ & \cpuregs[12]_t0 ;
  assign _0736_ = _0247_ & \cpuregs[14]_t0 ;
  assign _0738_ = _0247_ & \cpuregs[16]_t0 ;
  assign _0740_ = _0247_ & \cpuregs[18]_t0 ;
  assign _0742_ = _0248_ & _1911_;
  assign _0744_ = _0249_ & _1915_;
  assign _0746_ = _0249_ & _1919_;
  assign _0748_ = _0250_ & _1923_;
  assign _0750_ = _0250_ & _1927_;
  assign _0752_ = _0250_ & _1931_;
  assign _0754_ = _0250_ & _1935_;
  assign _0756_ = _0251_ & _1939_;
  assign _0758_ = _0251_ & _1943_;
  assign _0760_ = _0251_ & _1947_;
  assign _0762_ = _0251_ & _1951_;
  assign _0764_ = _0251_ & _1955_;
  assign _0766_ = _0251_ & _1959_;
  assign _0768_ = _0251_ & _1963_;
  assign _0770_ = _0251_ & _1967_;
  assign _0772_ = _0252_ & \cpuregs[0]_t0 ;
  assign _0774_ = _0252_ & \cpuregs[20]_t0 ;
  assign _0776_ = _0252_ & \cpuregs[22]_t0 ;
  assign _0778_ = _0252_ & \cpuregs[24]_t0 ;
  assign _0780_ = _0252_ & \cpuregs[26]_t0 ;
  assign _0782_ = _0252_ & \cpuregs[28]_t0 ;
  assign _0784_ = _0252_ & \cpuregs[30]_t0 ;
  assign _0786_ = _0252_ & \cpuregs[2]_t0 ;
  assign _0788_ = _0252_ & \cpuregs[4]_t0 ;
  assign _0790_ = _0252_ & \cpuregs[6]_t0 ;
  assign _0792_ = _0252_ & \cpuregs[8]_t0 ;
  assign _0794_ = _0252_ & \cpuregs[10]_t0 ;
  assign _0796_ = _0252_ & \cpuregs[12]_t0 ;
  assign _0798_ = _0252_ & \cpuregs[14]_t0 ;
  assign _0800_ = _0252_ & \cpuregs[16]_t0 ;
  assign _0802_ = _0252_ & \cpuregs[18]_t0 ;
  assign _0807_ = _0254_ & reg_next_pc_t0;
  assign _2084_ = _0259_ & dbg_rs2val_t0;
  assign _0809_ = _0260_ & cpuregs_rs2_t0;
  assign _0811_ = _0255_ & _2084_;
  assign _2088_ = _0259_ & dbg_rs1val_t0;
  assign _0813_ = _0261_ & cpuregs_rs1_t0;
  assign _0815_ = _0166_ & _2088_;
  assign _0817_ = _0255_ & _2088_;
  assign _2103_ = _0262_ & _0081_;
  assign _2107_ = _0263_ & _0081_;
  assign _0819_ = _0264_ & _1407_;
  assign _2113_ = _0257_ & _2111_;
  assign _0821_ = _0198_ & _0073_;
  assign _0823_ = _0265_ & _0047_;
  assign _2125_ = _0267_ & _2123_;
  assign _0825_ = _0268_ & _2125_;
  assign _0827_ = _0269_ & _2127_;
  assign _2132_ = _0270_ & mem_rdata_latched_t0[11];
  assign _0829_ = _0271_ & _2138_;
  assign _0831_ = _0272_ & _2140_;
  assign _0833_ = _0273_ & mem_rdata_latched_t0[19];
  assign _0835_ = _0273_ & mem_rdata_latched_t0[30];
  assign _0837_ = _0273_ & mem_rdata_latched_t0[27];
  assign _0839_ = _0273_ & mem_rdata_latched_t0[26];
  assign _0841_ = _0274_ & mem_rdata_latched_t0[23:21];
  assign _0843_ = _0273_ & mem_rdata_latched_t0[25];
  assign _0845_ = _0275_ & mem_rdata_latched_t0[29:28];
  assign _0847_ = _0276_ & { mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31], mem_rdata_latched_t0[31] };
  assign _0849_ = _0273_ & mem_rdata_latched_t0[24];
  assign _0851_ = _0273_ & mem_rdata_latched_t0[20];
  assign _2176_ = _0277_ & _2174_;
  assign _0853_ = _0278_ & _2176_;
  assign _0855_ = _0279_ & _2178_;
  assign _2183_ = _0280_ & mem_rdata_latched_t0[10:7];
  assign _0857_ = _0281_ & _2185_;
  assign _0859_ = _0282_ & _2187_;
  assign _0861_ = _0283_ & mem_rdata_latched_t0[18:15];
  assign _0863_ = _0285_ & _2223_;
  assign _2227_ = _0286_ & mem_rdata_latched_t0[6:2];
  assign _0865_ = _0287_ & _2229_;
  assign _0867_ = _0288_ & mem_rdata_latched_t0[24:20];
  assign _0869_ = _0289_ & mem_rdata_latched_t0[19:12];
  assign _2243_ = _0290_ & _2241_;
  assign _0871_ = _0285_ & _2243_;
  assign _2249_ = _0286_ & mem_rdata_latched_t0[11:7];
  assign _0873_ = _0291_ & _2251_;
  assign _0875_ = _0287_ & _2253_;
  assign _0877_ = _0288_ & mem_rdata_latched_t0[11:7];
  assign _0879_ = _0292_ & decoded_rs2_t0;
  assign _0881_ = _0292_ & decoded_rs1_t0;
  assign _0883_ = _0293_ & _0049_;
  assign _0885_ = _0294_ & q_insn_rs2_t0;
  assign _0887_ = _0294_ & q_insn_rs1_t0;
  assign _0889_ = _0295_ & { rvfi_insn_t0[31:25], 5'h00, rvfi_insn_t0[19:15], 3'h0, rvfi_insn_t0[11:0] };
  assign _0891_ = _0296_ & { 16'h0000, next_insn_opcode_t0[15:0] };
  assign _2281_ = _0297_ & _2279_;
  assign _2283_ = _0298_ & mem_rdata_t0[31:16];
  assign _0893_ = _0299_ & _2281_;
  assign _0895_ = _0301_ & mem_wstrb_t0;
  assign _2299_ = _0302_ & _2297_;
  assign _0897_ = _0303_ & _2297_;
  assign _0899_ = _0122_ & mem_rdata_q_t0[31];
  assign _2311_ = _0304_ & _2309_;
  assign _2313_ = _0267_ & _2311_;
  assign _2315_ = _0268_ & _2313_;
  assign _2317_ = _0269_ & _2315_;
  assign _2319_ = _0305_ & _2309_;
  assign _2321_ = _0306_ & _2319_;
  assign _0901_ = _0271_ & _2321_;
  assign _2325_ = _0272_ & _2323_;
  assign _2327_ = _0211_ & _2309_;
  assign _0903_ = _0307_ & _2309_;
  assign _0905_ = _0122_ & mem_rdata_q_t0[7];
  assign _2331_ = _0284_ & _2329_;
  assign _0907_ = _0183_ & _2329_;
  assign _0909_ = _0307_ & _2329_;
  assign _0911_ = _0308_ & mem_rdata_q_t0[24:20];
  assign _2337_ = _0309_ & _2335_;
  assign _2339_ = _0290_ & _2337_;
  assign _0913_ = _0291_ & _2335_;
  assign _0915_ = _0310_ & { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] };
  assign _0917_ = _0311_ & _2335_;
  assign _0919_ = _0308_ & mem_rdata_q_t0[19:15];
  assign _0921_ = _0310_ & { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[6:5] };
  assign _0923_ = _0312_ & _2345_;
  assign _0925_ = _0313_ & _2345_;
  assign _0927_ = _0311_ & _2345_;
  assign _0929_ = _0314_ & mem_rdata_q_t0[14:12];
  assign _2355_ = _0315_ & _2353_;
  assign _2357_ = _0316_ & _2355_;
  assign _2359_ = _0317_ & _2357_;
  assign _2361_ = _0318_ & _2359_;
  assign _2363_ = _0319_ & _2353_;
  assign _2365_ = _0320_ & _2363_;
  assign _2367_ = _0321_ & _2365_;
  assign _2369_ = _0322_ & _2367_;
  assign _2371_ = _0323_ & _2369_;
  assign _2373_ = _0324_ & _2371_;
  assign _2375_ = _0325_ & _2373_;
  assign _0931_ = _0326_ & _2367_;
  assign _2379_ = _0327_ & mem_rdata_latched_t0[4:2];
  assign _0933_ = _0328_ & _2353_;
  assign _0935_ = _0329_ & mem_rdata_q_t0[11:8];
  assign _0937_ = _0186_ & _2381_;
  assign _0939_ = _0192_ & _2381_;
  assign _0942_ = _0330_ & _2381_;
  assign _0944_ = _0331_ & mem_rdata_q_t0[30:25];
  assign _2391_ = _0332_ & _2389_;
  assign _2393_ = _0333_ & _2391_;
  assign _2395_ = _0334_ & _2393_;
  assign _2397_ = _0335_ & _2395_;
  assign _2399_ = _0336_ & _2389_;
  assign _2401_ = _0337_ & _2399_;
  assign _0946_ = _0338_ & _2401_;
  assign _2405_ = _0339_ & _2403_;
  assign _0948_ = _0340_ & { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] };
  assign _0950_ = _0341_ & _2389_;
  assign _0952_ = _0342_ & _0041_;
  assign _0954_ = _0343_ & _0038_;
  assign _0958_ = _0344_ & reg_next_pc_t0;
  assign _0960_ = _0345_ & _0067_;
  assign _0962_ = _0346_ & reg_next_pc_t0;
  assign _0964_ = _0347_ & reg_out_t0;
  assign _2437_ = _0348_ & reg_pc_t0;
  assign _0966_ = _0349_ & { pcpi_rs1_t0[31:2], 2'h0 };
  assign _0968_ = _0350_ & mem_rdata_q_t0;
  assign _0970_ = _0351_ & _2444_;
  assign _0972_ = _0352_ & mem_rdata_latched_noshuffle_t0;
  assign _0974_ = _0353_ & _2442_;
  assign _0482_ = { _1692_, _1692_, _1692_, _1692_, _1692_ } & _2237_;
  assign _0484_ = { latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh, latched_is_lh } & { mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15], mem_rdata_word_t0[15:0] };
  assign _0486_ = { latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb, latched_is_lb } & { mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7], mem_rdata_word_t0[7:0] };
  assign _0488_ = { _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_ } & _2042_;
  assign _0490_ = { _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_ } & _2048_;
  assign _0492_ = { _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_, _1631_ } & _0079_;
  assign _0494_ = { _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_, _1177_ } & _1322_;
  assign _0496_ = { is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_rdcycle_rdcycleh_rdinstr_rdinstrh } & _1336_;
  assign _0498_ = { instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh, instr_rdinstrh } & count_instr_t0[63:32];
  assign _0500_ = { instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh, instr_rdcycleh } & count_cycle_t0[63:32];
  assign _0502_ = { _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_, _1178_ } & _1332_;
  assign _0504_ = { _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_ } & _2086_;
  assign _0506_ = { _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_, _1630_ } & cpuregs_rs2_t0;
  assign _0509_ = { _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_, _0443_ } & decoded_imm_t0;
  assign _0511_ = { _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_, _1634_ } & _2105_;
  assign _0513_ = { _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_, _1632_ } & _2113_;
  assign _0515_ = { _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_, _1184_ } & _1399_;
  assign _0517_ = { _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_ } & { 1'h0, pcpi_rs1_t0[31:1] };
  assign _0519_ = { _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_ } & { 1'h0, pcpi_rs1_t0[31:1] };
  assign _0521_ = { _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_, _1828_ } & { 4'h0, pcpi_rs1_t0[31:4] };
  assign _0523_ = { _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_, _1823_ } & { 1'h0, pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31], pcpi_rs1_t0[31:4] };
  assign _0525_ = { is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal, is_lui_auipc_jal } & _2437_;
  assign _0527_ = { _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_, _1687_ } & { _0093_[31:1], _2433_[0] };
  assign _0529_ = { _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_, _1826_ } & _0091_;
  assign _0531_ = { _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_, _1824_ } & _2449_;
  assign _0533_ = { _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_, _1185_ } & _1417_;
  assign _1427_ = _2133_ & _2132_;
  assign _0535_ = _2130_ & _2129_;
  assign _0537_ = _2134_ & _1429_;
  assign _1433_ = _2152_ & _2150_;
  assign _0539_ = _1186_ & _1431_;
  assign _0541_ = _0442_ & _0089_[4];
  assign _1439_ = _2133_ & mem_rdata_latched_t0[11];
  assign _0543_ = _2147_ & _2146_;
  assign _0545_ = _1187_ & _1437_;
  assign _1447_ = { _2133_, _2133_, _2133_, _2133_ } & _2183_;
  assign _0547_ = { _1188_, _1188_, _1188_, _1188_ } & _1445_;
  assign _0549_ = { _2134_, _2134_, _2134_, _2134_ } & _1451_;
  assign _1455_ = { _2152_, _2152_, _2152_, _2152_ } & _1468_;
  assign _0551_ = { _1186_, _1186_, _1186_, _1186_ } & _1453_;
  assign _0553_ = { _0442_, _0442_, _0442_, _0442_ } & _0089_[3:0];
  assign _1461_ = { _2133_, _2133_, _2133_, _2133_ } & mem_rdata_latched_t0[10:7];
  assign _0555_ = { _2147_, _2147_, _2147_, _2147_ } & _2193_;
  assign _0557_ = { _1187_, _1187_, _1187_, _1187_ } & _1459_;
  assign _1468_ = { _0441_, _0441_, _0441_, _0441_ } & _0089_[3:0];
  assign _0559_ = { is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu, is_beq_bne_blt_bge_bltu_bgeu } & { mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[7], mem_rdata_q_t0[30:25], mem_rdata_q_t0[11:8], 1'h0 };
  assign _0561_ = { is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw, is_sb_sh_sw } & { mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31], mem_rdata_q_t0[31:25], mem_rdata_q_t0[11:7] };
  assign _1484_ = { instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal } & { decoded_imm_j_t0[31:1], 1'h0 };
  assign _0563_ = { _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_, _2221_ } & { mem_rdata_q_t0[31:12], 12'h000 };
  assign _0565_ = { _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_, _0366_ } & _1482_;
  assign _0567_ = { _2136_, _2136_, _2136_, _2136_, _2136_ } & mem_rdata_latched_t0[6:2];
  assign _1492_ = { _2133_, _2133_, _2133_, _2133_, _2133_ } & _2227_;
  assign _0569_ = { _1188_, _1188_, _1188_, _1188_, _1188_ } & _1490_;
  assign _0571_ = { _2134_, _2134_, _2134_, _2134_, _2134_ } & _1494_;
  assign _1498_ = { _2152_, _2152_, _2152_, _2152_, _2152_ } & _2235_;
  assign _0573_ = { _1186_, _1186_, _1186_, _1186_, _1186_ } & _1496_;
  assign _0575_ = { _2130_, _2130_, _2130_, _2130_, _2130_ } & _2245_;
  assign _1504_ = { _2133_, _2133_, _2133_, _2133_, _2133_ } & _2249_;
  assign _0577_ = { _1190_, _1190_, _1190_, _1190_, _1190_ } & _1502_;
  assign _0579_ = { _2134_, _2134_, _2134_, _2134_, _2134_ } & _1506_;
  assign _1510_ = { _2152_, _2152_, _2152_, _2152_, _2152_ } & _2260_;
  assign _0581_ = { _1186_, _1186_, _1186_, _1186_, _1186_ } & _1508_;
  assign _0583_ = { _2130_, _2130_, _2130_, _2130_, _2130_ } & _2255_;
  assign _1517_ = { _0362_, _0362_, _0362_, _0362_, _0362_ } & mem_rdata_latched_t0[11:7];
  assign _0585_ = { _1189_, _1189_, _1189_, _1189_, _1189_ } & _1514_;
  assign _0587_ = _2130_ & _2317_;
  assign _0589_ = _2134_ & _1528_;
  assign _0591_ = _2152_ & _2327_;
  assign _0593_ = _1186_ & _1530_;
  assign _0594_ = _2130_ & _2325_;
  assign _0596_ = _0449_ & mem_rdata_latched_t0[12];
  assign _0598_ = _2148_ & _2333_;
  assign _0600_ = _0361_ & _2331_;
  assign _0602_ = { _2151_, _2151_, _2151_, _2151_, _2151_ } & { mem_rdata_latched_t0[6:4], 2'h0 };
  assign _0604_ = { _2130_, _2130_, _2130_, _2130_, _2130_ } & _2339_;
  assign _0606_ = { _2134_, _2134_, _2134_, _2134_, _2134_ } & _1546_;
  assign _0608_ = { _2152_, _2152_, _2152_, _2152_, _2152_ } & _1562_;
  assign _0610_ = { _1186_, _1186_, _1186_, _1186_, _1186_ } & _1548_;
  assign _0612_ = { _2130_, _2130_, _2130_, _2130_, _2130_ } & _2341_;
  assign _0614_ = { _0362_, _0362_, _0362_, _0362_, _0362_ } & mem_rdata_latched_t0[6:2];
  assign _0616_ = { _1189_, _1189_, _1189_, _1189_, _1189_ } & _1554_;
  assign _0618_ = { _2133_, _2133_, _2133_, _2133_, _2133_ } & { mem_rdata_latched_t0[11], mem_rdata_latched_t0[5], mem_rdata_latched_t0[6], 2'h0 };
  assign _0620_ = { _2151_, _2151_, _2151_, _2151_, _2151_ } & { mem_rdata_latched_t0[11:10], mem_rdata_latched_t0[6], 2'h0 };
  assign _0622_ = { _1192_, _1192_, _1192_ } & _1564_;
  assign _0624_ = { _2134_, _2134_, _2134_ } & _1568_;
  assign _0626_ = { _2152_, _2152_, _2152_ } & _1584_;
  assign _0628_ = { _1186_, _1186_, _1186_ } & _1570_;
  assign _0630_ = { _2147_, _2147_, _2147_ } & _2379_;
  assign _0632_ = { _2130_, _2130_, _2130_ } & _2377_;
  assign _0634_ = { _2134_, _2134_, _2134_, _2134_ } & _2383_;
  assign _0636_ = { _2152_, _2152_, _2152_, _2152_ } & _2387_;
  assign _0638_ = { _1186_, _1186_, _1186_, _1186_ } & _1586_;
  assign _0640_ = { _2136_, _2136_, _2136_, _2136_, _2136_, _2136_ } & { 3'h0, mem_rdata_latched_t0[8:7], mem_rdata_latched_t0[12] };
  assign _0642_ = { _2151_, _2151_, _2151_, _2151_, _2151_, _2151_ } & { 3'h0, mem_rdata_latched_t0[3:2], mem_rdata_latched_t0[12] };
  assign _0644_ = { _1188_, _1188_, _1188_, _1188_, _1188_, _1188_ } & _1592_;
  assign _0646_ = { _2134_, _2134_, _2134_, _2134_, _2134_, _2134_ } & _1598_;
  assign _0648_ = { _2152_, _2152_, _2152_, _2152_, _2152_, _2152_ } & _1616_;
  assign _0650_ = { _1186_, _1186_, _1186_, _1186_, _1186_, _1186_ } & _1600_;
  assign _0652_ = { _0442_, _0442_, _0442_, _0442_, _0442_, _0442_ } & { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[6:5], mem_rdata_latched_t0[2] };
  assign _0654_ = { _0362_, _0362_, _0362_, _0362_, _0362_, _0362_ } & { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] };
  assign _0656_ = { _2147_, _2147_, _2147_, _2147_, _2147_, _2147_ } & _2407_;
  assign _0658_ = { _1187_, _1187_, _1187_, _1187_, _1187_, _1187_ } & _1606_;
  assign _0659_ = { _2133_, _2133_, _2133_, _2133_, _2133_, _2133_ } & { 1'h0, mem_rdata_latched_t0[10:7], mem_rdata_latched_t0[12] };
  assign _0661_ = { _0441_, _0441_, _0441_, _0441_, _0441_, _0441_ } & { 4'h0, mem_rdata_latched_t0[5], mem_rdata_latched_t0[12] };
  assign _0663_ = { _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_, _2408_ } & { 24'h000000, mem_rdata_t0[31:24] };
  assign _0665_ = { _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_, _2410_ } & { 24'h000000, mem_rdata_t0[15:8] };
  assign _0667_ = { _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_ } & _1618_;
  assign _0669_ = { pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1], pcpi_rs1[1] } & { 16'h0000, mem_rdata_t0[31:16] };
  assign _0671_ = { _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_ } & _0036_;
  assign _0673_ = { _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_ } & _0051_;
  assign mem_la_wstrb_t0 = { _2411_, _2411_, _2411_, _2411_ } & _2426_;
  assign _0675_ = { _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_, _1637_ } & { pcpi_rs2_t0[15:0], pcpi_rs2_t0[15:0] };
  assign _0677_ = { _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_, _2411_ } & { pcpi_rs2_t0[7:0], pcpi_rs2_t0[7:0], pcpi_rs2_t0[7:0], pcpi_rs2_t0[7:0] };
  assign _0679_ = { pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready, pcpi_div_ready } & pcpi_div_rd_t0;
  assign _0681_ = { _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4], _0064_[4] } & _1853_;
  assign _0683_ = { _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3] } & _1857_;
  assign _0685_ = { _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3], _0064_[3] } & _1861_;
  assign _0687_ = { _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2] } & _1865_;
  assign _0689_ = { _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2] } & _1869_;
  assign _0691_ = { _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2] } & _1873_;
  assign _0693_ = { _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2], _0064_[2] } & _1877_;
  assign _0695_ = { _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1] } & _1881_;
  assign _0697_ = { _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1] } & _1885_;
  assign _0699_ = { _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1] } & _1889_;
  assign _0701_ = { _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1] } & _1893_;
  assign _0703_ = { _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1] } & _1897_;
  assign _0705_ = { _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1] } & _1901_;
  assign _0707_ = { _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1] } & _1905_;
  assign _0709_ = { _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1], _0064_[1] } & _1909_;
  assign _0711_ = { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] } & \cpuregs[1]_t0 ;
  assign _0713_ = { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] } & \cpuregs[21]_t0 ;
  assign _0715_ = { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] } & \cpuregs[23]_t0 ;
  assign _0717_ = { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] } & \cpuregs[25]_t0 ;
  assign _0719_ = { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] } & \cpuregs[27]_t0 ;
  assign _0721_ = { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] } & \cpuregs[29]_t0 ;
  assign _0723_ = { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] } & \cpuregs[31]_t0 ;
  assign _0725_ = { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] } & \cpuregs[3]_t0 ;
  assign _0727_ = { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] } & \cpuregs[5]_t0 ;
  assign _0729_ = { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] } & \cpuregs[7]_t0 ;
  assign _0731_ = { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] } & \cpuregs[9]_t0 ;
  assign _0733_ = { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] } & \cpuregs[11]_t0 ;
  assign _0735_ = { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] } & \cpuregs[13]_t0 ;
  assign _0737_ = { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] } & \cpuregs[15]_t0 ;
  assign _0739_ = { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] } & \cpuregs[17]_t0 ;
  assign _0741_ = { _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0], _0064_[0] } & \cpuregs[19]_t0 ;
  assign _0743_ = { _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4], _0065_[4] } & _1913_;
  assign _0745_ = { _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3] } & _1917_;
  assign _0747_ = { _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3], _0065_[3] } & _1921_;
  assign _0749_ = { _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2] } & _1925_;
  assign _0751_ = { _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2] } & _1929_;
  assign _0753_ = { _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2] } & _1933_;
  assign _0755_ = { _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2], _0065_[2] } & _1937_;
  assign _0757_ = { _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1] } & _1941_;
  assign _0759_ = { _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1] } & _1945_;
  assign _0761_ = { _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1] } & _1949_;
  assign _0763_ = { _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1] } & _1953_;
  assign _0765_ = { _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1] } & _1957_;
  assign _0767_ = { _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1] } & _1961_;
  assign _0769_ = { _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1] } & _1965_;
  assign _0771_ = { _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1], _0065_[1] } & _1969_;
  assign _0773_ = { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] } & \cpuregs[1]_t0 ;
  assign _0775_ = { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] } & \cpuregs[21]_t0 ;
  assign _0777_ = { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] } & \cpuregs[23]_t0 ;
  assign _0779_ = { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] } & \cpuregs[25]_t0 ;
  assign _0781_ = { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] } & \cpuregs[27]_t0 ;
  assign _0783_ = { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] } & \cpuregs[29]_t0 ;
  assign _0785_ = { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] } & \cpuregs[31]_t0 ;
  assign _0787_ = { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] } & \cpuregs[3]_t0 ;
  assign _0789_ = { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] } & \cpuregs[5]_t0 ;
  assign _0791_ = { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] } & \cpuregs[7]_t0 ;
  assign _0793_ = { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] } & \cpuregs[9]_t0 ;
  assign _0795_ = { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] } & \cpuregs[11]_t0 ;
  assign _0797_ = { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] } & \cpuregs[13]_t0 ;
  assign _0799_ = { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] } & \cpuregs[15]_t0 ;
  assign _0801_ = { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] } & \cpuregs[17]_t0 ;
  assign _0803_ = { _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0], _0065_[0] } & \cpuregs[19]_t0 ;
  assign rvfi_csr_minstret_rdata_t0 = { _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_ } & _0056_;
  assign rvfi_csr_mcycle_rdata_t0 = { _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_, _1706_ } & _0053_;
  assign _2015_ = { _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_ } & mem_wdata_t0;
  assign _2017_ = { _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_ } & mem_rdata_t0;
  assign _2019_ = { _1704_, _1704_, _1704_, _1704_ } & mem_wstrb_t0;
  assign _2022_ = { _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_, _1704_ } & mem_addr_t0;
  assign _2025_ = { cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write } & _2439_;
  assign _2029_ = { cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write, cpuregs_write } & latched_rd_t0;
  assign _0808_ = { latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch, latched_branch } & _2435_;
  assign _2033_ = { _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_ } & _2031_;
  assign _0047_ = { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn } & _2033_;
  assign _2040_ = { _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_, _1697_ } & _1320_;
  assign _2042_ = { _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_ } & _2040_;
  assign _2044_ = { _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_, _1635_ } & pcpi_rs1_t0;
  assign _2048_ = { instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap, instr_trap } & _2046_;
  assign _2046_ = { pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready, pcpi_int_ready } & pcpi_int_rd_t0;
  assign _0019_ = { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn } & _1328_;
  assign _0810_ = { _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_, _0357_ } & _2084_;
  assign _0812_ = { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn } & _1373_;
  assign _0814_ = { _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_, _0359_ } & _2088_;
  assign _0816_ = { _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_, _1629_ } & _2090_;
  assign _0818_ = { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn } & _2092_;
  assign _2105_ = { _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_ } & _2103_;
  assign _2109_ = { _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_, _1831_ } & _2107_;
  assign _0820_ = { _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_, _1685_ } & _1411_;
  assign _0822_ = { instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal, instr_jal } & _0077_;
  assign _0824_ = { decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger, decoder_trigger } & _2115_;
  assign _0002_ = { _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_, _1689_ } & cpuregs_wrdata_t0;
  assign cpuregs_wrdata_t0 = { _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_ } & _0027_;
  assign _2123_ = _1732_ & mem_rdata_latched_t0[11];
  assign _0826_ = _1726_ & mem_rdata_latched_t0[11];
  assign _0828_ = _1727_ & mem_rdata_latched_t0[11];
  assign _2138_ = _1730_ & _0089_[4];
  assign _0830_ = _1647_ & _0089_[4];
  assign _0832_ = _1648_ & _0089_[4];
  assign _2144_ = _1644_ & mem_rdata_latched_t0[11];
  assign _2146_ = _1847_ & _2144_;
  assign _2150_ = _0441_ & _0089_[4];
  assign _0834_ = _1729_ & _1435_;
  assign _0836_ = _1729_ & mem_rdata_latched_t0[8];
  assign _0838_ = _1729_ & mem_rdata_latched_t0[6];
  assign _0840_ = _1729_ & mem_rdata_latched_t0[7];
  assign _0842_ = { _1729_, _1729_, _1729_ } & mem_rdata_latched_t0[5:3];
  assign _0844_ = _1729_ & mem_rdata_latched_t0[2];
  assign _0846_ = { _1729_, _1729_ } & mem_rdata_latched_t0[10:9];
  assign _0848_ = { _1729_, _1729_, _1729_, _1729_, _1729_, _1729_, _1729_, _1729_, _1729_, _1729_, _1729_, _1729_ } & { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] };
  assign _0850_ = _1729_ & mem_rdata_latched_t0[11];
  assign _0852_ = _1729_ & mem_rdata_latched_t0[12];
  assign _2174_ = { _1732_, _1732_, _1732_, _1732_ } & mem_rdata_latched_t0[10:7];
  assign _0854_ = { _1726_, _1726_, _1726_, _1726_ } & mem_rdata_latched_t0[10:7];
  assign _0856_ = { _1727_, _1727_, _1727_, _1727_ } & mem_rdata_latched_t0[10:7];
  assign _2185_ = { _1730_, _1730_, _1730_, _1730_ } & _0089_[3:0];
  assign _0858_ = { _1647_, _1647_, _1647_, _1647_ } & _0089_[3:0];
  assign _0860_ = { _1648_, _1648_, _1648_, _1648_ } & _0089_[3:0];
  assign _2191_ = { _1644_, _1644_, _1644_, _1644_ } & mem_rdata_latched_t0[10:7];
  assign _2193_ = { _1847_, _1847_, _1847_, _1847_ } & _2191_;
  assign _0862_ = { _1729_, _1729_, _1729_, _1729_ } & _1457_;
  assign _2223_ = { _1724_, _1724_, _1724_, _1724_, _1724_ } & mem_rdata_latched_t0[6:2];
  assign _0864_ = { _1727_, _1727_, _1727_, _1727_, _1727_ } & mem_rdata_latched_t0[6:2];
  assign _2229_ = { _1730_, _1730_, _1730_, _1730_, _1730_ } & mem_rdata_latched_t0[6:2];
  assign _0866_ = { _1648_, _1648_, _1648_, _1648_, _1648_ } & _0087_[4:0];
  assign _2233_ = { _2130_, _2130_, _2130_, _2130_, _2130_ } & _2231_;
  assign _2235_ = { _2136_, _2136_, _2136_, _2136_, _2136_ } & _0087_[4:0];
  assign _0868_ = { _1729_, _1729_, _1729_, _1729_, _1729_ } & _1500_;
  assign _0870_ = { _1729_, _1729_, _1729_, _1729_, _1729_, _1729_, _1729_, _1729_ } & { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] };
  assign _2241_ = { _1724_, _1724_, _1724_, _1724_, _1724_ } & mem_rdata_latched_t0[11:7];
  assign _0872_ = { _1727_, _1727_, _1727_, _1727_, _1727_ } & mem_rdata_latched_t0[11:7];
  assign _2247_ = { _2008_, _2008_, _2008_, _2008_, _2008_ } & mem_rdata_latched_t0[11:7];
  assign _2251_ = { _1730_, _1730_, _1730_, _1730_, _1730_ } & _0089_[4:0];
  assign _0874_ = { _1647_, _1647_, _1647_, _1647_, _1647_ } & _0089_[4:0];
  assign _0876_ = { _1648_, _1648_, _1648_, _1648_, _1648_ } & _0089_[4:0];
  assign _2257_ = { _1847_, _1847_, _1847_, _1847_, _1847_ } & mem_rdata_latched_t0[11:7];
  assign _2260_ = { _0362_, _0362_, _0362_, _0362_, _0362_ } & _0087_[4:0];
  assign _0878_ = { _1729_, _1729_, _1729_, _1729_, _1729_ } & _1512_;
  assign _0880_ = { decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q } & cached_insn_rs2_t0;
  assign _0882_ = { decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q } & cached_insn_rs1_t0;
  assign _0884_ = { decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q, decoder_pseudo_trigger_q } & cached_insn_opcode_t0;
  assign _0886_ = { dbg_next, dbg_next, dbg_next, dbg_next, dbg_next } & _0034_;
  assign _0888_ = { dbg_next, dbg_next, dbg_next, dbg_next, dbg_next } & _0032_;
  assign _0890_ = { dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next, dbg_next } & _0030_;
  assign _0892_ = { _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_, _2277_ } & next_insn_opcode_t0;
  assign _2279_ = { _1846_, _1846_, _1846_, _1846_, _1846_, _1846_, _1846_, _1846_, _1846_, _1846_, _1846_, _1846_, _1846_, _1846_, _1846_, _1846_ } & mem_rdata_t0[31:16];
  assign _0894_ = { mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read } & _2283_;
  assign _0896_ = { _1845_, _1845_, _1845_, _1845_ } & _0095_;
  assign _0898_ = { _1814_, _1814_, _1814_, _1814_ } & _2299_;
  assign _0900_ = mem_xfer & mem_rdata_latched_t0[31];
  assign _0902_ = _1647_ & mem_rdata_latched_t0[12];
  assign _0904_ = _1722_ & _1534_;
  assign _0906_ = mem_xfer & mem_rdata_latched_t0[7];
  assign _0908_ = _0442_ & mem_rdata_latched_t0[12];
  assign _0910_ = _1722_ & _1542_;
  assign _0912_ = { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer } & mem_rdata_latched_t0[24:20];
  assign _0914_ = { _1647_, _1647_, _1647_, _1647_, _1647_ } & mem_rdata_latched_t0[6:2];
  assign _0916_ = { _1644_, _1644_, _1644_, _1644_, _1644_ } & { mem_rdata_latched_t0[6], 4'h0 };
  assign _0918_ = { _1722_, _1722_, _1722_, _1722_, _1722_ } & _1552_;
  assign _0920_ = { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer } & mem_rdata_latched_t0[19:15];
  assign _0922_ = { _1644_, _1644_, _1644_, _1644_, _1644_ } & _2345_;
  assign _0924_ = { _2147_, _2147_, _2147_, _2147_, _2147_ } & _2347_;
  assign _0926_ = { _2148_, _2148_, _2148_, _2148_, _2148_ } & _2349_;
  assign _0928_ = { _1722_, _1722_, _1722_, _1722_, _1722_ } & _2351_;
  assign _0930_ = { mem_xfer, mem_xfer, mem_xfer } & mem_rdata_latched_t0[14:12];
  assign _0932_ = { _1648_, _1648_, _1648_ } & _2375_;
  assign _0934_ = { _1722_, _1722_, _1722_ } & _1574_;
  assign _0936_ = { mem_xfer, mem_xfer, mem_xfer, mem_xfer } & mem_rdata_latched_t0[11:8];
  assign _0938_ = { _2136_, _2136_, _2136_, _2136_ } & { mem_rdata_latched_t0[11:9], 1'h0 };
  assign _0940_ = { _0442_, _0442_, _0442_, _0442_ } & { mem_rdata_latched_t0[11:10], mem_rdata_latched_t0[4:3] };
  assign _0941_ = { _2136_, _2136_, _2136_, _2136_ } & { mem_rdata_latched_t0[11:10], mem_rdata_latched_t0[6], 1'h0 };
  assign _0943_ = { _1722_, _1722_, _1722_, _1722_ } & _1590_;
  assign _0945_ = { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer } & mem_rdata_latched_t0[30:25];
  assign _0947_ = { _1647_, _1647_, _1647_, _1647_, _1647_, _1647_ } & { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[12] };
  assign _0949_ = { _1644_, _1644_, _1644_, _1644_, _1644_, _1644_ } & { mem_rdata_latched_t0[12], mem_rdata_latched_t0[12], mem_rdata_latched_t0[4:3], mem_rdata_latched_t0[5], mem_rdata_latched_t0[2] };
  assign _0951_ = { _1722_, _1722_, _1722_, _1722_, _1722_, _1722_ } & _1604_;
  assign _0953_ = { _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_, _1643_ } & { rvfi_rd_wdata_t0, 32'h00000000 };
  assign _0041_ = { _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_, _1642_ } & { 32'h00000000, rvfi_rd_wdata_t0 };
  assign _0955_ = { _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_, _1641_ } & { rvfi_rd_wdata_t0, 32'h00000000 };
  assign _0038_ = { _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_, _1640_ } & { 32'h00000000, rvfi_rd_wdata_t0 };
  assign _0959_ = { _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_, _1686_ } & { reg_out_t0[31:1], 1'h0 };
  assign _0961_ = { instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub, instr_sub } & _2428_;
  assign cpuregs_rs1_t0 = { _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_, _2416_ } & _2003_;
  assign cpuregs_rs2_t0 = { _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_, _2417_ } & _2005_;
  assign _0963_ = { latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store, latched_store } & { _0093_[31:1], 1'h0 };
  assign _0965_ = { latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu, latched_stalu } & alu_out_q_t0;
  assign _2439_ = { _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_, _2418_ } & cpuregs_wrdata_t0;
  assign _0967_ = { _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_, _1707_ } & { _0085_, 2'h0 };
  assign _0969_ = { mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer, mem_xfer } & mem_rdata_t0;
  assign _0971_ = { mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word, mem_la_use_prefetched_high_word } & { 16'h0000, mem_16bit_buffer_t0 };
  assign _0973_ = { mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword, mem_la_firstword } & { 16'h0000, mem_rdata_latched_noshuffle_t0[31:16] };
  assign _0975_ = { mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword, mem_la_secondword } & { mem_rdata_latched_noshuffle_t0[15:0], mem_16bit_buffer_t0 };
  assign _1318_ = _0483_ | _0484_;
  assign _1320_ = _0485_ | _0486_;
  assign _1322_ = _0487_ | _0488_;
  assign _1324_ = _0489_ | _0490_;
  assign _1326_ = _0491_ | _0492_;
  assign _1328_ = _0493_ | _0494_;
  assign _1330_ = _0495_ | _0496_;
  assign _1332_ = _0497_ | _0498_;
  assign _1334_ = _0499_ | _0500_;
  assign _1336_ = _0501_ | _0502_;
  assign _1371_ = _0503_ | _0504_;
  assign _1373_ = _0505_ | _0506_;
  assign _1393_ = _0507_ | _0506_;
  assign _1397_ = _0508_ | _0509_;
  assign _1399_ = _0510_ | _0511_;
  assign _1401_ = _0512_ | _0513_;
  assign _1403_ = _0514_ | _0515_;
  assign _1405_ = _0516_ | _0517_;
  assign _1407_ = _0518_ | _0519_;
  assign _1409_ = _0520_ | _0521_;
  assign _1411_ = _0522_ | _0523_;
  assign _1415_ = _0524_ | _0525_;
  assign _0027_ = _0526_ | _0527_;
  assign _1417_ = _0528_ | _0529_;
  assign _1421_ = _0530_ | _0531_;
  assign alu_out_t0 = _0532_ | _0533_;
  assign _1429_ = _0534_ | _0535_;
  assign _1431_ = _0536_ | _0537_;
  assign _1435_ = _0538_ | _0539_;
  assign _1437_ = _0540_ | _0541_;
  assign _1441_ = _0542_ | _0543_;
  assign _1443_ = _0544_ | _0545_;
  assign _1451_ = _0546_ | _0547_;
  assign _1453_ = _0548_ | _0549_;
  assign _1457_ = _0550_ | _0551_;
  assign _1459_ = _0552_ | _0553_;
  assign _1463_ = _0554_ | _0555_;
  assign _1465_ = _0556_ | _0557_;
  assign _1480_ = _0558_ | _0559_;
  assign _1482_ = _0560_ | _0561_;
  assign _1486_ = _0562_ | _0563_;
  assign _1488_ = _0564_ | _0565_;
  assign _1490_ = _0566_ | _0567_;
  assign _1494_ = _0568_ | _0569_;
  assign _1496_ = _0570_ | _0571_;
  assign _1500_ = _0572_ | _0573_;
  assign _1502_ = _0574_ | _0575_;
  assign _1506_ = _0576_ | _0577_;
  assign _1508_ = _0578_ | _0579_;
  assign _1512_ = _0580_ | _0581_;
  assign _1514_ = _0582_ | _0583_;
  assign _1519_ = _0584_ | _0585_;
  assign _1526_ = _0586_ | _0587_;
  assign _1530_ = _0588_ | _0589_;
  assign _1532_ = _0590_ | _0591_;
  assign _1534_ = _0592_ | _0593_;
  assign _1536_ = _0586_ | _0594_;
  assign _1538_ = _0595_ | _0596_;
  assign _1540_ = _0597_ | _0598_;
  assign _1542_ = _0599_ | _0600_;
  assign _1544_ = _0601_ | _0602_;
  assign _1546_ = _0603_ | _0604_;
  assign _1548_ = _0605_ | _0606_;
  assign _1550_ = _0607_ | _0608_;
  assign _1552_ = _0609_ | _0610_;
  assign _1554_ = _0611_ | _0612_;
  assign _1556_ = _0613_ | _0614_;
  assign _1558_ = _0615_ | _0616_;
  assign _1560_ = _0617_ | _0618_;
  assign _1562_ = _0619_ | _0620_;
  assign _1568_ = _0621_ | _0622_;
  assign _1570_ = _0623_ | _0624_;
  assign _1572_ = _0625_ | _0626_;
  assign _1574_ = _0627_ | _0628_;
  assign _1577_ = _0629_ | _0630_;
  assign _1579_ = _0631_ | _0632_;
  assign _1586_ = _0633_ | _0634_;
  assign _1588_ = _0635_ | _0636_;
  assign _1590_ = _0637_ | _0638_;
  assign _1592_ = _0639_ | _0640_;
  assign _1596_ = _0641_ | _0642_;
  assign _1598_ = _0643_ | _0644_;
  assign _1600_ = _0645_ | _0646_;
  assign _1602_ = _0647_ | _0648_;
  assign _1604_ = _0649_ | _0650_;
  assign _1606_ = _0651_ | _0652_;
  assign _1608_ = _0653_ | _0654_;
  assign _1610_ = _0655_ | _0656_;
  assign _1612_ = _0657_ | _0658_;
  assign _1614_ = _1594_ | _0659_;
  assign _1616_ = _0660_ | _0661_;
  assign _1618_ = _0662_ | _0663_;
  assign _1620_ = _0664_ | _0665_;
  assign _0051_ = _0666_ | _0667_;
  assign _0036_ = _0668_ | _0669_;
  assign _1622_ = _0670_ | _0671_;
  assign mem_rdata_word_t0 = _0672_ | _0673_;
  assign _1625_ = _0674_ | _0675_;
  assign mem_la_wdata_t0 = _0676_ | _0677_;
  assign pcpi_int_rd_t0 = _0678_ | _0679_;
  assign _2005_ = _0680_ | _0681_;
  assign _1851_ = _0682_ | _0683_;
  assign _1853_ = _0684_ | _0685_;
  assign _1855_ = _0686_ | _0687_;
  assign _1857_ = _0688_ | _0689_;
  assign _1859_ = _0690_ | _0691_;
  assign _1861_ = _0692_ | _0693_;
  assign _1863_ = _0694_ | _0695_;
  assign _1865_ = _0696_ | _0697_;
  assign _1867_ = _0698_ | _0699_;
  assign _1869_ = _0700_ | _0701_;
  assign _1871_ = _0702_ | _0703_;
  assign _1873_ = _0704_ | _0705_;
  assign _1875_ = _0706_ | _0707_;
  assign _1877_ = _0708_ | _0709_;
  assign _1879_ = _0710_ | _0711_;
  assign _1899_ = _0712_ | _0713_;
  assign _1901_ = _0714_ | _0715_;
  assign _1903_ = _0716_ | _0717_;
  assign _1905_ = _0718_ | _0719_;
  assign _1907_ = _0720_ | _0721_;
  assign _1909_ = _0722_ | _0723_;
  assign _1881_ = _0724_ | _0725_;
  assign _1883_ = _0726_ | _0727_;
  assign _1885_ = _0728_ | _0729_;
  assign _1887_ = _0730_ | _0731_;
  assign _1889_ = _0732_ | _0733_;
  assign _1891_ = _0734_ | _0735_;
  assign _1893_ = _0736_ | _0737_;
  assign _1895_ = _0738_ | _0739_;
  assign _1897_ = _0740_ | _0741_;
  assign _2003_ = _0742_ | _0743_;
  assign _1911_ = _0744_ | _0745_;
  assign _1913_ = _0746_ | _0747_;
  assign _1915_ = _0748_ | _0749_;
  assign _1917_ = _0750_ | _0751_;
  assign _1919_ = _0752_ | _0753_;
  assign _1921_ = _0754_ | _0755_;
  assign _1923_ = _0756_ | _0757_;
  assign _1925_ = _0758_ | _0759_;
  assign _1927_ = _0760_ | _0761_;
  assign _1929_ = _0762_ | _0763_;
  assign _1931_ = _0764_ | _0765_;
  assign _1933_ = _0766_ | _0767_;
  assign _1935_ = _0768_ | _0769_;
  assign _1937_ = _0770_ | _0771_;
  assign _1939_ = _0772_ | _0773_;
  assign _1959_ = _0774_ | _0775_;
  assign _1961_ = _0776_ | _0777_;
  assign _1963_ = _0778_ | _0779_;
  assign _1965_ = _0780_ | _0781_;
  assign _1967_ = _0782_ | _0783_;
  assign _1969_ = _0784_ | _0785_;
  assign _1941_ = _0786_ | _0787_;
  assign _1943_ = _0788_ | _0789_;
  assign _1945_ = _0790_ | _0791_;
  assign _1947_ = _0792_ | _0793_;
  assign _1949_ = _0794_ | _0795_;
  assign _1951_ = _0796_ | _0797_;
  assign _1953_ = _0798_ | _0799_;
  assign _1955_ = _0800_ | _0801_;
  assign _1957_ = _0802_ | _0803_;
  assign _2031_ = _0807_ | _0808_;
  assign _2086_ = _0809_ | _0810_;
  assign _0008_ = _0811_ | _0812_;
  assign _2090_ = _0813_ | _0814_;
  assign _2092_ = _0815_ | _0816_;
  assign _0005_ = _0817_ | _0818_;
  assign _2111_ = _0819_ | _0820_;
  assign _2115_ = _0821_ | _0822_;
  assign _2117_ = _0823_ | _0824_;
  assign _2127_ = _0825_ | _0826_;
  assign _2129_ = _0827_ | _0828_;
  assign _2140_ = _0829_ | _0830_;
  assign _2142_ = _0831_ | _0832_;
  assign _2154_ = _0833_ | _0834_;
  assign _2156_ = _0835_ | _0836_;
  assign _2158_ = _0837_ | _0838_;
  assign _2160_ = _0839_ | _0840_;
  assign _2162_ = _0841_ | _0842_;
  assign _2164_ = _0843_ | _0844_;
  assign _2166_ = _0845_ | _0846_;
  assign _2168_ = _0847_ | _0848_;
  assign _2170_ = _0849_ | _0850_;
  assign _2172_ = _0851_ | _0852_;
  assign _2178_ = _0853_ | _0854_;
  assign _2180_ = _0855_ | _0856_;
  assign _2187_ = _0857_ | _0858_;
  assign _2189_ = _0859_ | _0860_;
  assign _2195_ = _0861_ | _0862_;
  assign _2225_ = _0863_ | _0864_;
  assign _2231_ = _0865_ | _0866_;
  assign _2237_ = _0867_ | _0868_;
  assign _2239_ = _0869_ | _0870_;
  assign _2245_ = _0871_ | _0872_;
  assign _2253_ = _0873_ | _0874_;
  assign _2255_ = _0875_ | _0876_;
  assign _2262_ = _0877_ | _0878_;
  assign _0034_ = _0879_ | _0880_;
  assign _0032_ = _0881_ | _0882_;
  assign _0030_ = _0883_ | _0884_;
  assign dbg_insn_rs2_t0 = _0885_ | _0886_;
  assign dbg_insn_rs1_t0 = _0887_ | _0888_;
  assign dbg_insn_opcode_t0 = _0889_ | _0890_;
  assign _0049_ = _0891_ | _0892_;
  assign _2285_ = _0893_ | _0894_;
  assign _2297_ = _0895_ | _0896_;
  assign _2301_ = _0897_ | _0898_;
  assign _2309_ = _0899_ | _0900_;
  assign _2323_ = _0901_ | _0902_;
  assign _0015_[31] = _0903_ | _0904_;
  assign _2329_ = _0905_ | _0906_;
  assign _2333_ = _0907_ | _0908_;
  assign _0015_[7] = _0909_ | _0910_;
  assign _2335_ = _0911_ | _0912_;
  assign _2341_ = _0913_ | _0914_;
  assign _2343_ = _0915_ | _0916_;
  assign _0015_[24:20] = _0917_ | _0918_;
  assign _2345_ = _0919_ | _0920_;
  assign _2347_ = _0921_ | _0922_;
  assign _2349_ = _0923_ | _0924_;
  assign _2351_ = _0925_ | _0926_;
  assign _0015_[19:15] = _0927_ | _0928_;
  assign _2353_ = _0929_ | _0930_;
  assign _2377_ = _0931_ | _0932_;
  assign _0015_[14:12] = _0933_ | _0934_;
  assign _2381_ = _0935_ | _0936_;
  assign _2383_ = _0937_ | _0938_;
  assign _2385_ = _0939_ | _0940_;
  assign _2387_ = _0937_ | _0941_;
  assign _0015_[11:8] = _0942_ | _0943_;
  assign _2389_ = _0944_ | _0945_;
  assign _2403_ = _0946_ | _0947_;
  assign _2407_ = _0948_ | _0949_;
  assign _0015_[30:25] = _0950_ | _0951_;
  assign _0056_ = _0952_ | _0953_;
  assign _0053_ = _0954_ | _0955_;
  assign next_pc_t0 = _0958_ | _0959_;
  assign alu_add_sub_t0 = _0960_ | _0961_;
  assign _2435_ = _0962_ | _0963_;
  assign { _0093_[31:1], _2433_[0] } = _0964_ | _0965_;
  assign mem_la_addr_t0 = _0966_ | _0967_;
  assign mem_rdata_latched_noshuffle_t0 = _0968_ | _0969_;
  assign mem_rdata_latched_t0 = _0970_ | _0971_;
  assign _2442_ = _0972_ | _0973_;
  assign _2444_ = _0974_ | _0975_;
  assign _0372_ = | { _1846_, mem_la_read, mem_do_rdata };
  assign _0373_ = { mem_la_read, mem_do_rdata } != 2'h1;
  assign _0374_ = { mem_la_read, mem_la_use_prefetched_high_word } != 2'h3;
  assign _0375_ = { _1843_, resetn } != 2'h3;
  assign _0376_ = { _1655_, _1843_, mem_do_rinst } != 3'h4;
  assign _0377_ = { _1814_, _1843_, _1841_, mem_do_wdata } != 4'h8;
  assign _0378_ = { _2286_, _1843_, mem_xfer } != 3'h4;
  assign _0379_ = { _1654_, _1843_, mem_xfer } != 3'h4;
  assign _0380_ = { _2286_, _1843_, mem_la_read, mem_xfer } != 4'hb;
  assign _0381_ = | { _1814_, _1654_, _1655_, _2286_, _1843_ };
  assign _0382_ = | { _1841_, mem_do_wdata };
  assign _0383_ = { _1843_, _1844_ } != 2'h2;
  assign _0384_ = | { _1814_, _1654_, _2286_, _1843_ };
  assign _0385_ = | { _1629_, _1630_ };
  assign _0386_ = | { _1704_, mem_instr };
  assign _0387_ = { _1631_, is_beq_bne_blt_bge_bltu_bgeu } != 2'h2;
  assign _0388_ = | { _1628_, _1631_ };
  assign _0389_ = { _1634_, _1831_, mem_do_rdata } != 3'h7;
  assign _0390_ = { _1634_, _1831_ } != 2'h2;
  assign _0391_ = | { _1628_, _1634_ };
  assign _0392_ = { _1631_, is_beq_bne_blt_bge_bltu_bgeu } != 2'h3;
  assign _0393_ = { _1629_, is_rdcycle_rdcycleh_rdinstr_rdinstrh, instr_trap } != 3'h4;
  assign _0394_ = { _1630_, instr_trap } != 2'h2;
  assign _0395_ = | { _1629_, _1630_, _1628_, _1631_, _0444_ };
  assign _0396_ = | { _1835_, resetn };
  assign _0397_ = { _0443_, _1629_, _0450_, _1835_, _1696_, instr_trap, is_sll_srl_sra, resetn } != 8'h43;
  assign _0398_ = { _1630_, _1835_, is_sll_srl_sra, resetn } != 4'hb;
  assign _0399_ = { _1632_, _1835_, _1635_, resetn } != 4'h9;
  assign _0400_ = { _1629_, _0450_, _1835_, resetn } != 4'hd;
  assign _0401_ = { _1629_, _1630_, _1628_, _1632_, _1835_, resetn } != 6'h01;
  assign _0402_ = { _1633_, _1831_, mem_do_wdata } != 3'h7;
  assign _0403_ = { _1632_, _1823_, _1828_, _1827_, _1685_, _1635_ } != 6'h20;
  assign _0404_ = { _1632_, _1823_, _1685_, _1635_ } != 4'hc;
  assign _0405_ = { _1632_, _1823_, _1828_, _1827_, _1685_, _1635_ } != 6'h22;
  assign _0406_ = { _1632_, _1823_, _1685_, _1635_ } != 4'he;
  assign _0407_ = { _1632_, _1635_ } != 2'h3;
  assign _0408_ = { _1633_, _1831_ } != 2'h2;
  assign _0409_ = | { _1629_, _1632_, _1633_, _1634_ };
  assign _0410_ = { _1634_, _1833_, _1832_, _1831_, instr_lw, mem_do_rdata } != 6'h24;
  assign _0411_ = { _1633_, _1831_, instr_sw, instr_sh, instr_sb, mem_do_wdata } != 6'h30;
  assign _0412_ = | { _1628_, _1633_, _1634_ };
  assign _0413_ = | { cpuregs_write, rvfi_valid };
  assign _0414_ = { _0358_, instr_trap } != 2'h2;
  assign _0415_ = & { _2286_, _0373_, _0372_, _0374_, _0124_, mem_xfer };
  assign _0416_ = & { _0300_, _0253_, _2286_, mem_xfer };
  assign _0417_ = & { _2286_, mem_xfer };
  assign _0418_ = & { _0376_, _0375_, _0380_, _0381_, _0377_, _0378_, _0379_ };
  assign _0419_ = & { _0382_, _0124_, _1814_ };
  assign _0420_ = & { _0124_, _1845_ };
  assign _0421_ = & { _0377_, _0378_, _0379_, _0384_, _0383_ };
  assign _0422_ = & { _0124_, mem_la_write };
  assign _0423_ = & { _0388_, _0387_, resetn };
  assign _0424_ = & { _0391_, _0390_, _0389_ };
  assign _0425_ = & { _1628_, resetn };
  assign _0426_ = & { _0392_, _0388_ };
  assign _0427_ = & { _0395_, _0394_, _0393_ };
  assign _0428_ = & { _0401_, _0400_, _0399_, _0398_, _0397_, _0396_ };
  assign _0429_ = & { _0385_, resetn };
  assign _0430_ = & { _0409_, _0408_, _0407_, _0406_, _0405_, _0404_, _0403_, _0402_, _0390_, _0389_, resetn };
  assign _0431_ = & { _0409_, _0408_, _0407_, _0405_, _0403_, _0402_, _0390_, _0389_, resetn };
  assign _0432_ = & { _0412_, _0411_, _0410_, _0408_, _0402_, _0390_, _0389_, resetn };
  assign _0433_ = & { _0258_, _1628_, decoder_trigger, resetn };
  assign _0434_ = & { _1628_, decoder_trigger };
  assign _0435_ = & { _0414_, _0385_ };
  assign _0354_ = ~ dbg_rs1val_valid;
  assign _0436_ = | { _1843_, clear_prefetched_high_word };
  assign _0437_ = | { _0256_, _1733_ };
  assign _0438_ = | { _0256_, _2026_ };
  assign _0439_ = | { _0354_, _2013_, _2012_ };
  assign _0440_ = & { _1831_, _0453_, resetn };
  assign _0443_ = | { is_jalr_addi_slti_sltiu_xori_ori_andi, is_lui_auipc_jal };
  assign _0444_ = | { _1634_, _1632_ };
  assign _0445_ = | { _1696_, is_jalr_addi_slti_sltiu_xori_ori_andi, is_lui_auipc_jal, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle };
  assign _0446_ = | { _1634_, _1633_, _1632_, _1630_, _1629_, _1628_, _1627_ };
  assign _0447_ = | { _1634_, _1632_, _1631_, _1630_, _1629_, _1628_, _1627_ };
  assign _0448_ = | { _2269_, _2258_ };
  assign _0441_ = | { _2151_, _2136_ };
  assign _0442_ = | { _2136_, _2135_ };
  assign _0449_ = | { _2151_, _2147_, _2136_, _2135_, _2133_ };
  assign _0450_ = | { is_slli_srli_srai, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle };
  assign _0451_ = | { _1687_, latched_branch };
  assign _0452_ = | { _1696_, is_slli_srli_srai, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle };
  assign _0453_ = | { _1634_, _1633_ };
  assign _0355_ = ~ pcpi_rs1;
  assign _0356_ = ~ pcpi_rs2;
  assign _0804_ = pcpi_rs1_t0 & _0356_;
  assign _0805_ = pcpi_rs2_t0 & _0355_;
  assign _1173_ = _0804_ | _0805_;
  assign _2011_ = _1173_ | _0806_;
  assign _0358_ = | { _1630_, _1629_ };
  assign _0357_ = | { _1696_, is_jalr_addi_slti_sltiu_xori_ori_andi, is_slli_srli_srai, is_lui_auipc_jal, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle };
  assign _0359_ = | { is_lui_auipc_jal, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle };
  assign _0361_ = | { _2152_, _2134_ };
  assign _0362_ = | { _2151_, _2133_ };
  assign _0360_ = | { _2151_, _2136_, _2133_ };
  assign pcpi_int_ready = | { pcpi_div_ready, pcpi_mul_ready };
  assign _1177_ = _1632_ | _1634_;
  assign _1178_ = instr_rdinstr | instr_rdinstrh;
  assign _1179_ = _1631_ | _0444_;
  assign _1180_ = _1629_ | _1630_;
  assign _1182_ = _1630_ | _1632_;
  assign _1181_ = is_sb_sh_sw | is_sll_srl_sra;
  assign _1183_ = _0450_ | _0443_;
  assign _1184_ = _1633_ | _1634_;
  assign _1185_ = _1825_ | _1826_;
  assign _1190_ = _2151_ | _2130_;
  assign _1191_ = _1654_ | _1655_;
  assign _1189_ = _2147_ | _2130_;
  assign _1192_ = _2130_ | _0441_;
  assign _1193_ = _0360_ | _2135_;
  assign _1188_ = _2130_ | _2136_;
  assign _1186_ = _2148_ | _2134_;
  assign _1187_ = _2130_ | _0442_;
  assign _1194_ = _2409_ | _2408_;
  assign _0363_ = | { _1634_, _1633_, _1632_, _1631_ };
  assign _0364_ = | { _1696_, is_jalr_addi_slti_sltiu_xori_ori_andi, is_slli_srli_srai, is_lui_auipc_jal };
  assign _0365_ = | { is_sltiu_bltu_sltu, is_slti_blt_slt, instr_bgeu };
  assign _0366_ = | { is_alu_reg_imm, is_beq_bne_blt_bge_bltu_bgeu, is_sb_sh_sw, is_lb_lh_lw_lbu_lhu, instr_jalr };
  assign _0045_ = _0447_ ? 1'h0 : _0060_;
  assign _0043_ = _1634_ ? _0058_ : 1'h0;
  assign _0044_ = _0446_ ? 1'h0 : _0059_;
  assign _1315_ = _1631_ ? _2038_ : _1692_;
  assign _1316_ = _0453_ ? _2036_ : _1315_;
  assign _1317_ = latched_is_lh ? { mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15], mem_rdata_word[15:0] } : mem_rdata_word;
  assign _1319_ = latched_is_lb ? { mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7], mem_rdata_word[7:0] } : _1317_;
  assign _1321_ = _1634_ ? _2041_ : _2043_;
  assign _1323_ = _1630_ ? _2047_ : _1329_;
  assign _1325_ = _1631_ ? _0078_ : _1323_;
  assign _1327_ = _1177_ ? _1321_ : _1325_;
  assign _1329_ = is_rdcycle_rdcycleh_rdinstr_rdinstrh ? _1335_ : _2045_;
  assign _1331_ = instr_rdinstrh ? count_instr[63:32] : count_instr[31:0];
  assign _1333_ = instr_rdcycleh ? count_cycle[63:32] : count_cycle[31:0];
  assign _1335_ = _1178_ ? _1331_ : _1333_;
  assign _1337_ = _1630_ ? cpuregs_rs2[4:0] : _1340_;
  assign _1338_ = _1632_ ? _2050_ : _1337_;
  assign _1339_ = is_slli_srli_srai ? decoded_rs2 : cpuregs_rs2[4:0];
  assign _1340_ = _0445_ ? 5'hxx : _1339_;
  assign _1341_ = _1631_ ? _2053_ : decoded_rd;
  assign _1343_ = _1634_ ? _2055_ : 1'h0;
  assign _1344_ = _1634_ ? _2057_ : 1'h0;
  assign _1345_ = _1631_ ? _2058_ : _2060_;
  assign _1346_ = _1631_ ? _2061_ : 1'h0;
  assign _1347_ = _0444_ ? 1'h1 : _2062_;
  assign _1348_ = _1629_ ? _1351_ : 1'h0;
  assign _1349_ = _1630_ ? _2064_ : _1348_;
  assign _1350_ = _1179_ ? _1347_ : _1349_;
  assign _1351_ = is_rdcycle_rdcycleh_rdinstr_rdinstrh ? 1'h1 : _2063_;
  assign _1352_ = _1632_ ? _2067_ : _2069_;
  assign _1353_ = _0453_ ? _2066_ : _1352_;
  assign _1354_ = _1630_ ? _1360_ : _1367_;
  assign _1355_ = _1628_ ? _2073_ : cpu_state;
  assign _1356_ = _1180_ ? _1354_ : _1355_;
  assign _1357_ = _0363_ ? _1353_ : _1356_;
  assign _1358_ = is_sll_srl_sra ? 8'h04 : 8'h02;
  assign _1359_ = instr_trap ? _2071_ : 8'h08;
  assign _1360_ = _1181_ ? _1358_ : _1359_;
  assign _1361_ = is_sb_sh_sw ? 8'h02 : 8'h08;
  assign _1362_ = is_sll_srl_sra ? 8'h04 : _1361_;
  assign _1363_ = is_slli_srli_srai ? 8'h04 : 8'h01;
  assign _1364_ = _0443_ ? 8'h08 : _1363_;
  assign _1365_ = instr_trap ? _2071_ : _1362_;
  assign _1366_ = is_rdcycle_rdcycleh_rdinstr_rdinstrh ? 8'h40 : _1365_;
  assign _1367_ = _0364_ ? _1364_ : _1366_;
  assign _1368_ = _1629_ ? _2079_ : _2078_;
  assign _1369_ = _1630_ ? 1'h1 : _1368_;
  assign _1370_ = _1629_ ? _2085_ : _2083_;
  assign _1372_ = _1630_ ? cpuregs_rs2 : _1370_;
  assign _1374_ = _1632_ ? _2093_ : _1379_;
  assign _1375_ = _1629_ ? _1385_ : _2095_;
  assign _1376_ = _1182_ ? _1374_ : _1375_;
  assign _1377_ = is_sll_srl_sra ? 1'hx : 1'h1;
  assign _1378_ = instr_trap ? _2094_ : mem_do_prefetch;
  assign _1379_ = _1181_ ? _1377_ : _1378_;
  assign _1380_ = is_sb_sh_sw ? 1'h1 : mem_do_prefetch;
  assign _1381_ = is_sll_srl_sra ? 1'hx : _1380_;
  assign _1382_ = _0443_ ? mem_do_prefetch : 1'hx;
  assign _1383_ = instr_trap ? _2094_ : _1381_;
  assign _1384_ = _1696_ ? 1'h1 : _1383_;
  assign _1385_ = _1183_ ? _1382_ : _1384_;
  assign _1386_ = _1833_ ? 2'h1 : 2'h2;
  assign _1387_ = instr_lw ? 2'h0 : _1386_;
  assign _1388_ = _1633_ ? _2101_ : 2'h0;
  assign _1389_ = _1634_ ? _2099_ : _1388_;
  assign _1390_ = instr_sh ? 2'h1 : 2'h2;
  assign _1391_ = instr_sw ? 2'h0 : _1390_;
  assign _1392_ = _1630_ ? cpuregs_rs2 : _1396_;
  assign _1394_ = _0452_ ? 32'hxxxxxxxx : cpuregs_rs2;
  assign _1396_ = _0443_ ? decoded_imm : _1394_;
  assign _1398_ = _1634_ ? _2104_ : _2108_;
  assign _1400_ = _1632_ ? _2112_ : _1414_;
  assign _1402_ = _1184_ ? _1398_ : _1400_;
  assign _1404_ = _1828_ ? { 1'h0, pcpi_rs1[31:1] } : { pcpi_rs1[30:0], 1'h0 };
  assign _1406_ = _1823_ ? { 1'hx, pcpi_rs1[31:1] } : _1404_;
  assign _1408_ = _1828_ ? { 4'h0, pcpi_rs1[31:4] } : { pcpi_rs1[27:0], 4'h0 };
  assign _1410_ = _1823_ ? { 1'hx, pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31:4] } : _1408_;
  assign _1412_ = is_rdcycle_rdcycleh_rdinstr_rdinstrh ? 32'hxxxxxxxx : cpuregs_rs1;
  assign _1414_ = is_lui_auipc_jal ? _2436_ : _1412_;
  assign _0026_ = _1687_ ? { _0092_[31:1], _2432_[0] } : _0068_;
  assign _1416_ = _1826_ ? _0090_ : _2010_;
  assign _1418_ = is_compare ? { 31'h00000000, alu_out_0 } : alu_add_sub;
  assign _1420_ = _1824_ ? _2448_ : _1418_;
  assign alu_out = _1185_ ? _1416_ : _1420_;
  assign _1422_ = is_slti_blt_slt ? alu_lts : _1805_;
  assign _1423_ = is_sltiu_bltu_sltu ? alu_ltu : _1422_;
  assign _1424_ = instr_bne ? _1803_ : alu_eq;
  assign _1425_ = instr_bge ? _1804_ : _1424_;
  assign alu_out_0 = _0365_ ? _1423_ : _1425_;
  assign _1426_ = _2133_ ? _2131_ : 1'h0;
  assign _1428_ = _2130_ ? _2128_ : _1426_;
  assign _1430_ = _2134_ ? _1428_ : _1442_;
  assign _1432_ = _2152_ ? _2149_ : 1'h0;
  assign _1434_ = _1186_ ? _1430_ : _1432_;
  assign _1436_ = _0442_ ? _0088_[4] : _2141_;
  assign _1438_ = _2133_ ? mem_rdata_latched[11] : 1'h0;
  assign _1440_ = _2147_ ? _2145_ : _1438_;
  assign _1442_ = _1187_ ? _1436_ : _1440_;
  assign _1444_ = _2136_ ? 4'h2 : _2179_;
  assign _1446_ = _2133_ ? _2182_ : 4'h0;
  assign _1448_ = _2151_ ? _2181_ : _1446_;
  assign _1450_ = _1188_ ? _1444_ : _1448_;
  assign _1452_ = _2134_ ? _1450_ : _1464_;
  assign _1454_ = _2152_ ? _1467_ : 4'h0;
  assign _1456_ = _1186_ ? _1452_ : _1454_;
  assign _1458_ = _0442_ ? _0088_[3:0] : _2188_;
  assign _1460_ = _2133_ ? mem_rdata_latched[10:7] : 4'h0;
  assign _1462_ = _2147_ ? _2192_ : _1460_;
  assign _1464_ = _1187_ ? _1458_ : _1462_;
  assign _1466_ = _2133_ ? 4'h2 : 4'h0;
  assign _1467_ = _0441_ ? _0088_[3:0] : _1466_;
  assign _1469_ = _2148_ ? _2200_ : _1665_;
  assign _1470_ = _2134_ ? _2198_ : _1469_;
  assign _1471_ = _2134_ ? _2203_ : _1476_;
  assign _1472_ = _2152_ ? _2208_ : _1664_;
  assign _1473_ = _1186_ ? _1471_ : _1472_;
  assign _1474_ = _2130_ ? _2205_ : _2207_;
  assign _1475_ = _0362_ ? 1'h1 : _1664_;
  assign _1476_ = _1189_ ? _1474_ : _1475_;
  assign _1477_ = _2152_ ? _2218_ : _1662_;
  assign _1478_ = _2134_ ? _2217_ : _1477_;
  assign _1479_ = is_beq_bne_blt_bge_bltu_bgeu ? { mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[7], mem_rdata_q[30:25], mem_rdata_q[11:8], 1'h0 } : { mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31:20] };
  assign _1481_ = is_sb_sh_sw ? { mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31], mem_rdata_q[31:25], mem_rdata_q[11:7] } : _1479_;
  assign _1483_ = instr_jal ? { decoded_imm_j[31:1], 1'h0 } : 32'b0000000000000000000000000000000x;
  assign _1485_ = _2221_ ? { mem_rdata_q[31:12], 12'h000 } : _1483_;
  assign _1487_ = _0366_ ? _1481_ : _1485_;
  assign _1489_ = _2136_ ? mem_rdata_latched[6:2] : _2224_;
  assign _1491_ = _2133_ ? _2226_ : 5'h00;
  assign _1493_ = _1188_ ? _1489_ : _1491_;
  assign _1495_ = _2134_ ? _1493_ : _2232_;
  assign _1497_ = _2152_ ? _2234_ : 5'h00;
  assign _1499_ = _1186_ ? _1495_ : _1497_;
  assign _1501_ = _2130_ ? _2244_ : _2246_;
  assign _1503_ = _2133_ ? _2248_ : 5'h00;
  assign _1505_ = _1190_ ? _1501_ : _1503_;
  assign _1507_ = _2134_ ? _1505_ : _1518_;
  assign _1509_ = _2152_ ? _2259_ : 5'h00;
  assign _1511_ = _1186_ ? _1507_ : _1509_;
  assign _1513_ = _2130_ ? _2254_ : _2256_;
  assign _1515_ = _2258_ ? 5'h01 : 5'h00;
  assign _1516_ = _0362_ ? mem_rdata_latched[11:7] : _1515_;
  assign _1518_ = _1189_ ? _1513_ : _1516_;
  assign _1520_ = _1655_ ? _2289_ : _2290_;
  assign _1521_ = _2286_ ? _2292_ : _2294_;
  assign _1522_ = _1191_ ? _1520_ : _1521_;
  assign _1523_ = _2286_ ? _2304_ : _2306_;
  assign _1524_ = _1654_ ? _2303_ : _1523_;
  assign _1525_ = _2130_ ? _2316_ : _2308_;
  assign _1527_ = _0360_ ? 1'h0 : _1525_;
  assign _1529_ = _2134_ ? _1527_ : _1537_;
  assign _1531_ = _2152_ ? _2326_ : _2308_;
  assign _1533_ = _1186_ ? _1529_ : _1531_;
  assign _1535_ = _2130_ ? _2324_ : _2308_;
  assign _1537_ = _0449_ ? mem_rdata_latched[12] : _1535_;
  assign _1539_ = _2148_ ? _2332_ : _2328_;
  assign _1541_ = _0361_ ? _2330_ : _1539_;
  assign _1543_ = _2151_ ? { mem_rdata_latched[6:4], 2'h0 } : _2334_;
  assign _1545_ = _2130_ ? _2338_ : _1543_;
  assign _1547_ = _2134_ ? _1545_ : _1557_;
  assign _1549_ = _2152_ ? _1561_ : _2334_;
  assign _1551_ = _1186_ ? _1547_ : _1549_;
  assign _1553_ = _2130_ ? _2340_ : _2342_;
  assign _1555_ = _0362_ ? mem_rdata_latched[6:2] : _2334_;
  assign _1557_ = _1189_ ? _1553_ : _1555_;
  assign _1559_ = _2133_ ? { mem_rdata_latched[11], mem_rdata_latched[5], mem_rdata_latched[6], 2'h0 } : _2334_;
  assign _1561_ = _2151_ ? { mem_rdata_latched[11:10], mem_rdata_latched[6], 2'h0 } : _1559_;
  assign _1563_ = _0441_ ? 3'h2 : _2360_;
  assign _1565_ = _2133_ ? 3'h1 : _2352_;
  assign _1567_ = _1192_ ? _1563_ : _1565_;
  assign _1569_ = _2134_ ? _1567_ : _1580_;
  assign _1571_ = _2152_ ? _1583_ : _2352_;
  assign _1573_ = _1186_ ? _1569_ : _1571_;
  assign _1575_ = _2135_ ? 3'h1 : 3'h0;
  assign _1576_ = _2147_ ? _2378_ : _2352_;
  assign _1578_ = _2130_ ? _2376_ : _1576_;
  assign _1580_ = _1193_ ? _1575_ : _1578_;
  assign _1582_ = _2133_ ? 3'h0 : _2352_;
  assign _1583_ = _0441_ ? 3'h2 : _1582_;
  assign _1585_ = _2134_ ? _2382_ : _2384_;
  assign _1587_ = _2152_ ? _2386_ : _2380_;
  assign _1589_ = _1186_ ? _1585_ : _1587_;
  assign _1591_ = _2136_ ? { 3'h0, mem_rdata_latched[8:7], mem_rdata_latched[12] } : _2396_;
  assign _1593_ = _2133_ ? 6'h00 : _2388_;
  assign _1595_ = _2151_ ? { 3'h0, mem_rdata_latched[3:2], mem_rdata_latched[12] } : _1593_;
  assign _1597_ = _1188_ ? _1591_ : _1595_;
  assign _1599_ = _2134_ ? _1597_ : _1611_;
  assign _1601_ = _2152_ ? _1615_ : _2388_;
  assign _1603_ = _1186_ ? _1599_ : _1601_;
  assign _1605_ = _0442_ ? { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[6:5], mem_rdata_latched[2] } : _2404_;
  assign _1607_ = _0362_ ? { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] } : _2388_;
  assign _1609_ = _2147_ ? _2406_ : _1607_;
  assign _1611_ = _1187_ ? _1605_ : _1609_;
  assign _1613_ = _2133_ ? { 1'h0, mem_rdata_latched[10:7], mem_rdata_latched[12] } : _2388_;
  assign _1615_ = _0441_ ? { 4'h0, mem_rdata_latched[5], mem_rdata_latched[12] } : _1613_;
  assign _1617_ = _2408_ ? { 24'h000000, mem_rdata[31:24] } : { 24'h000000, mem_rdata[23:16] };
  assign _1619_ = _2410_ ? { 24'h000000, mem_rdata[15:8] } : { 24'h000000, mem_rdata[7:0] };
  assign _0050_ = _1194_ ? _1617_ : _1619_;
  assign _0035_ = pcpi_rs1[1] ? { 16'h0000, mem_rdata[31:16] } : { 16'h0000, mem_rdata[15:0] };
  assign _1621_ = _1637_ ? _0035_ : mem_rdata;
  assign mem_rdata_word = _2411_ ? _0050_ : _1621_;
  assign _1623_ = _1637_ ? _2445_ : 4'hf;
  assign mem_la_wstrb = _2411_ ? _2425_ : _1623_;
  assign _1624_ = _1637_ ? { pcpi_rs2[15:0], pcpi_rs2[15:0] } : pcpi_rs2;
  assign mem_la_wdata = _2411_ ? { pcpi_rs2[7:0], pcpi_rs2[7:0], pcpi_rs2[7:0], pcpi_rs2[7:0] } : _1624_;
  assign pcpi_int_rd = pcpi_div_ready ? pcpi_div_rd : pcpi_mul_rd;
  assign _1626_ = pcpi_mul_ready ? pcpi_mul_wr : 1'h0;
  assign pcpi_int_wr = pcpi_div_ready ? pcpi_div_wr : _1626_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME count_cycle_t0 */
  always_ff @(posedge clk)
    if (!resetn) count_cycle_t0 <= 64'h0000000000000000;
    else count_cycle_t0 <= _0071_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rs2_rdata_t0 */
  always_ff @(posedge clk)
    if (!dbg_rs2val_valid) rvfi_rs2_rdata_t0 <= 32'd0;
    else rvfi_rs2_rdata_t0 <= dbg_rs2val_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rs1_rdata_t0 */
  always_ff @(posedge clk)
    if (_0439_) rvfi_rs1_rdata_t0 <= 32'd0;
    else rvfi_rs1_rdata_t0 <= dbg_rs1val_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rs2_addr_t0 */
  always_ff @(posedge clk)
    if (!dbg_rs2val_valid) rvfi_rs2_addr_t0 <= 5'h00;
    else rvfi_rs2_addr_t0 <= dbg_insn_rs2_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rs1_addr_t0 */
  always_ff @(posedge clk)
    if (_0439_) rvfi_rs1_addr_t0 <= 5'h00;
    else rvfi_rs1_addr_t0 <= dbg_insn_rs1_t0;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_order_t0 */
  always_ff @(posedge clk)
    if (!resetn) rvfi_order_t0 <= 64'h0000000000000000;
    else rvfi_order_t0 <= _0083_;
  assign _0367_ = ~ _0419_;
  assign _0368_ = ~ _0386_;
  assign _1079_ = { _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_ } & _2015_;
  assign _1097_ = { _0386_, _0386_, _0386_, _0386_ } & _2019_;
  assign _1106_ = { _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_ } & _2017_;
  assign _1108_ = { _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_, _0386_ } & _2022_;
  assign _1119_ = launch_next_insn & reg_next_pc_t0[0];
  assign _1046_ = _0367_ & mem_instr_t0;
  assign _1080_ = { _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_ } & rvfi_mem_wdata_t0;
  assign _1098_ = { _0368_, _0368_, _0368_, _0368_ } & rvfi_mem_wmask_t0;
  assign _1099_ = { _0368_, _0368_, _0368_, _0368_ } & rvfi_mem_rmask_t0;
  assign _1107_ = { _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_ } & rvfi_mem_rdata_t0;
  assign _1109_ = { _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_, _0368_ } & rvfi_mem_addr_t0;
  assign _1120_ = _0136_ & rvfi_pc_wdata_t0[0];
  assign _1232_ = _1079_ | _1080_;
  assign _1241_ = _1097_ | _1098_;
  assign _1245_ = _1106_ | _1107_;
  assign _1246_ = _1108_ | _1109_;
  assign _1251_ = _1119_ | _1120_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME mem_instr_t0 */
  always_ff @(posedge clk)
    if (mem_do_wdata) mem_instr_t0 <= 1'h0;
    else mem_instr_t0 <= _1046_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_wdata_t0 */
  always_ff @(posedge clk)
    if (mem_instr) rvfi_mem_wdata_t0 <= 32'd0;
    else rvfi_mem_wdata_t0 <= _1232_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_wmask_t0 */
  always_ff @(posedge clk)
    if (mem_instr) rvfi_mem_wmask_t0 <= 4'h0;
    else rvfi_mem_wmask_t0 <= _1241_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_rmask_t0 */
  always_ff @(posedge clk)
    if (mem_instr) rvfi_mem_rmask_t0 <= 4'h0;
    else rvfi_mem_rmask_t0 <= _1099_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_rdata_t0 */
  always_ff @(posedge clk)
    if (mem_instr) rvfi_mem_rdata_t0 <= 32'd0;
    else rvfi_mem_rdata_t0 <= _1245_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_mem_addr_t0 */
  always_ff @(posedge clk)
    if (mem_instr) rvfi_mem_addr_t0 <= 32'd0;
    else rvfi_mem_addr_t0 <= _1246_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_pc_wdata_t0[0] */
  always_ff @(posedge clk)
    if (_1686_) rvfi_pc_wdata_t0[0] <= 1'h0;
    else rvfi_pc_wdata_t0[0] <= _1251_;
  assign _0369_ = ~ _0413_;
  assign _0370_ = ~ _0434_;
  assign _0371_ = ~ _0435_;
  assign _1093_ = { _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_ } & _0047_;
  assign _1095_ = { _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_, _1628_ } & _2117_;
  assign _1110_ = { _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_ } & _2025_;
  assign _1112_ = { _0413_, _0413_, _0413_, _0413_, _0413_ } & _2029_;
  assign _1116_ = { _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_ } & _0075_;
  assign _1094_ = { _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_ } & reg_pc_t0;
  assign _1096_ = { _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_, _0266_ } & reg_next_pc_t0;
  assign _1111_ = { _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_, _0369_ } & rvfi_rd_wdata_t0;
  assign _1113_ = { _0369_, _0369_, _0369_, _0369_, _0369_ } & rvfi_rd_addr_t0;
  assign _1117_ = { _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_, _0370_ } & count_instr_t0;
  assign _1118_ = _0371_ & pcpi_valid_t0;
  assign _1239_ = _1093_ | _1094_;
  assign _1240_ = _1095_ | _1096_;
  assign _1247_ = _1110_ | _1111_;
  assign _1248_ = _1112_ | _1113_;
  assign _1250_ = _1116_ | _1117_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME reg_pc_t0 */
  always_ff @(posedge clk)
    if (!resetn) reg_pc_t0 <= 32'd0;
    else reg_pc_t0 <= _1239_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME reg_next_pc_t0 */
  always_ff @(posedge clk)
    if (!resetn) reg_next_pc_t0 <= 32'd0;
    else reg_next_pc_t0 <= _1240_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rd_wdata_t0 */
  always_ff @(posedge clk)
    if (_0438_) rvfi_rd_wdata_t0 <= 32'd0;
    else rvfi_rd_wdata_t0 <= _1247_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_rd_addr_t0 */
  always_ff @(posedge clk)
    if (_0438_) rvfi_rd_addr_t0 <= 5'h00;
    else rvfi_rd_addr_t0 <= _1248_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME count_instr_t0 */
  always_ff @(posedge clk)
    if (!resetn) count_instr_t0 <= 64'h0000000000000000;
    else count_instr_t0 <= _1250_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME pcpi_valid_t0 */
  always_ff @(posedge clk)
    if (!resetn) pcpi_valid_t0 <= 1'h0;
    else pcpi_valid_t0 <= _1118_;
  assign _2426_ = 4'h0 << pcpi_rs1[1:0];
  assign _1311_ = _1174_ - _0957_;
  assign _1312_ = _0956_ - _1175_;
  assign _1271_ = _1311_ ^ _1312_;
  assign _1176_ = _1271_ | pcpi_rs1_t0;
  assign _2428_ = _1176_ | pcpi_rs2_t0;
  assign _2449_ = pcpi_rs1_t0 | pcpi_rs2_t0;
  assign alu_eq = pcpi_rs1 == /* src = "generated/out/vanilla.sv:1111.14-1111.32" */ pcpi_rs2;
  assign _1635_ = ! /* src = "generated/out/vanilla.sv:1579.10-1579.21" */ reg_sh;
  assign _1638_ = rvfi_insn[6:0] == /* src = "generated/out/vanilla.sv:1792.23-1792.51" */ 7'h73;
  assign _1639_ = rvfi_insn[13:12] == /* src = "generated/out/vanilla.sv:1792.58-1792.84" */ 2'h2;
  assign _1640_ = rvfi_insn[31:20] == /* src = "generated/out/vanilla.sv:1793.8-1793.35" */ 12'hc00;
  assign _1641_ = rvfi_insn[31:20] == /* src = "generated/out/vanilla.sv:1797.8-1797.35" */ 12'hc80;
  assign _1642_ = rvfi_insn[31:20] == /* src = "generated/out/vanilla.sv:1801.8-1801.35" */ 12'hc02;
  assign _1643_ = rvfi_insn[31:20] == /* src = "generated/out/vanilla.sv:1805.8-1805.35" */ 12'hc82;
  assign _1645_ = ! /* src = "generated/out/vanilla.sv:379.12-379.45" */ mem_rdata_latched[11:10];
  assign _1646_ = mem_rdata_latched[11:10] == /* src = "generated/out/vanilla.sv:383.12-383.45" */ 2'h1;
  assign _1650_ = mem_rdata_latched[6:5] == /* src = "generated/out/vanilla.sv:394.13-394.44" */ 2'h1;
  assign _1651_ = mem_rdata_latched[6:5] == /* src = "generated/out/vanilla.sv:396.13-396.44" */ 2'h2;
  assign _1652_ = mem_rdata_latched[6:5] == /* src = "generated/out/vanilla.sv:398.13-398.44" */ 2'h3;
  assign _1649_ = ! /* src = "generated/out/vanilla.sv:400.32-400.63" */ mem_rdata_latched[6:5];
  assign _1656_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:797.17-797.53" */ 7'h37;
  assign _1657_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:798.19-798.55" */ 7'h17;
  assign _1658_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:799.17-799.53" */ 7'h6f;
  assign _1659_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:800.19-800.55" */ 7'h67;
  assign _1660_ = ! /* src = "generated/out/vanilla.sv:800.61-800.95" */ mem_rdata_latched[14:12];
  assign _1661_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:803.36-803.72" */ 7'h63;
  assign _1662_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:804.27-804.63" */ 7'h03;
  assign _1663_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:805.19-805.55" */ 7'h23;
  assign _1664_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:806.22-806.58" */ 7'h13;
  assign _1665_ = mem_rdata_latched[6:0] == /* src = "generated/out/vanilla.sv:807.22-807.58" */ 7'h33;
  assign _1644_ = mem_rdata_latched[11:7] == /* src = "generated/out/vanilla.sv:860.14-860.42" */ 5'h02;
  assign _1647_ = mem_rdata_latched[11:10] == /* src = "generated/out/vanilla.sv:877.13-877.46" */ 2'h2;
  assign _1648_ = mem_rdata_latched[12:10] == /* src = "generated/out/vanilla.sv:882.13-882.47" */ 3'h3;
  assign _1653_ = ! /* src = "generated/out/vanilla.sv:928.82-928.109" */ mem_rdata_latched[6:2];
  assign _1677_ = mem_rdata_q[31:20] == /* src = "generated/out/vanilla.sv:984.61-984.97" */ 12'hb00;
  assign _1678_ = mem_rdata_q[31:20] == /* src = "generated/out/vanilla.sv:984.174-984.210" */ 12'hb01;
  assign _1679_ = mem_rdata_q[31:20] == /* src = "generated/out/vanilla.sv:985.63-985.99" */ 12'hb80;
  assign _1680_ = mem_rdata_q[31:20] == /* src = "generated/out/vanilla.sv:985.176-985.212" */ 12'hb81;
  assign _1681_ = mem_rdata_q[31:20] == /* src = "generated/out/vanilla.sv:986.60-986.96" */ 12'hb02;
  assign _1682_ = mem_rdata_q[31:20] == /* src = "generated/out/vanilla.sv:987.62-987.98" */ 12'hb82;
  assign _1676_ = mem_rdata_q[6:0] == /* src = "generated/out/vanilla.sv:988.29-988.59" */ 7'h73;
  assign _1683_ = mem_rdata_q[15:0] == /* src = "generated/out/vanilla.sv:988.131-988.160" */ 16'h9002;
  assign _1684_ = mem_rdata_q[6:0] == /* src = "generated/out/vanilla.sv:989.20-989.50" */ 7'h0f;
  assign _1671_ = mem_rdata_q[14:12] == /* src = "generated/out/vanilla.sv:995.230-995.258" */ 3'h7;
  assign _1670_ = mem_rdata_q[14:12] == /* src = "generated/out/vanilla.sv:995.200-995.228" */ 3'h6;
  assign _1668_ = mem_rdata_q[14:12] == /* src = "generated/out/vanilla.sv:995.170-995.198" */ 3'h4;
  assign _1673_ = mem_rdata_q[14:12] == /* src = "generated/out/vanilla.sv:995.140-995.168" */ 3'h3;
  assign _1672_ = mem_rdata_q[14:12] == /* src = "generated/out/vanilla.sv:995.110-995.138" */ 3'h2;
  assign _1666_ = ! /* src = "generated/out/vanilla.sv:995.80-995.108" */ mem_rdata_q[14:12];
  assign _1675_ = mem_rdata_q[31:25] == /* src = "generated/out/vanilla.sv:996.217-996.249" */ 7'h20;
  assign _1669_ = mem_rdata_q[14:12] == /* src = "generated/out/vanilla.sv:996.113-996.141" */ 3'h5;
  assign _1667_ = mem_rdata_q[14:12] == /* src = "generated/out/vanilla.sv:996.43-996.71" */ 3'h1;
  assign _1674_ = ! /* src = "generated/out/vanilla.sv:996.77-996.109" */ mem_rdata_q[31:25];
  assign _1685_ = reg_sh >= /* src = "generated/out/vanilla.sv:1584.35-1584.46" */ 32'd4;
  assign _1686_ = latched_store && /* src = "generated/out/vanilla.sv:1080.20-1080.51" */ latched_branch;
  assign _1688_ = resetn && /* src = "generated/out/vanilla.sv:1181.8-1181.31" */ cpuregs_write;
  assign _1689_ = _1688_ && /* src = "generated/out/vanilla.sv:1181.7-1181.46" */ latched_rd;
  assign launch_next_insn = _1628_ && /* src = "generated/out/vanilla.sv:1195.29-1195.78" */ decoder_trigger;
  assign _1690_ = resetn && /* src = "generated/out/vanilla.sv:1214.9-1214.29" */ pcpi_valid;
  assign _1691_ = _1690_ && /* src = "generated/out/vanilla.sv:1214.8-1214.48" */ _1807_;
  assign _1692_ = mem_do_rinst && /* src = "generated/out/vanilla.sv:1234.22-1234.46" */ mem_done;
  assign _1687_ = latched_store && /* src = "generated/out/vanilla.sv:1281.7-1281.39" */ _1806_;
  assign _1696_ = is_lb_lh_lw_lbu_lhu && /* src = "generated/out/vanilla.sv:1454.7-1454.41" */ _1809_;
  assign _1697_ = _1810_ && /* src = "generated/out/vanilla.sv:1648.11-1648.39" */ mem_done;
  assign _1698_ = resetn && /* src = "generated/out/vanilla.sv:1668.7-1668.67" */ _1834_;
  assign _1699_ = _1636_ && /* src = "generated/out/vanilla.sv:1669.8-1669.50" */ _2006_;
  assign _1700_ = _1637_ && /* src = "generated/out/vanilla.sv:1674.8-1674.48" */ pcpi_rs1[0];
  assign _1701_ = resetn && /* src = "generated/out/vanilla.sv:1680.8-1680.50" */ mem_do_rinst;
  assign _1702_ = _1701_ && /* src = "generated/out/vanilla.sv:1680.7-1680.98" */ reg_pc[0];
  assign _1703_ = resetn && /* src = "generated/out/vanilla.sv:1715.18-1715.54" */ _1836_;
  assign _0021_ = _1703_ && /* src = "generated/out/vanilla.sv:1715.17-1715.73" */ dbg_valid_insn;
  assign _1704_ = mem_valid && /* src = "generated/out/vanilla.sv:1774.13-1774.43" */ mem_ready;
  assign _1705_ = rvfi_valid && /* src = "generated/out/vanilla.sv:1792.8-1792.52" */ _1638_;
  assign _1706_ = _1705_ && /* src = "generated/out/vanilla.sv:1792.7-1792.85" */ _1639_;
  assign _1708_ = _1707_ && /* src = "generated/out/vanilla.sv:286.27-286.94" */ next_pc[1];
  assign mem_la_firstword = _1708_ && /* src = "generated/out/vanilla.sv:286.26-286.117" */ _1811_;
  assign _1709_ = mem_la_firstword && /* src = "generated/out/vanilla.sv:293.42-293.102" */ prefetched_high_word;
  assign mem_la_use_prefetched_high_word = _1709_ && /* src = "generated/out/vanilla.sv:293.41-293.134" */ _1812_;
  assign _1710_ = mem_la_use_prefetched_high_word && /* src = "generated/out/vanilla.sv:294.49-294.96" */ mem_do_rinst;
  assign _1711_ = mem_xfer && /* src = "generated/out/vanilla.sv:296.32-296.54" */ _2420_;
  assign _1712_ = _1711_ && /* src = "generated/out/vanilla.sv:296.31-296.107" */ _1838_;
  assign _1713_ = _2413_ && /* src = "generated/out/vanilla.sv:296.113-296.139" */ mem_do_rinst;
  assign _1714_ = resetn && /* src = "generated/out/vanilla.sv:296.19-296.141" */ _1839_;
  assign _1715_ = _1801_ && /* src = "generated/out/vanilla.sv:296.169-296.205" */ mem_xfer;
  assign mem_done = _1714_ && /* src = "generated/out/vanilla.sv:296.18-296.207" */ _1840_;
  assign _1716_ = resetn && /* src = "generated/out/vanilla.sv:297.25-297.45" */ _1814_;
  assign mem_la_write = _1716_ && /* src = "generated/out/vanilla.sv:297.24-297.62" */ mem_do_wdata;
  assign _1717_ = _1815_ && /* src = "generated/out/vanilla.sv:298.36-298.82" */ _1814_;
  assign _1718_ = _1717_ && /* src = "generated/out/vanilla.sv:298.35-298.138" */ _1841_;
  assign mem_la_firstword_xfer = mem_xfer && /* src = "generated/out/vanilla.sv:298.146-298.237" */ _2412_;
  assign _1719_ = mem_la_firstword_xfer && /* src = "generated/out/vanilla.sv:298.145-298.260" */ _1811_;
  assign _1720_ = _1719_ && /* src = "generated/out/vanilla.sv:298.144-298.288" */ _2414_;
  assign mem_la_read = resetn && /* src = "generated/out/vanilla.sv:298.23-298.290" */ _1842_;
  assign _1721_ = mem_valid && /* src = "generated/out/vanilla.sv:310.22-310.45" */ _1816_;
  assign _1722_ = mem_done && /* src = "generated/out/vanilla.sv:344.7-344.72" */ _1707_;
  assign _1723_ = _0270_ && /* src = "generated/out/vanilla.sv:423.12-423.73" */ _1653_;
  assign _1728_ = _1659_ && /* src = "generated/out/vanilla.sv:800.18-800.96" */ _1660_;
  assign _1730_ = _1817_ && /* src = "generated/out/vanilla.sv:871.13-871.61" */ _1818_;
  assign _1731_ = _0270_ && /* src = "generated/out/vanilla.sv:917.14-917.76" */ _2008_;
  assign _1732_ = _1731_ && /* src = "generated/out/vanilla.sv:917.13-917.110" */ _1653_;
  assign _1724_ = _0270_ && /* src = "generated/out/vanilla.sv:922.13-922.74" */ _2007_;
  assign _1725_ = mem_rdata_latched[12] && /* src = "generated/out/vanilla.sv:928.14-928.76" */ _2008_;
  assign _1726_ = _1725_ && /* src = "generated/out/vanilla.sv:928.13-928.110" */ _1653_;
  assign _1727_ = mem_rdata_latched[12] && /* src = "generated/out/vanilla.sv:933.13-933.74" */ _2007_;
  assign _1733_ = decoder_trigger && /* src = "generated/out/vanilla.sv:949.7-949.49" */ _1819_;
  assign _1734_ = is_beq_bne_blt_bge_bltu_bgeu && /* src = "generated/out/vanilla.sv:951.17-951.79" */ _1666_;
  assign _1735_ = is_beq_bne_blt_bge_bltu_bgeu && /* src = "generated/out/vanilla.sv:952.17-952.79" */ _1667_;
  assign _1736_ = is_beq_bne_blt_bge_bltu_bgeu && /* src = "generated/out/vanilla.sv:953.17-953.79" */ _1668_;
  assign _1737_ = is_beq_bne_blt_bge_bltu_bgeu && /* src = "generated/out/vanilla.sv:954.17-954.79" */ _1669_;
  assign _1738_ = is_beq_bne_blt_bge_bltu_bgeu && /* src = "generated/out/vanilla.sv:955.18-955.80" */ _1670_;
  assign _1739_ = is_beq_bne_blt_bge_bltu_bgeu && /* src = "generated/out/vanilla.sv:956.18-956.80" */ _1671_;
  assign _1740_ = is_lb_lh_lw_lbu_lhu && /* src = "generated/out/vanilla.sv:957.16-957.69" */ _1666_;
  assign _1741_ = is_lb_lh_lw_lbu_lhu && /* src = "generated/out/vanilla.sv:958.16-958.69" */ _1667_;
  assign _1742_ = is_lb_lh_lw_lbu_lhu && /* src = "generated/out/vanilla.sv:959.16-959.69" */ _1672_;
  assign _1743_ = is_lb_lh_lw_lbu_lhu && /* src = "generated/out/vanilla.sv:960.17-960.70" */ _1668_;
  assign _1744_ = is_lb_lh_lw_lbu_lhu && /* src = "generated/out/vanilla.sv:961.17-961.70" */ _1669_;
  assign _1745_ = is_sb_sh_sw && /* src = "generated/out/vanilla.sv:962.16-962.61" */ _1666_;
  assign _1746_ = is_sb_sh_sw && /* src = "generated/out/vanilla.sv:963.16-963.61" */ _1667_;
  assign _1747_ = is_sb_sh_sw && /* src = "generated/out/vanilla.sv:964.16-964.61" */ _1672_;
  assign _1748_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:965.18-965.66" */ _1666_;
  assign _1749_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:966.18-966.66" */ _1672_;
  assign _1750_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:967.19-967.67" */ _1673_;
  assign _1751_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:968.18-968.66" */ _1668_;
  assign _1752_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:969.17-969.65" */ _1670_;
  assign _1753_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:970.18-970.66" */ _1671_;
  assign _1754_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:971.19-971.67" */ _1667_;
  assign _1755_ = _1754_ && /* src = "generated/out/vanilla.sv:971.18-971.106" */ _1674_;
  assign _1757_ = _1756_ && /* src = "generated/out/vanilla.sv:972.18-972.106" */ _1674_;
  assign _1756_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:973.19-973.67" */ _1669_;
  assign _1758_ = _1756_ && /* src = "generated/out/vanilla.sv:973.18-973.106" */ _1675_;
  assign _1760_ = _1759_ && /* src = "generated/out/vanilla.sv:974.17-974.105" */ _1674_;
  assign _1759_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:975.18-975.66" */ _1666_;
  assign _1761_ = _1759_ && /* src = "generated/out/vanilla.sv:975.17-975.105" */ _1675_;
  assign _1762_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:976.18-976.66" */ _1667_;
  assign _1763_ = _1762_ && /* src = "generated/out/vanilla.sv:976.17-976.105" */ _1674_;
  assign _1764_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:977.18-977.66" */ _1672_;
  assign _1765_ = _1764_ && /* src = "generated/out/vanilla.sv:977.17-977.105" */ _1674_;
  assign _1766_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:978.19-978.67" */ _1673_;
  assign _1767_ = _1766_ && /* src = "generated/out/vanilla.sv:978.18-978.106" */ _1674_;
  assign _1768_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:979.18-979.66" */ _1668_;
  assign _1769_ = _1768_ && /* src = "generated/out/vanilla.sv:979.17-979.105" */ _1674_;
  assign _1771_ = _1770_ && /* src = "generated/out/vanilla.sv:980.17-980.105" */ _1674_;
  assign _1770_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:981.18-981.66" */ _1669_;
  assign _1772_ = _1770_ && /* src = "generated/out/vanilla.sv:981.17-981.105" */ _1675_;
  assign _1773_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:982.17-982.65" */ _1670_;
  assign _1774_ = _1773_ && /* src = "generated/out/vanilla.sv:982.16-982.104" */ _1674_;
  assign _1775_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:983.18-983.66" */ _1671_;
  assign _1776_ = _1775_ && /* src = "generated/out/vanilla.sv:983.17-983.105" */ _1674_;
  assign _1777_ = _1676_ && /* src = "generated/out/vanilla.sv:984.24-984.98" */ _1677_;
  assign _1778_ = _1777_ && /* src = "generated/out/vanilla.sv:984.23-984.130" */ _2009_;
  assign _1779_ = _1676_ && /* src = "generated/out/vanilla.sv:984.137-984.211" */ _1678_;
  assign _1780_ = _1779_ && /* src = "generated/out/vanilla.sv:984.136-984.243" */ _2009_;
  assign _1782_ = _1676_ && /* src = "generated/out/vanilla.sv:985.26-985.100" */ _1679_;
  assign _1783_ = _1782_ && /* src = "generated/out/vanilla.sv:985.25-985.132" */ _2009_;
  assign _1784_ = _1676_ && /* src = "generated/out/vanilla.sv:985.139-985.213" */ _1680_;
  assign _1785_ = _1784_ && /* src = "generated/out/vanilla.sv:985.138-985.245" */ _2009_;
  assign _1787_ = _1676_ && /* src = "generated/out/vanilla.sv:986.23-986.97" */ _1681_;
  assign _1788_ = _1787_ && /* src = "generated/out/vanilla.sv:986.22-986.129" */ _2009_;
  assign _1789_ = _1676_ && /* src = "generated/out/vanilla.sv:987.25-987.99" */ _1682_;
  assign _1790_ = _1789_ && /* src = "generated/out/vanilla.sv:987.24-987.131" */ _2009_;
  assign _1791_ = _1676_ && /* src = "generated/out/vanilla.sv:988.28-988.83" */ _1820_;
  assign _1792_ = _1791_ && /* src = "generated/out/vanilla.sv:988.27-988.106" */ _1821_;
  assign _1793_ = _1684_ && /* src = "generated/out/vanilla.sv:989.19-989.74" */ _1822_;
  assign _1797_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:994.25-994.254" */ _2423_;
  assign _1798_ = is_alu_reg_imm && /* src = "generated/out/vanilla.sv:995.60-995.259" */ _2424_;
  assign _1794_ = _1669_ && /* src = "generated/out/vanilla.sv:996.182-996.250" */ _1675_;
  assign _1795_ = _1669_ && /* src = "generated/out/vanilla.sv:996.112-996.180" */ _1674_;
  assign _1796_ = _1667_ && /* src = "generated/out/vanilla.sv:996.42-996.110" */ _1674_;
  assign _1799_ = is_alu_reg_reg && /* src = "generated/out/vanilla.sv:996.22-996.251" */ _2423_;
  assign _1800_ = ! /* src = "generated/out/vanilla.sv:0.0-0.0" */ _2415_;
  assign _1801_ = ! /* src = "generated/out/vanilla.sv:0.0-0.0" */ _2414_;
  assign _1803_ = ! /* src = "generated/out/vanilla.sv:1124.27-1124.34" */ alu_eq;
  assign _1804_ = ! /* src = "generated/out/vanilla.sv:1125.27-1125.35" */ alu_lts;
  assign _1805_ = ! /* src = "generated/out/vanilla.sv:1126.28-1126.36" */ alu_ltu;
  assign _1807_ = ! /* src = "generated/out/vanilla.sv:1214.34-1214.48" */ pcpi_int_wait;
  assign _1808_ = ! /* src = "generated/out/vanilla.sv:1220.20-1220.41" */ pcpi_timeout_counter;
  assign _1693_ = ! /* src = "generated/out/vanilla.sv:1275.22-1275.38" */ decoder_trigger;
  assign _1806_ = ! /* src = "generated/out/vanilla.sv:1281.24-1281.39" */ latched_branch;
  assign _1694_ = ! /* src = "generated/out/vanilla.sv:1346.27-1346.38" */ instr_jalr;
  assign _1809_ = ! /* src = "generated/out/vanilla.sv:1454.30-1454.41" */ instr_trap;
  assign _1810_ = ! /* src = "generated/out/vanilla.sv:1648.11-1648.27" */ mem_do_prefetch;
  assign _1802_ = ! /* src = "generated/out/vanilla.sv:1740.7-1740.14" */ resetn;
  assign _1812_ = ! /* src = "generated/out/vanilla.sv:293.107-293.134" */ clear_prefetched_high_word;
  assign _1813_ = ! /* src = "generated/out/vanilla.sv:296.147-296.164" */ mem_la_firstword;
  assign _1811_ = ! /* src = "generated/out/vanilla.sv:298.242-298.260" */ mem_la_secondword;
  assign _1816_ = ! /* src = "generated/out/vanilla.sv:310.35-310.45" */ mem_ready;
  assign _1815_ = ! /* src = "generated/out/vanilla.sv:499.12-499.44" */ mem_la_use_prefetched_high_word;
  assign instr_trap = ! /* src = "generated/out/vanilla.sv:608.54-608.626" */ { instr_lui, instr_auipc, instr_jal, instr_jalr, instr_beq, instr_bne, instr_blt, instr_bge, instr_bltu, instr_bgeu, instr_lb, instr_lh, instr_lw, instr_lbu, instr_lhu, instr_sb, instr_sh, instr_sw, instr_addi, instr_slti, instr_sltiu, instr_xori, instr_ori, instr_andi, instr_slli, instr_srli, instr_srai, instr_add, instr_sub, instr_sll, instr_slt, instr_sltu, instr_xor, instr_srl, instr_sra, instr_or, instr_and, instr_rdcycle, instr_rdcycleh, instr_rdinstr, instr_rdinstrh, instr_fence, 6'h00 };
  assign _1817_ = ! /* src = "generated/out/vanilla.sv:871.13-871.35" */ mem_rdata_latched[11];
  assign _1818_ = ! /* src = "generated/out/vanilla.sv:904.13-904.35" */ mem_rdata_latched[12];
  assign _1819_ = ! /* src = "generated/out/vanilla.sv:949.26-949.49" */ decoder_pseudo_trigger;
  assign _1820_ = ! /* src = "generated/out/vanilla.sv:988.64-988.83" */ mem_rdata_q[31:21];
  assign _1821_ = ! /* src = "generated/out/vanilla.sv:988.88-988.106" */ mem_rdata_q[19:7];
  assign _1822_ = ! /* src = "generated/out/vanilla.sv:989.55-989.74" */ mem_rdata_q[15:12];
  assign _1823_ = instr_sra || /* src = "generated/out/vanilla.sv:1115.25-1115.48" */ instr_srai;
  assign _1824_ = instr_xori || /* src = "generated/out/vanilla.sv:1135.4-1135.27" */ instr_xor;
  assign _1825_ = instr_ori || /* src = "generated/out/vanilla.sv:1136.4-1136.25" */ instr_or;
  assign _1826_ = instr_andi || /* src = "generated/out/vanilla.sv:1137.4-1137.27" */ instr_and;
  assign _1829_ = latched_branch || /* src = "generated/out/vanilla.sv:1148.8-1148.35" */ 2'h0;
  assign _1830_ = _1829_ || /* src = "generated/out/vanilla.sv:1148.7-1148.47" */ _1802_;
  assign _1695_ = pcpi_timeout || /* src = "generated/out/vanilla.sv:1527.35-1527.69" */ instr_ecall_ebreak;
  assign _1827_ = instr_slli || /* src = "generated/out/vanilla.sv:1596.8-1596.31" */ instr_sll;
  assign _1828_ = instr_srli || /* src = "generated/out/vanilla.sv:1597.8-1597.31" */ instr_srl;
  assign _1831_ = _1810_ || /* src = "generated/out/vanilla.sv:1630.10-1630.38" */ mem_done;
  assign _1832_ = instr_lb || /* src = "generated/out/vanilla.sv:1634.9-1634.30" */ instr_lbu;
  assign _1833_ = instr_lh || /* src = "generated/out/vanilla.sv:1635.9-1635.30" */ instr_lhu;
  assign _1834_ = mem_do_rdata || /* src = "generated/out/vanilla.sv:1668.38-1668.66" */ mem_do_wdata;
  assign _1835_ = _1802_ || /* src = "generated/out/vanilla.sv:1687.7-1687.26" */ mem_done;
  assign _1836_ = launch_next_insn || /* src = "generated/out/vanilla.sv:1715.29-1715.53" */ trap;
  assign mem_xfer = _1704_ || /* src = "generated/out/vanilla.sv:294.20-294.97" */ _1710_;
  assign _1838_ = _1837_ || /* src = "generated/out/vanilla.sv:296.60-296.106" */ mem_do_wdata;
  assign _1839_ = _1712_ || /* src = "generated/out/vanilla.sv:296.30-296.140" */ _1713_;
  assign _1840_ = _1813_ || /* src = "generated/out/vanilla.sv:296.147-296.206" */ _1715_;
  assign _1842_ = _1718_ || /* src = "generated/out/vanilla.sv:298.34-298.289" */ _1720_;
  assign _1844_ = _1802_ || /* src = "generated/out/vanilla.sv:464.8-464.28" */ mem_ready;
  assign _1845_ = mem_la_read || /* src = "generated/out/vanilla.sv:470.8-470.35" */ mem_la_write;
  assign _1841_ = _1707_ || /* src = "generated/out/vanilla.sv:478.10-478.59" */ mem_do_rdata;
  assign _1707_ = mem_do_prefetch || /* src = "generated/out/vanilla.sv:480.20-480.51" */ mem_do_rinst;
  assign _1846_ = _1800_ || /* src = "generated/out/vanilla.sv:506.13-506.50" */ mem_la_secondword;
  assign _1837_ = mem_do_rinst || /* src = "generated/out/vanilla.sv:512.22-512.50" */ mem_do_rdata;
  assign _1843_ = _1802_ || /* src = "generated/out/vanilla.sv:743.7-743.22" */ trap;
  assign _1847_ = mem_rdata_latched[12] || /* src = "generated/out/vanilla.sv:859.13-859.60" */ mem_rdata_latched[6:2];
  assign _1781_ = _1778_ || /* src = "generated/out/vanilla.sv:984.22-984.244" */ _1780_;
  assign _1786_ = _1783_ || /* src = "generated/out/vanilla.sv:985.24-985.246" */ _1785_;
  assign _1848_ = _1792_ || /* src = "generated/out/vanilla.sv:988.26-988.162" */ _1683_;
  assign _1849_ = instr_jalr || /* src = "generated/out/vanilla.sv:995.45-995.260" */ _1798_;
  assign alu_lts = $signed(pcpi_rs1) < /* src = "generated/out/vanilla.sv:1112.15-1112.50" */ $signed(pcpi_rs2);
  assign alu_ltu = pcpi_rs1 < /* src = "generated/out/vanilla.sv:1113.15-1113.32" */ pcpi_rs2;
  assign _2004_ = _0064_[4] ? _1852_ : _1850_;
  assign _1850_ = _0064_[3] ? _1856_ : _1854_;
  assign _1852_ = _0064_[3] ? _1860_ : _1858_;
  assign _1854_ = _0064_[2] ? _1864_ : _1862_;
  assign _1856_ = _0064_[2] ? _1868_ : _1866_;
  assign _1858_ = _0064_[2] ? _1872_ : _1870_;
  assign _1860_ = _0064_[2] ? _1876_ : _1874_;
  assign _1862_ = _0064_[1] ? _1880_ : _1878_;
  assign _1864_ = _0064_[1] ? _1884_ : _1882_;
  assign _1866_ = _0064_[1] ? _1888_ : _1886_;
  assign _1868_ = _0064_[1] ? _1892_ : _1890_;
  assign _1870_ = _0064_[1] ? _1896_ : _1894_;
  assign _1872_ = _0064_[1] ? _1900_ : _1898_;
  assign _1874_ = _0064_[1] ? _1904_ : _1902_;
  assign _1876_ = _0064_[1] ? _1908_ : _1906_;
  assign _1878_ = _0064_[0] ? \cpuregs[1]  : \cpuregs[0] ;
  assign _1898_ = _0064_[0] ? \cpuregs[21]  : \cpuregs[20] ;
  assign _1900_ = _0064_[0] ? \cpuregs[23]  : \cpuregs[22] ;
  assign _1902_ = _0064_[0] ? \cpuregs[25]  : \cpuregs[24] ;
  assign _1904_ = _0064_[0] ? \cpuregs[27]  : \cpuregs[26] ;
  assign _1906_ = _0064_[0] ? \cpuregs[29]  : \cpuregs[28] ;
  assign _1908_ = _0064_[0] ? \cpuregs[31]  : \cpuregs[30] ;
  assign _1880_ = _0064_[0] ? \cpuregs[3]  : \cpuregs[2] ;
  assign _1882_ = _0064_[0] ? \cpuregs[5]  : \cpuregs[4] ;
  assign _1884_ = _0064_[0] ? \cpuregs[7]  : \cpuregs[6] ;
  assign _1886_ = _0064_[0] ? \cpuregs[9]  : \cpuregs[8] ;
  assign _1888_ = _0064_[0] ? \cpuregs[11]  : \cpuregs[10] ;
  assign _1890_ = _0064_[0] ? \cpuregs[13]  : \cpuregs[12] ;
  assign _1892_ = _0064_[0] ? \cpuregs[15]  : \cpuregs[14] ;
  assign _1894_ = _0064_[0] ? \cpuregs[17]  : \cpuregs[16] ;
  assign _1896_ = _0064_[0] ? \cpuregs[19]  : \cpuregs[18] ;
  assign _2002_ = _0065_[4] ? _1912_ : _1910_;
  assign _1910_ = _0065_[3] ? _1916_ : _1914_;
  assign _1912_ = _0065_[3] ? _1920_ : _1918_;
  assign _1914_ = _0065_[2] ? _1924_ : _1922_;
  assign _1916_ = _0065_[2] ? _1928_ : _1926_;
  assign _1918_ = _0065_[2] ? _1932_ : _1930_;
  assign _1920_ = _0065_[2] ? _1936_ : _1934_;
  assign _1922_ = _0065_[1] ? _1940_ : _1938_;
  assign _1924_ = _0065_[1] ? _1944_ : _1942_;
  assign _1926_ = _0065_[1] ? _1948_ : _1946_;
  assign _1928_ = _0065_[1] ? _1952_ : _1950_;
  assign _1930_ = _0065_[1] ? _1956_ : _1954_;
  assign _1932_ = _0065_[1] ? _1960_ : _1958_;
  assign _1934_ = _0065_[1] ? _1964_ : _1962_;
  assign _1936_ = _0065_[1] ? _1968_ : _1966_;
  assign _1938_ = _0065_[0] ? \cpuregs[1]  : \cpuregs[0] ;
  assign _1958_ = _0065_[0] ? \cpuregs[21]  : \cpuregs[20] ;
  assign _1960_ = _0065_[0] ? \cpuregs[23]  : \cpuregs[22] ;
  assign _1962_ = _0065_[0] ? \cpuregs[25]  : \cpuregs[24] ;
  assign _1964_ = _0065_[0] ? \cpuregs[27]  : \cpuregs[26] ;
  assign _1966_ = _0065_[0] ? \cpuregs[29]  : \cpuregs[28] ;
  assign _1968_ = _0065_[0] ? \cpuregs[31]  : \cpuregs[30] ;
  assign _1940_ = _0065_[0] ? \cpuregs[3]  : \cpuregs[2] ;
  assign _1942_ = _0065_[0] ? \cpuregs[5]  : \cpuregs[4] ;
  assign _1944_ = _0065_[0] ? \cpuregs[7]  : \cpuregs[6] ;
  assign _1946_ = _0065_[0] ? \cpuregs[9]  : \cpuregs[8] ;
  assign _1948_ = _0065_[0] ? \cpuregs[11]  : \cpuregs[10] ;
  assign _1950_ = _0065_[0] ? \cpuregs[13]  : \cpuregs[12] ;
  assign _1952_ = _0065_[0] ? \cpuregs[15]  : \cpuregs[14] ;
  assign _1954_ = _0065_[0] ? \cpuregs[17]  : \cpuregs[16] ;
  assign _1956_ = _0065_[0] ? \cpuregs[19]  : \cpuregs[18] ;
  assign _1970_ = _0979_ & _0003_[31];
  assign _1971_ = _0995_ & _0003_[31];
  assign _1972_ = _0996_ & _0003_[31];
  assign _1973_ = _0998_ & _0003_[31];
  assign _1974_ = _0999_ & _0003_[31];
  assign _1975_ = _1000_ & _0003_[31];
  assign _1976_ = _1001_ & _0003_[31];
  assign _1977_ = _1004_ & _0003_[31];
  assign _1978_ = _1005_ & _0003_[31];
  assign _1979_ = _1006_ & _0003_[31];
  assign _1980_ = _1007_ & _0003_[31];
  assign _1981_ = _0981_ & _0003_[31];
  assign _1982_ = _1009_ & _0003_[31];
  assign _1983_ = _1010_ & _0003_[31];
  assign _1984_ = _1011_ & _0003_[31];
  assign _1985_ = _1012_ & _0003_[31];
  assign _1986_ = _1015_ & _0003_[31];
  assign _1987_ = _1016_ & _0003_[31];
  assign _1988_ = _1017_ & _0003_[31];
  assign _1989_ = _1018_ & _0003_[31];
  assign _1990_ = _1020_ & _0003_[31];
  assign _1991_ = _1021_ & _0003_[31];
  assign _1992_ = _0983_ & _0003_[31];
  assign _1993_ = _1022_ & _0003_[31];
  assign _1994_ = _1023_ & _0003_[31];
  assign _1995_ = _0985_ & _0003_[31];
  assign _1996_ = _0987_ & _0003_[31];
  assign _1997_ = _0988_ & _0003_[31];
  assign _1998_ = _0989_ & _0003_[31];
  assign _1999_ = _0990_ & _0003_[31];
  assign _2000_ = _0993_ & _0003_[31];
  assign _2001_ = _0994_ & _0003_[31];
  assign _2006_ = | /* src = "generated/out/vanilla.sv:1669.32-1669.49" */ pcpi_rs1[1:0];
  assign _1729_ = mem_rdata_latched[1:0] != /* src = "generated/out/vanilla.sv:817.27-817.58" */ 2'h3;
  assign _2008_ = | /* src = "generated/out/vanilla.sv:928.47-928.75" */ mem_rdata_latched[11:7];
  assign _2007_ = | /* src = "generated/out/vanilla.sv:933.46-933.73" */ mem_rdata_latched[6:2];
  assign _2009_ = | /* src = "generated/out/vanilla.sv:987.105-987.130" */ mem_rdata_q[13:12];
  assign _2010_ = pcpi_rs1 | /* src = "generated/out/vanilla.sv:1136.37-1136.54" */ pcpi_rs2;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_valid */
  always_ff @(posedge clk)
    rvfi_valid <= _0021_;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_halt */
  always_ff @(posedge clk)
    rvfi_halt <= trap;
  /* src = "generated/out/vanilla.sv:1714.2-1781.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME rvfi_pc_rdata */
  always_ff @(posedge clk)
    rvfi_pc_rdata <= rvfi_pc_wdata;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME reg_out */
  always_ff @(posedge clk)
    reg_out <= _0018_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME reg_sh */
  always_ff @(posedge clk)
    reg_sh <= _0020_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME decoder_trigger */
  always_ff @(posedge clk)
    decoder_trigger <= _0010_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME decoder_trigger_q */
  always_ff @(posedge clk)
    decoder_trigger_q <= decoder_trigger;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME decoder_pseudo_trigger_q */
  always_ff @(posedge clk)
    decoder_pseudo_trigger_q <= decoder_pseudo_trigger;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_rs1val */
  always_ff @(posedge clk)
    dbg_rs1val <= _0004_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_rs2val */
  always_ff @(posedge clk)
    dbg_rs2val <= _0007_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_rs1val_valid */
  always_ff @(posedge clk)
    dbg_rs1val_valid <= _0006_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_rs2val_valid */
  always_ff @(posedge clk)
    dbg_rs2val_valid <= _0009_;
  /* src = "generated/out/vanilla.sv:1196.2-1710.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME alu_out_q */
  always_ff @(posedge clk)
    alu_out_q <= alu_out;
  /* src = "generated/out/vanilla.sv:1143.2-1143.83" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME clear_prefetched_high_word_q */
  always_ff @(posedge clk)
    clear_prefetched_high_word_q <= clear_prefetched_high_word;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME is_lui_auipc_jal */
  always_ff @(posedge clk)
    is_lui_auipc_jal <= _0011_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME is_slti_blt_slt */
  always_ff @(posedge clk)
    is_slti_blt_slt <= _0012_;
  /* src = "generated/out/vanilla.sv:789.2-1036.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME is_sltiu_bltu_sltu */
  always_ff @(posedge clk)
    is_sltiu_bltu_sltu <= _0013_;
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME q_insn_rs1 */
  always_ff @(posedge clk)
    q_insn_rs1 <= dbg_insn_rs1;
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME q_insn_rs2 */
  always_ff @(posedge clk)
    q_insn_rs2 <= dbg_insn_rs2;
  /* src = "generated/out/vanilla.sv:735.2-760.5" */
/* PC_TAINT_INFO MODULE_NAME cellift_data_flow_picorv32  */
/* PC_TAINT_INFO STATE_NAME dbg_next */
  always_ff @(posedge clk)
    dbg_next <= launch_next_insn;
  assign _0039_ = _1640_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1793.8-1793.35|generated/out/vanilla.sv:1793.4-1796.7" */ 64'h00000000ffffffff : 64'h0000000000000000;
  assign rvfi_csr_minstret_rdata = _1706_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1792.7-1792.85|generated/out/vanilla.sv:1792.3-1809.6" */ _0055_ : 64'h0000000000000000;
  assign rvfi_csr_minstret_rmask = _1706_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1792.7-1792.85|generated/out/vanilla.sv:1792.3-1809.6" */ _0057_ : 64'h0000000000000000;
  assign rvfi_csr_mcycle_rdata = _1706_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1792.7-1792.85|generated/out/vanilla.sv:1792.3-1809.6" */ _0052_ : 64'h0000000000000000;
  assign rvfi_csr_mcycle_rmask = _1706_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1792.7-1792.85|generated/out/vanilla.sv:1792.3-1809.6" */ _0054_ : 64'h0000000000000000;
  assign _2012_ = { dbg_insn_opcode[31:25], dbg_insn_opcode[19:15], dbg_insn_opcode[11:0] } == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1752.3-1765.10" */ 24'h04000b;
  assign _2013_ = { dbg_insn_opcode[31:25], dbg_insn_opcode[19:17], dbg_insn_opcode[6:0] } == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1752.3-1765.10" */ 17'h0000b;
  assign _2014_ = _1704_ ? /* src = "generated/out/vanilla.sv:1774.13-1774.43|generated/out/vanilla.sv:1774.9-1780.7" */ mem_wdata : 32'hxxxxxxxx;
  assign _2016_ = _1704_ ? /* src = "generated/out/vanilla.sv:1774.13-1774.43|generated/out/vanilla.sv:1774.9-1780.7" */ mem_rdata : 32'hxxxxxxxx;
  assign _2018_ = _1704_ ? /* src = "generated/out/vanilla.sv:1774.13-1774.43|generated/out/vanilla.sv:1774.9-1780.7" */ mem_wstrb : 4'hx;
  assign _2020_ = _1704_ ? /* src = "generated/out/vanilla.sv:1774.13-1774.43|generated/out/vanilla.sv:1774.9-1780.7" */ _2440_[3:0] : 4'hx;
  assign _2021_ = _1704_ ? /* src = "generated/out/vanilla.sv:1774.13-1774.43|generated/out/vanilla.sv:1774.9-1780.7" */ mem_addr : 32'hxxxxxxxx;
  assign _2023_ = rvfi_valid ? /* src = "generated/out/vanilla.sv:1748.12-1748.22|generated/out/vanilla.sv:1748.8-1751.6" */ 32'd0 : 32'hxxxxxxxx;
  assign _2024_ = cpuregs_write ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1744.12-1744.39|generated/out/vanilla.sv:1744.8-1751.6" */ _2438_ : _2023_;
  assign _2027_ = rvfi_valid ? /* src = "generated/out/vanilla.sv:1748.12-1748.22|generated/out/vanilla.sv:1748.8-1751.6" */ 5'h00 : 5'hxx;
  assign _2028_ = cpuregs_write ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1744.12-1744.39|generated/out/vanilla.sv:1744.8-1751.6" */ latched_rd : _2027_;
  assign _2026_ = { dbg_insn_opcode[31:25], dbg_insn_opcode[11:9], dbg_insn_opcode[6:0] } == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1752.3-1765.10" */ 17'h0040b;
  assign _0058_ = _1831_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1630.10-1630.38|generated/out/vanilla.sv:1630.6-1659.9" */ _0061_ : 1'h0;
  assign _0060_ = _1831_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1606.10-1606.38|generated/out/vanilla.sv:1606.6-1626.9" */ _0062_ : 1'h0;
  assign _0059_ = is_beq_bne_blt_bge_bltu_bgeu ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1559.15-1559.43|generated/out/vanilla.sv:1559.11-1575.9" */ _0063_ : 1'h0;
  assign _0062_ = mem_do_wdata ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1607.11-1607.24|generated/out/vanilla.sv:1607.7-1620.10" */ 1'h0 : 1'h1;
  assign _0061_ = mem_do_rdata ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1631.11-1631.24|generated/out/vanilla.sv:1631.7-1647.10" */ 1'h0 : 1'h1;
  assign _0063_ = alu_out_0 ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1565.11-1565.56|generated/out/vanilla.sv:1565.7-1568.10" */ 1'h1 : 1'h0;
  assign _2030_ = latched_branch ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1279.6-1292.13" */ _2434_ : reg_next_pc;
  assign _2032_ = _1628_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ _2030_ : 32'hxxxxxxxx;
  assign _0046_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _2032_ : 32'hxxxxxxxx;
  assign _0024_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _0045_ : 1'h0;
  assign _0022_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _0043_ : 1'h0;
  assign _0023_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _0044_ : 1'h0;
  assign _2034_ = _1697_ ? /* src = "generated/out/vanilla.sv:1621.11-1621.39|generated/out/vanilla.sv:1621.7-1625.10" */ 1'h1 : 1'h0;
  assign _2035_ = _1697_ ? /* src = "generated/out/vanilla.sv:1621.11-1621.39|generated/out/vanilla.sv:1621.7-1625.10" */ 1'h1 : _1692_;
  assign _2036_ = _1831_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1606.10-1606.38|generated/out/vanilla.sv:1606.6-1626.9" */ _2035_ : _1692_;
  assign _2037_ = alu_out_0 ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1565.11-1565.56|generated/out/vanilla.sv:1565.7-1568.10" */ 1'h0 : _1692_;
  assign _2038_ = is_beq_bne_blt_bge_bltu_bgeu ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1559.15-1559.43|generated/out/vanilla.sv:1559.11-1575.9" */ _2037_ : _1692_;
  assign _0010_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _1316_ : _1692_;
  assign _2039_ = _1697_ ? /* src = "generated/out/vanilla.sv:1648.11-1648.39|generated/out/vanilla.sv:1648.7-1658.10" */ _1319_ : 32'hxxxxxxxx;
  assign _2041_ = _1831_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1630.10-1630.38|generated/out/vanilla.sv:1630.6-1659.9" */ _2039_ : 32'hxxxxxxxx;
  assign _2043_ = _1635_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1579.10-1579.21|generated/out/vanilla.sv:1579.6-1601.9" */ pcpi_rs1 : 32'hxxxxxxxx;
  assign _2047_ = instr_trap ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1517.6-1551.13" */ _2045_ : 32'hxxxxxxxx;
  assign _2045_ = pcpi_int_ready ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1367.14-1367.28|generated/out/vanilla.sv:1367.10-1382.13" */ pcpi_int_rd : 32'hxxxxxxxx;
  assign _0018_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _1327_ : 32'hxxxxxxxx;
  assign _2049_ = _1685_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1584.15-1584.47|generated/out/vanilla.sv:1584.11-1601.9" */ _2430_[4:0] : _2431_[4:0];
  assign _2050_ = _1635_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1579.10-1579.21|generated/out/vanilla.sv:1579.6-1601.9" */ 5'hxx : _2049_;
  assign _0020_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _1338_ : 5'hxx;
  assign _2051_ = _1627_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 1'h1 : 1'h0;
  assign _1627_ = cpu_state == /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 8'h80;
  assign _2053_ = is_beq_bne_blt_bge_bltu_bgeu ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1559.15-1559.43|generated/out/vanilla.sv:1559.11-1575.9" */ 5'h00 : 5'hxx;
  assign _2054_ = mem_do_rdata ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1631.11-1631.24|generated/out/vanilla.sv:1631.7-1647.10" */ 1'hx : instr_lb;
  assign _2055_ = _1831_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1630.10-1630.38|generated/out/vanilla.sv:1630.6-1659.9" */ _2054_ : 1'hx;
  assign _2056_ = mem_do_rdata ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1631.11-1631.24|generated/out/vanilla.sv:1631.7-1647.10" */ 1'hx : instr_lh;
  assign _2057_ = _1831_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1630.10-1630.38|generated/out/vanilla.sv:1630.6-1659.9" */ _2056_ : 1'hx;
  assign _2058_ = is_beq_bne_blt_bge_bltu_bgeu ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1559.15-1559.43|generated/out/vanilla.sv:1559.11-1575.9" */ alu_out_0 : instr_jalr;
  assign _2059_ = instr_jal ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1339.11-1339.20|generated/out/vanilla.sv:1339.7-1348.10" */ 1'h1 : 1'h0;
  assign _2060_ = decoder_trigger ? /* src = "generated/out/vanilla.sv:1329.15-1329.30|generated/out/vanilla.sv:1329.11-1349.9" */ _2059_ : 1'h0;
  assign _2061_ = is_beq_bne_blt_bge_bltu_bgeu ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1559.15-1559.43|generated/out/vanilla.sv:1559.11-1575.9" */ 1'hx : 1'h1;
  assign _2062_ = is_beq_bne_blt_bge_bltu_bgeu ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1559.15-1559.43|generated/out/vanilla.sv:1559.11-1575.9" */ alu_out_0 : 1'h1;
  assign _2064_ = instr_trap ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1517.6-1551.13" */ _2063_ : 1'hx;
  assign _2063_ = pcpi_int_ready ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1367.14-1367.28|generated/out/vanilla.sv:1367.10-1382.13" */ pcpi_int_wr : latched_store;
  assign _2065_ = _1697_ ? /* src = "generated/out/vanilla.sv:1621.11-1621.39|generated/out/vanilla.sv:1621.7-1625.10" */ 8'h40 : cpu_state;
  assign _2066_ = _1831_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1606.10-1606.38|generated/out/vanilla.sv:1606.6-1626.9" */ _2065_ : cpu_state;
  assign _2067_ = _1635_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1579.10-1579.21|generated/out/vanilla.sv:1579.6-1601.9" */ 8'h40 : cpu_state;
  assign _2068_ = mem_done ? /* src = "generated/out/vanilla.sv:1563.11-1563.19|generated/out/vanilla.sv:1563.7-1564.37" */ 8'h40 : cpu_state;
  assign _2069_ = is_beq_bne_blt_bge_bltu_bgeu ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1559.15-1559.43|generated/out/vanilla.sv:1559.11-1575.9" */ _2068_ : 8'h40;
  assign _2070_ = _1695_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1374.19-1374.72|generated/out/vanilla.sv:1374.15-1382.13" */ 8'h80 : cpu_state;
  assign _2071_ = pcpi_int_ready ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1367.14-1367.28|generated/out/vanilla.sv:1367.10-1382.13" */ 8'h40 : _2070_;
  assign _2072_ = instr_jal ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1339.11-1339.20|generated/out/vanilla.sv:1339.7-1348.10" */ cpu_state : 8'h20;
  assign _2073_ = decoder_trigger ? /* src = "generated/out/vanilla.sv:1329.15-1329.30|generated/out/vanilla.sv:1329.11-1349.9" */ _2072_ : cpu_state;
  assign _2074_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _1357_ : 8'h40;
  assign _2075_ = _1699_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1669.8-1669.50|generated/out/vanilla.sv:1669.4-1673.34" */ 8'h80 : _2074_;
  assign _2076_ = _1700_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1674.8-1674.48|generated/out/vanilla.sv:1674.4-1678.34" */ 8'h80 : _2075_;
  assign _2077_ = _1698_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1668.7-1668.67|generated/out/vanilla.sv:1668.3-1679.6" */ _2076_ : _2074_;
  assign _2078_ = launch_next_insn ? /* src = "generated/out/vanilla.sv:1207.7-1207.23|generated/out/vanilla.sv:1207.3-1212.6" */ 1'h0 : dbg_rs2val_valid;
  assign _2079_ = _0357_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1355.6-1509.13" */ _2078_ : 1'h1;
  assign _0009_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _1369_ : _2078_;
  assign _2080_ = launch_next_insn ? /* src = "generated/out/vanilla.sv:1207.7-1207.23|generated/out/vanilla.sv:1207.3-1212.6" */ 1'h0 : dbg_rs1val_valid;
  assign _2081_ = _0359_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1355.6-1509.13" */ _2080_ : 1'h1;
  assign _2082_ = _1629_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ _2081_ : _2080_;
  assign _0006_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _2082_ : _2080_;
  assign _2083_ = launch_next_insn ? /* src = "generated/out/vanilla.sv:1207.7-1207.23|generated/out/vanilla.sv:1207.3-1212.6" */ 32'hxxxxxxxx : dbg_rs2val;
  assign _2085_ = _0357_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1355.6-1509.13" */ _2083_ : cpuregs_rs2;
  assign _0007_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _1372_ : _2083_;
  assign _2087_ = launch_next_insn ? /* src = "generated/out/vanilla.sv:1207.7-1207.23|generated/out/vanilla.sv:1207.3-1212.6" */ 32'hxxxxxxxx : dbg_rs1val;
  assign _2089_ = _0359_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1355.6-1509.13" */ _2087_ : cpuregs_rs1;
  assign _2091_ = _1629_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ _2089_ : _2087_;
  assign _0004_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _2091_ : _2087_;
  assign _2093_ = _1635_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1579.10-1579.21|generated/out/vanilla.sv:1579.6-1601.9" */ mem_do_prefetch : 1'hx;
  assign _1631_ = cpu_state == /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 8'h08;
  assign _2094_ = pcpi_int_ready ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1367.14-1367.28|generated/out/vanilla.sv:1367.10-1382.13" */ 1'h1 : mem_do_rinst;
  assign _2095_ = decoder_trigger ? /* src = "generated/out/vanilla.sv:1329.15-1329.30|generated/out/vanilla.sv:1329.11-1349.9" */ _2059_ : _1693_;
  assign _2096_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1242.7-1242.14|generated/out/vanilla.sv:1242.3-1661.11" */ _1376_ : 1'hx;
  assign _2097_ = _1835_ ? /* src = "generated/out/vanilla.sv:1687.7-1687.26|generated/out/vanilla.sv:1687.3-1692.6" */ 1'h0 : _2096_;
  assign _2098_ = mem_do_rdata ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1631.11-1631.24|generated/out/vanilla.sv:1631.7-1647.10" */ 2'hx : _1387_;
  assign _2099_ = _1831_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1630.10-1630.38|generated/out/vanilla.sv:1630.6-1659.9" */ _2098_ : 2'hx;
  assign _2100_ = mem_do_wdata ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1607.11-1607.24|generated/out/vanilla.sv:1607.7-1620.10" */ 2'hx : _1391_;
  assign _2101_ = _1831_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1606.10-1606.38|generated/out/vanilla.sv:1606.6-1626.9" */ _2100_ : 2'hx;
  assign _2102_ = mem_do_rdata ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1631.11-1631.24|generated/out/vanilla.sv:1631.7-1647.10" */ 32'hxxxxxxxx : _0080_;
  assign _2104_ = _1831_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1630.10-1630.38|generated/out/vanilla.sv:1630.6-1659.9" */ _2102_ : 32'hxxxxxxxx;
  assign _1634_ = cpu_state == /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 8'h01;
  assign _2106_ = mem_do_wdata ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1607.11-1607.24|generated/out/vanilla.sv:1607.7-1620.10" */ 32'hxxxxxxxx : _0080_;
  assign _2108_ = _1831_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1606.10-1606.38|generated/out/vanilla.sv:1606.6-1626.9" */ _2106_ : 32'hxxxxxxxx;
  assign _1633_ = cpu_state == /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 8'h02;
  assign _2110_ = _1685_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1584.15-1584.47|generated/out/vanilla.sv:1584.11-1601.9" */ _1410_ : _1406_;
  assign _2112_ = _1635_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1579.10-1579.21|generated/out/vanilla.sv:1579.6-1601.9" */ 32'hxxxxxxxx : _2110_;
  assign _1632_ = cpu_state == /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 8'h04;
  assign _2114_ = instr_jal ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1339.11-1339.20|generated/out/vanilla.sv:1339.7-1348.10" */ _0076_ : _0072_;
  assign _2116_ = decoder_trigger ? /* src = "generated/out/vanilla.sv:1329.15-1329.30|generated/out/vanilla.sv:1329.11-1349.9" */ _2114_ : _0046_;
  assign _1628_ = cpu_state == /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 8'h40;
  assign _2121_ = _0358_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ _2120_ : 1'hx;
  assign _1630_ = cpu_state == /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 8'h10;
  assign _2118_ = _1695_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1374.19-1374.72|generated/out/vanilla.sv:1374.15-1382.13" */ 1'h0 : 1'h1;
  assign _2119_ = pcpi_int_ready ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1367.14-1367.28|generated/out/vanilla.sv:1367.10-1382.13" */ 1'h0 : _2118_;
  assign _2120_ = instr_trap ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1355.6-1509.13" */ _2119_ : 1'hx;
  assign _1629_ = cpu_state == /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1272.4-1661.11" */ 8'h20;
  assign _0003_[31] = _1689_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1181.7-1181.46|generated/out/vanilla.sv:1181.3-1182.42" */ 1'h1 : 1'h0;
  assign _0001_ = _1689_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1181.7-1181.46|generated/out/vanilla.sv:1181.3-1182.42" */ cpuregs_wrdata : 32'hxxxxxxxx;
  assign _0000_ = _1689_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1181.7-1181.46|generated/out/vanilla.sv:1181.3-1182.42" */ latched_rd : 5'hxx;
  assign _0028_ = _0451_ ? /* full_case = 32'd1 */ /* parallel_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1161.4-1178.11" */ 1'h1 : 1'h0;
  assign cpuregs_wrdata = _1628_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1159.7-1159.35|generated/out/vanilla.sv:1159.3-1178.11" */ _0026_ : 32'hxxxxxxxx;
  assign cpuregs_write = _1628_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1159.7-1159.35|generated/out/vanilla.sv:1159.3-1178.11" */ _0028_ : 1'h0;
  assign clear_prefetched_high_word = _1830_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1148.7-1148.47|generated/out/vanilla.sv:1148.3-1149.48" */ 1'h1 : _0025_;
  assign _0025_ = prefetched_high_word ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1146.7-1146.28|generated/out/vanilla.sv:1146.3-1147.35" */ clear_prefetched_high_word_q : 1'h0;
  assign _2122_ = _1732_ ? /* src = "generated/out/vanilla.sv:917.13-917.110|generated/out/vanilla.sv:917.9-921.12" */ mem_rdata_latched[11] : 1'h0;
  assign _2124_ = _1724_ ? /* src = "generated/out/vanilla.sv:922.13-922.74|generated/out/vanilla.sv:922.9-927.12" */ 1'h0 : _2122_;
  assign _2126_ = _1726_ ? /* src = "generated/out/vanilla.sv:928.13-928.110|generated/out/vanilla.sv:928.9-932.12" */ mem_rdata_latched[11] : _2124_;
  assign _2128_ = _1727_ ? /* src = "generated/out/vanilla.sv:933.13-933.74|generated/out/vanilla.sv:933.9-938.12" */ mem_rdata_latched[11] : _2126_;
  assign _2131_ = mem_rdata_latched[12] ? /* src = "generated/out/vanilla.sv:904.13-904.35|generated/out/vanilla.sv:904.9-909.12" */ 1'h0 : mem_rdata_latched[11];
  assign _2137_ = _1730_ ? /* src = "generated/out/vanilla.sv:871.13-871.61|generated/out/vanilla.sv:871.9-876.12" */ _0088_[4] : 1'h0;
  assign _2139_ = _1647_ ? /* src = "generated/out/vanilla.sv:877.13-877.46|generated/out/vanilla.sv:877.9-881.12" */ _0088_[4] : _2137_;
  assign _2141_ = _1648_ ? /* src = "generated/out/vanilla.sv:882.13-882.47|generated/out/vanilla.sv:882.9-887.12" */ _0088_[4] : _2139_;
  assign _2143_ = _1644_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:860.14-860.42|generated/out/vanilla.sv:860.10-869.13" */ mem_rdata_latched[11] : 1'h0;
  assign _2145_ = _1847_ ? /* src = "generated/out/vanilla.sv:859.13-859.60|generated/out/vanilla.sv:859.9-869.13" */ _2143_ : 1'h0;
  assign _2149_ = _0441_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ _0088_[4] : 1'h0;
  assign _2153_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _1434_ : mem_rdata_latched[19];
  assign _2155_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ mem_rdata_latched[8] : mem_rdata_latched[30];
  assign _2157_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ mem_rdata_latched[6] : mem_rdata_latched[27];
  assign _2159_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ mem_rdata_latched[7] : mem_rdata_latched[26];
  assign _2161_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ mem_rdata_latched[5:3] : mem_rdata_latched[23:21];
  assign _2163_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ mem_rdata_latched[2] : mem_rdata_latched[25];
  assign _2165_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ mem_rdata_latched[10:9] : mem_rdata_latched[29:28];
  assign _2167_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] } : { mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31], mem_rdata_latched[31] };
  assign _2169_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ mem_rdata_latched[11] : mem_rdata_latched[24];
  assign _2171_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ mem_rdata_latched[12] : mem_rdata_latched[20];
  assign _2173_ = _1732_ ? /* src = "generated/out/vanilla.sv:917.13-917.110|generated/out/vanilla.sv:917.9-921.12" */ mem_rdata_latched[10:7] : 4'h0;
  assign _2175_ = _1724_ ? /* src = "generated/out/vanilla.sv:922.13-922.74|generated/out/vanilla.sv:922.9-927.12" */ 4'h0 : _2173_;
  assign _2177_ = _1726_ ? /* src = "generated/out/vanilla.sv:928.13-928.110|generated/out/vanilla.sv:928.9-932.12" */ mem_rdata_latched[10:7] : _2175_;
  assign _2179_ = _1727_ ? /* src = "generated/out/vanilla.sv:933.13-933.74|generated/out/vanilla.sv:933.9-938.12" */ mem_rdata_latched[10:7] : _2177_;
  assign _2181_ = _2008_ ? /* src = "generated/out/vanilla.sv:911.13-911.36|generated/out/vanilla.sv:911.9-915.12" */ 4'h2 : 4'h0;
  assign _2182_ = mem_rdata_latched[12] ? /* src = "generated/out/vanilla.sv:904.13-904.35|generated/out/vanilla.sv:904.9-909.12" */ 4'h0 : mem_rdata_latched[10:7];
  assign _2184_ = _1730_ ? /* src = "generated/out/vanilla.sv:871.13-871.61|generated/out/vanilla.sv:871.9-876.12" */ _0088_[3:0] : 4'h0;
  assign _2186_ = _1647_ ? /* src = "generated/out/vanilla.sv:877.13-877.46|generated/out/vanilla.sv:877.9-881.12" */ _0088_[3:0] : _2184_;
  assign _2188_ = _1648_ ? /* src = "generated/out/vanilla.sv:882.13-882.47|generated/out/vanilla.sv:882.9-887.12" */ _0088_[3:0] : _2186_;
  assign _2190_ = _1644_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:860.14-860.42|generated/out/vanilla.sv:860.10-869.13" */ mem_rdata_latched[10:7] : 4'h0;
  assign _2192_ = _1847_ ? /* src = "generated/out/vanilla.sv:859.13-859.60|generated/out/vanilla.sv:859.9-869.13" */ _2190_ : 4'h0;
  assign _2194_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _1456_ : mem_rdata_latched[18:15];
  assign _2196_ = _1724_ ? /* src = "generated/out/vanilla.sv:922.13-922.74|generated/out/vanilla.sv:922.9-927.12" */ 1'h1 : _1665_;
  assign _2197_ = _1727_ ? /* src = "generated/out/vanilla.sv:933.13-933.74|generated/out/vanilla.sv:933.9-938.12" */ 1'h1 : _2196_;
  assign _2198_ = _2130_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:902.7-945.14" */ _2197_ : _1665_;
  assign _2199_ = _1648_ ? /* src = "generated/out/vanilla.sv:882.13-882.47|generated/out/vanilla.sv:882.9-887.12" */ 1'h1 : _1665_;
  assign _2200_ = _2130_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:843.7-900.14" */ _2199_ : _1665_;
  assign _2201_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _1470_ : _1665_;
  assign _2202_ = mem_rdata_latched[12] ? /* src = "generated/out/vanilla.sv:904.13-904.35|generated/out/vanilla.sv:904.9-909.12" */ _1664_ : 1'h1;
  assign _2203_ = _2133_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:902.7-945.14" */ _2202_ : _1664_;
  assign _2204_ = _1730_ ? /* src = "generated/out/vanilla.sv:871.13-871.61|generated/out/vanilla.sv:871.9-876.12" */ 1'h1 : _1664_;
  assign _2205_ = _1647_ ? /* src = "generated/out/vanilla.sv:877.13-877.46|generated/out/vanilla.sv:877.9-881.12" */ 1'h1 : _2204_;
  assign _2206_ = _1644_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:860.14-860.42|generated/out/vanilla.sv:860.10-869.13" */ 1'h1 : _1664_;
  assign _2207_ = _1847_ ? /* src = "generated/out/vanilla.sv:859.13-859.60|generated/out/vanilla.sv:859.9-869.13" */ _2206_ : _1664_;
  assign _2208_ = _2133_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ _2422_ : _1664_;
  assign _2209_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _1473_ : _1664_;
  assign _2210_ = _0442_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:843.7-900.14" */ 1'h1 : _1661_;
  assign _2211_ = _2148_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:823.5-946.12" */ _2210_ : _1661_;
  assign _2212_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _2211_ : _1661_;
  assign _2214_ = _0361_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:823.5-946.12" */ _2213_ : _1663_;
  assign _2213_ = _2136_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ 1'h1 : _1663_;
  assign _2215_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _2214_ : _1663_;
  assign _2216_ = _2008_ ? /* src = "generated/out/vanilla.sv:911.13-911.36|generated/out/vanilla.sv:911.9-915.12" */ 1'h1 : _1662_;
  assign _2217_ = _2151_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:902.7-945.14" */ _2216_ : _1662_;
  assign _2218_ = _2151_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ 1'h1 : _1662_;
  assign _2219_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _1478_ : _1662_;
  assign _2220_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ 1'h1 : 1'h0;
  assign _2222_ = _1724_ ? /* src = "generated/out/vanilla.sv:922.13-922.74|generated/out/vanilla.sv:922.9-927.12" */ mem_rdata_latched[6:2] : 5'h00;
  assign _2224_ = _1727_ ? /* src = "generated/out/vanilla.sv:933.13-933.74|generated/out/vanilla.sv:933.9-938.12" */ mem_rdata_latched[6:2] : _2222_;
  assign _2226_ = mem_rdata_latched[12] ? /* src = "generated/out/vanilla.sv:904.13-904.35|generated/out/vanilla.sv:904.9-909.12" */ 5'h00 : mem_rdata_latched[6:2];
  assign _2228_ = _1730_ ? /* src = "generated/out/vanilla.sv:871.13-871.61|generated/out/vanilla.sv:871.9-876.12" */ mem_rdata_latched[6:2] : 5'h00;
  assign _2230_ = _1648_ ? /* src = "generated/out/vanilla.sv:882.13-882.47|generated/out/vanilla.sv:882.9-887.12" */ _0086_[4:0] : _2228_;
  assign _2232_ = _2130_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:843.7-900.14" */ _2230_ : 5'h00;
  assign _2234_ = _2136_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ _0086_[4:0] : 5'h00;
  assign _2136_ = mem_rdata_latched[15:13] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ 3'h6;
  assign _2236_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _1499_ : mem_rdata_latched[24:20];
  assign _2238_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] } : mem_rdata_latched[19:12];
  assign _2240_ = _1724_ ? /* src = "generated/out/vanilla.sv:922.13-922.74|generated/out/vanilla.sv:922.9-927.12" */ mem_rdata_latched[11:7] : 5'h00;
  assign _2242_ = _1726_ ? /* src = "generated/out/vanilla.sv:928.13-928.110|generated/out/vanilla.sv:928.9-932.12" */ 5'h01 : _2240_;
  assign _2244_ = _1727_ ? /* src = "generated/out/vanilla.sv:933.13-933.74|generated/out/vanilla.sv:933.9-938.12" */ mem_rdata_latched[11:7] : _2242_;
  assign _2246_ = _2008_ ? /* src = "generated/out/vanilla.sv:911.13-911.36|generated/out/vanilla.sv:911.9-915.12" */ mem_rdata_latched[11:7] : 5'h00;
  assign _2248_ = mem_rdata_latched[12] ? /* src = "generated/out/vanilla.sv:904.13-904.35|generated/out/vanilla.sv:904.9-909.12" */ 5'h00 : mem_rdata_latched[11:7];
  assign _2250_ = _1730_ ? /* src = "generated/out/vanilla.sv:871.13-871.61|generated/out/vanilla.sv:871.9-876.12" */ _0088_[4:0] : 5'h00;
  assign _2252_ = _1647_ ? /* src = "generated/out/vanilla.sv:877.13-877.46|generated/out/vanilla.sv:877.9-881.12" */ _0088_[4:0] : _2250_;
  assign _2254_ = _1648_ ? /* src = "generated/out/vanilla.sv:882.13-882.47|generated/out/vanilla.sv:882.9-887.12" */ _0088_[4:0] : _2252_;
  assign _2256_ = _1847_ ? /* src = "generated/out/vanilla.sv:859.13-859.60|generated/out/vanilla.sv:859.9-869.13" */ mem_rdata_latched[11:7] : 5'h00;
  assign _2259_ = _0362_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ _0086_[4:0] : 5'h00;
  assign _2151_ = mem_rdata_latched[15:13] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ 3'h2;
  assign _2133_ = ! /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:825.7-841.14" */ mem_rdata_latched[15:13];
  assign _2152_ = ! /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:823.5-946.12" */ mem_rdata_latched[1:0];
  assign _2261_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _1511_ : mem_rdata_latched[11:7];
  assign _2263_ = _1732_ ? /* src = "generated/out/vanilla.sv:917.13-917.110|generated/out/vanilla.sv:917.9-921.12" */ 1'h1 : _1728_;
  assign _2264_ = _1726_ ? /* src = "generated/out/vanilla.sv:928.13-928.110|generated/out/vanilla.sv:928.9-932.12" */ 1'h1 : _2263_;
  assign _2265_ = _2130_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:902.7-945.14" */ _2264_ : _1728_;
  assign _2130_ = mem_rdata_latched[15:13] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:902.7-945.14" */ 3'h4;
  assign _2266_ = _2134_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:823.5-946.12" */ _2265_ : _1728_;
  assign _2134_ = mem_rdata_latched[1:0] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:823.5-946.12" */ 2'h2;
  assign _2267_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _2266_ : _1728_;
  assign _2268_ = _0448_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:843.7-900.14" */ 1'h1 : _1658_;
  assign _2269_ = mem_rdata_latched[15:13] == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:843.7-900.14" */ 3'h5;
  assign _2258_ = mem_rdata_latched[15:13] == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:843.7-900.14" */ 3'h1;
  assign _2270_ = _2148_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:823.5-946.12" */ _2268_ : _1658_;
  assign _2271_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _2270_ : _1658_;
  assign _2272_ = _1644_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:860.14-860.42|generated/out/vanilla.sv:860.10-869.13" */ _1656_ : 1'h1;
  assign _2273_ = _1847_ ? /* src = "generated/out/vanilla.sv:859.13-859.60|generated/out/vanilla.sv:859.9-869.13" */ _2272_ : _1656_;
  assign _2274_ = _2147_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:843.7-900.14" */ _2273_ : _1656_;
  assign _2147_ = mem_rdata_latched[15:13] == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:843.7-900.14" */ 3'h3;
  assign _2275_ = _2148_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:823.5-946.12" */ _2274_ : _1656_;
  assign _2148_ = mem_rdata_latched[1:0] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:823.5-946.12" */ 2'h1;
  assign _2276_ = _1729_ ? /* src = "generated/out/vanilla.sv:817.8-817.59|generated/out/vanilla.sv:817.4-947.7" */ _2275_ : _1656_;
  assign _0033_ = decoder_pseudo_trigger_q ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:769.8-769.32|generated/out/vanilla.sv:769.4-787.7" */ cached_insn_rs2 : decoded_rs2;
  assign _0031_ = decoder_pseudo_trigger_q ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:769.8-769.32|generated/out/vanilla.sv:769.4-787.7" */ cached_insn_rs1 : decoded_rs1;
  assign _0029_ = decoder_pseudo_trigger_q ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:769.8-769.32|generated/out/vanilla.sv:769.4-787.7" */ cached_insn_opcode : _0048_;
  assign dbg_insn_rs2 = dbg_next ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:768.7-768.15|generated/out/vanilla.sv:768.3-787.7" */ _0033_ : q_insn_rs2;
  assign dbg_insn_rs1 = dbg_next ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:768.7-768.15|generated/out/vanilla.sv:768.3-787.7" */ _0031_ : q_insn_rs1;
  assign dbg_insn_opcode = dbg_next ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:768.7-768.15|generated/out/vanilla.sv:768.3-787.7" */ _0029_ : { rvfi_insn[31:25], 5'hxx, rvfi_insn[19:15], 3'hx, rvfi_insn[11:0] };
  assign _0048_ = _2277_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:750.8-750.30|generated/out/vanilla.sv:750.4-753.74" */ next_insn_opcode : { 16'h0000, next_insn_opcode[15:0] };
  assign _2278_ = _1846_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:506.13-506.50|generated/out/vanilla.sv:506.9-511.36" */ mem_rdata[31:16] : 16'hxxxx;
  assign _2280_ = mem_do_rdata ? /* src = "generated/out/vanilla.sv:505.12-505.43|generated/out/vanilla.sv:505.8-511.36" */ 16'hxxxx : _2278_;
  assign _2282_ = mem_la_use_prefetched_high_word ? /* src = "generated/out/vanilla.sv:499.12-499.44|generated/out/vanilla.sv:499.8-500.46" */ 16'hxxxx : mem_rdata[31:16];
  assign _2284_ = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:496.11-496.40|generated/out/vanilla.sv:496.7-513.10" */ _2282_ : _2280_;
  assign _2286_ = mem_state == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:476.4-529.11" */ 2'h1;
  assign _2287_ = _1846_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:506.13-506.50|generated/out/vanilla.sv:506.9-511.36" */ 1'h1 : 1'h0;
  assign _2288_ = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:496.11-496.40|generated/out/vanilla.sv:496.7-513.10" */ 1'h1 : 1'h0;
  assign _2289_ = mem_do_rinst ? /* src = "generated/out/vanilla.sv:526.10-526.22|generated/out/vanilla.sv:526.6-527.22" */ 2'h0 : 2'hx;
  assign _1655_ = mem_state == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:476.4-529.11" */ 2'h3;
  assign _2290_ = mem_xfer ? /* src = "generated/out/vanilla.sv:518.10-518.18|generated/out/vanilla.sv:518.6-521.9" */ 2'h0 : 2'hx;
  assign _1654_ = mem_state == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:476.4-529.11" */ 2'h2;
  assign _2291_ = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:496.11-496.40|generated/out/vanilla.sv:496.7-513.10" */ 2'hx : _2447_[1:0];
  assign _2292_ = mem_xfer ? /* src = "generated/out/vanilla.sv:495.10-495.18|generated/out/vanilla.sv:495.6-513.10" */ _2291_ : 2'hx;
  assign _2293_ = _1841_ ? /* src = "generated/out/vanilla.sv:478.10-478.59|generated/out/vanilla.sv:478.6-483.9" */ 2'h1 : 2'hx;
  assign _2294_ = mem_do_wdata ? /* src = "generated/out/vanilla.sv:484.10-484.22|generated/out/vanilla.sv:484.6-488.9" */ 2'h2 : _2293_;
  assign _2295_ = resetn ? /* src = "generated/out/vanilla.sv:462.8-462.15|generated/out/vanilla.sv:462.4-463.20" */ 2'hx : 2'h0;
  assign _0016_ = _1843_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:461.7-461.22|generated/out/vanilla.sv:461.3-530.6" */ _2295_ : _1522_;
  assign _2296_ = _1845_ ? /* src = "generated/out/vanilla.sv:470.8-470.35|generated/out/vanilla.sv:470.4-473.7" */ _0094_ : mem_wstrb;
  assign _2298_ = _1841_ ? /* src = "generated/out/vanilla.sv:478.10-478.59|generated/out/vanilla.sv:478.6-483.9" */ 4'h0 : _2296_;
  assign _2300_ = _1814_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:476.4-529.11" */ _2298_ : _2296_;
  assign _1814_ = ! /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:476.4-529.11" */ mem_state;
  assign _2302_ = _1841_ ? /* src = "generated/out/vanilla.sv:478.10-478.59|generated/out/vanilla.sv:478.6-483.9" */ _1707_ : 1'hx;
  assign _2303_ = mem_xfer ? /* src = "generated/out/vanilla.sv:518.10-518.18|generated/out/vanilla.sv:518.6-521.9" */ 1'h0 : 1'hx;
  assign _2304_ = mem_xfer ? /* src = "generated/out/vanilla.sv:495.10-495.18|generated/out/vanilla.sv:495.6-513.10" */ _2288_ : 1'hx;
  assign _2305_ = _1841_ ? /* src = "generated/out/vanilla.sv:478.10-478.59|generated/out/vanilla.sv:478.6-483.9" */ _1815_ : 1'hx;
  assign _2306_ = mem_do_wdata ? /* src = "generated/out/vanilla.sv:484.10-484.22|generated/out/vanilla.sv:484.6-488.9" */ 1'h1 : _2305_;
  assign _2307_ = _1844_ ? /* src = "generated/out/vanilla.sv:464.8-464.28|generated/out/vanilla.sv:464.4-465.20" */ 1'h0 : 1'hx;
  assign _0017_ = _1843_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:461.7-461.22|generated/out/vanilla.sv:461.3-530.6" */ _2307_ : _1524_;
  assign _2308_ = mem_xfer ? /* src = "generated/out/vanilla.sv:340.7-340.15|generated/out/vanilla.sv:340.3-343.6" */ mem_rdata_latched[31] : mem_rdata_q[31];
  assign _2310_ = _1723_ ? /* src = "generated/out/vanilla.sv:423.12-423.73|generated/out/vanilla.sv:423.8-426.11" */ 1'h0 : _2308_;
  assign _2312_ = _1724_ ? /* src = "generated/out/vanilla.sv:427.12-427.73|generated/out/vanilla.sv:427.8-430.11" */ 1'h0 : _2310_;
  assign _2314_ = _1726_ ? /* src = "generated/out/vanilla.sv:431.12-431.109|generated/out/vanilla.sv:431.8-434.11" */ 1'h0 : _2312_;
  assign _2316_ = _1727_ ? /* src = "generated/out/vanilla.sv:435.12-435.73|generated/out/vanilla.sv:435.8-438.11" */ 1'h0 : _2314_;
  assign _2318_ = _1645_ ? /* src = "generated/out/vanilla.sv:379.12-379.45|generated/out/vanilla.sv:379.8-382.11" */ 1'h0 : _2308_;
  assign _2320_ = _1646_ ? /* src = "generated/out/vanilla.sv:383.12-383.45|generated/out/vanilla.sv:383.8-386.11" */ 1'h0 : _2318_;
  assign _2322_ = _1647_ ? /* src = "generated/out/vanilla.sv:387.12-387.45|generated/out/vanilla.sv:387.8-390.11" */ mem_rdata_latched[12] : _2320_;
  assign _2324_ = _1648_ ? /* src = "generated/out/vanilla.sv:391.12-391.46|generated/out/vanilla.sv:391.8-401.11" */ _2446_[6] : _2322_;
  assign _2326_ = _0360_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:347.6-360.13" */ 1'h0 : _2308_;
  assign _0014_[31] = _1722_ ? /* src = "generated/out/vanilla.sv:344.7-344.72|generated/out/vanilla.sv:344.3-445.11" */ _1533_ : _2308_;
  assign _2328_ = mem_xfer ? /* src = "generated/out/vanilla.sv:340.7-340.15|generated/out/vanilla.sv:340.3-343.6" */ mem_rdata_latched[7] : mem_rdata_q[7];
  assign _2330_ = _2136_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:413.6-444.13" */ 1'h0 : _2328_;
  assign _2332_ = _0442_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:362.6-411.13" */ mem_rdata_latched[12] : _2328_;
  assign _2135_ = mem_rdata_latched[15:13] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:362.6-411.13" */ 3'h7;
  assign _0014_[7] = _1722_ ? /* src = "generated/out/vanilla.sv:344.7-344.72|generated/out/vanilla.sv:344.3-445.11" */ _1541_ : _2328_;
  assign _2334_ = mem_xfer ? /* src = "generated/out/vanilla.sv:340.7-340.15|generated/out/vanilla.sv:340.3-343.6" */ mem_rdata_latched[24:20] : mem_rdata_q[24:20];
  assign _2336_ = _1723_ ? /* src = "generated/out/vanilla.sv:423.12-423.73|generated/out/vanilla.sv:423.8-426.11" */ 5'h00 : _2334_;
  assign _2338_ = _1726_ ? /* src = "generated/out/vanilla.sv:431.12-431.109|generated/out/vanilla.sv:431.8-434.11" */ 5'h00 : _2336_;
  assign _2340_ = _1647_ ? /* src = "generated/out/vanilla.sv:387.12-387.45|generated/out/vanilla.sv:387.8-390.11" */ mem_rdata_latched[6:2] : _2334_;
  assign _2342_ = _1644_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:372.12-372.40|generated/out/vanilla.sv:372.8-377.88" */ { mem_rdata_latched[6], 4'h0 } : { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] };
  assign _0014_[24:20] = _1722_ ? /* src = "generated/out/vanilla.sv:344.7-344.72|generated/out/vanilla.sv:344.3-445.11" */ _1551_ : _2334_;
  assign _2344_ = mem_xfer ? /* src = "generated/out/vanilla.sv:340.7-340.15|generated/out/vanilla.sv:340.3-343.6" */ mem_rdata_latched[19:15] : mem_rdata_q[19:15];
  assign _2346_ = _1644_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:372.12-372.40|generated/out/vanilla.sv:372.8-377.88" */ _2344_ : { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[6:5] };
  assign _2348_ = _2147_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:362.6-411.13" */ _2346_ : _2344_;
  assign _2350_ = _2148_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:345.4-445.11" */ _2348_ : _2344_;
  assign _0014_[19:15] = _1722_ ? /* src = "generated/out/vanilla.sv:344.7-344.72|generated/out/vanilla.sv:344.3-445.11" */ _2350_ : _2344_;
  assign _2352_ = mem_xfer ? /* src = "generated/out/vanilla.sv:340.7-340.15|generated/out/vanilla.sv:340.3-343.6" */ mem_rdata_latched[14:12] : mem_rdata_q[14:12];
  assign _2354_ = _1723_ ? /* src = "generated/out/vanilla.sv:423.12-423.73|generated/out/vanilla.sv:423.8-426.11" */ 3'h0 : _2352_;
  assign _2356_ = _1724_ ? /* src = "generated/out/vanilla.sv:427.12-427.73|generated/out/vanilla.sv:427.8-430.11" */ 3'h0 : _2354_;
  assign _2358_ = _1726_ ? /* src = "generated/out/vanilla.sv:431.12-431.109|generated/out/vanilla.sv:431.8-434.11" */ 3'h0 : _2356_;
  assign _2360_ = _1727_ ? /* src = "generated/out/vanilla.sv:435.12-435.73|generated/out/vanilla.sv:435.8-438.11" */ 3'h0 : _2358_;
  assign _2362_ = _1645_ ? /* src = "generated/out/vanilla.sv:379.12-379.45|generated/out/vanilla.sv:379.8-382.11" */ 3'h5 : _2352_;
  assign _2364_ = _1646_ ? /* src = "generated/out/vanilla.sv:383.12-383.45|generated/out/vanilla.sv:383.8-386.11" */ 3'h5 : _2362_;
  assign _2366_ = _1647_ ? /* src = "generated/out/vanilla.sv:387.12-387.45|generated/out/vanilla.sv:387.8-390.11" */ 3'h7 : _2364_;
  assign _2368_ = _1649_ ? /* src = "generated/out/vanilla.sv:392.13-392.44|generated/out/vanilla.sv:392.9-393.39" */ 3'h0 : _2366_;
  assign _2370_ = _1650_ ? /* src = "generated/out/vanilla.sv:394.13-394.44|generated/out/vanilla.sv:394.9-395.39" */ 3'h4 : _2368_;
  assign _2372_ = _1651_ ? /* src = "generated/out/vanilla.sv:396.13-396.44|generated/out/vanilla.sv:396.9-397.39" */ 3'h6 : _2370_;
  assign _2374_ = _1652_ ? /* src = "generated/out/vanilla.sv:398.13-398.44|generated/out/vanilla.sv:398.9-399.39" */ 3'h7 : _2372_;
  assign _2376_ = _1648_ ? /* src = "generated/out/vanilla.sv:391.12-391.46|generated/out/vanilla.sv:391.8-401.11" */ _2374_ : _2366_;
  assign _2378_ = _1644_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:372.12-372.40|generated/out/vanilla.sv:372.8-377.88" */ 3'h0 : mem_rdata_latched[4:2];
  assign _0014_[14:12] = _1722_ ? /* src = "generated/out/vanilla.sv:344.7-344.72|generated/out/vanilla.sv:344.3-445.11" */ _1573_ : _2352_;
  assign _2380_ = mem_xfer ? /* src = "generated/out/vanilla.sv:340.7-340.15|generated/out/vanilla.sv:340.3-343.6" */ mem_rdata_latched[11:8] : mem_rdata_q[11:8];
  assign _2382_ = _2136_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:413.6-444.13" */ { mem_rdata_latched[11:9], 1'h0 } : _2380_;
  assign _2384_ = _0442_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:362.6-411.13" */ { mem_rdata_latched[11:10], mem_rdata_latched[4:3] } : _2380_;
  assign _2386_ = _2136_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:347.6-360.13" */ { mem_rdata_latched[11:10], mem_rdata_latched[6], 1'h0 } : _2380_;
  assign _0014_[11:8] = _1722_ ? /* src = "generated/out/vanilla.sv:344.7-344.72|generated/out/vanilla.sv:344.3-445.11" */ _1589_ : _2380_;
  assign _2388_ = mem_xfer ? /* src = "generated/out/vanilla.sv:340.7-340.15|generated/out/vanilla.sv:340.3-343.6" */ mem_rdata_latched[30:25] : mem_rdata_q[30:25];
  assign _2390_ = _1723_ ? /* src = "generated/out/vanilla.sv:423.12-423.73|generated/out/vanilla.sv:423.8-426.11" */ 6'h00 : _2388_;
  assign _2392_ = _1724_ ? /* src = "generated/out/vanilla.sv:427.12-427.73|generated/out/vanilla.sv:427.8-430.11" */ 6'h00 : _2390_;
  assign _2394_ = _1726_ ? /* src = "generated/out/vanilla.sv:431.12-431.109|generated/out/vanilla.sv:431.8-434.11" */ 6'h00 : _2392_;
  assign _2396_ = _1727_ ? /* src = "generated/out/vanilla.sv:435.12-435.73|generated/out/vanilla.sv:435.8-438.11" */ 6'h00 : _2394_;
  assign _2398_ = _1645_ ? /* src = "generated/out/vanilla.sv:379.12-379.45|generated/out/vanilla.sv:379.8-382.11" */ 6'h00 : _2388_;
  assign _2400_ = _1646_ ? /* src = "generated/out/vanilla.sv:383.12-383.45|generated/out/vanilla.sv:383.8-386.11" */ 6'h20 : _2398_;
  assign _2402_ = _1647_ ? /* src = "generated/out/vanilla.sv:387.12-387.45|generated/out/vanilla.sv:387.8-390.11" */ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] } : _2400_;
  assign _2404_ = _1648_ ? /* src = "generated/out/vanilla.sv:391.12-391.46|generated/out/vanilla.sv:391.8-401.11" */ _2446_[5:0] : _2402_;
  assign _2406_ = _1644_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:372.12-372.40|generated/out/vanilla.sv:372.8-377.88" */ { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[4:3], mem_rdata_latched[5], mem_rdata_latched[2] } : { mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12], mem_rdata_latched[12] };
  assign _0014_[30:25] = _1722_ ? /* src = "generated/out/vanilla.sv:344.7-344.72|generated/out/vanilla.sv:344.3-445.11" */ _1603_ : _2388_;
  assign _2408_ = pcpi_rs1[1:0] == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:331.5-336.12" */ 2'h3;
  assign _2409_ = pcpi_rs1[1:0] == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:331.5-336.12" */ 2'h2;
  assign _2410_ = pcpi_rs1[1:0] == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:331.5-336.12" */ 2'h1;
  assign _2411_ = mem_wordsize == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:314.3-338.10" */ 2'h2;
  assign _1637_ = mem_wordsize == /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:314.3-338.10" */ 2'h1;
  assign _1636_ = ! /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:314.3-338.10" */ mem_wordsize;
  assign _2412_ = last_mem_valid ? /* src = "generated/out/vanilla.sv:308.8-308.23|generated/out/vanilla.sv:308.4-309.46" */ mem_la_firstword_reg : mem_la_firstword;
  assign _0055_ = _1643_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1805.8-1805.35|generated/out/vanilla.sv:1805.4-1808.7" */ { rvfi_rd_wdata, 32'h00000000 } : _0040_;
  assign _0057_ = _1643_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1805.8-1805.35|generated/out/vanilla.sv:1805.4-1808.7" */ 64'hffffffff00000000 : _0042_;
  assign _0040_ = _1642_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1801.8-1801.35|generated/out/vanilla.sv:1801.4-1804.7" */ { 32'h00000000, rvfi_rd_wdata } : 64'h0000000000000000;
  assign _0042_ = _1642_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1801.8-1801.35|generated/out/vanilla.sv:1801.4-1804.7" */ 64'h00000000ffffffff : 64'h0000000000000000;
  assign _0052_ = _1641_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1797.8-1797.35|generated/out/vanilla.sv:1797.4-1800.7" */ { rvfi_rd_wdata, 32'h00000000 } : _0037_;
  assign _0054_ = _1641_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1797.8-1797.35|generated/out/vanilla.sv:1797.4-1800.7" */ 64'hffffffff00000000 : _0039_;
  assign _0037_ = _1640_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1793.8-1793.35|generated/out/vanilla.sv:1793.4-1796.7" */ { 32'h00000000, rvfi_rd_wdata } : 64'h0000000000000000;
  assign _2413_ = & /* src = "generated/out/vanilla.sv:296.113-296.123" */ mem_state;
  assign _2414_ = & /* src = "generated/out/vanilla.sv:298.265-298.288" */ mem_rdata_latched[1:0];
  assign _2415_ = & /* src = "generated/out/vanilla.sv:506.13-506.29" */ mem_rdata[1:0];
  assign _2277_ = & /* src = "generated/out/vanilla.sv:779.9-779.31" */ next_insn_opcode[1:0];
  assign _2052_ = | /* src = "generated/out/vanilla.sv:0.0-0.0" */ pcpi_timeout_counter;
  assign _2416_ = | /* src = "generated/out/vanilla.sv:1186.19-1186.57" */ decoded_rs1;
  assign _2417_ = | /* src = "generated/out/vanilla.sv:1187.19-1187.57" */ decoded_rs2;
  assign _2418_ = | /* src = "generated/out/vanilla.sv:1746.22-1746.53" */ latched_rd;
  assign _2419_ = | /* src = "generated/out/vanilla.sv:1776.24-1776.46" */ mem_wstrb;
  assign _2221_ = | /* src = "generated/out/vanilla.sv:1002.5-1002.30" */ { instr_auipc, instr_lui };
  assign pcpi_int_wait = | /* src = "generated/out/vanilla.sv:256.19-256.125" */ { pcpi_div_wait, pcpi_mul_wait };
  assign _2420_ = | /* src = "generated/out/vanilla.sv:296.44-296.54" */ mem_state;
  assign is_rdcycle_rdcycleh_rdinstr_rdinstrh = | /* src = "generated/out/vanilla.sv:610.48-610.111" */ { instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle };
  assign _0011_ = | /* src = "generated/out/vanilla.sv:790.23-790.59" */ { instr_jal, instr_auipc, instr_lui };
  assign _0012_ = | /* src = "generated/out/vanilla.sv:792.22-792.57" */ { instr_slt, instr_slti, instr_blt };
  assign _0013_ = | /* src = "generated/out/vanilla.sv:793.25-793.63" */ { instr_sltu, instr_sltiu, instr_bltu };
  assign _2421_ = | /* src = "generated/out/vanilla.sv:795.17-795.96" */ { is_beq_bne_blt_bge_bltu_bgeu, instr_sltu, instr_slt, instr_sltiu, instr_slti };
  assign _2422_ = | /* src = "generated/out/vanilla.sv:827.27-827.51" */ mem_rdata_latched[12:5];
  assign _2424_ = | /* src = "generated/out/vanilla.sv:995.78-995.259" */ { _1673_, _1672_, _1671_, _1670_, _1668_, _1666_ };
  assign _2423_ = | /* src = "generated/out/vanilla.sv:996.40-996.251" */ { _1796_, _1795_, _1794_ };
  assign _2425_ = 4'h1 << /* src = "generated/out/vanilla.sv:330.20-330.43" */ pcpi_rs1[1:0];
  assign _2427_ = pcpi_rs1 - /* src = "generated/out/vanilla.sv:1110.32-1110.49" */ pcpi_rs2;
  assign _2429_ = pcpi_timeout_counter - /* src = "generated/out/vanilla.sv:1216.30-1216.54" */ 32'd1;
  assign _2430_ = reg_sh - /* src = "generated/out/vanilla.sv:1591.17-1591.27" */ 32'd4;
  assign _2431_ = reg_sh - /* src = "generated/out/vanilla.sv:1600.17-1600.27" */ 32'd1;
  assign next_pc = _1686_ ? /* src = "generated/out/vanilla.sv:1080.20-1080.80" */ { reg_out[31:1], 1'h0 } : reg_next_pc;
  assign alu_add_sub = instr_sub ? /* src = "generated/out/vanilla.sv:1110.20-1110.69" */ _2427_ : _0066_;
  assign _1025_ = latched_compr ? /* src = "generated/out/vanilla.sv:1163.33-1163.54" */ 32'd2 : 32'd4;
  assign cpuregs_rs1 = _2416_ ? /* src = "generated/out/vanilla.sv:1186.19-1186.57" */ _2002_ : 32'd0;
  assign cpuregs_rs2 = _2417_ ? /* src = "generated/out/vanilla.sv:1187.19-1187.57" */ _2004_ : 32'd0;
  assign _2434_ = latched_store ? /* src = "generated/out/vanilla.sv:1280.37-1280.109" */ { _0092_[31:1], 1'h0 } : reg_next_pc;
  assign { _0092_[31:1], _2432_[0] } = latched_stalu ? /* src = "generated/out/vanilla.sv:1299.54-1299.89" */ alu_out_q : reg_out;
  assign _1028_ = compressed_instr ? /* src = "generated/out/vanilla.sv:1331.36-1331.60" */ 32'd2 : 32'd4;
  assign _2436_ = instr_lui ? /* src = "generated/out/vanilla.sv:1405.20-1405.42" */ 32'd0 : reg_pc;
  assign _2438_ = _2418_ ? /* src = "generated/out/vanilla.sv:1746.22-1746.53" */ cpuregs_wrdata : 32'd0;
  assign _2440_ = _2419_ ? /* src = "generated/out/vanilla.sv:1776.24-1776.46" */ 32'd0 : 32'd4294967295;
  assign mem_la_addr = _1707_ ? /* src = "generated/out/vanilla.sv:299.24-299.129" */ { _0084_, 2'h0 } : { pcpi_rs1[31:2], 2'h0 };
  assign mem_rdata_latched_noshuffle = mem_xfer ? /* src = "generated/out/vanilla.sv:300.40-300.95" */ mem_rdata : mem_rdata_q;
  assign mem_rdata_latched = mem_la_use_prefetched_high_word ? /* src = "generated/out/vanilla.sv:301.30-301.348" */ { 16'hxxxx, mem_16bit_buffer } : _2443_;
  assign _2441_ = mem_la_firstword ? /* src = "generated/out/vanilla.sv:301.221-301.346" */ { 16'hxxxx, mem_rdata_latched_noshuffle[31:16] } : mem_rdata_latched_noshuffle;
  assign _2443_ = mem_la_secondword ? /* src = "generated/out/vanilla.sv:301.126-301.347" */ { mem_rdata_latched_noshuffle[15:0], mem_16bit_buffer } : _2441_;
  assign _2445_ = pcpi_rs1[1] ? /* src = "generated/out/vanilla.sv:322.21-322.51" */ 4'hc : 4'h3;
  assign _2446_ = _1649_ ? /* src = "generated/out/vanilla.sv:400.32-400.89" */ 7'h20 : 7'h00;
  assign _2447_ = _1837_ ? /* src = "generated/out/vanilla.sv:512.22-512.58" */ 32'd0 : 32'd3;
  assign _2448_ = pcpi_rs1 ^ /* src = "generated/out/vanilla.sv:1135.39-1135.56" */ pcpi_rs2;
  /* module_not_derived = 32'd1 */
  /* src = "generated/out/vanilla.sv:213.22-224.5" */
  picorv32_pcpi_mul \genblk1.genblk1.pcpi_mul  (
    .clk(clk),
    .pcpi_insn(pcpi_insn),
    .pcpi_insn_t0(pcpi_insn_t0),
    .pcpi_rd(pcpi_mul_rd),
    .pcpi_rd_t0(pcpi_mul_rd_t0),
    .pcpi_ready(pcpi_mul_ready),
    .pcpi_ready_t0(pcpi_mul_ready_t0),
    .pcpi_rs1(pcpi_rs1),
    .pcpi_rs1_t0(pcpi_rs1_t0),
    .pcpi_rs2(pcpi_rs2),
    .pcpi_rs2_t0(pcpi_rs2_t0),
    .pcpi_valid(pcpi_valid),
    .pcpi_valid_t0(pcpi_valid_t0),
    .pcpi_wait(pcpi_mul_wait),
    .pcpi_wait_t0(pcpi_mul_wait_t0),
    .pcpi_wr(pcpi_mul_wr),
    .pcpi_wr_t0(pcpi_mul_wr_t0),
    .resetn(resetn)
  );
  /* module_not_derived = 32'd1 */
  /* src = "generated/out/vanilla.sv:233.22-244.5" */
  picorv32_pcpi_div \genblk2.pcpi_div  (
    .clk(clk),
    .pcpi_insn(pcpi_insn),
    .pcpi_insn_t0(pcpi_insn_t0),
    .pcpi_rd(pcpi_div_rd),
    .pcpi_rd_t0(pcpi_div_rd_t0),
    .pcpi_ready(pcpi_div_ready),
    .pcpi_ready_t0(pcpi_div_ready_t0),
    .pcpi_rs1(pcpi_rs1),
    .pcpi_rs1_t0(pcpi_rs1_t0),
    .pcpi_rs2(pcpi_rs2),
    .pcpi_rs2_t0(pcpi_rs2_t0),
    .pcpi_valid(pcpi_valid),
    .pcpi_valid_t0(pcpi_valid_t0),
    .pcpi_wait(pcpi_div_wait),
    .pcpi_wait_t0(pcpi_div_wait_t0),
    .pcpi_wr(pcpi_div_wr),
    .pcpi_wr_t0(pcpi_div_wr_t0),
    .resetn(resetn)
  );
  assign _0003_[30:0] = { _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31], _0003_[31] };
  assign _0092_[0] = 1'h0;
  assign _0093_[0] = 1'h0;
  assign _2432_[31:1] = _0092_[31:1];
  assign _2433_[31:1] = _0093_[31:1];
  assign decoded_imm_j[0] = 1'h0;
  assign decoded_imm_j_t0[0] = 1'h0;
  assign eoi = 32'd0;
  assign eoi_t0 = 32'd0;
  assign mem_la_read_t0 = 1'h0;
  assign mem_la_write_t0 = 1'h0;
  assign rvfi_csr_mcycle_rmask_t0 = 64'h0000000000000000;
  assign rvfi_csr_mcycle_wdata = 64'h0000000000000000;
  assign rvfi_csr_mcycle_wdata_t0 = 64'h0000000000000000;
  assign rvfi_csr_mcycle_wmask = 64'h0000000000000000;
  assign rvfi_csr_mcycle_wmask_t0 = 64'h0000000000000000;
  assign rvfi_csr_minstret_rmask_t0 = 64'h0000000000000000;
  assign rvfi_csr_minstret_wdata = 64'h0000000000000000;
  assign rvfi_csr_minstret_wdata_t0 = 64'h0000000000000000;
  assign rvfi_csr_minstret_wmask = 64'h0000000000000000;
  assign rvfi_csr_minstret_wmask_t0 = 64'h0000000000000000;
  assign rvfi_halt_t0 = 1'h0;
  assign rvfi_intr = 1'h0;
  assign rvfi_intr_t0 = 1'h0;
  assign rvfi_ixl = 2'h1;
  assign rvfi_ixl_t0 = 2'h0;
  assign rvfi_mode = 2'h3;
  assign rvfi_mode_t0 = 2'h0;
  assign rvfi_trap = rvfi_halt;
  assign rvfi_trap_t0 = 1'h0;
  assign rvfi_valid_t0 = 1'h0;
  assign trace_data = 36'hxxxxxxxxx;
  assign trace_data_t0 = 36'h000000000;
  assign trace_valid = 1'h0;
  assign trace_valid_t0 = 1'h0;
  assign trap_t0 = 1'h0;
endmodule

/* cellift =  1  */
/* hdlname = "\\picorv32_mem_top" */
/* top =  1  */
/* src = "generated/out/vanilla.sv:2703.1-2890.10" */
module picorv32_mem_top(clk, resetn, trap, instr_mem_req, instr_mem_gnt, instr_mem_addr, instr_mem_wdata, instr_mem_strb, instr_mem_we, instr_mem_rdata, data_mem_req, data_mem_gnt, data_mem_addr, data_mem_wdata, data_mem_strb, data_mem_we, data_mem_rdata, mem_la_read, mem_la_write, mem_la_addr, mem_la_wdata
, mem_la_wstrb, pcpi_valid, pcpi_insn, pcpi_rs1, pcpi_rs2, pcpi_wr, pcpi_rd, pcpi_wait, pcpi_ready, irq, eoi, trace_valid, trace_data, trap_t0, trace_valid_t0, trace_data_t0, mem_la_wstrb_t0, mem_la_write_t0, mem_la_wdata_t0, mem_la_read_t0, mem_la_addr_t0
, irq_t0, eoi_t0, pcpi_insn_t0, pcpi_rd_t0, pcpi_ready_t0, pcpi_rs1_t0, pcpi_rs2_t0, pcpi_valid_t0, pcpi_wait_t0, pcpi_wr_t0, data_mem_addr_t0, data_mem_gnt_t0, data_mem_rdata_t0, data_mem_req_t0, data_mem_strb_t0, data_mem_wdata_t0, data_mem_we_t0, instr_mem_addr_t0, instr_mem_gnt_t0, instr_mem_rdata_t0, instr_mem_req_t0
, instr_mem_strb_t0, instr_mem_wdata_t0, instr_mem_we_t0);
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _00_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _01_;
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire _02_;
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [3:0] _03_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [3:0] _04_;
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _05_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _06_;
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _07_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _08_;
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _09_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _10_;
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _11_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2781.2-2817.5" */
  wire [31:0] _12_;
  wire [31:0] _13_;
  wire [31:0] _14_;
  wire [3:0] _15_;
  wire [31:0] _16_;
  wire [31:0] _17_;
  wire [31:0] _18_;
  wire [3:0] _19_;
  wire [31:0] _20_;
  wire [31:0] _21_;
  /* src = "generated/out/vanilla.sv:2739.8-2739.11" */
  input clk;
  wire clk;
  /* src = "generated/out/vanilla.sv:2751.20-2751.33" */
  output [31:0] data_mem_addr;
  wire [31:0] data_mem_addr;
  /* cellift = 32'd1 */
  output [31:0] data_mem_addr_t0;
  wire [31:0] data_mem_addr_t0;
  /* src = "generated/out/vanilla.sv:2750.13-2750.25" */
  input data_mem_gnt;
  wire data_mem_gnt;
  /* cellift = 32'd1 */
  input data_mem_gnt_t0;
  wire data_mem_gnt_t0;
  /* src = "generated/out/vanilla.sv:2755.20-2755.34" */
  input [31:0] data_mem_rdata;
  wire [31:0] data_mem_rdata;
  /* cellift = 32'd1 */
  input [31:0] data_mem_rdata_t0;
  wire [31:0] data_mem_rdata_t0;
  /* src = "generated/out/vanilla.sv:2749.13-2749.25" */
  output data_mem_req;
  wire data_mem_req;
  /* cellift = 32'd1 */
  output data_mem_req_t0;
  wire data_mem_req_t0;
  /* src = "generated/out/vanilla.sv:2753.19-2753.32" */
  output [3:0] data_mem_strb;
  wire [3:0] data_mem_strb;
  /* cellift = 32'd1 */
  output [3:0] data_mem_strb_t0;
  wire [3:0] data_mem_strb_t0;
  /* src = "generated/out/vanilla.sv:2752.20-2752.34" */
  output [31:0] data_mem_wdata;
  wire [31:0] data_mem_wdata;
  /* cellift = 32'd1 */
  output [31:0] data_mem_wdata_t0;
  wire [31:0] data_mem_wdata_t0;
  /* src = "generated/out/vanilla.sv:2754.13-2754.24" */
  output data_mem_we;
  wire data_mem_we;
  /* cellift = 32'd1 */
  output data_mem_we_t0;
  wire data_mem_we_t0;
  /* src = "generated/out/vanilla.sv:2770.20-2770.23" */
  output [31:0] eoi;
  wire [31:0] eoi;
  /* cellift = 32'd1 */
  output [31:0] eoi_t0;
  wire [31:0] eoi_t0;
  /* src = "generated/out/vanilla.sv:2744.20-2744.34" */
  output [31:0] instr_mem_addr;
  wire [31:0] instr_mem_addr;
  /* cellift = 32'd1 */
  output [31:0] instr_mem_addr_t0;
  wire [31:0] instr_mem_addr_t0;
  /* src = "generated/out/vanilla.sv:2743.13-2743.26" */
  input instr_mem_gnt;
  wire instr_mem_gnt;
  /* cellift = 32'd1 */
  input instr_mem_gnt_t0;
  wire instr_mem_gnt_t0;
  /* src = "generated/out/vanilla.sv:2748.20-2748.35" */
  input [31:0] instr_mem_rdata;
  wire [31:0] instr_mem_rdata;
  /* cellift = 32'd1 */
  input [31:0] instr_mem_rdata_t0;
  wire [31:0] instr_mem_rdata_t0;
  /* src = "generated/out/vanilla.sv:2742.13-2742.26" */
  output instr_mem_req;
  wire instr_mem_req;
  /* cellift = 32'd1 */
  output instr_mem_req_t0;
  wire instr_mem_req_t0;
  /* src = "generated/out/vanilla.sv:2746.19-2746.33" */
  output [3:0] instr_mem_strb;
  wire [3:0] instr_mem_strb;
  /* cellift = 32'd1 */
  output [3:0] instr_mem_strb_t0;
  wire [3:0] instr_mem_strb_t0;
  /* src = "generated/out/vanilla.sv:2745.20-2745.35" */
  output [31:0] instr_mem_wdata;
  wire [31:0] instr_mem_wdata;
  /* cellift = 32'd1 */
  output [31:0] instr_mem_wdata_t0;
  wire [31:0] instr_mem_wdata_t0;
  /* src = "generated/out/vanilla.sv:2747.13-2747.25" */
  output instr_mem_we;
  wire instr_mem_we;
  /* cellift = 32'd1 */
  output instr_mem_we_t0;
  wire instr_mem_we_t0;
  /* src = "generated/out/vanilla.sv:2769.15-2769.18" */
  input [31:0] irq;
  wire [31:0] irq;
  /* cellift = 32'd1 */
  input [31:0] irq_t0;
  wire [31:0] irq_t0;
  /* src = "generated/out/vanilla.sv:2776.14-2776.22" */
  /* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] mem_addr;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2776.14-2776.22" */
  /* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] mem_addr_t0;
  /* src = "generated/out/vanilla.sv:2774.7-2774.16" */
  wire mem_instr;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2774.7-2774.16" */
  /* unused_bits = "0" */
  wire mem_instr_t0;
  /* src = "generated/out/vanilla.sv:2758.21-2758.32" */
  output [31:0] mem_la_addr;
  wire [31:0] mem_la_addr;
  /* cellift = 32'd1 */
  output [31:0] mem_la_addr_t0;
  wire [31:0] mem_la_addr_t0;
  /* src = "generated/out/vanilla.sv:2756.14-2756.25" */
  output mem_la_read;
  wire mem_la_read;
  /* cellift = 32'd1 */
  output mem_la_read_t0;
  wire mem_la_read_t0;
  /* src = "generated/out/vanilla.sv:2759.20-2759.32" */
  output [31:0] mem_la_wdata;
  wire [31:0] mem_la_wdata;
  /* cellift = 32'd1 */
  output [31:0] mem_la_wdata_t0;
  wire [31:0] mem_la_wdata_t0;
  /* src = "generated/out/vanilla.sv:2757.14-2757.26" */
  output mem_la_write;
  wire mem_la_write;
  /* cellift = 32'd1 */
  output mem_la_write_t0;
  wire mem_la_write_t0;
  /* src = "generated/out/vanilla.sv:2760.19-2760.31" */
  output [3:0] mem_la_wstrb;
  wire [3:0] mem_la_wstrb;
  /* cellift = 32'd1 */
  output [3:0] mem_la_wstrb_t0;
  wire [3:0] mem_la_wstrb_t0;
  /* src = "generated/out/vanilla.sv:2779.13-2779.22" */
  wire [31:0] mem_rdata;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2779.13-2779.22" */
  wire [31:0] mem_rdata_t0;
  /* src = "generated/out/vanilla.sv:2775.7-2775.16" */
  wire mem_ready;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2775.7-2775.16" */
  wire mem_ready_t0;
  /* src = "generated/out/vanilla.sv:2777.14-2777.23" */
  /* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] mem_wdata;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2777.14-2777.23" */
  /* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] mem_wdata_t0;
  /* src = "generated/out/vanilla.sv:2778.13-2778.22" */
  /* unused_bits = "0 1 2 3" */
  wire [3:0] mem_wstrb;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2778.13-2778.22" */
  /* unused_bits = "0 1 2 3" */
  wire [3:0] mem_wstrb_t0;
  /* src = "generated/out/vanilla.sv:2762.20-2762.29" */
  output [31:0] pcpi_insn;
  wire [31:0] pcpi_insn;
  /* cellift = 32'd1 */
  output [31:0] pcpi_insn_t0;
  wire [31:0] pcpi_insn_t0;
  /* src = "generated/out/vanilla.sv:2766.15-2766.22" */
  input [31:0] pcpi_rd;
  wire [31:0] pcpi_rd;
  /* cellift = 32'd1 */
  input [31:0] pcpi_rd_t0;
  wire [31:0] pcpi_rd_t0;
  /* src = "generated/out/vanilla.sv:2768.8-2768.18" */
  input pcpi_ready;
  wire pcpi_ready;
  /* cellift = 32'd1 */
  input pcpi_ready_t0;
  wire pcpi_ready_t0;
  /* src = "generated/out/vanilla.sv:2763.21-2763.29" */
  output [31:0] pcpi_rs1;
  wire [31:0] pcpi_rs1;
  /* cellift = 32'd1 */
  output [31:0] pcpi_rs1_t0;
  wire [31:0] pcpi_rs1_t0;
  /* src = "generated/out/vanilla.sv:2764.21-2764.29" */
  output [31:0] pcpi_rs2;
  wire [31:0] pcpi_rs2;
  /* cellift = 32'd1 */
  output [31:0] pcpi_rs2_t0;
  wire [31:0] pcpi_rs2_t0;
  /* src = "generated/out/vanilla.sv:2761.13-2761.23" */
  output pcpi_valid;
  wire pcpi_valid;
  /* cellift = 32'd1 */
  output pcpi_valid_t0;
  wire pcpi_valid_t0;
  /* src = "generated/out/vanilla.sv:2767.8-2767.17" */
  input pcpi_wait;
  wire pcpi_wait;
  /* cellift = 32'd1 */
  input pcpi_wait_t0;
  wire pcpi_wait_t0;
  /* src = "generated/out/vanilla.sv:2765.8-2765.15" */
  input pcpi_wr;
  wire pcpi_wr;
  /* cellift = 32'd1 */
  input pcpi_wr_t0;
  wire pcpi_wr_t0;
  /* src = "generated/out/vanilla.sv:2740.8-2740.14" */
  input resetn;
  wire resetn;
  /* src = "generated/out/vanilla.sv:2772.20-2772.30" */
  output [35:0] trace_data;
  wire [35:0] trace_data;
  /* cellift = 32'd1 */
  output [35:0] trace_data_t0;
  wire [35:0] trace_data_t0;
  /* src = "generated/out/vanilla.sv:2771.13-2771.24" */
  output trace_valid;
  wire trace_valid;
  /* cellift = 32'd1 */
  output trace_valid_t0;
  wire trace_valid_t0;
  /* src = "generated/out/vanilla.sv:2741.13-2741.17" */
  output trap;
  wire trap;
  /* cellift = 32'd1 */
  output trap_t0;
  wire trap_t0;
  assign _13_ = ~ { mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr };
  assign _14_ = ~ { mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write };
  assign _16_ = ~ { mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read };
  assign _15_ = ~ { mem_la_read, mem_la_read, mem_la_read, mem_la_read };
  assign _17_ = _13_ & data_mem_rdata_t0;
  assign _08_ = _14_ & _10_;
  assign _19_ = _15_ & _04_;
  assign _20_ = _16_ & _06_;
  assign _21_ = _16_ & _01_;
  assign mem_rdata_t0 = _16_ & _08_;
  assign _18_ = { mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr, mem_instr } & instr_mem_rdata_t0;
  assign _10_ = { mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready, mem_ready } & _12_;
  assign _04_ = { mem_la_write, mem_la_write, mem_la_write, mem_la_write } & mem_la_wstrb_t0;
  assign _06_ = { mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write } & mem_la_wdata_t0;
  assign _01_ = { mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write, mem_la_write } & mem_la_addr_t0;
  assign instr_mem_strb_t0 = { mem_la_read, mem_la_read, mem_la_read, mem_la_read } & mem_la_wstrb_t0;
  assign instr_mem_wdata_t0 = { mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read } & mem_la_wdata_t0;
  assign instr_mem_addr_t0 = { mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read, mem_la_read } & mem_la_addr_t0;
  assign _12_ = _17_ | _18_;
  assign data_mem_strb_t0 = _19_ | instr_mem_strb_t0;
  assign data_mem_wdata_t0 = _20_ | instr_mem_wdata_t0;
  assign data_mem_addr_t0 = _21_ | instr_mem_addr_t0;
  assign _11_ = mem_instr ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2813.8-2813.17|generated/out/vanilla.sv:2813.4-2816.32" */ instr_mem_rdata : data_mem_rdata;
  assign _09_ = mem_ready ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2812.12-2812.21|generated/out/vanilla.sv:2812.8-2816.32" */ _11_ : 32'd0;
  assign _03_ = mem_la_write ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2805.12-2805.24|generated/out/vanilla.sv:2805.8-2816.32" */ mem_la_wstrb : 4'h0;
  assign _05_ = mem_la_write ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2805.12-2805.24|generated/out/vanilla.sv:2805.8-2816.32" */ mem_la_wdata : 32'd0;
  assign _00_ = mem_la_write ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2805.12-2805.24|generated/out/vanilla.sv:2805.8-2816.32" */ mem_la_addr : 32'd0;
  assign _02_ = mem_la_write ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2805.12-2805.24|generated/out/vanilla.sv:2805.8-2816.32" */ 1'h1 : 1'h0;
  assign _07_ = mem_la_write ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2805.12-2805.24|generated/out/vanilla.sv:2805.8-2816.32" */ 32'd0 : _09_;
  assign data_mem_we = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ 1'h0 : _02_;
  assign data_mem_strb = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ mem_la_wstrb : _03_;
  assign data_mem_wdata = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ mem_la_wdata : _05_;
  assign data_mem_addr = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ mem_la_addr : _00_;
  assign data_mem_req = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ 1'h1 : _02_;
  assign instr_mem_strb = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ mem_la_wstrb : 4'h0;
  assign instr_mem_wdata = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ mem_la_wdata : 32'd0;
  assign instr_mem_addr = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ mem_la_addr : 32'd0;
  assign instr_mem_req = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ 1'h1 : 1'h0;
  assign mem_rdata = mem_la_read ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2793.7-2793.18|generated/out/vanilla.sv:2793.3-2816.32" */ 32'd0 : _07_;
  /* module_not_derived = 32'd1 */
  /* src = "generated/out/vanilla.sv:2861.4-2889.3" */
  cellift_data_flow_picorv32  i_picorv32 (
    .clk(clk),
    .eoi(eoi),
    .eoi_t0(eoi_t0),
    .irq(irq),
    .irq_t0(irq_t0),
    .mem_addr(mem_addr),
    .mem_addr_t0(mem_addr_t0),
    .mem_instr(mem_instr),
    .mem_instr_t0(mem_instr_t0),
    .mem_la_addr(mem_la_addr),
    .mem_la_addr_t0(mem_la_addr_t0),
    .mem_la_read(mem_la_read),
    .mem_la_read_t0(mem_la_read_t0),
    .mem_la_wdata(mem_la_wdata),
    .mem_la_wdata_t0(mem_la_wdata_t0),
    .mem_la_write(mem_la_write),
    .mem_la_write_t0(mem_la_write_t0),
    .mem_la_wstrb(mem_la_wstrb),
    .mem_la_wstrb_t0(mem_la_wstrb_t0),
    .mem_rdata(mem_rdata),
    .mem_rdata_t0(mem_rdata_t0),
    .mem_ready(mem_ready),
    .mem_ready_t0(mem_ready_t0),
    .mem_valid(mem_ready),
    .mem_valid_t0(mem_ready_t0),
    .mem_wdata(mem_wdata),
    .mem_wdata_t0(mem_wdata_t0),
    .mem_wstrb(mem_wstrb),
    .mem_wstrb_t0(mem_wstrb_t0),
    .pcpi_insn(pcpi_insn),
    .pcpi_insn_t0(pcpi_insn_t0),
    .pcpi_rd(pcpi_rd),
    .pcpi_rd_t0(pcpi_rd_t0),
    .pcpi_ready(pcpi_ready),
    .pcpi_ready_t0(pcpi_ready_t0),
    .pcpi_rs1(pcpi_rs1),
    .pcpi_rs1_t0(pcpi_rs1_t0),
    .pcpi_rs2(pcpi_rs2),
    .pcpi_rs2_t0(pcpi_rs2_t0),
    .pcpi_valid(pcpi_valid),
    .pcpi_valid_t0(pcpi_valid_t0),
    .pcpi_wait(pcpi_wait),
    .pcpi_wait_t0(pcpi_wait_t0),
    .pcpi_wr(pcpi_wr),
    .pcpi_wr_t0(pcpi_wr_t0),
    .resetn(resetn),
    .trace_data(trace_data),
    .trace_data_t0(trace_data_t0),
    .trace_valid(trace_valid),
    .trace_valid_t0(trace_valid_t0),
    .trap(trap),
    .trap_t0(trap_t0)
  );
  assign data_mem_req_t0 = 1'h0;
  assign data_mem_we_t0 = 1'h0;
  assign instr_mem_req_t0 = 1'h0;
  assign instr_mem_we = 1'h0;
  assign instr_mem_we_t0 = 1'h0;
endmodule

/* cellift =  1  */
/* hdlname = "\\picorv32_pcpi_div" */
/* src = "generated/out/vanilla.sv:2055.1-2137.10" */
module picorv32_pcpi_div(clk, resetn, pcpi_valid, pcpi_insn, pcpi_rs1, pcpi_rs2, pcpi_wr, pcpi_rd, pcpi_wait, pcpi_ready, pcpi_insn_t0, pcpi_rd_t0, pcpi_ready_t0, pcpi_rs1_t0, pcpi_rs2_t0, pcpi_valid_t0, pcpi_wait_t0, pcpi_wr_t0);
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
  wire [31:0] _000_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
  wire [31:0] _001_;
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
  wire _002_;
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
  wire _003_;
  wire _004_;
  wire _005_;
  wire [31:0] _006_;
  wire [31:0] _007_;
  wire [31:0] _008_;
  wire [62:0] _009_;
  wire [62:0] _010_;
  wire [31:0] _011_;
  wire [62:0] _012_;
  wire [31:0] _013_;
  wire [31:0] _014_;
  wire [62:0] _015_;
  wire [31:0] _016_;
  wire [31:0] _017_;
  wire [31:0] _018_;
  wire [62:0] _019_;
  wire [31:0] _020_;
  wire [31:0] _021_;
  wire [31:0] _022_;
  wire [62:0] _023_;
  wire [31:0] _024_;
  wire [31:0] _025_;
  wire _026_;
  wire [31:0] _027_;
  wire [31:0] _028_;
  wire [62:0] _029_;
  wire [62:0] _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire [31:0] _038_;
  wire [31:0] _039_;
  wire [31:0] _040_;
  wire [31:0] _041_;
  wire [31:0] _042_;
  wire [31:0] _043_;
  wire [30:0] _044_;
  wire [30:0] _045_;
  wire [31:0] _046_;
  wire [31:0] _047_;
  wire [31:0] _048_;
  wire [62:0] _049_;
  wire [31:0] _050_;
  wire [31:0] _051_;
  wire [31:0] _052_;
  wire [31:0] _053_;
  wire [31:0] _054_;
  wire [31:0] _055_;
  wire [31:0] _056_;
  wire [62:0] _057_;
  wire [62:0] _058_;
  wire [31:0] _059_;
  wire [31:0] _060_;
  wire [62:0] _061_;
  wire [62:0] _062_;
  wire [31:0] _063_;
  wire [31:0] _064_;
  wire [62:0] _065_;
  wire [62:0] _066_;
  wire [31:0] _067_;
  wire [31:0] _068_;
  wire [31:0] _069_;
  wire [31:0] _070_;
  wire [31:0] _071_;
  wire [31:0] _072_;
  wire [31:0] _073_;
  wire [30:0] _074_;
  wire [31:0] _075_;
  wire [31:0] _076_;
  wire [62:0] _077_;
  wire [31:0] _078_;
  wire [31:0] _079_;
  wire [31:0] _080_;
  wire [62:0] _081_;
  wire [62:0] _082_;
  wire [62:0] _083_;
  wire [31:0] _084_;
  wire [62:0] _085_;
  wire [31:0] _086_;
  wire [31:0] _087_;
  wire [62:0] _088_;
  wire [62:0] _089_;
  wire [62:0] _090_;
  /* src = "generated/out/vanilla.sv:2089.52-2089.80" */
  wire _091_;
  /* src = "generated/out/vanilla.sv:2089.87-2089.117" */
  wire _092_;
  /* src = "generated/out/vanilla.sv:2129.8-2129.27" */
  wire _093_;
  /* src = "generated/out/vanilla.sv:2089.10-2089.30" */
  wire _094_;
  /* src = "generated/out/vanilla.sv:2089.9-2089.46" */
  wire _095_;
  /* src = "generated/out/vanilla.sv:2089.8-2089.81" */
  wire _096_;
  /* src = "generated/out/vanilla.sv:2089.7-2089.118" */
  wire _097_;
  /* src = "generated/out/vanilla.sv:2113.17-2113.57" */
  wire _098_;
  /* src = "generated/out/vanilla.sv:2114.16-2114.56" */
  wire _099_;
  /* src = "generated/out/vanilla.sv:2115.17-2115.60" */
  wire _100_;
  /* src = "generated/out/vanilla.sv:2115.16-2115.74" */
  wire _101_;
  /* src = "generated/out/vanilla.sv:2115.80-2115.105" */
  wire _102_;
  /* src = "generated/out/vanilla.sv:2119.12-2119.36" */
  wire _103_;
  /* src = "generated/out/vanilla.sv:2083.28-2083.40" */
  wire _104_;
  /* src = "generated/out/vanilla.sv:2089.35-2089.46" */
  wire _105_;
  /* src = "generated/out/vanilla.sv:2119.12-2119.25" */
  wire _106_;
  /* src = "generated/out/vanilla.sv:2113.18-2113.40" */
  wire _107_;
  /* src = "generated/out/vanilla.sv:2115.15-2115.106" */
  wire _108_;
  /* src = "generated/out/vanilla.sv:2123.8-2123.31" */
  wire _109_;
  /* src = "generated/out/vanilla.sv:2115.31-2115.59" */
  wire _110_;
  /* src = "generated/out/vanilla.sv:2113.60-2113.69" */
  wire [31:0] _111_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2113.60-2113.69" */
  wire [31:0] _112_;
  /* src = "generated/out/vanilla.sv:2114.59-2114.68" */
  wire [62:0] _113_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2114.59-2114.68" */
  wire [62:0] _114_;
  /* src = "generated/out/vanilla.sv:2124.27-2124.36" */
  wire [31:0] _115_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2124.27-2124.36" */
  wire [31:0] _116_;
  /* src = "generated/out/vanilla.sv:2126.27-2126.36" */
  wire [31:0] _117_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2126.27-2126.36" */
  wire [31:0] _118_;
  /* src = "generated/out/vanilla.sv:2131.17-2131.40" */
  wire [31:0] _119_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2131.17-2131.40" */
  wire [31:0] _120_;
  wire [31:0] _121_;
  /* cellift = 32'd1 */
  wire [31:0] _122_;
  wire [31:0] _123_;
  /* cellift = 32'd1 */
  wire [31:0] _124_;
  wire [31:0] _125_;
  /* cellift = 32'd1 */
  wire [31:0] _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire [31:0] _130_;
  /* cellift = 32'd1 */
  wire [31:0] _131_;
  wire [31:0] _132_;
  /* cellift = 32'd1 */
  wire [31:0] _133_;
  wire [31:0] _134_;
  /* cellift = 32'd1 */
  wire [31:0] _135_;
  wire [62:0] _136_;
  /* cellift = 32'd1 */
  wire [62:0] _137_;
  /* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30" */
  wire [62:0] _138_;
  /* cellift = 32'd1 */
  /* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30" */
  wire [62:0] _139_;
  wire [31:0] _140_;
  /* cellift = 32'd1 */
  wire [31:0] _141_;
  wire [31:0] _142_;
  /* cellift = 32'd1 */
  wire [31:0] _143_;
  wire [31:0] _144_;
  /* cellift = 32'd1 */
  wire [31:0] _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  /* src = "generated/out/vanilla.sv:2115.65-2115.74" */
  wire _154_;
  /* src = "generated/out/vanilla.sv:2114.15-2114.86" */
  wire [62:0] _155_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2114.15-2114.86" */
  wire [62:0] _156_;
  /* src = "generated/out/vanilla.sv:2130.17-2130.35" */
  /* unused_bits = "32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62" */
  wire [62:0] _157_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2130.17-2130.35" */
  /* unused_bits = "32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62" */
  wire [62:0] _158_;
  /* src = "generated/out/vanilla.sv:2113.17-2113.80" */
  wire [31:0] _159_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2113.17-2113.80" */
  wire [31:0] _160_;
  /* src = "generated/out/vanilla.sv:2114.16-2114.79" */
  /* unused_bits = "32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62" */
  wire [62:0] _161_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2114.16-2114.79" */
  /* unused_bits = "32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62" */
  wire [62:0] _162_;
  /* src = "generated/out/vanilla.sv:2124.17-2124.47" */
  wire [31:0] _163_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2124.17-2124.47" */
  wire [31:0] _164_;
  /* src = "generated/out/vanilla.sv:2126.17-2126.47" */
  wire [31:0] _165_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2126.17-2126.47" */
  wire [31:0] _166_;
  /* src = "generated/out/vanilla.sv:2067.8-2067.11" */
  input clk;
  wire clk;
  /* src = "generated/out/vanilla.sv:2099.13-2099.21" */
  reg [31:0] dividend;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2099.13-2099.21" */
  reg [31:0] dividend_t0;
  /* src = "generated/out/vanilla.sv:2100.13-2100.20" */
  reg [62:0] divisor;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2100.13-2100.20" */
  reg [62:0] divisor_t0;
  /* src = "generated/out/vanilla.sv:2081.7-2081.24" */
  wire instr_any_div_rem;
  /* src = "generated/out/vanilla.sv:2077.6-2077.15" */
  reg instr_div;
  /* src = "generated/out/vanilla.sv:2078.6-2078.16" */
  reg instr_divu;
  /* src = "generated/out/vanilla.sv:2079.6-2079.15" */
  reg instr_rem;
  /* src = "generated/out/vanilla.sv:2080.6-2080.16" */
  reg instr_remu;
  /* src = "generated/out/vanilla.sv:2104.6-2104.13" */
  reg outsign;
  /* src = "generated/out/vanilla.sv:2070.15-2070.24" */
  input [31:0] pcpi_insn;
  wire [31:0] pcpi_insn;
  /* cellift = 32'd1 */
  input [31:0] pcpi_insn_t0;
  wire [31:0] pcpi_insn_t0;
  /* src = "generated/out/vanilla.sv:2074.20-2074.27" */
  output [31:0] pcpi_rd;
  reg [31:0] pcpi_rd;
  /* cellift = 32'd1 */
  output [31:0] pcpi_rd_t0;
  reg [31:0] pcpi_rd_t0;
  /* src = "generated/out/vanilla.sv:2076.13-2076.23" */
  output pcpi_ready;
  reg pcpi_ready;
  /* cellift = 32'd1 */
  output pcpi_ready_t0;
  wire pcpi_ready_t0;
  /* src = "generated/out/vanilla.sv:2071.15-2071.23" */
  input [31:0] pcpi_rs1;
  wire [31:0] pcpi_rs1;
  /* cellift = 32'd1 */
  input [31:0] pcpi_rs1_t0;
  wire [31:0] pcpi_rs1_t0;
  /* src = "generated/out/vanilla.sv:2072.15-2072.23" */
  input [31:0] pcpi_rs2;
  wire [31:0] pcpi_rs2;
  /* cellift = 32'd1 */
  input [31:0] pcpi_rs2_t0;
  wire [31:0] pcpi_rs2_t0;
  /* src = "generated/out/vanilla.sv:2069.8-2069.18" */
  input pcpi_valid;
  wire pcpi_valid;
  /* cellift = 32'd1 */
  input pcpi_valid_t0;
  wire pcpi_valid_t0;
  /* src = "generated/out/vanilla.sv:2075.13-2075.22" */
  output pcpi_wait;
  reg pcpi_wait;
  /* src = "generated/out/vanilla.sv:2082.6-2082.17" */
  reg pcpi_wait_q;
  /* cellift = 32'd1 */
  output pcpi_wait_t0;
  wire pcpi_wait_t0;
  /* src = "generated/out/vanilla.sv:2073.13-2073.20" */
  output pcpi_wr;
  wire pcpi_wr;
  /* cellift = 32'd1 */
  output pcpi_wr_t0;
  wire pcpi_wr_t0;
  /* src = "generated/out/vanilla.sv:2101.13-2101.21" */
  reg [31:0] quotient;
  /* src = "generated/out/vanilla.sv:2102.13-2102.25" */
  reg [31:0] quotient_msk;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2102.13-2102.25" */
  reg [31:0] quotient_msk_t0;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:2101.13-2101.21" */
  reg [31:0] quotient_t0;
  /* src = "generated/out/vanilla.sv:2068.8-2068.14" */
  input resetn;
  wire resetn;
  /* src = "generated/out/vanilla.sv:2103.6-2103.13" */
  reg running;
  /* src = "generated/out/vanilla.sv:2083.7-2083.12" */
  wire start;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME pcpi_rd_t0 */
  always_ff @(posedge clk)
    pcpi_rd_t0 <= _001_;
  assign _004_ = ~ _036_;
  assign _005_ = ~ _035_;
  assign _040_ = { _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_ } & _145_;
  assign _046_ = { _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_ } & _139_[62:31];
  assign _041_ = { _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_ } & dividend_t0;
  assign _047_ = { _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_ } & divisor_t0[62:31];
  assign _072_ = _040_ | _041_;
  assign _075_ = _046_ | _047_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME dividend_t0 */
  always_ff @(posedge clk)
    dividend_t0 <= _072_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME divisor_t0[62:31] */
  always_ff @(posedge clk)
    divisor_t0[62:31] <= _075_;
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME instr_div */
  always_ff @(posedge clk)
    if (!_097_) instr_div <= 1'h0;
    else instr_div <= _152_;
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME instr_divu */
  always_ff @(posedge clk)
    if (!_097_) instr_divu <= 1'h0;
    else instr_divu <= _150_;
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME instr_remu */
  always_ff @(posedge clk)
    if (!_097_) instr_remu <= 1'h0;
    else instr_remu <= _146_;
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME instr_rem */
  always_ff @(posedge clk)
    if (!_097_) instr_rem <= 1'h0;
    else instr_rem <= _148_;
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME outsign */
  always_ff @(posedge clk)
    if (_034_) outsign <= _108_;
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME running */
  always_ff @(posedge clk)
    if (!resetn) running <= 1'h0;
    else if (_031_) running <= _129_;
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME quotient_msk */
  always_ff @(posedge clk)
    if (_035_)
      if (start) quotient_msk <= 32'd2147483648;
      else quotient_msk <= _130_;
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME pcpi_ready */
  always_ff @(posedge clk)
    if (_037_) pcpi_ready <= 1'h0;
    else pcpi_ready <= _127_;
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME dividend */
  always_ff @(posedge clk)
    if (_036_) dividend <= _144_;
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME quotient */
  always_ff @(posedge clk)
    if (_036_)
      if (start) quotient <= 32'd0;
      else quotient <= _134_;
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME divisor[30:0] */
  always_ff @(posedge clk)
    if (_035_)
      if (start) divisor[30:0] <= 31'h00000000;
      else divisor[30:0] <= _136_[30:0];
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME divisor[62:31] */
  always_ff @(posedge clk)
    if (_035_) divisor[62:31] <= _138_[62:31];
  assign _006_ = ~ { _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_ };
  assign _009_ = ~ { _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_ };
  assign _010_ = ~ { start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start };
  assign _007_ = ~ { _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_ };
  assign _008_ = ~ { start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start };
  assign _011_ = ~ { _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_ };
  assign _012_ = ~ { _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_ };
  assign _013_ = ~ { outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign };
  assign _055_ = _006_ & _166_;
  assign _126_ = _008_ & _124_;
  assign _131_ = _007_ & { 1'h0, quotient_msk_t0[31:1] };
  assign _135_ = _007_ & _133_;
  assign _137_ = _009_ & { 1'h0, divisor_t0[62:1] };
  assign _057_ = _010_ & _137_;
  assign _143_ = _007_ & _141_;
  assign _059_ = _008_ & _143_;
  assign _063_ = _011_ & pcpi_rs1_t0;
  assign _065_ = _012_ & { 31'h00000000, pcpi_rs2_t0 };
  assign _067_ = _013_ & quotient_t0;
  assign _069_ = _013_ & dividend_t0;
  assign _056_ = { _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_ } & _164_;
  assign _124_ = { _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_, _103_ } & _122_;
  assign _001_ = { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn } & _126_;
  assign _133_ = { _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_ } & _120_;
  assign _058_ = { start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start } & { _156_[62:31], 31'h00000000 };
  assign _141_ = { _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_ } & _158_[31:0];
  assign _060_ = { start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start, start } & _160_;
  assign _064_ = { _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_, _098_ } & _112_;
  assign _066_ = { _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_, _099_ } & _114_;
  assign _068_ = { outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign } & _116_;
  assign _070_ = { outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign, outsign } & _118_;
  assign _122_ = _055_ | _056_;
  assign _139_ = _057_ | _058_;
  assign _145_ = _059_ | _060_;
  assign _160_ = _063_ | _064_;
  assign { _162_[62:32], _156_[62:31] } = _065_ | _066_;
  assign _164_ = _067_ | _068_;
  assign _166_ = _069_ | _070_;
  assign _014_ = ~ pcpi_rs1_t0;
  assign _015_ = ~ { 31'h00000000, pcpi_rs2_t0 };
  assign _016_ = ~ quotient_t0;
  assign _017_ = ~ dividend_t0;
  assign _048_ = pcpi_rs1 & _014_;
  assign _049_ = { 31'h00000000, pcpi_rs2 } & _015_;
  assign _050_ = quotient & _016_;
  assign _051_ = dividend & _017_;
  assign _076_ = pcpi_rs1 | pcpi_rs1_t0;
  assign _077_ = { 31'h00000000, pcpi_rs2 } | { 31'h00000000, pcpi_rs2_t0 };
  assign _078_ = quotient | quotient_t0;
  assign _079_ = dividend | dividend_t0;
  assign _018_ = - _048_;
  assign _019_ = - _049_;
  assign _020_ = - _050_;
  assign _021_ = - _051_;
  assign _022_ = - _076_;
  assign _023_ = - _077_;
  assign _024_ = - _078_;
  assign _025_ = - _079_;
  assign _084_ = _018_ ^ _022_;
  assign _085_ = _019_ ^ _023_;
  assign _086_ = _020_ ^ _024_;
  assign _087_ = _021_ ^ _025_;
  assign _112_ = _084_ | pcpi_rs1_t0;
  assign _114_ = _085_ | { 31'h00000000, pcpi_rs2_t0 };
  assign _116_ = _086_ | quotient_t0;
  assign _118_ = _087_ | dividend_t0;
  assign _031_ = | { _103_, start };
  assign _032_ = { _103_, start } != 2'h2;
  assign _033_ = | { _093_, _103_, start };
  assign _034_ = & { start, resetn };
  assign _035_ = & { _032_, resetn };
  assign _036_ = & { _032_, _033_, resetn };
  assign _026_ = ~ resetn;
  assign _037_ = | { _026_, start };
  assign _027_ = ~ quotient;
  assign _028_ = ~ quotient_msk;
  assign _052_ = quotient_t0 & _028_;
  assign _053_ = quotient_msk_t0 & _027_;
  assign _054_ = quotient_t0 & quotient_msk_t0;
  assign _080_ = _052_ | _053_;
  assign _120_ = _080_ | _054_;
  assign _038_ = { _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_ } & _131_;
  assign _042_ = { _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_, _036_ } & _135_;
  assign _044_ = { _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_ } & _137_[30:0];
  assign _039_ = { _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_ } & quotient_msk_t0;
  assign _043_ = { _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_ } & quotient_t0;
  assign _045_ = { _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_, _005_ } & divisor_t0[30:0];
  assign _071_ = _038_ | _039_;
  assign _073_ = _042_ | _043_;
  assign _074_ = _044_ | _045_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME quotient_msk_t0 */
  always_ff @(posedge clk)
    if (start) quotient_msk_t0 <= 32'd0;
    else quotient_msk_t0 <= _071_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME quotient_t0 */
  always_ff @(posedge clk)
    if (start) quotient_t0 <= 32'd0;
    else quotient_t0 <= _073_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME divisor_t0[30:0] */
  always_ff @(posedge clk)
    if (start) divisor_t0[30:0] <= 31'h00000000;
    else divisor_t0[30:0] <= _074_;
  assign _029_ = ~ { 31'h00000000, dividend_t0 };
  assign _030_ = ~ divisor_t0;
  assign _061_ = { 31'h00000000, dividend } & _029_;
  assign _062_ = divisor & _030_;
  assign _081_ = { 31'h00000000, dividend } | { 31'h00000000, dividend_t0 };
  assign _082_ = divisor | divisor_t0;
  assign _089_ = _081_ - _062_;
  assign _090_ = _061_ - _082_;
  assign _088_ = _089_ ^ _090_;
  assign _083_ = _088_ | { 31'h00000000, dividend_t0 };
  assign _158_ = _083_ | divisor_t0;
  assign _091_ = pcpi_insn[6:0] == /* src = "generated/out/vanilla.sv:2089.52-2089.80" */ 7'h33;
  assign _092_ = pcpi_insn[31:25] == /* src = "generated/out/vanilla.sv:2089.87-2089.117" */ 7'h01;
  assign _093_ = divisor <= /* src = "generated/out/vanilla.sv:2129.8-2129.27" */ dividend;
  assign start = pcpi_wait && /* src = "generated/out/vanilla.sv:2083.15-2083.40" */ _104_;
  assign _094_ = resetn && /* src = "generated/out/vanilla.sv:2089.10-2089.30" */ pcpi_valid;
  assign _095_ = _094_ && /* src = "generated/out/vanilla.sv:2089.9-2089.46" */ _105_;
  assign _096_ = _095_ && /* src = "generated/out/vanilla.sv:2089.8-2089.81" */ _091_;
  assign _097_ = _096_ && /* src = "generated/out/vanilla.sv:2089.7-2089.118" */ _092_;
  assign _002_ = instr_any_div_rem && /* src = "generated/out/vanilla.sv:2096.16-2096.43" */ resetn;
  assign _003_ = pcpi_wait && /* src = "generated/out/vanilla.sv:2097.18-2097.37" */ resetn;
  assign _098_ = _107_ && /* src = "generated/out/vanilla.sv:2113.17-2113.57" */ pcpi_rs1[31];
  assign _099_ = _107_ && /* src = "generated/out/vanilla.sv:2114.16-2114.56" */ pcpi_rs2[31];
  assign _100_ = instr_div && /* src = "generated/out/vanilla.sv:2115.17-2115.60" */ _110_;
  assign _101_ = _100_ && /* src = "generated/out/vanilla.sv:2115.16-2115.74" */ _154_;
  assign _102_ = instr_rem && /* src = "generated/out/vanilla.sv:2115.80-2115.105" */ pcpi_rs1[31];
  assign _103_ = _106_ && /* src = "generated/out/vanilla.sv:2119.12-2119.36" */ running;
  assign _104_ = ! /* src = "generated/out/vanilla.sv:2083.28-2083.40" */ pcpi_wait_q;
  assign _105_ = ! /* src = "generated/out/vanilla.sv:2089.35-2089.46" */ pcpi_ready;
  assign _106_ = ! /* src = "generated/out/vanilla.sv:2119.12-2119.25" */ quotient_msk;
  assign _107_ = instr_div || /* src = "generated/out/vanilla.sv:2114.17-2114.39" */ instr_rem;
  assign _108_ = _101_ || /* src = "generated/out/vanilla.sv:2115.15-2115.106" */ _102_;
  assign _109_ = instr_div || /* src = "generated/out/vanilla.sv:2123.8-2123.31" */ instr_divu;
  assign _110_ = pcpi_rs1[31] != /* src = "generated/out/vanilla.sv:2115.31-2115.59" */ pcpi_rs2[31];
  assign _111_ = - /* src = "generated/out/vanilla.sv:2113.60-2113.69" */ pcpi_rs1;
  assign _113_ = - /* src = "generated/out/vanilla.sv:2114.59-2114.68" */ { 31'h00000000, pcpi_rs2 };
  assign _115_ = - /* src = "generated/out/vanilla.sv:2124.27-2124.36" */ quotient;
  assign _117_ = - /* src = "generated/out/vanilla.sv:2126.27-2126.36" */ dividend;
  assign _119_ = quotient | /* src = "generated/out/vanilla.sv:2131.17-2131.40" */ quotient_msk;
  /* src = "generated/out/vanilla.sv:2105.2-2136.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME pcpi_rd */
  always_ff @(posedge clk)
    pcpi_rd <= _000_;
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME pcpi_wait */
  always_ff @(posedge clk)
    pcpi_wait <= _002_;
  /* src = "generated/out/vanilla.sv:2084.2-2098.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_div */
/* PC_TAINT_INFO STATE_NAME pcpi_wait_q */
  always_ff @(posedge clk)
    pcpi_wait_q <= _003_;
  assign _121_ = _109_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2123.8-2123.31|generated/out/vanilla.sv:2123.4-2126.49" */ _163_ : _165_;
  assign _123_ = _103_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2119.12-2119.36|generated/out/vanilla.sv:2119.8-2135.6" */ _121_ : 32'hxxxxxxxx;
  assign _125_ = start ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2111.12-2111.17|generated/out/vanilla.sv:2111.8-2135.6" */ 32'hxxxxxxxx : _123_;
  assign _000_ = resetn ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2109.7-2109.14|generated/out/vanilla.sv:2109.3-2135.6" */ _125_ : 32'hxxxxxxxx;
  assign _127_ = _103_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2119.12-2119.36|generated/out/vanilla.sv:2119.8-2135.6" */ 1'h1 : 1'h0;
  assign _128_ = _103_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2119.12-2119.36|generated/out/vanilla.sv:2119.8-2135.6" */ 1'h0 : 1'hx;
  assign _129_ = start ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2111.12-2111.17|generated/out/vanilla.sv:2111.8-2135.6" */ 1'h1 : _128_;
  assign _130_ = _103_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2119.12-2119.36|generated/out/vanilla.sv:2119.8-2135.6" */ 32'hxxxxxxxx : { 1'h0, quotient_msk[31:1] };
  assign _132_ = _093_ ? /* src = "generated/out/vanilla.sv:2129.8-2129.27|generated/out/vanilla.sv:2129.4-2132.7" */ _119_ : 32'hxxxxxxxx;
  assign _134_ = _103_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2119.12-2119.36|generated/out/vanilla.sv:2119.8-2135.6" */ 32'hxxxxxxxx : _132_;
  assign _136_ = _103_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2119.12-2119.36|generated/out/vanilla.sv:2119.8-2135.6" */ 63'hxxxxxxxxxxxxxxxx : { 1'h0, divisor[62:1] };
  assign _138_ = start ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2111.12-2111.17|generated/out/vanilla.sv:2111.8-2135.6" */ { _155_[62:31], 31'h00000000 } : _136_;
  assign _140_ = _093_ ? /* src = "generated/out/vanilla.sv:2129.8-2129.27|generated/out/vanilla.sv:2129.4-2132.7" */ _157_[31:0] : 32'hxxxxxxxx;
  assign _142_ = _103_ ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2119.12-2119.36|generated/out/vanilla.sv:2119.8-2135.6" */ 32'hxxxxxxxx : _140_;
  assign _144_ = start ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:2111.12-2111.17|generated/out/vanilla.sv:2111.8-2135.6" */ _159_ : _142_;
  assign _146_ = _147_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:2090.4-2095.11" */ 1'h1 : 1'h0;
  assign _147_ = pcpi_insn[14:12] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:2090.4-2095.11" */ 3'h7;
  assign _148_ = _149_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:2090.4-2095.11" */ 1'h1 : 1'h0;
  assign _149_ = pcpi_insn[14:12] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:2090.4-2095.11" */ 3'h6;
  assign _150_ = _151_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:2090.4-2095.11" */ 1'h1 : 1'h0;
  assign _151_ = pcpi_insn[14:12] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:2090.4-2095.11" */ 3'h5;
  assign _152_ = _153_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:2090.4-2095.11" */ 1'h1 : 1'h0;
  assign _153_ = pcpi_insn[14:12] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:2090.4-2095.11" */ 3'h4;
  assign instr_any_div_rem = | /* src = "generated/out/vanilla.sv:2081.27-2081.74" */ { instr_remu, instr_rem, instr_divu, instr_div };
  assign _154_ = | /* src = "generated/out/vanilla.sv:2115.65-2115.74" */ pcpi_rs2;
  assign _157_ = dividend - /* src = "generated/out/vanilla.sv:2130.17-2130.35" */ divisor;
  assign _159_ = _098_ ? /* src = "generated/out/vanilla.sv:2113.17-2113.80" */ _111_ : pcpi_rs1;
  assign { _161_[62:32], _155_[62:31] } = _099_ ? /* src = "generated/out/vanilla.sv:2114.16-2114.79" */ _113_ : { 31'h00000000, pcpi_rs2 };
  assign _163_ = outsign ? /* src = "generated/out/vanilla.sv:2124.17-2124.47" */ _115_ : quotient;
  assign _165_ = outsign ? /* src = "generated/out/vanilla.sv:2126.17-2126.47" */ _117_ : dividend;
  assign _155_[30:0] = 31'h00000000;
  assign _156_[30:0] = 31'h00000000;
  assign _161_[31:0] = _155_[62:31];
  assign _162_[31:0] = _156_[62:31];
  assign pcpi_ready_t0 = 1'h0;
  assign pcpi_wait_t0 = 1'h0;
  assign pcpi_wr = pcpi_ready;
  assign pcpi_wr_t0 = 1'h0;
endmodule

/* cellift =  1  */
/* hdlname = "\\picorv32_pcpi_mul" */
/* src = "generated/out/vanilla.sv:1837.1-1963.10" */
module picorv32_pcpi_mul(clk, resetn, pcpi_valid, pcpi_insn, pcpi_rs1, pcpi_rs2, pcpi_wr, pcpi_rd, pcpi_wait, pcpi_ready, pcpi_insn_t0, pcpi_rd_t0, pcpi_ready_t0, pcpi_rs1_t0, pcpi_rs2_t0, pcpi_valid_t0, pcpi_wait_t0, pcpi_wr_t0);
  /* src = "generated/out/vanilla.sv:1954.2-1962.5" */
  wire _000_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _001_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _002_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _003_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _004_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _005_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _006_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _007_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _008_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _009_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _010_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _011_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _012_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _013_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _014_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _015_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _016_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _017_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _018_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _019_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _020_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _021_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _022_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _023_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _024_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _025_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _026_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _027_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _028_;
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _029_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1917.69-1917.119" */
  wire [4:0] _030_;
  wire [4:0] _031_;
  wire [4:0] _032_;
  wire [4:0] _033_;
  wire [4:0] _034_;
  wire [4:0] _035_;
  wire [4:0] _036_;
  wire [4:0] _037_;
  wire [4:0] _038_;
  wire [4:0] _039_;
  wire [4:0] _040_;
  wire [4:0] _041_;
  wire [4:0] _042_;
  wire [4:0] _043_;
  wire [4:0] _044_;
  wire [4:0] _045_;
  wire [4:0] _046_;
  wire [4:0] _047_;
  wire [4:0] _048_;
  wire [4:0] _049_;
  wire [4:0] _050_;
  wire [4:0] _051_;
  wire [4:0] _052_;
  wire [4:0] _053_;
  wire [4:0] _054_;
  wire [4:0] _055_;
  wire [4:0] _056_;
  wire [4:0] _057_;
  wire [4:0] _058_;
  wire [4:0] _059_;
  wire [4:0] _060_;
  wire [4:0] _061_;
  wire [4:0] _062_;
  wire [4:0] _063_;
  wire [4:0] _064_;
  wire [4:0] _065_;
  wire [4:0] _066_;
  wire [4:0] _067_;
  wire [4:0] _068_;
  wire [4:0] _069_;
  wire [4:0] _070_;
  wire [4:0] _071_;
  wire [4:0] _072_;
  wire [4:0] _073_;
  wire [4:0] _074_;
  wire [4:0] _075_;
  wire [4:0] _076_;
  wire [4:0] _077_;
  wire [4:0] _078_;
  wire [4:0] _079_;
  wire [4:0] _080_;
  wire [4:0] _081_;
  wire [4:0] _082_;
  wire [4:0] _083_;
  wire [4:0] _084_;
  wire [4:0] _085_;
  wire [4:0] _086_;
  wire [4:0] _087_;
  wire [4:0] _088_;
  wire [4:0] _089_;
  wire [4:0] _090_;
  wire [4:0] _091_;
  wire [4:0] _092_;
  wire _093_;
  wire _094_;
  wire [63:0] _095_;
  wire [63:0] _096_;
  wire [63:0] _097_;
  wire _098_;
  wire _099_;
  wire [4:0] _100_;
  wire [4:0] _101_;
  wire [4:0] _102_;
  wire [4:0] _103_;
  wire [4:0] _104_;
  wire [4:0] _105_;
  wire [4:0] _106_;
  wire [4:0] _107_;
  wire [4:0] _108_;
  wire [4:0] _109_;
  wire [4:0] _110_;
  wire [4:0] _111_;
  wire [4:0] _112_;
  wire [4:0] _113_;
  wire [4:0] _114_;
  wire [4:0] _115_;
  wire [4:0] _116_;
  wire [4:0] _117_;
  wire [4:0] _118_;
  wire [4:0] _119_;
  wire [4:0] _120_;
  wire [4:0] _121_;
  wire [4:0] _122_;
  wire [4:0] _123_;
  wire [4:0] _124_;
  wire [4:0] _125_;
  wire [4:0] _126_;
  wire [4:0] _127_;
  wire [4:0] _128_;
  wire [4:0] _129_;
  wire [4:0] _130_;
  wire [4:0] _131_;
  wire [4:0] _132_;
  wire [4:0] _133_;
  wire [4:0] _134_;
  wire [4:0] _135_;
  wire [4:0] _136_;
  wire [4:0] _137_;
  wire [4:0] _138_;
  wire [4:0] _139_;
  wire [4:0] _140_;
  wire [4:0] _141_;
  wire [4:0] _142_;
  wire [4:0] _143_;
  wire [4:0] _144_;
  wire [4:0] _145_;
  wire [4:0] _146_;
  wire [4:0] _147_;
  wire [4:0] _148_;
  wire [4:0] _149_;
  wire [4:0] _150_;
  wire [4:0] _151_;
  wire [4:0] _152_;
  wire [4:0] _153_;
  wire [4:0] _154_;
  wire [4:0] _155_;
  wire [4:0] _156_;
  wire [4:0] _157_;
  wire [4:0] _158_;
  wire [4:0] _159_;
  wire [4:0] _160_;
  wire [4:0] _161_;
  wire [31:0] _162_;
  wire [31:0] _163_;
  wire [63:0] _164_;
  wire [63:0] _165_;
  wire _166_;
  wire _167_;
  wire [62:0] _168_;
  wire [62:0] _169_;
  wire [14:0] _170_;
  wire [14:0] _171_;
  wire [63:0] _172_;
  wire [63:0] _173_;
  wire [63:0] _174_;
  wire [63:0] _175_;
  wire [63:0] _176_;
  wire [63:0] _177_;
  wire [4:0] _178_;
  wire [4:0] _179_;
  wire [4:0] _180_;
  wire [4:0] _181_;
  wire [4:0] _182_;
  wire [4:0] _183_;
  wire [4:0] _184_;
  wire [4:0] _185_;
  wire [4:0] _186_;
  wire [4:0] _187_;
  wire [4:0] _188_;
  wire [4:0] _189_;
  wire [4:0] _190_;
  wire [4:0] _191_;
  wire [4:0] _192_;
  wire [4:0] _193_;
  wire [4:0] _194_;
  wire [4:0] _195_;
  wire [4:0] _196_;
  wire [4:0] _197_;
  wire [4:0] _198_;
  wire [4:0] _199_;
  wire [4:0] _200_;
  wire [4:0] _201_;
  wire [4:0] _202_;
  wire [4:0] _203_;
  wire [4:0] _204_;
  wire [4:0] _205_;
  wire [4:0] _206_;
  wire [4:0] _207_;
  wire [4:0] _208_;
  wire [4:0] _209_;
  wire [4:0] _210_;
  wire [4:0] _211_;
  wire [4:0] _212_;
  wire [4:0] _213_;
  wire [4:0] _214_;
  wire [4:0] _215_;
  wire [4:0] _216_;
  wire [4:0] _217_;
  wire [4:0] _218_;
  wire [4:0] _219_;
  wire [4:0] _220_;
  wire [4:0] _221_;
  wire [4:0] _222_;
  wire [4:0] _223_;
  wire [4:0] _224_;
  wire [4:0] _225_;
  wire [4:0] _226_;
  wire [4:0] _227_;
  wire [4:0] _228_;
  wire [4:0] _229_;
  wire [4:0] _230_;
  wire [4:0] _231_;
  wire [4:0] _232_;
  wire [4:0] _233_;
  wire [4:0] _234_;
  wire [4:0] _235_;
  wire [4:0] _236_;
  wire [4:0] _237_;
  wire [4:0] _238_;
  wire [4:0] _239_;
  wire [4:0] _240_;
  wire [4:0] _241_;
  wire [4:0] _242_;
  wire [4:0] _243_;
  wire [4:0] _244_;
  wire [4:0] _245_;
  wire [4:0] _246_;
  wire [4:0] _247_;
  wire [4:0] _248_;
  wire [4:0] _249_;
  wire [4:0] _250_;
  wire [4:0] _251_;
  wire [4:0] _252_;
  wire [4:0] _253_;
  wire [4:0] _254_;
  wire [4:0] _255_;
  wire [4:0] _256_;
  wire [4:0] _257_;
  wire [4:0] _258_;
  wire [4:0] _259_;
  wire [4:0] _260_;
  wire [4:0] _261_;
  wire [4:0] _262_;
  wire [4:0] _263_;
  wire [4:0] _264_;
  wire [4:0] _265_;
  wire [4:0] _266_;
  wire [4:0] _267_;
  wire [4:0] _268_;
  wire [4:0] _269_;
  wire [4:0] _270_;
  wire [31:0] _271_;
  wire [63:0] _272_;
  wire _273_;
  wire [62:0] _274_;
  wire [14:0] _275_;
  wire [4:0] _276_;
  wire [4:0] _277_;
  wire [4:0] _278_;
  wire [4:0] _279_;
  wire [4:0] _280_;
  wire [4:0] _281_;
  wire [4:0] _282_;
  wire [4:0] _283_;
  wire [4:0] _284_;
  wire [4:0] _285_;
  wire [4:0] _286_;
  wire [4:0] _287_;
  wire [4:0] _288_;
  wire [4:0] _289_;
  wire [4:0] _290_;
  wire [4:0] _291_;
  wire [4:0] _292_;
  wire [4:0] _293_;
  wire [4:0] _294_;
  wire [4:0] _295_;
  wire [4:0] _296_;
  wire [4:0] _297_;
  wire [4:0] _298_;
  wire [4:0] _299_;
  wire [4:0] _300_;
  wire [4:0] _301_;
  wire [4:0] _302_;
  wire [4:0] _303_;
  wire [4:0] _304_;
  wire [4:0] _305_;
  wire [4:0] _306_;
  wire [4:0] _307_;
  wire [4:0] _308_;
  wire [4:0] _309_;
  wire [4:0] _310_;
  wire [4:0] _311_;
  wire [4:0] _312_;
  wire [4:0] _313_;
  wire [4:0] _314_;
  wire [4:0] _315_;
  wire [4:0] _316_;
  wire [4:0] _317_;
  wire [4:0] _318_;
  wire [4:0] _319_;
  wire [4:0] _320_;
  wire [4:0] _321_;
  wire [4:0] _322_;
  wire [4:0] _323_;
  wire [4:0] _324_;
  wire [4:0] _325_;
  wire [4:0] _326_;
  wire [4:0] _327_;
  wire [4:0] _328_;
  wire [4:0] _329_;
  wire [4:0] _330_;
  wire [4:0] _331_;
  wire [4:0] _332_;
  wire [4:0] _333_;
  wire [4:0] _334_;
  wire [4:0] _335_;
  wire [4:0] _336_;
  wire [4:0] _337_;
  wire [4:0] _338_;
  wire [4:0] _339_;
  wire [4:0] _340_;
  wire [4:0] _341_;
  wire [4:0] _342_;
  wire [4:0] _343_;
  wire [4:0] _344_;
  wire [4:0] _345_;
  wire [4:0] _346_;
  wire [4:0] _347_;
  wire [4:0] _348_;
  wire [4:0] _349_;
  wire [4:0] _350_;
  wire [4:0] _351_;
  wire [4:0] _352_;
  wire [4:0] _353_;
  wire [4:0] _354_;
  wire [4:0] _355_;
  wire [4:0] _356_;
  wire [4:0] _357_;
  wire [4:0] _358_;
  wire [4:0] _359_;
  wire [4:0] _360_;
  wire [4:0] _361_;
  wire [4:0] _362_;
  wire [4:0] _363_;
  wire [4:0] _364_;
  wire [4:0] _365_;
  wire [4:0] _366_;
  wire [4:0] _367_;
  wire [4:0] _368_;
  /* src = "generated/out/vanilla.sv:1876.35-1876.63" */
  wire _369_;
  /* src = "generated/out/vanilla.sv:1876.70-1876.100" */
  wire _370_;
  /* src = "generated/out/vanilla.sv:1876.9-1876.29" */
  wire _371_;
  /* src = "generated/out/vanilla.sv:1876.8-1876.64" */
  wire _372_;
  /* src = "generated/out/vanilla.sv:1876.7-1876.101" */
  wire _373_;
  /* src = "generated/out/vanilla.sv:1957.7-1957.27" */
  wire _374_;
  /* src = "generated/out/vanilla.sv:1870.32-1870.44" */
  wire _375_;
  /* src = "generated/out/vanilla.sv:1940.19-1940.29" */
  wire _376_;
  wire _377_;
  wire _378_;
  wire [6:0] _379_;
  wire [63:0] _380_;
  /* cellift = 32'd1 */
  wire [63:0] _381_;
  /* unused_bits = "0" */
  wire [63:0] _382_;
  /* cellift = 32'd1 */
  /* unused_bits = "0" */
  wire [63:0] _383_;
  wire [63:0] _384_;
  /* unused_bits = "63" */
  wire [63:0] _385_;
  wire _386_;
  wire _387_;
  wire _388_;
  wire _389_;
  wire _390_;
  wire _391_;
  wire _392_;
  wire _393_;
  /* src = "generated/out/vanilla.sv:1947.19-1947.46" */
  /* unused_bits = "7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _394_;
  /* src = "generated/out/vanilla.sv:1939.20-1939.76" */
  /* unused_bits = "7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
  wire [31:0] _395_;
  /* src = "generated/out/vanilla.sv:1960.16-1960.46" */
  /* unused_bits = "32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63" */
  wire [63:0] _396_;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1960.16-1960.46" */
  /* unused_bits = "32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63" */
  wire [63:0] _397_;
  /* src = "generated/out/vanilla.sv:1851.8-1851.11" */
  input clk;
  wire clk;
  /* src = "generated/out/vanilla.sv:1865.7-1865.20" */
  wire instr_any_mul;
  /* src = "generated/out/vanilla.sv:1866.7-1866.21" */
  wire instr_any_mulh;
  /* src = "generated/out/vanilla.sv:1861.6-1861.15" */
  reg instr_mul;
  /* src = "generated/out/vanilla.sv:1862.6-1862.16" */
  reg instr_mulh;
  /* src = "generated/out/vanilla.sv:1863.6-1863.18" */
  reg instr_mulhsu;
  /* src = "generated/out/vanilla.sv:1864.6-1864.17" */
  reg instr_mulhu;
  /* src = "generated/out/vanilla.sv:1867.7-1867.23" */
  wire instr_rs1_signed;
  /* src = "generated/out/vanilla.sv:1896.12-1896.23" */
  reg [6:0] mul_counter;
  /* src = "generated/out/vanilla.sv:1898.6-1898.16" */
  reg mul_finish;
  /* src = "generated/out/vanilla.sv:1870.7-1870.16" */
  wire mul_start;
  /* src = "generated/out/vanilla.sv:1897.6-1897.17" */
  reg mul_waiting;
  /* src = "generated/out/vanilla.sv:1893.13-1893.20" */
  wire [63:0] next_rd;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1893.13-1893.20" */
  wire [63:0] next_rd_t0;
  /* src = "generated/out/vanilla.sv:1895.13-1895.21" */
  /* unused_bits = "63" */
  wire [63:0] next_rdt;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1895.13-1895.21" */
  /* unused_bits = "63" */
  wire [63:0] next_rdt_t0;
  /* src = "generated/out/vanilla.sv:1854.15-1854.24" */
  input [31:0] pcpi_insn;
  wire [31:0] pcpi_insn;
  /* cellift = 32'd1 */
  input [31:0] pcpi_insn_t0;
  wire [31:0] pcpi_insn_t0;
  /* src = "generated/out/vanilla.sv:1858.20-1858.27" */
  output [31:0] pcpi_rd;
  reg [31:0] pcpi_rd;
  /* cellift = 32'd1 */
  output [31:0] pcpi_rd_t0;
  reg [31:0] pcpi_rd_t0;
  /* src = "generated/out/vanilla.sv:1860.13-1860.23" */
  output pcpi_ready;
  reg pcpi_ready;
  /* cellift = 32'd1 */
  output pcpi_ready_t0;
  wire pcpi_ready_t0;
  /* src = "generated/out/vanilla.sv:1855.15-1855.23" */
  input [31:0] pcpi_rs1;
  wire [31:0] pcpi_rs1;
  /* cellift = 32'd1 */
  input [31:0] pcpi_rs1_t0;
  wire [31:0] pcpi_rs1_t0;
  /* src = "generated/out/vanilla.sv:1856.15-1856.23" */
  input [31:0] pcpi_rs2;
  wire [31:0] pcpi_rs2;
  /* cellift = 32'd1 */
  input [31:0] pcpi_rs2_t0;
  wire [31:0] pcpi_rs2_t0;
  /* src = "generated/out/vanilla.sv:1853.8-1853.18" */
  input pcpi_valid;
  wire pcpi_valid;
  /* cellift = 32'd1 */
  input pcpi_valid_t0;
  wire pcpi_valid_t0;
  /* src = "generated/out/vanilla.sv:1859.13-1859.22" */
  output pcpi_wait;
  reg pcpi_wait;
  /* src = "generated/out/vanilla.sv:1869.6-1869.17" */
  reg pcpi_wait_q;
  /* cellift = 32'd1 */
  output pcpi_wait_t0;
  wire pcpi_wait_t0;
  /* src = "generated/out/vanilla.sv:1857.13-1857.20" */
  output pcpi_wr;
  wire pcpi_wr;
  /* cellift = 32'd1 */
  output pcpi_wr_t0;
  wire pcpi_wr_t0;
  /* src = "generated/out/vanilla.sv:1888.13-1888.15" */
  reg [63:0] rd;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1888.13-1888.15" */
  reg [63:0] rd_t0;
  /* src = "generated/out/vanilla.sv:1889.13-1889.16" */
  wire [63:0] rdx;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1889.13-1889.16" */
  wire [63:0] rdx_t0;
  /* src = "generated/out/vanilla.sv:1852.8-1852.14" */
  input resetn;
  wire resetn;
  /* src = "generated/out/vanilla.sv:1886.13-1886.16" */
  reg [63:0] rs1;
  /* src = "generated/out/vanilla.sv:1887.13-1887.16" */
  reg [63:0] rs2;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1887.13-1887.16" */
  reg [63:0] rs2_t0;
  /* src = "generated/out/vanilla.sv:1892.13-1892.21" */
  wire [63:0] this_rs2;
  /* cellift = 32'd1 */
  /* src = "generated/out/vanilla.sv:1892.13-1892.21" */
  wire [63:0] this_rs2_t0;
  assign { next_rdt[3], next_rd[3:0] } = { 1'h0, rd[3:0] } + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[3:0];
  assign _001_ = rd[7:4] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[4] };
  assign { next_rdt[7], next_rd[7:4] } = _001_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[7:4];
  assign _003_ = rd[11:8] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[8] };
  assign { next_rdt[11], next_rd[11:8] } = _003_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[11:8];
  assign _005_ = rd[15:12] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[12] };
  assign { next_rdt[15], next_rd[15:12] } = _005_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[15:12];
  assign _007_ = rd[19:16] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[16] };
  assign { next_rdt[19], next_rd[19:16] } = _007_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[19:16];
  assign _009_ = rd[23:20] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[20] };
  assign { next_rdt[23], next_rd[23:20] } = _009_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[23:20];
  assign _011_ = rd[27:24] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[24] };
  assign { next_rdt[27], next_rd[27:24] } = _011_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[27:24];
  assign _013_ = rd[31:28] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[28] };
  assign { next_rdt[31], next_rd[31:28] } = _013_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[31:28];
  assign _015_ = rd[35:32] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[32] };
  assign { next_rdt[35], next_rd[35:32] } = _015_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[35:32];
  assign _017_ = rd[39:36] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[36] };
  assign { next_rdt[39], next_rd[39:36] } = _017_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[39:36];
  assign _019_ = rd[43:40] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[40] };
  assign { next_rdt[43], next_rd[43:40] } = _019_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[43:40];
  assign _021_ = rd[47:44] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[44] };
  assign { next_rdt[47], next_rd[47:44] } = _021_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[47:44];
  assign _023_ = rd[51:48] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[48] };
  assign { next_rdt[51], next_rd[51:48] } = _023_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[51:48];
  assign _025_ = rd[55:52] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[52] };
  assign { next_rdt[55], next_rd[55:52] } = _025_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[55:52];
  assign _027_ = rd[59:56] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[56] };
  assign { next_rdt[59], next_rd[59:56] } = _027_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[59:56];
  assign _029_ = rd[63:60] + /* src = "generated/out/vanilla.sv:1917.69-1917.119" */ { 3'h0, rdx[60] };
  assign { next_rdt[63], next_rd[63:60] } = _029_ + /* src = "generated/out/vanilla.sv:1917.68-1917.147" */ this_rs2[63:60];
  assign _031_ = ~ { 1'h0, rd_t0[3:0] };
  assign _032_ = ~ { 1'h0, rd_t0[7:4] };
  assign _033_ = ~ _002_;
  assign _034_ = ~ { 1'h0, rd_t0[11:8] };
  assign _035_ = ~ _004_;
  assign _036_ = ~ { 1'h0, rd_t0[15:12] };
  assign _037_ = ~ _006_;
  assign _038_ = ~ { 1'h0, rd_t0[19:16] };
  assign _039_ = ~ _008_;
  assign _040_ = ~ { 1'h0, rd_t0[23:20] };
  assign _041_ = ~ _010_;
  assign _042_ = ~ { 1'h0, rd_t0[27:24] };
  assign _043_ = ~ _012_;
  assign _044_ = ~ { 1'h0, rd_t0[31:28] };
  assign _045_ = ~ _014_;
  assign _046_ = ~ { 1'h0, rd_t0[35:32] };
  assign _047_ = ~ _016_;
  assign _048_ = ~ { 1'h0, rd_t0[39:36] };
  assign _049_ = ~ _018_;
  assign _050_ = ~ { 1'h0, rd_t0[43:40] };
  assign _051_ = ~ _020_;
  assign _052_ = ~ { 1'h0, rd_t0[47:44] };
  assign _053_ = ~ _022_;
  assign _054_ = ~ { 1'h0, rd_t0[51:48] };
  assign _055_ = ~ _024_;
  assign _056_ = ~ { 1'h0, rd_t0[55:52] };
  assign _057_ = ~ _026_;
  assign _058_ = ~ { 1'h0, rd_t0[59:56] };
  assign _059_ = ~ _028_;
  assign _060_ = ~ { 1'h0, rd_t0[63:60] };
  assign _061_ = ~ _030_;
  assign _062_ = ~ { 1'h0, this_rs2_t0[3:0] };
  assign _063_ = ~ { 4'h0, rdx_t0[4] };
  assign _064_ = ~ { 1'h0, this_rs2_t0[7:4] };
  assign _065_ = ~ { 4'h0, rdx_t0[8] };
  assign _066_ = ~ { 1'h0, this_rs2_t0[11:8] };
  assign _067_ = ~ { 4'h0, rdx_t0[12] };
  assign _068_ = ~ { 1'h0, this_rs2_t0[15:12] };
  assign _069_ = ~ { 4'h0, rdx_t0[16] };
  assign _070_ = ~ { 1'h0, this_rs2_t0[19:16] };
  assign _071_ = ~ { 4'h0, rdx_t0[20] };
  assign _072_ = ~ { 1'h0, this_rs2_t0[23:20] };
  assign _073_ = ~ { 4'h0, rdx_t0[24] };
  assign _074_ = ~ { 1'h0, this_rs2_t0[27:24] };
  assign _075_ = ~ { 4'h0, rdx_t0[28] };
  assign _076_ = ~ { 1'h0, this_rs2_t0[31:28] };
  assign _077_ = ~ { 4'h0, rdx_t0[32] };
  assign _078_ = ~ { 1'h0, this_rs2_t0[35:32] };
  assign _079_ = ~ { 4'h0, rdx_t0[36] };
  assign _080_ = ~ { 1'h0, this_rs2_t0[39:36] };
  assign _081_ = ~ { 4'h0, rdx_t0[40] };
  assign _082_ = ~ { 1'h0, this_rs2_t0[43:40] };
  assign _083_ = ~ { 4'h0, rdx_t0[44] };
  assign _084_ = ~ { 1'h0, this_rs2_t0[47:44] };
  assign _085_ = ~ { 4'h0, rdx_t0[48] };
  assign _086_ = ~ { 1'h0, this_rs2_t0[51:48] };
  assign _087_ = ~ { 4'h0, rdx_t0[52] };
  assign _088_ = ~ { 1'h0, this_rs2_t0[55:52] };
  assign _089_ = ~ { 4'h0, rdx_t0[56] };
  assign _090_ = ~ { 1'h0, this_rs2_t0[59:56] };
  assign _091_ = ~ { 4'h0, rdx_t0[60] };
  assign _092_ = ~ { 1'h0, this_rs2_t0[63:60] };
  assign _100_ = { 1'h0, rd[3:0] } & _031_;
  assign _102_ = { 1'h0, rd[7:4] } & _032_;
  assign _104_ = _001_ & _033_;
  assign _106_ = { 1'h0, rd[11:8] } & _034_;
  assign _108_ = _003_ & _035_;
  assign _110_ = { 1'h0, rd[15:12] } & _036_;
  assign _112_ = _005_ & _037_;
  assign _114_ = { 1'h0, rd[19:16] } & _038_;
  assign _116_ = _007_ & _039_;
  assign _118_ = { 1'h0, rd[23:20] } & _040_;
  assign _120_ = _009_ & _041_;
  assign _122_ = { 1'h0, rd[27:24] } & _042_;
  assign _124_ = _011_ & _043_;
  assign _126_ = { 1'h0, rd[31:28] } & _044_;
  assign _128_ = _013_ & _045_;
  assign _130_ = { 1'h0, rd[35:32] } & _046_;
  assign _132_ = _015_ & _047_;
  assign _134_ = { 1'h0, rd[39:36] } & _048_;
  assign _136_ = _017_ & _049_;
  assign _138_ = { 1'h0, rd[43:40] } & _050_;
  assign _140_ = _019_ & _051_;
  assign _142_ = { 1'h0, rd[47:44] } & _052_;
  assign _144_ = _021_ & _053_;
  assign _146_ = { 1'h0, rd[51:48] } & _054_;
  assign _148_ = _023_ & _055_;
  assign _150_ = { 1'h0, rd[55:52] } & _056_;
  assign _152_ = _025_ & _057_;
  assign _154_ = { 1'h0, rd[59:56] } & _058_;
  assign _156_ = _027_ & _059_;
  assign _158_ = { 1'h0, rd[63:60] } & _060_;
  assign _160_ = _029_ & _061_;
  assign _101_ = { 1'h0, this_rs2[3:0] } & _062_;
  assign _103_ = { 4'h0, rdx[4] } & _063_;
  assign _105_ = { 1'h0, this_rs2[7:4] } & _064_;
  assign _107_ = { 4'h0, rdx[8] } & _065_;
  assign _109_ = { 1'h0, this_rs2[11:8] } & _066_;
  assign _111_ = { 4'h0, rdx[12] } & _067_;
  assign _113_ = { 1'h0, this_rs2[15:12] } & _068_;
  assign _115_ = { 4'h0, rdx[16] } & _069_;
  assign _117_ = { 1'h0, this_rs2[19:16] } & _070_;
  assign _119_ = { 4'h0, rdx[20] } & _071_;
  assign _121_ = { 1'h0, this_rs2[23:20] } & _072_;
  assign _123_ = { 4'h0, rdx[24] } & _073_;
  assign _125_ = { 1'h0, this_rs2[27:24] } & _074_;
  assign _127_ = { 4'h0, rdx[28] } & _075_;
  assign _129_ = { 1'h0, this_rs2[31:28] } & _076_;
  assign _131_ = { 4'h0, rdx[32] } & _077_;
  assign _133_ = { 1'h0, this_rs2[35:32] } & _078_;
  assign _135_ = { 4'h0, rdx[36] } & _079_;
  assign _137_ = { 1'h0, this_rs2[39:36] } & _080_;
  assign _139_ = { 4'h0, rdx[40] } & _081_;
  assign _141_ = { 1'h0, this_rs2[43:40] } & _082_;
  assign _143_ = { 4'h0, rdx[44] } & _083_;
  assign _145_ = { 1'h0, this_rs2[47:44] } & _084_;
  assign _147_ = { 4'h0, rdx[48] } & _085_;
  assign _149_ = { 1'h0, this_rs2[51:48] } & _086_;
  assign _151_ = { 4'h0, rdx[52] } & _087_;
  assign _153_ = { 1'h0, this_rs2[55:52] } & _088_;
  assign _155_ = { 4'h0, rdx[56] } & _089_;
  assign _157_ = { 1'h0, this_rs2[59:56] } & _090_;
  assign _159_ = { 4'h0, rdx[60] } & _091_;
  assign _161_ = { 1'h0, this_rs2[63:60] } & _092_;
  assign _307_ = _100_ + _101_;
  assign _309_ = _102_ + _103_;
  assign _311_ = _104_ + _105_;
  assign _313_ = _106_ + _107_;
  assign _315_ = _108_ + _109_;
  assign _317_ = _110_ + _111_;
  assign _319_ = _112_ + _113_;
  assign _321_ = _114_ + _115_;
  assign _323_ = _116_ + _117_;
  assign _325_ = _118_ + _119_;
  assign _327_ = _120_ + _121_;
  assign _329_ = _122_ + _123_;
  assign _331_ = _124_ + _125_;
  assign _333_ = _126_ + _127_;
  assign _335_ = _128_ + _129_;
  assign _337_ = _130_ + _131_;
  assign _339_ = _132_ + _133_;
  assign _341_ = _134_ + _135_;
  assign _343_ = _136_ + _137_;
  assign _345_ = _138_ + _139_;
  assign _347_ = _140_ + _141_;
  assign _349_ = _142_ + _143_;
  assign _351_ = _144_ + _145_;
  assign _353_ = _146_ + _147_;
  assign _355_ = _148_ + _149_;
  assign _357_ = _150_ + _151_;
  assign _359_ = _152_ + _153_;
  assign _361_ = _154_ + _155_;
  assign _363_ = _156_ + _157_;
  assign _365_ = _158_ + _159_;
  assign _367_ = _160_ + _161_;
  assign _178_ = { 1'h0, rd[3:0] } | { 1'h0, rd_t0[3:0] };
  assign _181_ = { 1'h0, rd[7:4] } | { 1'h0, rd_t0[7:4] };
  assign _184_ = _001_ | _002_;
  assign _187_ = { 1'h0, rd[11:8] } | { 1'h0, rd_t0[11:8] };
  assign _190_ = _003_ | _004_;
  assign _193_ = { 1'h0, rd[15:12] } | { 1'h0, rd_t0[15:12] };
  assign _196_ = _005_ | _006_;
  assign _199_ = { 1'h0, rd[19:16] } | { 1'h0, rd_t0[19:16] };
  assign _202_ = _007_ | _008_;
  assign _205_ = { 1'h0, rd[23:20] } | { 1'h0, rd_t0[23:20] };
  assign _208_ = _009_ | _010_;
  assign _211_ = { 1'h0, rd[27:24] } | { 1'h0, rd_t0[27:24] };
  assign _214_ = _011_ | _012_;
  assign _217_ = { 1'h0, rd[31:28] } | { 1'h0, rd_t0[31:28] };
  assign _220_ = _013_ | _014_;
  assign _223_ = { 1'h0, rd[35:32] } | { 1'h0, rd_t0[35:32] };
  assign _226_ = _015_ | _016_;
  assign _229_ = { 1'h0, rd[39:36] } | { 1'h0, rd_t0[39:36] };
  assign _232_ = _017_ | _018_;
  assign _235_ = { 1'h0, rd[43:40] } | { 1'h0, rd_t0[43:40] };
  assign _238_ = _019_ | _020_;
  assign _241_ = { 1'h0, rd[47:44] } | { 1'h0, rd_t0[47:44] };
  assign _244_ = _021_ | _022_;
  assign _247_ = { 1'h0, rd[51:48] } | { 1'h0, rd_t0[51:48] };
  assign _250_ = _023_ | _024_;
  assign _253_ = { 1'h0, rd[55:52] } | { 1'h0, rd_t0[55:52] };
  assign _256_ = _025_ | _026_;
  assign _259_ = { 1'h0, rd[59:56] } | { 1'h0, rd_t0[59:56] };
  assign _262_ = _027_ | _028_;
  assign _265_ = { 1'h0, rd[63:60] } | { 1'h0, rd_t0[63:60] };
  assign _268_ = _029_ | _030_;
  assign _179_ = { 1'h0, this_rs2[3:0] } | { 1'h0, this_rs2_t0[3:0] };
  assign _182_ = { 4'h0, rdx[4] } | { 4'h0, rdx_t0[4] };
  assign _185_ = { 1'h0, this_rs2[7:4] } | { 1'h0, this_rs2_t0[7:4] };
  assign _188_ = { 4'h0, rdx[8] } | { 4'h0, rdx_t0[8] };
  assign _191_ = { 1'h0, this_rs2[11:8] } | { 1'h0, this_rs2_t0[11:8] };
  assign _194_ = { 4'h0, rdx[12] } | { 4'h0, rdx_t0[12] };
  assign _197_ = { 1'h0, this_rs2[15:12] } | { 1'h0, this_rs2_t0[15:12] };
  assign _200_ = { 4'h0, rdx[16] } | { 4'h0, rdx_t0[16] };
  assign _203_ = { 1'h0, this_rs2[19:16] } | { 1'h0, this_rs2_t0[19:16] };
  assign _206_ = { 4'h0, rdx[20] } | { 4'h0, rdx_t0[20] };
  assign _209_ = { 1'h0, this_rs2[23:20] } | { 1'h0, this_rs2_t0[23:20] };
  assign _212_ = { 4'h0, rdx[24] } | { 4'h0, rdx_t0[24] };
  assign _215_ = { 1'h0, this_rs2[27:24] } | { 1'h0, this_rs2_t0[27:24] };
  assign _218_ = { 4'h0, rdx[28] } | { 4'h0, rdx_t0[28] };
  assign _221_ = { 1'h0, this_rs2[31:28] } | { 1'h0, this_rs2_t0[31:28] };
  assign _224_ = { 4'h0, rdx[32] } | { 4'h0, rdx_t0[32] };
  assign _227_ = { 1'h0, this_rs2[35:32] } | { 1'h0, this_rs2_t0[35:32] };
  assign _230_ = { 4'h0, rdx[36] } | { 4'h0, rdx_t0[36] };
  assign _233_ = { 1'h0, this_rs2[39:36] } | { 1'h0, this_rs2_t0[39:36] };
  assign _236_ = { 4'h0, rdx[40] } | { 4'h0, rdx_t0[40] };
  assign _239_ = { 1'h0, this_rs2[43:40] } | { 1'h0, this_rs2_t0[43:40] };
  assign _242_ = { 4'h0, rdx[44] } | { 4'h0, rdx_t0[44] };
  assign _245_ = { 1'h0, this_rs2[47:44] } | { 1'h0, this_rs2_t0[47:44] };
  assign _248_ = { 4'h0, rdx[48] } | { 4'h0, rdx_t0[48] };
  assign _251_ = { 1'h0, this_rs2[51:48] } | { 1'h0, this_rs2_t0[51:48] };
  assign _254_ = { 4'h0, rdx[52] } | { 4'h0, rdx_t0[52] };
  assign _257_ = { 1'h0, this_rs2[55:52] } | { 1'h0, this_rs2_t0[55:52] };
  assign _260_ = { 4'h0, rdx[56] } | { 4'h0, rdx_t0[56] };
  assign _263_ = { 1'h0, this_rs2[59:56] } | { 1'h0, this_rs2_t0[59:56] };
  assign _266_ = { 4'h0, rdx[60] } | { 4'h0, rdx_t0[60] };
  assign _269_ = { 1'h0, this_rs2[63:60] } | { 1'h0, this_rs2_t0[63:60] };
  assign _308_ = _178_ + _179_;
  assign _310_ = _181_ + _182_;
  assign _312_ = _184_ + _185_;
  assign _314_ = _187_ + _188_;
  assign _316_ = _190_ + _191_;
  assign _318_ = _193_ + _194_;
  assign _320_ = _196_ + _197_;
  assign _322_ = _199_ + _200_;
  assign _324_ = _202_ + _203_;
  assign _326_ = _205_ + _206_;
  assign _328_ = _208_ + _209_;
  assign _330_ = _211_ + _212_;
  assign _332_ = _214_ + _215_;
  assign _334_ = _217_ + _218_;
  assign _336_ = _220_ + _221_;
  assign _338_ = _223_ + _224_;
  assign _340_ = _226_ + _227_;
  assign _342_ = _229_ + _230_;
  assign _344_ = _232_ + _233_;
  assign _346_ = _235_ + _236_;
  assign _348_ = _238_ + _239_;
  assign _350_ = _241_ + _242_;
  assign _352_ = _244_ + _245_;
  assign _354_ = _247_ + _248_;
  assign _356_ = _250_ + _251_;
  assign _358_ = _253_ + _254_;
  assign _360_ = _256_ + _257_;
  assign _362_ = _259_ + _260_;
  assign _364_ = _262_ + _263_;
  assign _366_ = _265_ + _266_;
  assign _368_ = _268_ + _269_;
  assign _276_ = _307_ ^ _308_;
  assign _277_ = _309_ ^ _310_;
  assign _278_ = _311_ ^ _312_;
  assign _279_ = _313_ ^ _314_;
  assign _280_ = _315_ ^ _316_;
  assign _281_ = _317_ ^ _318_;
  assign _282_ = _319_ ^ _320_;
  assign _283_ = _321_ ^ _322_;
  assign _284_ = _323_ ^ _324_;
  assign _285_ = _325_ ^ _326_;
  assign _286_ = _327_ ^ _328_;
  assign _287_ = _329_ ^ _330_;
  assign _288_ = _331_ ^ _332_;
  assign _289_ = _333_ ^ _334_;
  assign _290_ = _335_ ^ _336_;
  assign _291_ = _337_ ^ _338_;
  assign _292_ = _339_ ^ _340_;
  assign _293_ = _341_ ^ _342_;
  assign _294_ = _343_ ^ _344_;
  assign _295_ = _345_ ^ _346_;
  assign _296_ = _347_ ^ _348_;
  assign _297_ = _349_ ^ _350_;
  assign _298_ = _351_ ^ _352_;
  assign _299_ = _353_ ^ _354_;
  assign _300_ = _355_ ^ _356_;
  assign _301_ = _357_ ^ _358_;
  assign _302_ = _359_ ^ _360_;
  assign _303_ = _361_ ^ _362_;
  assign _304_ = _363_ ^ _364_;
  assign _305_ = _365_ ^ _366_;
  assign _306_ = _367_ ^ _368_;
  assign _180_ = _276_ | { 1'h0, rd_t0[3:0] };
  assign _183_ = _277_ | { 1'h0, rd_t0[7:4] };
  assign _186_ = _278_ | _002_;
  assign _189_ = _279_ | { 1'h0, rd_t0[11:8] };
  assign _192_ = _280_ | _004_;
  assign _195_ = _281_ | { 1'h0, rd_t0[15:12] };
  assign _198_ = _282_ | _006_;
  assign _201_ = _283_ | { 1'h0, rd_t0[19:16] };
  assign _204_ = _284_ | _008_;
  assign _207_ = _285_ | { 1'h0, rd_t0[23:20] };
  assign _210_ = _286_ | _010_;
  assign _213_ = _287_ | { 1'h0, rd_t0[27:24] };
  assign _216_ = _288_ | _012_;
  assign _219_ = _289_ | { 1'h0, rd_t0[31:28] };
  assign _222_ = _290_ | _014_;
  assign _225_ = _291_ | { 1'h0, rd_t0[35:32] };
  assign _228_ = _292_ | _016_;
  assign _231_ = _293_ | { 1'h0, rd_t0[39:36] };
  assign _234_ = _294_ | _018_;
  assign _237_ = _295_ | { 1'h0, rd_t0[43:40] };
  assign _240_ = _296_ | _020_;
  assign _243_ = _297_ | { 1'h0, rd_t0[47:44] };
  assign _246_ = _298_ | _022_;
  assign _249_ = _299_ | { 1'h0, rd_t0[51:48] };
  assign _252_ = _300_ | _024_;
  assign _255_ = _301_ | { 1'h0, rd_t0[55:52] };
  assign _258_ = _302_ | _026_;
  assign _261_ = _303_ | { 1'h0, rd_t0[59:56] };
  assign _264_ = _304_ | _028_;
  assign _267_ = _305_ | { 1'h0, rd_t0[63:60] };
  assign _270_ = _306_ | _030_;
  assign { next_rdt_t0[3], next_rd_t0[3:0] } = _180_ | { 1'h0, this_rs2_t0[3:0] };
  assign _002_ = _183_ | { 4'h0, rdx_t0[4] };
  assign { next_rdt_t0[7], next_rd_t0[7:4] } = _186_ | { 1'h0, this_rs2_t0[7:4] };
  assign _004_ = _189_ | { 4'h0, rdx_t0[8] };
  assign { next_rdt_t0[11], next_rd_t0[11:8] } = _192_ | { 1'h0, this_rs2_t0[11:8] };
  assign _006_ = _195_ | { 4'h0, rdx_t0[12] };
  assign { next_rdt_t0[15], next_rd_t0[15:12] } = _198_ | { 1'h0, this_rs2_t0[15:12] };
  assign _008_ = _201_ | { 4'h0, rdx_t0[16] };
  assign { next_rdt_t0[19], next_rd_t0[19:16] } = _204_ | { 1'h0, this_rs2_t0[19:16] };
  assign _010_ = _207_ | { 4'h0, rdx_t0[20] };
  assign { next_rdt_t0[23], next_rd_t0[23:20] } = _210_ | { 1'h0, this_rs2_t0[23:20] };
  assign _012_ = _213_ | { 4'h0, rdx_t0[24] };
  assign { next_rdt_t0[27], next_rd_t0[27:24] } = _216_ | { 1'h0, this_rs2_t0[27:24] };
  assign _014_ = _219_ | { 4'h0, rdx_t0[28] };
  assign { next_rdt_t0[31], next_rd_t0[31:28] } = _222_ | { 1'h0, this_rs2_t0[31:28] };
  assign _016_ = _225_ | { 4'h0, rdx_t0[32] };
  assign { next_rdt_t0[35], next_rd_t0[35:32] } = _228_ | { 1'h0, this_rs2_t0[35:32] };
  assign _018_ = _231_ | { 4'h0, rdx_t0[36] };
  assign { next_rdt_t0[39], next_rd_t0[39:36] } = _234_ | { 1'h0, this_rs2_t0[39:36] };
  assign _020_ = _237_ | { 4'h0, rdx_t0[40] };
  assign { next_rdt_t0[43], next_rd_t0[43:40] } = _240_ | { 1'h0, this_rs2_t0[43:40] };
  assign _022_ = _243_ | { 4'h0, rdx_t0[44] };
  assign { next_rdt_t0[47], next_rd_t0[47:44] } = _246_ | { 1'h0, this_rs2_t0[47:44] };
  assign _024_ = _249_ | { 4'h0, rdx_t0[48] };
  assign { next_rdt_t0[51], next_rd_t0[51:48] } = _252_ | { 1'h0, this_rs2_t0[51:48] };
  assign _026_ = _255_ | { 4'h0, rdx_t0[52] };
  assign { next_rdt_t0[55], next_rd_t0[55:52] } = _258_ | { 1'h0, this_rs2_t0[55:52] };
  assign _028_ = _261_ | { 4'h0, rdx_t0[56] };
  assign { next_rdt_t0[59], next_rd_t0[59:56] } = _264_ | { 1'h0, this_rs2_t0[59:56] };
  assign _030_ = _267_ | { 4'h0, rdx_t0[60] };
  assign { next_rdt_t0[63], next_rd_t0[63:60] } = _270_ | { 1'h0, this_rs2_t0[63:60] };
  assign _093_ = ~ resetn;
  assign _094_ = ~ _374_;
  assign _162_ = { _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_, _374_ } & _397_[31:0];
  assign _168_ = { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn } & _383_[63:1];
  assign _163_ = { _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_, _094_ } & pcpi_rd_t0;
  assign _169_ = { _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_ } & rs2_t0[63:1];
  assign _271_ = _162_ | _163_;
  assign _274_ = _168_ | _169_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME pcpi_rd_t0 */
  always_ff @(posedge clk)
    pcpi_rd_t0 <= _271_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rs2_t0[63:1] */
  always_ff @(posedge clk)
    rs2_t0[63:1] <= _274_;
  /* src = "generated/out/vanilla.sv:1871.2-1885.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME instr_mulhu */
  always_ff @(posedge clk)
    if (!_373_) instr_mulhu <= 1'h0;
    else instr_mulhu <= _386_;
  /* src = "generated/out/vanilla.sv:1871.2-1885.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME instr_mulhsu */
  always_ff @(posedge clk)
    if (!_373_) instr_mulhsu <= 1'h0;
    else instr_mulhsu <= _388_;
  /* src = "generated/out/vanilla.sv:1871.2-1885.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME instr_mulh */
  always_ff @(posedge clk)
    if (!_373_) instr_mulh <= 1'h0;
    else instr_mulh <= _390_;
  /* src = "generated/out/vanilla.sv:1871.2-1885.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME instr_mul */
  always_ff @(posedge clk)
    if (!_373_) instr_mul <= 1'h0;
    else instr_mul <= _392_;
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME mul_waiting */
  always_ff @(posedge clk)
    if (!resetn) mul_waiting <= 1'h1;
    else mul_waiting <= _378_;
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME mul_finish */
  always_ff @(posedge clk)
    if (_098_) mul_finish <= 1'h0;
    else mul_finish <= _377_;
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME mul_counter */
  always_ff @(posedge clk)
    if (resetn) mul_counter <= _379_;
  /* src = "generated/out/vanilla.sv:1954.2-1962.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME pcpi_rd */
  always_ff @(posedge clk)
    if (_374_) pcpi_rd <= _396_[31:0];
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rd */
  always_ff @(posedge clk)
    if (resetn)
      if (mul_waiting) rd <= 64'h0000000000000000;
      else rd <= next_rd;
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rs2[0] */
  always_ff @(posedge clk)
    if (resetn)
      if (!mul_waiting) rs2[0] <= 1'h0;
      else rs2[0] <= _380_[0];
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rs2[63:1] */
  always_ff @(posedge clk)
    if (resetn) rs2[63:1] <= _382_[63:1];
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rs1[63] */
  always_ff @(posedge clk)
    if (resetn)
      if (!_099_) rs1[63] <= 1'h0;
      else rs1[63] <= pcpi_rs1[31];
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rs1[62:0] */
  always_ff @(posedge clk)
    if (resetn) rs1[62:0] <= _385_[62:0];
  reg [14:0] _793_;
  /* src = "generated/out/vanilla.sv:1924.2-1953.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME _793_ */
  always_ff @(posedge clk)
    if (resetn)
      if (mul_waiting) _793_ <= 15'h0000;
      else _793_ <= { next_rdt[59], next_rdt[55], next_rdt[51], next_rdt[47], next_rdt[43], next_rdt[39], next_rdt[35], next_rdt[31], next_rdt[27], next_rdt[23], next_rdt[19], next_rdt[15], next_rdt[11], next_rdt[7], next_rdt[3] };
  assign { rdx[60], rdx[56], rdx[52], rdx[48], rdx[44], rdx[40], rdx[36], rdx[32], rdx[28], rdx[24], rdx[20], rdx[16], rdx[12], rdx[8], rdx[4] } = _793_;
  assign _095_ = ~ { instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh };
  assign _096_ = ~ { mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting };
  assign _097_ = ~ { instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh };
  assign _172_ = _095_ & { 32'h00000000, pcpi_rs2_t0 };
  assign _174_ = _096_ & { rs2_t0[62:0], 1'h0 };
  assign _176_ = _097_ & rd_t0;
  assign _173_ = { instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh, instr_mulh } & { pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0[31], pcpi_rs2_t0 };
  assign _175_ = { mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting, mul_waiting } & _381_;
  assign this_rs2_t0 = { rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0], rs1[0] } & rs2_t0;
  assign _177_ = { instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh, instr_any_mulh } & { 32'h00000000, rd_t0[63:32] };
  assign _381_ = _172_ | _173_;
  assign _383_ = _174_ | _175_;
  assign _397_ = _176_ | _177_;
  assign _098_ = | { _093_, mul_waiting };
  assign _099_ = & { mul_waiting, instr_rs1_signed };
  assign _164_ = { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn } & next_rd_t0;
  assign _166_ = resetn & _381_[0];
  assign _170_ = { resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn, resetn } & { next_rdt_t0[59], next_rdt_t0[55], next_rdt_t0[51], next_rdt_t0[47], next_rdt_t0[43], next_rdt_t0[39], next_rdt_t0[35], next_rdt_t0[31], next_rdt_t0[27], next_rdt_t0[23], next_rdt_t0[19], next_rdt_t0[15], next_rdt_t0[11], next_rdt_t0[7], next_rdt_t0[3] };
  assign _165_ = { _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_ } & rd_t0;
  assign _167_ = _093_ & rs2_t0[0];
  assign _171_ = { _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_ } & { rdx_t0[60], rdx_t0[56], rdx_t0[52], rdx_t0[48], rdx_t0[44], rdx_t0[40], rdx_t0[36], rdx_t0[32], rdx_t0[28], rdx_t0[24], rdx_t0[20], rdx_t0[16], rdx_t0[12], rdx_t0[8], rdx_t0[4] };
  assign _272_ = _164_ | _165_;
  assign _273_ = _166_ | _167_;
  assign _275_ = _170_ | _171_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rd_t0 */
  always_ff @(posedge clk)
    if (mul_waiting) rd_t0 <= 64'h0000000000000000;
    else rd_t0 <= _272_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME rs2_t0[0] */
  always_ff @(posedge clk)
    if (!mul_waiting) rs2_t0[0] <= 1'h0;
    else rs2_t0[0] <= _273_;
  reg [14:0] _820_;
  /* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME _820_ */
  always_ff @(posedge clk)
    if (mul_waiting) _820_ <= 15'h0000;
    else _820_ <= _275_;
  assign { rdx_t0[60], rdx_t0[56], rdx_t0[52], rdx_t0[48], rdx_t0[44], rdx_t0[40], rdx_t0[36], rdx_t0[32], rdx_t0[28], rdx_t0[24], rdx_t0[20], rdx_t0[16], rdx_t0[12], rdx_t0[8], rdx_t0[4] } = _820_;
  assign _369_ = pcpi_insn[6:0] == /* src = "generated/out/vanilla.sv:1876.35-1876.63" */ 7'h33;
  assign _370_ = pcpi_insn[31:25] == /* src = "generated/out/vanilla.sv:1876.70-1876.100" */ 7'h01;
  assign mul_start = pcpi_wait && /* src = "generated/out/vanilla.sv:1870.19-1870.44" */ _375_;
  assign _371_ = resetn && /* src = "generated/out/vanilla.sv:1876.9-1876.29" */ pcpi_valid;
  assign _372_ = _371_ && /* src = "generated/out/vanilla.sv:1876.8-1876.64" */ _369_;
  assign _373_ = _372_ && /* src = "generated/out/vanilla.sv:1876.7-1876.101" */ _370_;
  assign _374_ = mul_finish && /* src = "generated/out/vanilla.sv:1957.7-1957.27" */ resetn;
  assign _375_ = ! /* src = "generated/out/vanilla.sv:1870.32-1870.44" */ pcpi_wait_q;
  assign _376_ = ! /* src = "generated/out/vanilla.sv:1940.19-1940.29" */ mul_start;
  /* src = "generated/out/vanilla.sv:1954.2-1962.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME pcpi_ready */
  always_ff @(posedge clk)
    pcpi_ready <= _000_;
  /* src = "generated/out/vanilla.sv:1871.2-1885.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME pcpi_wait */
  always_ff @(posedge clk)
    pcpi_wait <= instr_any_mul;
  /* src = "generated/out/vanilla.sv:1871.2-1885.5" */
/* PC_TAINT_INFO MODULE_NAME picorv32_pcpi_mul */
/* PC_TAINT_INFO STATE_NAME pcpi_wait_q */
  always_ff @(posedge clk)
    pcpi_wait_q <= pcpi_wait;
  assign _000_ = _374_ ? /* src = "generated/out/vanilla.sv:1957.7-1957.27|generated/out/vanilla.sv:1957.3-1961.6" */ 1'h1 : 1'h0;
  assign _377_ = mul_counter[6] ? /* src = "generated/out/vanilla.sv:1948.8-1948.22|generated/out/vanilla.sv:1948.4-1951.7" */ 1'h1 : 1'h0;
  assign _378_ = mul_waiting ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1928.12-1928.23|generated/out/vanilla.sv:1928.8-1952.6" */ _376_ : _377_;
  assign _379_ = mul_waiting ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1928.12-1928.23|generated/out/vanilla.sv:1928.8-1952.6" */ _395_[6:0] : _394_[6:0];
  assign _380_ = instr_mulh ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1933.8-1933.24|generated/out/vanilla.sv:1933.4-1936.32" */ { pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2[31], pcpi_rs2 } : { 32'h00000000, pcpi_rs2 };
  assign _382_ = mul_waiting ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1928.12-1928.23|generated/out/vanilla.sv:1928.8-1952.6" */ _380_ : { rs2[62:0], 1'h0 };
  assign _384_ = instr_rs1_signed ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1929.8-1929.24|generated/out/vanilla.sv:1929.4-1932.32" */ { pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1[31], pcpi_rs1 } : { 32'h00000000, pcpi_rs1 };
  assign _385_ = mul_waiting ? /* full_case = 32'd1 */ /* src = "generated/out/vanilla.sv:1928.12-1928.23|generated/out/vanilla.sv:1928.8-1952.6" */ _384_ : { 1'h0, rs1[63:1] };
  assign _386_ = _387_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1877.4-1882.11" */ 1'h1 : 1'h0;
  assign _387_ = pcpi_insn[14:12] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1877.4-1882.11" */ 3'h3;
  assign _388_ = _389_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1877.4-1882.11" */ 1'h1 : 1'h0;
  assign _389_ = pcpi_insn[14:12] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1877.4-1882.11" */ 3'h2;
  assign _390_ = _391_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1877.4-1882.11" */ 1'h1 : 1'h0;
  assign _391_ = pcpi_insn[14:12] == /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1877.4-1882.11" */ 3'h1;
  assign _392_ = _393_ ? /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1877.4-1882.11" */ 1'h1 : 1'h0;
  assign _393_ = ! /* src = "generated/out/vanilla.sv:0.0-0.0|generated/out/vanilla.sv:1877.4-1882.11" */ pcpi_insn[14:12];
  assign instr_any_mul = | /* src = "generated/out/vanilla.sv:1865.23-1865.74" */ { instr_mulhu, instr_mulhsu, instr_mulh, instr_mul };
  assign instr_any_mulh = | /* src = "generated/out/vanilla.sv:1866.24-1866.64" */ { instr_mulhu, instr_mulhsu, instr_mulh };
  assign instr_rs1_signed = | /* src = "generated/out/vanilla.sv:1867.26-1867.53" */ { instr_mulhsu, instr_mulh };
  assign _394_ = mul_counter - /* src = "generated/out/vanilla.sv:1947.19-1947.46" */ 32'd1;
  assign this_rs2 = rs1[0] ? /* src = "generated/out/vanilla.sv:1908.17-1908.43" */ rs2 : 64'h0000000000000000;
  assign _395_ = instr_any_mulh ? /* src = "generated/out/vanilla.sv:1939.20-1939.76" */ 32'd62 : 32'd30;
  assign _396_ = instr_any_mulh ? /* src = "generated/out/vanilla.sv:1960.16-1960.46" */ { 32'h00000000, rd[63:32] } : rd;
  assign { next_rdt[62:60], next_rdt[58:56], next_rdt[54:52], next_rdt[50:48], next_rdt[46:44], next_rdt[42:40], next_rdt[38:36], next_rdt[34:32], next_rdt[30:28], next_rdt[26:24], next_rdt[22:20], next_rdt[18:16], next_rdt[14:12], next_rdt[10:8], next_rdt[6:4], next_rdt[2:0] } = 48'h000000000000;
  assign { next_rdt_t0[62:60], next_rdt_t0[58:56], next_rdt_t0[54:52], next_rdt_t0[50:48], next_rdt_t0[46:44], next_rdt_t0[42:40], next_rdt_t0[38:36], next_rdt_t0[34:32], next_rdt_t0[30:28], next_rdt_t0[26:24], next_rdt_t0[22:20], next_rdt_t0[18:16], next_rdt_t0[14:12], next_rdt_t0[10:8], next_rdt_t0[6:4], next_rdt_t0[2:0] } = 48'h000000000000;
  assign pcpi_ready_t0 = 1'h0;
  assign pcpi_wait_t0 = 1'h0;
  assign pcpi_wr = pcpi_ready;
  assign pcpi_wr_t0 = 1'h0;
  assign { rdx[63:61], rdx[59:57], rdx[55:53], rdx[51:49], rdx[47:45], rdx[43:41], rdx[39:37], rdx[35:33], rdx[31:29], rdx[27:25], rdx[23:21], rdx[19:17], rdx[15:13], rdx[11:9], rdx[7:5], rdx[3:0] } = 49'h0000000000000;
  assign { rdx_t0[63:61], rdx_t0[59:57], rdx_t0[55:53], rdx_t0[51:49], rdx_t0[47:45], rdx_t0[43:41], rdx_t0[39:37], rdx_t0[35:33], rdx_t0[31:29], rdx_t0[27:25], rdx_t0[23:21], rdx_t0[19:17], rdx_t0[15:13], rdx_t0[11:9], rdx_t0[7:5], rdx_t0[3:0] } = 49'h0000000000000;
endmodule
