  asm_declass_cpuregs_wrdata: assume property (!cpuregs_wrdata_t0);