bit gen_instr_word_sampling_cond;
assign gen_instr_word_sampling_cond = (mem_do_rinst &&  mem_done);