bit gen_regrd_rs2;
assign gen_regrd_rs2 = 
 ((|  decoded_rs2));
;