bit gen_regrd_rs1;
assign gen_regrd_rs1 = 
 ((|  decoded_rs1));
;