asm_declass_rf_wdata_fwd_wb: assume property (!u_ibex_core__rf_wdata_fwd_wb_t0);
asm_declass_rf_wdata_wb: assume property (!u_ibex_core__rf_wdata_wb_ecc_o_t0);