asm_declass_u_ex__regwr_data_t0: assume property(!u_ex__regwr_data_t0);
