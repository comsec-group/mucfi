bind frv_core frv_core_fpv frv_core_fpv_bind (
.g_clk(
  g_clk),
.g_resetn(
  g_resetn),
.trs_pc(
  trs_pc),
.trs_instr(
  trs_instr),
.trs_valid(
  trs_valid),
.leak_prng(
  leak_prng),
.leak_fence_unc0(
  leak_fence_unc0),
.leak_fence_unc1(
  leak_fence_unc1),
.leak_fence_unc2(
  leak_fence_unc2),
.rng_req_valid(
  rng_req_valid),
.rng_req_op(
  rng_req_op),
.rng_req_data(
  rng_req_data),
.rng_req_ready(
  rng_req_ready),
.rng_rsp_valid(
  rng_rsp_valid),
.rng_rsp_status(
  rng_rsp_status),
.rng_rsp_data(
  rng_rsp_data),
.rng_rsp_ready(
  rng_rsp_ready),
.int_nmi(
  int_nmi),
.int_external(
  int_external),
.int_extern_cause(
  int_extern_cause),
.int_software(
  int_software),
.int_mtime(
  int_mtime),
.imem_req(
  imem_req),
.imem_wen(
  imem_wen),
.imem_strb(
  imem_strb),
.imem_wdata(
  imem_wdata),
.imem_addr(
  imem_addr),
.imem_gnt(
  imem_gnt),
.imem_recv(
  imem_recv),
.imem_ack(
  imem_ack),
.imem_error(
  imem_error),
.imem_rdata(
  imem_rdata),
.dmem_req(
  dmem_req),
.dmem_wen(
  dmem_wen),
.dmem_strb(
  dmem_strb),
.dmem_wdata(
  dmem_wdata),
.dmem_addr(
  dmem_addr),
.dmem_gnt(
  dmem_gnt),
.dmem_recv(
  dmem_recv),
.dmem_ack(
  dmem_ack),
.dmem_error(
  dmem_error),
.dmem_rdata(
  dmem_rdata),
.leak_prng_t0(
  leak_prng_t0),
.imem_wen_t0(
  imem_wen_t0),
.imem_wdata_t0(
  imem_wdata_t0),
.imem_strb_t0(
  imem_strb_t0),
.imem_req_t0(
  imem_req_t0),
.imem_recv_t0(
  imem_recv_t0),
.imem_rdata_t0(
  imem_rdata_t0),
.imem_gnt_t0(
  imem_gnt_t0),
.imem_error_t0(
  imem_error_t0),
.imem_addr_t0(
  imem_addr_t0),
.imem_ack_t0(
  imem_ack_t0),
.rng_req_data_t0(
  rng_req_data_t0),
.rng_req_op_t0(
  rng_req_op_t0),
.rng_req_ready_t0(
  rng_req_ready_t0),
.rng_req_valid_t0(
  rng_req_valid_t0),
.rng_rsp_data_t0(
  rng_rsp_data_t0),
.rng_rsp_ready_t0(
  rng_rsp_ready_t0),
.rng_rsp_status_t0(
  rng_rsp_status_t0),
.rng_rsp_valid_t0(
  rng_rsp_valid_t0),
.dmem_addr_t0(
  dmem_addr_t0),
.dmem_gnt_t0(
  dmem_gnt_t0),
.dmem_req_t0(
  dmem_req_t0),
.dmem_strb_t0(
  dmem_strb_t0),
.dmem_wdata_t0(
  dmem_wdata_t0),
.dmem_wen_t0(
  dmem_wen_t0),
.leak_fence_unc0_t0(
  leak_fence_unc0_t0),
.leak_fence_unc1_t0(
  leak_fence_unc1_t0),
.leak_fence_unc2_t0(
  leak_fence_unc2_t0),
.dmem_ack_t0(
  dmem_ack_t0),
.dmem_error_t0(
  dmem_error_t0),
.dmem_rdata_t0(
  dmem_rdata_t0),
.dmem_recv_t0(
  dmem_recv_t0),
.trs_instr_t0(
  trs_instr_t0),
.trs_pc_t0(
  trs_pc_t0),
.trs_valid_t0(
  trs_valid_t0),
.int_extern_cause_t0(
  int_extern_cause_t0),
.int_external_t0(
  int_external_t0),
.int_mtime_t0(
  int_mtime_t0),
.int_nmi_t0(
  int_nmi_t0),
.int_software_t0(
  int_software_t0),
.ctr_cycle(
  ctr_cycle),
.ctr_cycle_t0(
  ctr_cycle_t0),
.ctr_instret(
  ctr_instret),
.ctr_instret_t0(
  ctr_instret_t0),
.ctr_time(
  ctr_time),
.ctr_time_t0(
  ctr_time_t0),
.inhibit_cy(
  inhibit_cy),
.inhibit_cy_t0(
  inhibit_cy_t0),
.inhibit_ir(
  inhibit_ir),
.inhibit_ir_t0(
  inhibit_ir_t0),
.inhibit_tm(
  inhibit_tm),
.inhibit_tm_t0(
  inhibit_tm_t0),
.instr_ret(
  instr_ret),
.instr_ret_t0(
  instr_ret_t0),
.int_trap_ack(
  int_trap_ack),
.int_trap_ack_t0(
  int_trap_ack_t0),
.int_trap_cause(
  int_trap_cause),
.int_trap_cause_t0(
  int_trap_cause_t0),
.int_trap_req(
  int_trap_req),
.int_trap_req_t0(
  int_trap_req_t0),
.mie_meie(
  mie_meie),
.mie_meie_t0(
  mie_meie_t0),
.mie_msie(
  mie_msie),
.mie_msie_t0(
  mie_msie_t0),
.mie_mtie(
  mie_mtie),
.mie_mtie_t0(
  mie_mtie_t0),
.mip_meip(
  mip_meip),
.mip_meip_t0(
  mip_meip_t0),
.mip_msip(
  mip_msip),
.mip_msip_t0(
  mip_msip_t0),
.mmio_addr(
  mmio_addr),
.mmio_addr_t0(
  mmio_addr_t0),
.mmio_en(
  mmio_en),
.mmio_en_t0(
  mmio_en_t0),
.mmio_error(
  mmio_error),
.mmio_error_t0(
  mmio_error_t0),
.mmio_rdata(
  mmio_rdata),
.mmio_rdata_t0(
  mmio_rdata_t0),
.mmio_wdata(
  mmio_wdata),
.mmio_wdata_t0(
  mmio_wdata_t0),
.mmio_wen(
  mmio_wen),
.mmio_wen_t0(
  mmio_wen_t0),
.mstatus_mie(
  mstatus_mie),
.mstatus_mie_t0(
  mstatus_mie_t0),
.ti_pending(
  ti_pending),
.ti_pending_t0(
  ti_pending_t0),
.i_counters__g_clk(
  i_counters.g_clk),
.i_counters__g_resetn(
  i_counters.g_resetn),
.i_counters__instr_ret(
  i_counters.instr_ret),
.i_counters__timer_interrupt(
  i_counters.timer_interrupt),
.i_counters__ctr_time(
  i_counters.ctr_time),
.i_counters__ctr_cycle(
  i_counters.ctr_cycle),
.i_counters__ctr_instret(
  i_counters.ctr_instret),
.i_counters__inhibit_cy(
  i_counters.inhibit_cy),
.i_counters__inhibit_tm(
  i_counters.inhibit_tm),
.i_counters__inhibit_ir(
  i_counters.inhibit_ir),
.i_counters__mmio_en(
  i_counters.mmio_en),
.i_counters__mmio_wen(
  i_counters.mmio_wen),
.i_counters__mmio_addr(
  i_counters.mmio_addr),
.i_counters__mmio_wdata(
  i_counters.mmio_wdata),
.i_counters__mmio_rdata(
  i_counters.mmio_rdata),
.i_counters__mmio_error(
  i_counters.mmio_error),
.i_counters__timer_interrupt_t0(
  i_counters.timer_interrupt_t0),
.i_counters__mmio_wen_t0(
  i_counters.mmio_wen_t0),
.i_counters__mmio_wdata_t0(
  i_counters.mmio_wdata_t0),
.i_counters__mmio_rdata_t0(
  i_counters.mmio_rdata_t0),
.i_counters__mmio_error_t0(
  i_counters.mmio_error_t0),
.i_counters__mmio_en_t0(
  i_counters.mmio_en_t0),
.i_counters__mmio_addr_t0(
  i_counters.mmio_addr_t0),
.i_counters__instr_ret_t0(
  i_counters.instr_ret_t0),
.i_counters__inhibit_tm_t0(
  i_counters.inhibit_tm_t0),
.i_counters__inhibit_ir_t0(
  i_counters.inhibit_ir_t0),
.i_counters__inhibit_cy_t0(
  i_counters.inhibit_cy_t0),
.i_counters__ctr_time_t0(
  i_counters.ctr_time_t0),
.i_counters__ctr_instret_t0(
  i_counters.ctr_instret_t0),
.i_counters__ctr_cycle_t0(
  i_counters.ctr_cycle_t0),
.i_counters__addr_mtime_hi(
  i_counters.addr_mtime_hi),
.i_counters__addr_mtime_lo(
  i_counters.addr_mtime_lo),
.i_counters__addr_mtimecmp_hi(
  i_counters.addr_mtimecmp_hi),
.i_counters__addr_mtimecmp_lo(
  i_counters.addr_mtimecmp_lo),
.i_counters__mapped_mtimecmp(
  i_counters.mapped_mtimecmp),
.i_counters__mapped_mtimecmp_t0(
  i_counters.mapped_mtimecmp_t0),
.i_counters__n_ctr_cycle(
  i_counters.n_ctr_cycle),
.i_counters__n_ctr_cycle_t0(
  i_counters.n_ctr_cycle_t0),
.i_counters__n_ctr_instret(
  i_counters.n_ctr_instret),
.i_counters__n_ctr_instret_t0(
  i_counters.n_ctr_instret_t0),
.i_counters__n_mapped_mtime(
  i_counters.n_mapped_mtime),
.i_counters__n_mapped_mtime_t0(
  i_counters.n_mapped_mtime_t0),
.i_counters__n_mmio_error(
  i_counters.n_mmio_error),
.i_counters__n_mmio_rdata(
  i_counters.n_mmio_rdata),
.i_counters__n_mmio_rdata_t0(
  i_counters.n_mmio_rdata_t0),
.i_counters__n_timer_interrupt(
  i_counters.n_timer_interrupt),
.i_counters__wr_mtime_hi(
  i_counters.wr_mtime_hi),
.i_counters__wr_mtime_lo(
  i_counters.wr_mtime_lo),
.i_counters__wr_mtimecmp_hi(
  i_counters.wr_mtimecmp_hi),
.i_counters__wr_mtimecmp_lo(
  i_counters.wr_mtimecmp_lo),
.i_interrupts__g_clk(
  i_interrupts.g_clk),
.i_interrupts__g_resetn(
  i_interrupts.g_resetn),
.i_interrupts__mstatus_mie(
  i_interrupts.mstatus_mie),
.i_interrupts__mie_meie(
  i_interrupts.mie_meie),
.i_interrupts__mie_mtie(
  i_interrupts.mie_mtie),
.i_interrupts__mie_msie(
  i_interrupts.mie_msie),
.i_interrupts__nmi_pending(
  i_interrupts.nmi_pending),
.i_interrupts__ex_pending(
  i_interrupts.ex_pending),
.i_interrupts__ex_cause(
  i_interrupts.ex_cause),
.i_interrupts__ti_pending(
  i_interrupts.ti_pending),
.i_interrupts__sw_pending(
  i_interrupts.sw_pending),
.i_interrupts__mip_meip(
  i_interrupts.mip_meip),
.i_interrupts__mip_mtip(
  i_interrupts.mip_mtip),
.i_interrupts__mip_msip(
  i_interrupts.mip_msip),
.i_interrupts__int_trap_req(
  i_interrupts.int_trap_req),
.i_interrupts__int_trap_cause(
  i_interrupts.int_trap_cause),
.i_interrupts__int_trap_ack(
  i_interrupts.int_trap_ack),
.i_interrupts__sw_pending_t0(
  i_interrupts.sw_pending_t0),
.i_interrupts__mip_mtip_t0(
  i_interrupts.mip_mtip_t0),
.i_interrupts__mstatus_mie_t0(
  i_interrupts.mstatus_mie_t0),
.i_interrupts__mie_msie_t0(
  i_interrupts.mie_msie_t0),
.i_interrupts__mie_mtie_t0(
  i_interrupts.mie_mtie_t0),
.i_interrupts__mip_meip_t0(
  i_interrupts.mip_meip_t0),
.i_interrupts__ti_pending_t0(
  i_interrupts.ti_pending_t0),
.i_interrupts__int_trap_req_t0(
  i_interrupts.int_trap_req_t0),
.i_interrupts__ex_cause_t0(
  i_interrupts.ex_cause_t0),
.i_interrupts__mip_msip_t0(
  i_interrupts.mip_msip_t0),
.i_interrupts__ex_pending_t0(
  i_interrupts.ex_pending_t0),
.i_interrupts__int_trap_cause_t0(
  i_interrupts.int_trap_cause_t0),
.i_interrupts__int_trap_ack_t0(
  i_interrupts.int_trap_ack_t0),
.i_interrupts__mie_meie_t0(
  i_interrupts.mie_meie_t0),
.i_interrupts__nmi_pending_t0(
  i_interrupts.nmi_pending_t0),
.i_interrupts__extern_cause(
  i_interrupts.extern_cause),
.i_interrupts__extern_cause_t0(
  i_interrupts.extern_cause_t0),
.i_interrupts__mip_nmi(
  i_interrupts.mip_nmi),
.i_interrupts__n_int_trap_cause(
  i_interrupts.n_int_trap_cause),
.i_interrupts__n_int_trap_cause_t0(
  i_interrupts.n_int_trap_cause_t0),
.i_interrupts__raise_mei(
  i_interrupts.raise_mei),
.i_interrupts__raise_msi(
  i_interrupts.raise_msi),
.i_interrupts__raise_mti(
  i_interrupts.raise_mti),
.i_interrupts__raise_nmi(
  i_interrupts.raise_nmi),
.i_interrupts__use_extern_cause(
  i_interrupts.use_extern_cause),
.i_pipeline__g_clk(
  i_pipeline.g_clk),
.i_pipeline__g_resetn(
  i_pipeline.g_resetn),
.i_pipeline__trs_pc(
  i_pipeline.trs_pc),
.i_pipeline__trs_instr(
  i_pipeline.trs_instr),
.i_pipeline__trs_valid(
  i_pipeline.trs_valid),
.i_pipeline__leak_prng(
  i_pipeline.leak_prng),
.i_pipeline__leak_fence_unc0(
  i_pipeline.leak_fence_unc0),
.i_pipeline__leak_fence_unc1(
  i_pipeline.leak_fence_unc1),
.i_pipeline__leak_fence_unc2(
  i_pipeline.leak_fence_unc2),
.i_pipeline__rng_req_valid(
  i_pipeline.rng_req_valid),
.i_pipeline__rng_req_op(
  i_pipeline.rng_req_op),
.i_pipeline__rng_req_data(
  i_pipeline.rng_req_data),
.i_pipeline__rng_req_ready(
  i_pipeline.rng_req_ready),
.i_pipeline__rng_rsp_valid(
  i_pipeline.rng_rsp_valid),
.i_pipeline__rng_rsp_status(
  i_pipeline.rng_rsp_status),
.i_pipeline__rng_rsp_data(
  i_pipeline.rng_rsp_data),
.i_pipeline__rng_rsp_ready(
  i_pipeline.rng_rsp_ready),
.i_pipeline__instr_ret(
  i_pipeline.instr_ret),
.i_pipeline__mstatus_mie(
  i_pipeline.mstatus_mie),
.i_pipeline__mie_meie(
  i_pipeline.mie_meie),
.i_pipeline__mie_mtie(
  i_pipeline.mie_mtie),
.i_pipeline__mie_msie(
  i_pipeline.mie_msie),
.i_pipeline__mip_meip(
  i_pipeline.mip_meip),
.i_pipeline__mip_mtip(
  i_pipeline.mip_mtip),
.i_pipeline__mip_msip(
  i_pipeline.mip_msip),
.i_pipeline__ctr_time(
  i_pipeline.ctr_time),
.i_pipeline__ctr_cycle(
  i_pipeline.ctr_cycle),
.i_pipeline__ctr_instret(
  i_pipeline.ctr_instret),
.i_pipeline__int_trap_req(
  i_pipeline.int_trap_req),
.i_pipeline__int_trap_cause(
  i_pipeline.int_trap_cause),
.i_pipeline__int_trap_ack(
  i_pipeline.int_trap_ack),
.i_pipeline__inhibit_cy(
  i_pipeline.inhibit_cy),
.i_pipeline__inhibit_tm(
  i_pipeline.inhibit_tm),
.i_pipeline__inhibit_ir(
  i_pipeline.inhibit_ir),
.i_pipeline__mmio_en(
  i_pipeline.mmio_en),
.i_pipeline__mmio_wen(
  i_pipeline.mmio_wen),
.i_pipeline__mmio_addr(
  i_pipeline.mmio_addr),
.i_pipeline__mmio_wdata(
  i_pipeline.mmio_wdata),
.i_pipeline__mmio_rdata(
  i_pipeline.mmio_rdata),
.i_pipeline__mmio_error(
  i_pipeline.mmio_error),
.i_pipeline__imem_req(
  i_pipeline.imem_req),
.i_pipeline__imem_wen(
  i_pipeline.imem_wen),
.i_pipeline__imem_strb(
  i_pipeline.imem_strb),
.i_pipeline__imem_wdata(
  i_pipeline.imem_wdata),
.i_pipeline__imem_addr(
  i_pipeline.imem_addr),
.i_pipeline__imem_gnt(
  i_pipeline.imem_gnt),
.i_pipeline__imem_recv(
  i_pipeline.imem_recv),
.i_pipeline__imem_ack(
  i_pipeline.imem_ack),
.i_pipeline__imem_error(
  i_pipeline.imem_error),
.i_pipeline__imem_rdata(
  i_pipeline.imem_rdata),
.i_pipeline__dmem_req(
  i_pipeline.dmem_req),
.i_pipeline__dmem_wen(
  i_pipeline.dmem_wen),
.i_pipeline__dmem_strb(
  i_pipeline.dmem_strb),
.i_pipeline__dmem_wdata(
  i_pipeline.dmem_wdata),
.i_pipeline__dmem_addr(
  i_pipeline.dmem_addr),
.i_pipeline__dmem_gnt(
  i_pipeline.dmem_gnt),
.i_pipeline__dmem_recv(
  i_pipeline.dmem_recv),
.i_pipeline__dmem_ack(
  i_pipeline.dmem_ack),
.i_pipeline__dmem_error(
  i_pipeline.dmem_error),
.i_pipeline__dmem_rdata(
  i_pipeline.dmem_rdata),
.i_pipeline__mip_mtip_t0(
  i_pipeline.mip_mtip_t0),
.i_pipeline__mstatus_mie_t0(
  i_pipeline.mstatus_mie_t0),
.i_pipeline__mie_msie_t0(
  i_pipeline.mie_msie_t0),
.i_pipeline__mie_mtie_t0(
  i_pipeline.mie_mtie_t0),
.i_pipeline__mip_meip_t0(
  i_pipeline.mip_meip_t0),
.i_pipeline__leak_prng_t0(
  i_pipeline.leak_prng_t0),
.i_pipeline__imem_wen_t0(
  i_pipeline.imem_wen_t0),
.i_pipeline__imem_wdata_t0(
  i_pipeline.imem_wdata_t0),
.i_pipeline__imem_strb_t0(
  i_pipeline.imem_strb_t0),
.i_pipeline__imem_req_t0(
  i_pipeline.imem_req_t0),
.i_pipeline__imem_recv_t0(
  i_pipeline.imem_recv_t0),
.i_pipeline__imem_rdata_t0(
  i_pipeline.imem_rdata_t0),
.i_pipeline__imem_gnt_t0(
  i_pipeline.imem_gnt_t0),
.i_pipeline__imem_error_t0(
  i_pipeline.imem_error_t0),
.i_pipeline__imem_addr_t0(
  i_pipeline.imem_addr_t0),
.i_pipeline__imem_ack_t0(
  i_pipeline.imem_ack_t0),
.i_pipeline__int_trap_req_t0(
  i_pipeline.int_trap_req_t0),
.i_pipeline__mmio_wen_t0(
  i_pipeline.mmio_wen_t0),
.i_pipeline__mmio_wdata_t0(
  i_pipeline.mmio_wdata_t0),
.i_pipeline__mmio_rdata_t0(
  i_pipeline.mmio_rdata_t0),
.i_pipeline__mmio_error_t0(
  i_pipeline.mmio_error_t0),
.i_pipeline__mmio_en_t0(
  i_pipeline.mmio_en_t0),
.i_pipeline__mmio_addr_t0(
  i_pipeline.mmio_addr_t0),
.i_pipeline__instr_ret_t0(
  i_pipeline.instr_ret_t0),
.i_pipeline__inhibit_tm_t0(
  i_pipeline.inhibit_tm_t0),
.i_pipeline__inhibit_ir_t0(
  i_pipeline.inhibit_ir_t0),
.i_pipeline__inhibit_cy_t0(
  i_pipeline.inhibit_cy_t0),
.i_pipeline__ctr_time_t0(
  i_pipeline.ctr_time_t0),
.i_pipeline__ctr_instret_t0(
  i_pipeline.ctr_instret_t0),
.i_pipeline__ctr_cycle_t0(
  i_pipeline.ctr_cycle_t0),
.i_pipeline__mip_msip_t0(
  i_pipeline.mip_msip_t0),
.i_pipeline__int_trap_cause_t0(
  i_pipeline.int_trap_cause_t0),
.i_pipeline__int_trap_ack_t0(
  i_pipeline.int_trap_ack_t0),
.i_pipeline__mie_meie_t0(
  i_pipeline.mie_meie_t0),
.i_pipeline__rng_req_data_t0(
  i_pipeline.rng_req_data_t0),
.i_pipeline__rng_req_op_t0(
  i_pipeline.rng_req_op_t0),
.i_pipeline__rng_req_ready_t0(
  i_pipeline.rng_req_ready_t0),
.i_pipeline__rng_req_valid_t0(
  i_pipeline.rng_req_valid_t0),
.i_pipeline__rng_rsp_data_t0(
  i_pipeline.rng_rsp_data_t0),
.i_pipeline__rng_rsp_ready_t0(
  i_pipeline.rng_rsp_ready_t0),
.i_pipeline__rng_rsp_status_t0(
  i_pipeline.rng_rsp_status_t0),
.i_pipeline__rng_rsp_valid_t0(
  i_pipeline.rng_rsp_valid_t0),
.i_pipeline__dmem_addr_t0(
  i_pipeline.dmem_addr_t0),
.i_pipeline__dmem_gnt_t0(
  i_pipeline.dmem_gnt_t0),
.i_pipeline__dmem_req_t0(
  i_pipeline.dmem_req_t0),
.i_pipeline__dmem_strb_t0(
  i_pipeline.dmem_strb_t0),
.i_pipeline__dmem_wdata_t0(
  i_pipeline.dmem_wdata_t0),
.i_pipeline__dmem_wen_t0(
  i_pipeline.dmem_wen_t0),
.i_pipeline__leak_fence_unc0_t0(
  i_pipeline.leak_fence_unc0_t0),
.i_pipeline__leak_fence_unc1_t0(
  i_pipeline.leak_fence_unc1_t0),
.i_pipeline__leak_fence_unc2_t0(
  i_pipeline.leak_fence_unc2_t0),
.i_pipeline__dmem_ack_t0(
  i_pipeline.dmem_ack_t0),
.i_pipeline__dmem_error_t0(
  i_pipeline.dmem_error_t0),
.i_pipeline__dmem_rdata_t0(
  i_pipeline.dmem_rdata_t0),
.i_pipeline__dmem_recv_t0(
  i_pipeline.dmem_recv_t0),
.i_pipeline__trs_instr_t0(
  i_pipeline.trs_instr_t0),
.i_pipeline__trs_pc_t0(
  i_pipeline.trs_pc_t0),
.i_pipeline__trs_valid_t0(
  i_pipeline.trs_valid_t0),
.i_pipeline__cf_ack(
  i_pipeline.cf_ack),
.i_pipeline__cf_ack_t0(
  i_pipeline.cf_ack_t0),
.i_pipeline__cf_req(
  i_pipeline.cf_req),
.i_pipeline__cf_req_t0(
  i_pipeline.cf_req_t0),
.i_pipeline__cf_target(
  i_pipeline.cf_target),
.i_pipeline__cf_target_t0(
  i_pipeline.cf_target_t0),
.i_pipeline__csr_addr(
  i_pipeline.csr_addr),
.i_pipeline__csr_addr_t0(
  i_pipeline.csr_addr_t0),
.i_pipeline__csr_en(
  i_pipeline.csr_en),
.i_pipeline__csr_en_t0(
  i_pipeline.csr_en_t0),
.i_pipeline__csr_error(
  i_pipeline.csr_error),
.i_pipeline__csr_error_t0(
  i_pipeline.csr_error_t0),
.i_pipeline__csr_mepc(
  i_pipeline.csr_mepc),
.i_pipeline__csr_mepc_t0(
  i_pipeline.csr_mepc_t0),
.i_pipeline__csr_mtvec(
  i_pipeline.csr_mtvec),
.i_pipeline__csr_mtvec_t0(
  i_pipeline.csr_mtvec_t0),
.i_pipeline__csr_rdata(
  i_pipeline.csr_rdata),
.i_pipeline__csr_rdata_t0(
  i_pipeline.csr_rdata_t0),
.i_pipeline__csr_wdata(
  i_pipeline.csr_wdata),
.i_pipeline__csr_wdata_t0(
  i_pipeline.csr_wdata_t0),
.i_pipeline__csr_wr(
  i_pipeline.csr_wr),
.i_pipeline__csr_wr_clr(
  i_pipeline.csr_wr_clr),
.i_pipeline__csr_wr_clr_t0(
  i_pipeline.csr_wr_clr_t0),
.i_pipeline__csr_wr_set(
  i_pipeline.csr_wr_set),
.i_pipeline__csr_wr_set_t0(
  i_pipeline.csr_wr_set_t0),
.i_pipeline__csr_wr_t0(
  i_pipeline.csr_wr_t0),
.i_pipeline__exec_mret(
  i_pipeline.exec_mret),
.i_pipeline__exec_mret_t0(
  i_pipeline.exec_mret_t0),
.i_pipeline__fwd_rs1_rdata(
  i_pipeline.fwd_rs1_rdata),
.i_pipeline__fwd_rs1_rdata_t0(
  i_pipeline.fwd_rs1_rdata_t0),
.i_pipeline__fwd_rs2_rdata(
  i_pipeline.fwd_rs2_rdata),
.i_pipeline__fwd_rs2_rdata_t0(
  i_pipeline.fwd_rs2_rdata_t0),
.i_pipeline__fwd_rs3_rdata(
  i_pipeline.fwd_rs3_rdata),
.i_pipeline__fwd_rs3_rdata_t0(
  i_pipeline.fwd_rs3_rdata_t0),
.i_pipeline__fwd_s2_csr(
  i_pipeline.fwd_s2_csr),
.i_pipeline__fwd_s2_csr_t0(
  i_pipeline.fwd_s2_csr_t0),
.i_pipeline__fwd_s2_load(
  i_pipeline.fwd_s2_load),
.i_pipeline__fwd_s2_load_t0(
  i_pipeline.fwd_s2_load_t0),
.i_pipeline__fwd_s2_rd(
  i_pipeline.fwd_s2_rd),
.i_pipeline__fwd_s2_rd_t0(
  i_pipeline.fwd_s2_rd_t0),
.i_pipeline__fwd_s2_rs1_hi(
  i_pipeline.fwd_s2_rs1_hi),
.i_pipeline__fwd_s2_rs2_hi(
  i_pipeline.fwd_s2_rs2_hi),
.i_pipeline__fwd_s2_rs3_hi(
  i_pipeline.fwd_s2_rs3_hi),
.i_pipeline__fwd_s2_wdata(
  i_pipeline.fwd_s2_wdata),
.i_pipeline__fwd_s2_wdata_hi(
  i_pipeline.fwd_s2_wdata_hi),
.i_pipeline__fwd_s2_wdata_hi_t0(
  i_pipeline.fwd_s2_wdata_hi_t0),
.i_pipeline__fwd_s2_wdata_t0(
  i_pipeline.fwd_s2_wdata_t0),
.i_pipeline__fwd_s2_wide(
  i_pipeline.fwd_s2_wide),
.i_pipeline__fwd_s2_wide_t0(
  i_pipeline.fwd_s2_wide_t0),
.i_pipeline__fwd_s3_csr(
  i_pipeline.fwd_s3_csr),
.i_pipeline__fwd_s3_csr_t0(
  i_pipeline.fwd_s3_csr_t0),
.i_pipeline__fwd_s3_load(
  i_pipeline.fwd_s3_load),
.i_pipeline__fwd_s3_load_t0(
  i_pipeline.fwd_s3_load_t0),
.i_pipeline__fwd_s3_rd(
  i_pipeline.fwd_s3_rd),
.i_pipeline__fwd_s3_rd_t0(
  i_pipeline.fwd_s3_rd_t0),
.i_pipeline__fwd_s3_rs1_hi(
  i_pipeline.fwd_s3_rs1_hi),
.i_pipeline__fwd_s3_rs2_hi(
  i_pipeline.fwd_s3_rs2_hi),
.i_pipeline__fwd_s3_rs3_hi(
  i_pipeline.fwd_s3_rs3_hi),
.i_pipeline__fwd_s3_wdata(
  i_pipeline.fwd_s3_wdata),
.i_pipeline__fwd_s3_wdata_hi(
  i_pipeline.fwd_s3_wdata_hi),
.i_pipeline__fwd_s3_wdata_hi_t0(
  i_pipeline.fwd_s3_wdata_hi_t0),
.i_pipeline__fwd_s3_wdata_t0(
  i_pipeline.fwd_s3_wdata_t0),
.i_pipeline__fwd_s3_wide(
  i_pipeline.fwd_s3_wide),
.i_pipeline__fwd_s3_wide_t0(
  i_pipeline.fwd_s3_wide_t0),
.i_pipeline__fwd_s4_csr(
  i_pipeline.fwd_s4_csr),
.i_pipeline__fwd_s4_csr_t0(
  i_pipeline.fwd_s4_csr_t0),
.i_pipeline__fwd_s4_load(
  i_pipeline.fwd_s4_load),
.i_pipeline__fwd_s4_load_t0(
  i_pipeline.fwd_s4_load_t0),
.i_pipeline__fwd_s4_rd(
  i_pipeline.fwd_s4_rd),
.i_pipeline__fwd_s4_rd_t0(
  i_pipeline.fwd_s4_rd_t0),
.i_pipeline__fwd_s4_rs1_hi(
  i_pipeline.fwd_s4_rs1_hi),
.i_pipeline__fwd_s4_rs2_hi(
  i_pipeline.fwd_s4_rs2_hi),
.i_pipeline__fwd_s4_rs3_hi(
  i_pipeline.fwd_s4_rs3_hi),
.i_pipeline__fwd_s4_wdata(
  i_pipeline.fwd_s4_wdata),
.i_pipeline__fwd_s4_wdata_t0(
  i_pipeline.fwd_s4_wdata_t0),
.i_pipeline__gpr_rd(
  i_pipeline.gpr_rd),
.i_pipeline__gpr_rd_t0(
  i_pipeline.gpr_rd_t0),
.i_pipeline__gpr_wdata(
  i_pipeline.gpr_wdata),
.i_pipeline__gpr_wdata_hi(
  i_pipeline.gpr_wdata_hi),
.i_pipeline__gpr_wdata_hi_t0(
  i_pipeline.gpr_wdata_hi_t0),
.i_pipeline__gpr_wdata_t0(
  i_pipeline.gpr_wdata_t0),
.i_pipeline__gpr_wen(
  i_pipeline.gpr_wen),
.i_pipeline__gpr_wen_t0(
  i_pipeline.gpr_wen_t0),
.i_pipeline__gpr_wide(
  i_pipeline.gpr_wide),
.i_pipeline__gpr_wide_t0(
  i_pipeline.gpr_wide_t0),
.i_pipeline__hold_lsu_req(
  i_pipeline.hold_lsu_req),
.i_pipeline__hold_lsu_req_t0(
  i_pipeline.hold_lsu_req_t0),
.i_pipeline__hzd_rs1_s2(
  i_pipeline.hzd_rs1_s2),
.i_pipeline__hzd_rs1_s3(
  i_pipeline.hzd_rs1_s3),
.i_pipeline__hzd_rs1_s4(
  i_pipeline.hzd_rs1_s4),
.i_pipeline__hzd_rs2_s2(
  i_pipeline.hzd_rs2_s2),
.i_pipeline__hzd_rs2_s3(
  i_pipeline.hzd_rs2_s3),
.i_pipeline__hzd_rs2_s4(
  i_pipeline.hzd_rs2_s4),
.i_pipeline__hzd_rs3_s2(
  i_pipeline.hzd_rs3_s2),
.i_pipeline__hzd_rs3_s3(
  i_pipeline.hzd_rs3_s3),
.i_pipeline__hzd_rs3_s4(
  i_pipeline.hzd_rs3_s4),
.i_pipeline__leak_lkgcfg(
  i_pipeline.leak_lkgcfg),
.i_pipeline__leak_lkgcfg_t0(
  i_pipeline.leak_lkgcfg_t0),
.i_pipeline__nz_s1_rs1(
  i_pipeline.nz_s1_rs1),
.i_pipeline__nz_s1_rs2(
  i_pipeline.nz_s1_rs2),
.i_pipeline__nz_s1_rs3(
  i_pipeline.nz_s1_rs3),
.i_pipeline__s0_flush(
  i_pipeline.s0_flush),
.i_pipeline__s1_bubble(
  i_pipeline.s1_bubble),
.i_pipeline__s1_bubble_from_s2(
  i_pipeline.s1_bubble_from_s2),
.i_pipeline__s1_bubble_from_s3(
  i_pipeline.s1_bubble_from_s3),
.i_pipeline__s1_bubble_from_s4(
  i_pipeline.s1_bubble_from_s4),
.i_pipeline__s1_bubble_no_instr(
  i_pipeline.s1_bubble_no_instr),
.i_pipeline__s1_busy(
  i_pipeline.s1_busy),
.i_pipeline__s1_busy_t0(
  i_pipeline.s1_busy_t0),
.i_pipeline__s1_data(
  i_pipeline.s1_data),
.i_pipeline__s1_data_t0(
  i_pipeline.s1_data_t0),
.i_pipeline__s1_error(
  i_pipeline.s1_error),
.i_pipeline__s1_error_t0(
  i_pipeline.s1_error_t0),
.i_pipeline__s1_leak_fence(
  i_pipeline.s1_leak_fence),
.i_pipeline__s1_leak_fence_t0(
  i_pipeline.s1_leak_fence_t0),
.i_pipeline__s1_rs1_addr(
  i_pipeline.s1_rs1_addr),
.i_pipeline__s1_rs1_addr_t0(
  i_pipeline.s1_rs1_addr_t0),
.i_pipeline__s1_rs1_rdata(
  i_pipeline.s1_rs1_rdata),
.i_pipeline__s1_rs1_rdata_t0(
  i_pipeline.s1_rs1_rdata_t0),
.i_pipeline__s1_rs2_addr(
  i_pipeline.s1_rs2_addr),
.i_pipeline__s1_rs2_addr_t0(
  i_pipeline.s1_rs2_addr_t0),
.i_pipeline__s1_rs2_rdata(
  i_pipeline.s1_rs2_rdata),
.i_pipeline__s1_rs2_rdata_t0(
  i_pipeline.s1_rs2_rdata_t0),
.i_pipeline__s1_rs3_addr(
  i_pipeline.s1_rs3_addr),
.i_pipeline__s1_rs3_addr_t0(
  i_pipeline.s1_rs3_addr_t0),
.i_pipeline__s1_rs3_rdata(
  i_pipeline.s1_rs3_rdata),
.i_pipeline__s1_rs3_rdata_t0(
  i_pipeline.s1_rs3_rdata_t0),
.i_pipeline__s1_valid(
  i_pipeline.s1_valid),
.i_pipeline__s1_valid_t0(
  i_pipeline.s1_valid_t0),
.i_pipeline__s2_busy(
  i_pipeline.s2_busy),
.i_pipeline__s2_busy_t0(
  i_pipeline.s2_busy_t0),
.i_pipeline__s2_fu(
  i_pipeline.s2_fu),
.i_pipeline__s2_fu_t0(
  i_pipeline.s2_fu_t0),
.i_pipeline__s2_instr(
  i_pipeline.s2_instr),
.i_pipeline__s2_instr_t0(
  i_pipeline.s2_instr_t0),
.i_pipeline__s2_opr_a(
  i_pipeline.s2_opr_a),
.i_pipeline__s2_opr_a_t0(
  i_pipeline.s2_opr_a_t0),
.i_pipeline__s2_opr_b(
  i_pipeline.s2_opr_b),
.i_pipeline__s2_opr_b_t0(
  i_pipeline.s2_opr_b_t0),
.i_pipeline__s2_opr_c(
  i_pipeline.s2_opr_c),
.i_pipeline__s2_opr_c_t0(
  i_pipeline.s2_opr_c_t0),
.i_pipeline__s2_pw(
  i_pipeline.s2_pw),
.i_pipeline__s2_pw_t0(
  i_pipeline.s2_pw_t0),
.i_pipeline__s2_rd(
  i_pipeline.s2_rd),
.i_pipeline__s2_rd_t0(
  i_pipeline.s2_rd_t0),
.i_pipeline__s2_size(
  i_pipeline.s2_size),
.i_pipeline__s2_size_t0(
  i_pipeline.s2_size_t0),
.i_pipeline__s2_trap(
  i_pipeline.s2_trap),
.i_pipeline__s2_trap_t0(
  i_pipeline.s2_trap_t0),
.i_pipeline__s2_uop(
  i_pipeline.s2_uop),
.i_pipeline__s2_uop_t0(
  i_pipeline.s2_uop_t0),
.i_pipeline__s2_valid(
  i_pipeline.s2_valid),
.i_pipeline__s2_valid_t0(
  i_pipeline.s2_valid_t0),
.i_pipeline__s3_busy(
  i_pipeline.s3_busy),
.i_pipeline__s3_busy_t0(
  i_pipeline.s3_busy_t0),
.i_pipeline__s3_fu(
  i_pipeline.s3_fu),
.i_pipeline__s3_fu_t0(
  i_pipeline.s3_fu_t0),
.i_pipeline__s3_instr(
  i_pipeline.s3_instr),
.i_pipeline__s3_instr_t0(
  i_pipeline.s3_instr_t0),
.i_pipeline__s3_opr_a(
  i_pipeline.s3_opr_a),
.i_pipeline__s3_opr_a_t0(
  i_pipeline.s3_opr_a_t0),
.i_pipeline__s3_opr_b(
  i_pipeline.s3_opr_b),
.i_pipeline__s3_opr_b_t0(
  i_pipeline.s3_opr_b_t0),
.i_pipeline__s3_rd(
  i_pipeline.s3_rd),
.i_pipeline__s3_rd_t0(
  i_pipeline.s3_rd_t0),
.i_pipeline__s3_size(
  i_pipeline.s3_size),
.i_pipeline__s3_size_t0(
  i_pipeline.s3_size_t0),
.i_pipeline__s3_trap(
  i_pipeline.s3_trap),
.i_pipeline__s3_trap_t0(
  i_pipeline.s3_trap_t0),
.i_pipeline__s3_uop(
  i_pipeline.s3_uop),
.i_pipeline__s3_uop_t0(
  i_pipeline.s3_uop_t0),
.i_pipeline__s3_valid(
  i_pipeline.s3_valid),
.i_pipeline__s3_valid_t0(
  i_pipeline.s3_valid_t0),
.i_pipeline__s4_busy(
  i_pipeline.s4_busy),
.i_pipeline__s4_busy_t0(
  i_pipeline.s4_busy_t0),
.i_pipeline__s4_fu(
  i_pipeline.s4_fu),
.i_pipeline__s4_fu_t0(
  i_pipeline.s4_fu_t0),
.i_pipeline__s4_instr(
  i_pipeline.s4_instr),
.i_pipeline__s4_instr_t0(
  i_pipeline.s4_instr_t0),
.i_pipeline__s4_opr_a(
  i_pipeline.s4_opr_a),
.i_pipeline__s4_opr_a_t0(
  i_pipeline.s4_opr_a_t0),
.i_pipeline__s4_opr_b(
  i_pipeline.s4_opr_b),
.i_pipeline__s4_opr_b_t0(
  i_pipeline.s4_opr_b_t0),
.i_pipeline__s4_rd(
  i_pipeline.s4_rd),
.i_pipeline__s4_rd_t0(
  i_pipeline.s4_rd_t0),
.i_pipeline__s4_size(
  i_pipeline.s4_size),
.i_pipeline__s4_size_t0(
  i_pipeline.s4_size_t0),
.i_pipeline__s4_trap(
  i_pipeline.s4_trap),
.i_pipeline__s4_trap_t0(
  i_pipeline.s4_trap_t0),
.i_pipeline__s4_uop(
  i_pipeline.s4_uop),
.i_pipeline__s4_uop_t0(
  i_pipeline.s4_uop_t0),
.i_pipeline__s4_valid(
  i_pipeline.s4_valid),
.i_pipeline__s4_valid_t0(
  i_pipeline.s4_valid_t0),
.i_pipeline__trap_cause(
  i_pipeline.trap_cause),
.i_pipeline__trap_cause_t0(
  i_pipeline.trap_cause_t0),
.i_pipeline__trap_cpu(
  i_pipeline.trap_cpu),
.i_pipeline__trap_cpu_t0(
  i_pipeline.trap_cpu_t0),
.i_pipeline__trap_int(
  i_pipeline.trap_int),
.i_pipeline__trap_int_t0(
  i_pipeline.trap_int_t0),
.i_pipeline__trap_mtval(
  i_pipeline.trap_mtval),
.i_pipeline__trap_mtval_t0(
  i_pipeline.trap_mtval_t0),
.i_pipeline__trap_pc(
  i_pipeline.trap_pc),
.i_pipeline__trap_pc_t0(
  i_pipeline.trap_pc_t0),
.i_pipeline__uxcrypto_b0(
  i_pipeline.uxcrypto_b0),
.i_pipeline__uxcrypto_b0_t0(
  i_pipeline.uxcrypto_b0_t0),
.i_pipeline__uxcrypto_b1(
  i_pipeline.uxcrypto_b1),
.i_pipeline__uxcrypto_b1_t0(
  i_pipeline.uxcrypto_b1_t0),
.i_pipeline__uxcrypto_ct(
  i_pipeline.uxcrypto_ct),
.i_pipeline__uxcrypto_ct_t0(
  i_pipeline.uxcrypto_ct_t0),
.i_pipeline__vector_intrs(
  i_pipeline.vector_intrs),
.i_pipeline__vector_intrs_t0(
  i_pipeline.vector_intrs_t0),
.i_pipeline__i_csrs__g_clk(
  i_pipeline.i_csrs.g_clk),
.i_pipeline__i_csrs__g_resetn(
  i_pipeline.i_csrs.g_resetn),
.i_pipeline__i_csrs__csr_en(
  i_pipeline.i_csrs.csr_en),
.i_pipeline__i_csrs__csr_wr(
  i_pipeline.i_csrs.csr_wr),
.i_pipeline__i_csrs__csr_wr_set(
  i_pipeline.i_csrs.csr_wr_set),
.i_pipeline__i_csrs__csr_wr_clr(
  i_pipeline.i_csrs.csr_wr_clr),
.i_pipeline__i_csrs__csr_addr(
  i_pipeline.i_csrs.csr_addr),
.i_pipeline__i_csrs__csr_wdata(
  i_pipeline.i_csrs.csr_wdata),
.i_pipeline__i_csrs__csr_rdata(
  i_pipeline.i_csrs.csr_rdata),
.i_pipeline__i_csrs__csr_error(
  i_pipeline.i_csrs.csr_error),
.i_pipeline__i_csrs__csr_mepc(
  i_pipeline.i_csrs.csr_mepc),
.i_pipeline__i_csrs__csr_mtvec(
  i_pipeline.i_csrs.csr_mtvec),
.i_pipeline__i_csrs__vector_intrs(
  i_pipeline.i_csrs.vector_intrs),
.i_pipeline__i_csrs__exec_mret(
  i_pipeline.i_csrs.exec_mret),
.i_pipeline__i_csrs__mstatus_mie(
  i_pipeline.i_csrs.mstatus_mie),
.i_pipeline__i_csrs__mie_meie(
  i_pipeline.i_csrs.mie_meie),
.i_pipeline__i_csrs__mie_mtie(
  i_pipeline.i_csrs.mie_mtie),
.i_pipeline__i_csrs__mie_msie(
  i_pipeline.i_csrs.mie_msie),
.i_pipeline__i_csrs__mip_meip(
  i_pipeline.i_csrs.mip_meip),
.i_pipeline__i_csrs__mip_mtip(
  i_pipeline.i_csrs.mip_mtip),
.i_pipeline__i_csrs__mip_msip(
  i_pipeline.i_csrs.mip_msip),
.i_pipeline__i_csrs__ctr_time(
  i_pipeline.i_csrs.ctr_time),
.i_pipeline__i_csrs__ctr_cycle(
  i_pipeline.i_csrs.ctr_cycle),
.i_pipeline__i_csrs__ctr_instret(
  i_pipeline.i_csrs.ctr_instret),
.i_pipeline__i_csrs__inhibit_cy(
  i_pipeline.i_csrs.inhibit_cy),
.i_pipeline__i_csrs__inhibit_tm(
  i_pipeline.i_csrs.inhibit_tm),
.i_pipeline__i_csrs__inhibit_ir(
  i_pipeline.i_csrs.inhibit_ir),
.i_pipeline__i_csrs__uxcrypto_ct(
  i_pipeline.i_csrs.uxcrypto_ct),
.i_pipeline__i_csrs__uxcrypto_b0(
  i_pipeline.i_csrs.uxcrypto_b0),
.i_pipeline__i_csrs__uxcrypto_b1(
  i_pipeline.i_csrs.uxcrypto_b1),
.i_pipeline__i_csrs__leak_lkgcfg(
  i_pipeline.i_csrs.leak_lkgcfg),
.i_pipeline__i_csrs__trap_cpu(
  i_pipeline.i_csrs.trap_cpu),
.i_pipeline__i_csrs__trap_int(
  i_pipeline.i_csrs.trap_int),
.i_pipeline__i_csrs__trap_cause(
  i_pipeline.i_csrs.trap_cause),
.i_pipeline__i_csrs__trap_mtval(
  i_pipeline.i_csrs.trap_mtval),
.i_pipeline__i_csrs__trap_pc(
  i_pipeline.i_csrs.trap_pc),
.i_pipeline__i_csrs__mip_mtip_t0(
  i_pipeline.i_csrs.mip_mtip_t0),
.i_pipeline__i_csrs__mstatus_mie_t0(
  i_pipeline.i_csrs.mstatus_mie_t0),
.i_pipeline__i_csrs__mie_msie_t0(
  i_pipeline.i_csrs.mie_msie_t0),
.i_pipeline__i_csrs__mie_mtie_t0(
  i_pipeline.i_csrs.mie_mtie_t0),
.i_pipeline__i_csrs__mip_meip_t0(
  i_pipeline.i_csrs.mip_meip_t0),
.i_pipeline__i_csrs__leak_lkgcfg_t0(
  i_pipeline.i_csrs.leak_lkgcfg_t0),
.i_pipeline__i_csrs__trap_cause_t0(
  i_pipeline.i_csrs.trap_cause_t0),
.i_pipeline__i_csrs__inhibit_tm_t0(
  i_pipeline.i_csrs.inhibit_tm_t0),
.i_pipeline__i_csrs__inhibit_ir_t0(
  i_pipeline.i_csrs.inhibit_ir_t0),
.i_pipeline__i_csrs__inhibit_cy_t0(
  i_pipeline.i_csrs.inhibit_cy_t0),
.i_pipeline__i_csrs__ctr_time_t0(
  i_pipeline.i_csrs.ctr_time_t0),
.i_pipeline__i_csrs__ctr_instret_t0(
  i_pipeline.i_csrs.ctr_instret_t0),
.i_pipeline__i_csrs__ctr_cycle_t0(
  i_pipeline.i_csrs.ctr_cycle_t0),
.i_pipeline__i_csrs__mip_msip_t0(
  i_pipeline.i_csrs.mip_msip_t0),
.i_pipeline__i_csrs__mie_meie_t0(
  i_pipeline.i_csrs.mie_meie_t0),
.i_pipeline__i_csrs__uxcrypto_b0_t0(
  i_pipeline.i_csrs.uxcrypto_b0_t0),
.i_pipeline__i_csrs__uxcrypto_b1_t0(
  i_pipeline.i_csrs.uxcrypto_b1_t0),
.i_pipeline__i_csrs__uxcrypto_ct_t0(
  i_pipeline.i_csrs.uxcrypto_ct_t0),
.i_pipeline__i_csrs__csr_addr_t0(
  i_pipeline.i_csrs.csr_addr_t0),
.i_pipeline__i_csrs__csr_en_t0(
  i_pipeline.i_csrs.csr_en_t0),
.i_pipeline__i_csrs__csr_error_t0(
  i_pipeline.i_csrs.csr_error_t0),
.i_pipeline__i_csrs__csr_mepc_t0(
  i_pipeline.i_csrs.csr_mepc_t0),
.i_pipeline__i_csrs__csr_mtvec_t0(
  i_pipeline.i_csrs.csr_mtvec_t0),
.i_pipeline__i_csrs__csr_rdata_t0(
  i_pipeline.i_csrs.csr_rdata_t0),
.i_pipeline__i_csrs__csr_wdata_t0(
  i_pipeline.i_csrs.csr_wdata_t0),
.i_pipeline__i_csrs__csr_wr_t0(
  i_pipeline.i_csrs.csr_wr_t0),
.i_pipeline__i_csrs__csr_wr_clr_t0(
  i_pipeline.i_csrs.csr_wr_clr_t0),
.i_pipeline__i_csrs__csr_wr_set_t0(
  i_pipeline.i_csrs.csr_wr_set_t0),
.i_pipeline__i_csrs__exec_mret_t0(
  i_pipeline.i_csrs.exec_mret_t0),
.i_pipeline__i_csrs__trap_cpu_t0(
  i_pipeline.i_csrs.trap_cpu_t0),
.i_pipeline__i_csrs__trap_int_t0(
  i_pipeline.i_csrs.trap_int_t0),
.i_pipeline__i_csrs__trap_mtval_t0(
  i_pipeline.i_csrs.trap_mtval_t0),
.i_pipeline__i_csrs__trap_pc_t0(
  i_pipeline.i_csrs.trap_pc_t0),
.i_pipeline__i_csrs__vector_intrs_t0(
  i_pipeline.i_csrs.vector_intrs_t0),
.i_pipeline__i_csrs__int_pulse(
  i_pipeline.i_csrs.int_pulse),
.i_pipeline__i_csrs__invalid_addr(
  i_pipeline.i_csrs.invalid_addr),
.i_pipeline__i_csrs__mtvec_bad_write(
  i_pipeline.i_csrs.mtvec_bad_write),
.i_pipeline__i_csrs__n_mcause_cause(
  i_pipeline.i_csrs.n_mcause_cause),
.i_pipeline__i_csrs__n_mcause_cause_t0(
  i_pipeline.i_csrs.n_mcause_cause_t0),
.i_pipeline__i_csrs__n_mepc(
  i_pipeline.i_csrs.n_mepc),
.i_pipeline__i_csrs__n_mepc_t0(
  i_pipeline.i_csrs.n_mepc_t0),
.i_pipeline__i_csrs__n_mstatus_mie(
  i_pipeline.i_csrs.n_mstatus_mie),
.i_pipeline__i_csrs__n_mstatus_mie_t0(
  i_pipeline.i_csrs.n_mstatus_mie_t0),
.i_pipeline__i_csrs__n_mstatus_mpie(
  i_pipeline.i_csrs.n_mstatus_mpie),
.i_pipeline__i_csrs__n_mstatus_mpie_t0(
  i_pipeline.i_csrs.n_mstatus_mpie_t0),
.i_pipeline__i_csrs__n_mtvec_base(
  i_pipeline.i_csrs.n_mtvec_base),
.i_pipeline__i_csrs__n_mtvec_base_t0(
  i_pipeline.i_csrs.n_mtvec_base_t0),
.i_pipeline__i_csrs__n_mtvec_mode(
  i_pipeline.i_csrs.n_mtvec_mode),
.i_pipeline__i_csrs__n_mtvec_mode_t0(
  i_pipeline.i_csrs.n_mtvec_mode_t0),
.i_pipeline__i_csrs__n_reg_lkgcfg(
  i_pipeline.i_csrs.n_reg_lkgcfg),
.i_pipeline__i_csrs__n_reg_lkgcfg_t0(
  i_pipeline.i_csrs.n_reg_lkgcfg_t0),
.i_pipeline__i_csrs__n_reg_mie(
  i_pipeline.i_csrs.n_reg_mie),
.i_pipeline__i_csrs__n_reg_mie_t0(
  i_pipeline.i_csrs.n_reg_mie_t0),
.i_pipeline__i_csrs__n_reg_mscratch(
  i_pipeline.i_csrs.n_reg_mscratch),
.i_pipeline__i_csrs__n_reg_mscratch_t0(
  i_pipeline.i_csrs.n_reg_mscratch_t0),
.i_pipeline__i_csrs__n_reg_mtval(
  i_pipeline.i_csrs.n_reg_mtval),
.i_pipeline__i_csrs__n_reg_mtval_t0(
  i_pipeline.i_csrs.n_reg_mtval_t0),
.i_pipeline__i_csrs__n_uxcrypto_b0(
  i_pipeline.i_csrs.n_uxcrypto_b0),
.i_pipeline__i_csrs__n_uxcrypto_b0_t0(
  i_pipeline.i_csrs.n_uxcrypto_b0_t0),
.i_pipeline__i_csrs__n_uxcrypto_b1(
  i_pipeline.i_csrs.n_uxcrypto_b1),
.i_pipeline__i_csrs__n_uxcrypto_b1_t0(
  i_pipeline.i_csrs.n_uxcrypto_b1_t0),
.i_pipeline__i_csrs__n_uxcrypto_ct(
  i_pipeline.i_csrs.n_uxcrypto_ct),
.i_pipeline__i_csrs__n_uxcrypto_ct_t0(
  i_pipeline.i_csrs.n_uxcrypto_ct_t0),
.i_pipeline__i_csrs__p_trap_int(
  i_pipeline.i_csrs.p_trap_int),
.i_pipeline__i_csrs__read_cycle(
  i_pipeline.i_csrs.read_cycle),
.i_pipeline__i_csrs__read_cycleh(
  i_pipeline.i_csrs.read_cycleh),
.i_pipeline__i_csrs__read_instret(
  i_pipeline.i_csrs.read_instret),
.i_pipeline__i_csrs__read_instreth(
  i_pipeline.i_csrs.read_instreth),
.i_pipeline__i_csrs__read_lkgcfg(
  i_pipeline.i_csrs.read_lkgcfg),
.i_pipeline__i_csrs__read_marchid(
  i_pipeline.i_csrs.read_marchid),
.i_pipeline__i_csrs__read_mcause(
  i_pipeline.i_csrs.read_mcause),
.i_pipeline__i_csrs__read_mcountin(
  i_pipeline.i_csrs.read_mcountin),
.i_pipeline__i_csrs__read_mcycle(
  i_pipeline.i_csrs.read_mcycle),
.i_pipeline__i_csrs__read_mcycleh(
  i_pipeline.i_csrs.read_mcycleh),
.i_pipeline__i_csrs__read_medeleg(
  i_pipeline.i_csrs.read_medeleg),
.i_pipeline__i_csrs__read_mepc(
  i_pipeline.i_csrs.read_mepc),
.i_pipeline__i_csrs__read_mhartid(
  i_pipeline.i_csrs.read_mhartid),
.i_pipeline__i_csrs__read_mideleg(
  i_pipeline.i_csrs.read_mideleg),
.i_pipeline__i_csrs__read_mie(
  i_pipeline.i_csrs.read_mie),
.i_pipeline__i_csrs__read_mimpid(
  i_pipeline.i_csrs.read_mimpid),
.i_pipeline__i_csrs__read_minstret(
  i_pipeline.i_csrs.read_minstret),
.i_pipeline__i_csrs__read_minstreth(
  i_pipeline.i_csrs.read_minstreth),
.i_pipeline__i_csrs__read_mip(
  i_pipeline.i_csrs.read_mip),
.i_pipeline__i_csrs__read_misa(
  i_pipeline.i_csrs.read_misa),
.i_pipeline__i_csrs__read_mscratch(
  i_pipeline.i_csrs.read_mscratch),
.i_pipeline__i_csrs__read_mstatus(
  i_pipeline.i_csrs.read_mstatus),
.i_pipeline__i_csrs__read_mtval(
  i_pipeline.i_csrs.read_mtval),
.i_pipeline__i_csrs__read_mtvec(
  i_pipeline.i_csrs.read_mtvec),
.i_pipeline__i_csrs__read_mvendorid(
  i_pipeline.i_csrs.read_mvendorid),
.i_pipeline__i_csrs__read_time(
  i_pipeline.i_csrs.read_time),
.i_pipeline__i_csrs__read_timeh(
  i_pipeline.i_csrs.read_timeh),
.i_pipeline__i_csrs__read_uxcrypto(
  i_pipeline.i_csrs.read_uxcrypto),
.i_pipeline__i_csrs__reg_mcause_cause(
  i_pipeline.i_csrs.reg_mcause_cause),
.i_pipeline__i_csrs__reg_mcause_cause_t0(
  i_pipeline.i_csrs.reg_mcause_cause_t0),
.i_pipeline__i_csrs__reg_mcause_interrupt(
  i_pipeline.i_csrs.reg_mcause_interrupt),
.i_pipeline__i_csrs__reg_mcause_interrupt_t0(
  i_pipeline.i_csrs.reg_mcause_interrupt_t0),
.i_pipeline__i_csrs__reg_mepc_mepc(
  i_pipeline.i_csrs.reg_mepc_mepc),
.i_pipeline__i_csrs__reg_mepc_mepc_t0(
  i_pipeline.i_csrs.reg_mepc_mepc_t0),
.i_pipeline__i_csrs__reg_mscratch(
  i_pipeline.i_csrs.reg_mscratch),
.i_pipeline__i_csrs__reg_mscratch_t0(
  i_pipeline.i_csrs.reg_mscratch_t0),
.i_pipeline__i_csrs__reg_mstatus_mpie(
  i_pipeline.i_csrs.reg_mstatus_mpie),
.i_pipeline__i_csrs__reg_mstatus_mpie_t0(
  i_pipeline.i_csrs.reg_mstatus_mpie_t0),
.i_pipeline__i_csrs__reg_mstatus_wpri1(
  i_pipeline.i_csrs.reg_mstatus_wpri1),
.i_pipeline__i_csrs__reg_mstatus_wpri1_t0(
  i_pipeline.i_csrs.reg_mstatus_wpri1_t0),
.i_pipeline__i_csrs__reg_mstatus_wpri2(
  i_pipeline.i_csrs.reg_mstatus_wpri2),
.i_pipeline__i_csrs__reg_mstatus_wpri2_t0(
  i_pipeline.i_csrs.reg_mstatus_wpri2_t0),
.i_pipeline__i_csrs__reg_mstatus_wpri3(
  i_pipeline.i_csrs.reg_mstatus_wpri3),
.i_pipeline__i_csrs__reg_mstatus_wpri3_t0(
  i_pipeline.i_csrs.reg_mstatus_wpri3_t0),
.i_pipeline__i_csrs__reg_mstatus_wpri4(
  i_pipeline.i_csrs.reg_mstatus_wpri4),
.i_pipeline__i_csrs__reg_mstatus_wpri4_t0(
  i_pipeline.i_csrs.reg_mstatus_wpri4_t0),
.i_pipeline__i_csrs__reg_mtval(
  i_pipeline.i_csrs.reg_mtval),
.i_pipeline__i_csrs__reg_mtval_t0(
  i_pipeline.i_csrs.reg_mtval_t0),
.i_pipeline__i_csrs__reg_mtvec_base(
  i_pipeline.i_csrs.reg_mtvec_base),
.i_pipeline__i_csrs__reg_mtvec_base_t0(
  i_pipeline.i_csrs.reg_mtvec_base_t0),
.i_pipeline__i_csrs__reg_mtvec_mode(
  i_pipeline.i_csrs.reg_mtvec_mode),
.i_pipeline__i_csrs__reg_mtvec_mode_t0(
  i_pipeline.i_csrs.reg_mtvec_mode_t0),
.i_pipeline__i_csrs__valid_addr(
  i_pipeline.i_csrs.valid_addr),
.i_pipeline__i_csrs__wen_lkgcfg(
  i_pipeline.i_csrs.wen_lkgcfg),
.i_pipeline__i_csrs__wen_mcause(
  i_pipeline.i_csrs.wen_mcause),
.i_pipeline__i_csrs__wen_mcountin(
  i_pipeline.i_csrs.wen_mcountin),
.i_pipeline__i_csrs__wen_mepc(
  i_pipeline.i_csrs.wen_mepc),
.i_pipeline__i_csrs__wen_mie(
  i_pipeline.i_csrs.wen_mie),
.i_pipeline__i_csrs__wen_mscratch(
  i_pipeline.i_csrs.wen_mscratch),
.i_pipeline__i_csrs__wen_mstatus(
  i_pipeline.i_csrs.wen_mstatus),
.i_pipeline__i_csrs__wen_mstatus_mie(
  i_pipeline.i_csrs.wen_mstatus_mie),
.i_pipeline__i_csrs__wen_mtval(
  i_pipeline.i_csrs.wen_mtval),
.i_pipeline__i_csrs__wen_mtvec(
  i_pipeline.i_csrs.wen_mtvec),
.i_pipeline__i_csrs__wen_uxcrypto(
  i_pipeline.i_csrs.wen_uxcrypto),
.i_pipeline__i_csrs__wen_valid_mcause(
  i_pipeline.i_csrs.wen_valid_mcause),
.i_pipeline__i_gprs__g_clk(
  i_pipeline.i_gprs.g_clk),
.i_pipeline__i_gprs__g_resetn(
  i_pipeline.i_gprs.g_resetn),
.i_pipeline__i_gprs__rs1_addr(
  i_pipeline.i_gprs.rs1_addr),
.i_pipeline__i_gprs__rs1_data(
  i_pipeline.i_gprs.rs1_data),
.i_pipeline__i_gprs__rs2_addr(
  i_pipeline.i_gprs.rs2_addr),
.i_pipeline__i_gprs__rs2_data(
  i_pipeline.i_gprs.rs2_data),
.i_pipeline__i_gprs__rs3_addr(
  i_pipeline.i_gprs.rs3_addr),
.i_pipeline__i_gprs__rs3_data(
  i_pipeline.i_gprs.rs3_data),
.i_pipeline__i_gprs__rd_wen(
  i_pipeline.i_gprs.rd_wen),
.i_pipeline__i_gprs__rd_wide(
  i_pipeline.i_gprs.rd_wide),
.i_pipeline__i_gprs__rd_addr(
  i_pipeline.i_gprs.rd_addr),
.i_pipeline__i_gprs__rd_wdata(
  i_pipeline.i_gprs.rd_wdata),
.i_pipeline__i_gprs__rd_wdata_hi(
  i_pipeline.i_gprs.rd_wdata_hi),
.i_pipeline__i_gprs__rs3_data_t0(
  i_pipeline.i_gprs.rs3_data_t0),
.i_pipeline__i_gprs__rs3_addr_t0(
  i_pipeline.i_gprs.rs3_addr_t0),
.i_pipeline__i_gprs__rs2_data_t0(
  i_pipeline.i_gprs.rs2_data_t0),
.i_pipeline__i_gprs__rs2_addr_t0(
  i_pipeline.i_gprs.rs2_addr_t0),
.i_pipeline__i_gprs__rs1_data_t0(
  i_pipeline.i_gprs.rs1_data_t0),
.i_pipeline__i_gprs__rs1_addr_t0(
  i_pipeline.i_gprs.rs1_addr_t0),
.i_pipeline__i_gprs__rd_wide_t0(
  i_pipeline.i_gprs.rd_wide_t0),
.i_pipeline__i_gprs__rd_wen_t0(
  i_pipeline.i_gprs.rd_wen_t0),
.i_pipeline__i_gprs__rd_wdata_hi_t0(
  i_pipeline.i_gprs.rd_wdata_hi_t0),
.i_pipeline__i_gprs__rd_wdata_t0(
  i_pipeline.i_gprs.rd_wdata_t0),
.i_pipeline__i_gprs__rd_addr_t0(
  i_pipeline.i_gprs.rd_addr_t0),
.i_pipeline__i_gprs__gprs_10_(
  i_pipeline.i_gprs.\gprs[10] ),
.i_pipeline__i_gprs__gprs_10__t0(
  i_pipeline.i_gprs.\gprs[10]_t0 ),
.i_pipeline__i_gprs__gprs_11_(
  i_pipeline.i_gprs.\gprs[11] ),
.i_pipeline__i_gprs__gprs_11__t0(
  i_pipeline.i_gprs.\gprs[11]_t0 ),
.i_pipeline__i_gprs__gprs_12_(
  i_pipeline.i_gprs.\gprs[12] ),
.i_pipeline__i_gprs__gprs_12__t0(
  i_pipeline.i_gprs.\gprs[12]_t0 ),
.i_pipeline__i_gprs__gprs_13_(
  i_pipeline.i_gprs.\gprs[13] ),
.i_pipeline__i_gprs__gprs_13__t0(
  i_pipeline.i_gprs.\gprs[13]_t0 ),
.i_pipeline__i_gprs__gprs_14_(
  i_pipeline.i_gprs.\gprs[14] ),
.i_pipeline__i_gprs__gprs_14__t0(
  i_pipeline.i_gprs.\gprs[14]_t0 ),
.i_pipeline__i_gprs__gprs_15_(
  i_pipeline.i_gprs.\gprs[15] ),
.i_pipeline__i_gprs__gprs_15__t0(
  i_pipeline.i_gprs.\gprs[15]_t0 ),
.i_pipeline__i_gprs__gprs_16_(
  i_pipeline.i_gprs.\gprs[16] ),
.i_pipeline__i_gprs__gprs_16__t0(
  i_pipeline.i_gprs.\gprs[16]_t0 ),
.i_pipeline__i_gprs__gprs_17_(
  i_pipeline.i_gprs.\gprs[17] ),
.i_pipeline__i_gprs__gprs_17__t0(
  i_pipeline.i_gprs.\gprs[17]_t0 ),
.i_pipeline__i_gprs__gprs_18_(
  i_pipeline.i_gprs.\gprs[18] ),
.i_pipeline__i_gprs__gprs_18__t0(
  i_pipeline.i_gprs.\gprs[18]_t0 ),
.i_pipeline__i_gprs__gprs_19_(
  i_pipeline.i_gprs.\gprs[19] ),
.i_pipeline__i_gprs__gprs_19__t0(
  i_pipeline.i_gprs.\gprs[19]_t0 ),
.i_pipeline__i_gprs__gprs_1_(
  i_pipeline.i_gprs.\gprs[1] ),
.i_pipeline__i_gprs__gprs_1__t0(
  i_pipeline.i_gprs.\gprs[1]_t0 ),
.i_pipeline__i_gprs__gprs_20_(
  i_pipeline.i_gprs.\gprs[20] ),
.i_pipeline__i_gprs__gprs_20__t0(
  i_pipeline.i_gprs.\gprs[20]_t0 ),
.i_pipeline__i_gprs__gprs_21_(
  i_pipeline.i_gprs.\gprs[21] ),
.i_pipeline__i_gprs__gprs_21__t0(
  i_pipeline.i_gprs.\gprs[21]_t0 ),
.i_pipeline__i_gprs__gprs_22_(
  i_pipeline.i_gprs.\gprs[22] ),
.i_pipeline__i_gprs__gprs_22__t0(
  i_pipeline.i_gprs.\gprs[22]_t0 ),
.i_pipeline__i_gprs__gprs_23_(
  i_pipeline.i_gprs.\gprs[23] ),
.i_pipeline__i_gprs__gprs_23__t0(
  i_pipeline.i_gprs.\gprs[23]_t0 ),
.i_pipeline__i_gprs__gprs_24_(
  i_pipeline.i_gprs.\gprs[24] ),
.i_pipeline__i_gprs__gprs_24__t0(
  i_pipeline.i_gprs.\gprs[24]_t0 ),
.i_pipeline__i_gprs__gprs_25_(
  i_pipeline.i_gprs.\gprs[25] ),
.i_pipeline__i_gprs__gprs_25__t0(
  i_pipeline.i_gprs.\gprs[25]_t0 ),
.i_pipeline__i_gprs__gprs_26_(
  i_pipeline.i_gprs.\gprs[26] ),
.i_pipeline__i_gprs__gprs_26__t0(
  i_pipeline.i_gprs.\gprs[26]_t0 ),
.i_pipeline__i_gprs__gprs_27_(
  i_pipeline.i_gprs.\gprs[27] ),
.i_pipeline__i_gprs__gprs_27__t0(
  i_pipeline.i_gprs.\gprs[27]_t0 ),
.i_pipeline__i_gprs__gprs_28_(
  i_pipeline.i_gprs.\gprs[28] ),
.i_pipeline__i_gprs__gprs_28__t0(
  i_pipeline.i_gprs.\gprs[28]_t0 ),
.i_pipeline__i_gprs__gprs_29_(
  i_pipeline.i_gprs.\gprs[29] ),
.i_pipeline__i_gprs__gprs_29__t0(
  i_pipeline.i_gprs.\gprs[29]_t0 ),
.i_pipeline__i_gprs__gprs_2_(
  i_pipeline.i_gprs.\gprs[2] ),
.i_pipeline__i_gprs__gprs_2__t0(
  i_pipeline.i_gprs.\gprs[2]_t0 ),
.i_pipeline__i_gprs__gprs_30_(
  i_pipeline.i_gprs.\gprs[30] ),
.i_pipeline__i_gprs__gprs_30__t0(
  i_pipeline.i_gprs.\gprs[30]_t0 ),
.i_pipeline__i_gprs__gprs_31_(
  i_pipeline.i_gprs.\gprs[31] ),
.i_pipeline__i_gprs__gprs_31__t0(
  i_pipeline.i_gprs.\gprs[31]_t0 ),
.i_pipeline__i_gprs__gprs_3_(
  i_pipeline.i_gprs.\gprs[3] ),
.i_pipeline__i_gprs__gprs_3__t0(
  i_pipeline.i_gprs.\gprs[3]_t0 ),
.i_pipeline__i_gprs__gprs_4_(
  i_pipeline.i_gprs.\gprs[4] ),
.i_pipeline__i_gprs__gprs_4__t0(
  i_pipeline.i_gprs.\gprs[4]_t0 ),
.i_pipeline__i_gprs__gprs_5_(
  i_pipeline.i_gprs.\gprs[5] ),
.i_pipeline__i_gprs__gprs_5__t0(
  i_pipeline.i_gprs.\gprs[5]_t0 ),
.i_pipeline__i_gprs__gprs_6_(
  i_pipeline.i_gprs.\gprs[6] ),
.i_pipeline__i_gprs__gprs_6__t0(
  i_pipeline.i_gprs.\gprs[6]_t0 ),
.i_pipeline__i_gprs__gprs_7_(
  i_pipeline.i_gprs.\gprs[7] ),
.i_pipeline__i_gprs__gprs_7__t0(
  i_pipeline.i_gprs.\gprs[7]_t0 ),
.i_pipeline__i_gprs__gprs_8_(
  i_pipeline.i_gprs.\gprs[8] ),
.i_pipeline__i_gprs__gprs_8__t0(
  i_pipeline.i_gprs.\gprs[8]_t0 ),
.i_pipeline__i_gprs__gprs_9_(
  i_pipeline.i_gprs.\gprs[9] ),
.i_pipeline__i_gprs__gprs_9__t0(
  i_pipeline.i_gprs.\gprs[9]_t0 ),
.i_pipeline__i_gprs__rd_even(
  i_pipeline.i_gprs.rd_even),
.i_pipeline__i_gprs__rd_wdata_odd(
  i_pipeline.i_gprs.rd_wdata_odd),
.i_pipeline__i_gprs__rd_wdata_odd_t0(
  i_pipeline.i_gprs.rd_wdata_odd_t0),
.i_pipeline__i_gprs__rd_wen_even(
  i_pipeline.i_gprs.rd_wen_even),
.i_pipeline__i_gprs__rd_wen_odd(
  i_pipeline.i_gprs.rd_wen_odd),
.i_pipeline__i_pipeline_s0_fetch__g_clk(
  i_pipeline.i_pipeline_s0_fetch.g_clk),
.i_pipeline__i_pipeline_s0_fetch__g_resetn(
  i_pipeline.i_pipeline_s0_fetch.g_resetn),
.i_pipeline__i_pipeline_s0_fetch__cf_req(
  i_pipeline.i_pipeline_s0_fetch.cf_req),
.i_pipeline__i_pipeline_s0_fetch__cf_target(
  i_pipeline.i_pipeline_s0_fetch.cf_target),
.i_pipeline__i_pipeline_s0_fetch__cf_ack(
  i_pipeline.i_pipeline_s0_fetch.cf_ack),
.i_pipeline__i_pipeline_s0_fetch__imem_req(
  i_pipeline.i_pipeline_s0_fetch.imem_req),
.i_pipeline__i_pipeline_s0_fetch__imem_wen(
  i_pipeline.i_pipeline_s0_fetch.imem_wen),
.i_pipeline__i_pipeline_s0_fetch__imem_strb(
  i_pipeline.i_pipeline_s0_fetch.imem_strb),
.i_pipeline__i_pipeline_s0_fetch__imem_wdata(
  i_pipeline.i_pipeline_s0_fetch.imem_wdata),
.i_pipeline__i_pipeline_s0_fetch__imem_addr(
  i_pipeline.i_pipeline_s0_fetch.imem_addr),
.i_pipeline__i_pipeline_s0_fetch__imem_gnt(
  i_pipeline.i_pipeline_s0_fetch.imem_gnt),
.i_pipeline__i_pipeline_s0_fetch__imem_ack(
  i_pipeline.i_pipeline_s0_fetch.imem_ack),
.i_pipeline__i_pipeline_s0_fetch__imem_recv(
  i_pipeline.i_pipeline_s0_fetch.imem_recv),
.i_pipeline__i_pipeline_s0_fetch__imem_error(
  i_pipeline.i_pipeline_s0_fetch.imem_error),
.i_pipeline__i_pipeline_s0_fetch__imem_rdata(
  i_pipeline.i_pipeline_s0_fetch.imem_rdata),
.i_pipeline__i_pipeline_s0_fetch__s0_flush(
  i_pipeline.i_pipeline_s0_fetch.s0_flush),
.i_pipeline__i_pipeline_s0_fetch__s1_busy(
  i_pipeline.i_pipeline_s0_fetch.s1_busy),
.i_pipeline__i_pipeline_s0_fetch__s1_valid(
  i_pipeline.i_pipeline_s0_fetch.s1_valid),
.i_pipeline__i_pipeline_s0_fetch__s1_data(
  i_pipeline.i_pipeline_s0_fetch.s1_data),
.i_pipeline__i_pipeline_s0_fetch__s1_error(
  i_pipeline.i_pipeline_s0_fetch.s1_error),
.i_pipeline__i_pipeline_s0_fetch__s1_valid_t0(
  i_pipeline.i_pipeline_s0_fetch.s1_valid_t0),
.i_pipeline__i_pipeline_s0_fetch__s1_error_t0(
  i_pipeline.i_pipeline_s0_fetch.s1_error_t0),
.i_pipeline__i_pipeline_s0_fetch__s1_data_t0(
  i_pipeline.i_pipeline_s0_fetch.s1_data_t0),
.i_pipeline__i_pipeline_s0_fetch__s1_busy_t0(
  i_pipeline.i_pipeline_s0_fetch.s1_busy_t0),
.i_pipeline__i_pipeline_s0_fetch__s0_flush_t0(
  i_pipeline.i_pipeline_s0_fetch.s0_flush_t0),
.i_pipeline__i_pipeline_s0_fetch__imem_wen_t0(
  i_pipeline.i_pipeline_s0_fetch.imem_wen_t0),
.i_pipeline__i_pipeline_s0_fetch__imem_wdata_t0(
  i_pipeline.i_pipeline_s0_fetch.imem_wdata_t0),
.i_pipeline__i_pipeline_s0_fetch__imem_strb_t0(
  i_pipeline.i_pipeline_s0_fetch.imem_strb_t0),
.i_pipeline__i_pipeline_s0_fetch__imem_req_t0(
  i_pipeline.i_pipeline_s0_fetch.imem_req_t0),
.i_pipeline__i_pipeline_s0_fetch__imem_recv_t0(
  i_pipeline.i_pipeline_s0_fetch.imem_recv_t0),
.i_pipeline__i_pipeline_s0_fetch__imem_rdata_t0(
  i_pipeline.i_pipeline_s0_fetch.imem_rdata_t0),
.i_pipeline__i_pipeline_s0_fetch__imem_gnt_t0(
  i_pipeline.i_pipeline_s0_fetch.imem_gnt_t0),
.i_pipeline__i_pipeline_s0_fetch__imem_error_t0(
  i_pipeline.i_pipeline_s0_fetch.imem_error_t0),
.i_pipeline__i_pipeline_s0_fetch__imem_addr_t0(
  i_pipeline.i_pipeline_s0_fetch.imem_addr_t0),
.i_pipeline__i_pipeline_s0_fetch__imem_ack_t0(
  i_pipeline.i_pipeline_s0_fetch.imem_ack_t0),
.i_pipeline__i_pipeline_s0_fetch__cf_target_t0(
  i_pipeline.i_pipeline_s0_fetch.cf_target_t0),
.i_pipeline__i_pipeline_s0_fetch__cf_req_t0(
  i_pipeline.i_pipeline_s0_fetch.cf_req_t0),
.i_pipeline__i_pipeline_s0_fetch__cf_ack_t0(
  i_pipeline.i_pipeline_s0_fetch.cf_ack_t0),
.i_pipeline__i_pipeline_s0_fetch__allow_new_mem_req(
  i_pipeline.i_pipeline_s0_fetch.allow_new_mem_req),
.i_pipeline__i_pipeline_s0_fetch__buf_16(
  i_pipeline.i_pipeline_s0_fetch.buf_16),
.i_pipeline__i_pipeline_s0_fetch__buf_16_t0(
  i_pipeline.i_pipeline_s0_fetch.buf_16_t0),
.i_pipeline__i_pipeline_s0_fetch__buf_32(
  i_pipeline.i_pipeline_s0_fetch.buf_32),
.i_pipeline__i_pipeline_s0_fetch__buf_32_t0(
  i_pipeline.i_pipeline_s0_fetch.buf_32_t0),
.i_pipeline__i_pipeline_s0_fetch__buf_depth(
  i_pipeline.i_pipeline_s0_fetch.buf_depth),
.i_pipeline__i_pipeline_s0_fetch__buf_depth_t0(
  i_pipeline.i_pipeline_s0_fetch.buf_depth_t0),
.i_pipeline__i_pipeline_s0_fetch__buf_out_2(
  i_pipeline.i_pipeline_s0_fetch.buf_out_2),
.i_pipeline__i_pipeline_s0_fetch__buf_out_2_t0(
  i_pipeline.i_pipeline_s0_fetch.buf_out_2_t0),
.i_pipeline__i_pipeline_s0_fetch__buf_out_4(
  i_pipeline.i_pipeline_s0_fetch.buf_out_4),
.i_pipeline__i_pipeline_s0_fetch__buf_out_4_t0(
  i_pipeline.i_pipeline_s0_fetch.buf_out_4_t0),
.i_pipeline__i_pipeline_s0_fetch__buf_ready(
  i_pipeline.i_pipeline_s0_fetch.buf_ready),
.i_pipeline__i_pipeline_s0_fetch__cf_change(
  i_pipeline.i_pipeline_s0_fetch.cf_change),
.i_pipeline__i_pipeline_s0_fetch__drop_response(
  i_pipeline.i_pipeline_s0_fetch.drop_response),
.i_pipeline__i_pipeline_s0_fetch__f_2byte(
  i_pipeline.i_pipeline_s0_fetch.f_2byte),
.i_pipeline__i_pipeline_s0_fetch__f_4byte(
  i_pipeline.i_pipeline_s0_fetch.f_4byte),
.i_pipeline__i_pipeline_s0_fetch__fetch_misaligned(
  i_pipeline.i_pipeline_s0_fetch.fetch_misaligned),
.i_pipeline__i_pipeline_s0_fetch__ignore_rsps(
  i_pipeline.i_pipeline_s0_fetch.ignore_rsps),
.i_pipeline__i_pipeline_s0_fetch__incomplete_instr(
  i_pipeline.i_pipeline_s0_fetch.incomplete_instr),
.i_pipeline__i_pipeline_s0_fetch__n_fetch_misaligned(
  i_pipeline.i_pipeline_s0_fetch.n_fetch_misaligned),
.i_pipeline__i_pipeline_s0_fetch__n_ignore_rsps(
  i_pipeline.i_pipeline_s0_fetch.n_ignore_rsps),
.i_pipeline__i_pipeline_s0_fetch__n_imem_addr(
  i_pipeline.i_pipeline_s0_fetch.n_imem_addr),
.i_pipeline__i_pipeline_s0_fetch__n_imem_addr_t0(
  i_pipeline.i_pipeline_s0_fetch.n_imem_addr_t0),
.i_pipeline__i_pipeline_s0_fetch__n_imem_req(
  i_pipeline.i_pipeline_s0_fetch.n_imem_req),
.i_pipeline__i_pipeline_s0_fetch__n_reqs_outstanding(
  i_pipeline.i_pipeline_s0_fetch.n_reqs_outstanding),
.i_pipeline__i_pipeline_s0_fetch__new_mem_req(
  i_pipeline.i_pipeline_s0_fetch.new_mem_req),
.i_pipeline__i_pipeline_s0_fetch__progress_imem_addr(
  i_pipeline.i_pipeline_s0_fetch.progress_imem_addr),
.i_pipeline__i_pipeline_s0_fetch__reqs_outstanding(
  i_pipeline.i_pipeline_s0_fetch.reqs_outstanding),
.i_pipeline__i_pipeline_s0_fetch__rsp_recv(
  i_pipeline.i_pipeline_s0_fetch.rsp_recv),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__g_clk(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.g_clk),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__g_resetn(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.g_resetn),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__flush(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.flush),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_4byte(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.f_4byte),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_2byte(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.f_2byte),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_err(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.f_err),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_in(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.f_in),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_ready(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.f_ready),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_depth(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_depth),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_16(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_16),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_32(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_32),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_out),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out_2(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_out_2),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out_4(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_out_4),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_err(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_err),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_valid(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_valid),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_ready(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_ready),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__flush_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.flush_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_ready_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.f_ready_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_in_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.f_in_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_err_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.f_err_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_4byte_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.f_4byte_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_2byte_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.f_2byte_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_valid_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_valid_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_ready_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_ready_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out_4_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_out_4_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out_2_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_out_2_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_out_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_err_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_err_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_depth_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_depth_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_32_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_32_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_16_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buf_16_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buffer(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buffer),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buffer_err(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buffer_err),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buffer_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.buffer_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__eat_2(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.eat_2),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__eat_4(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.eat_4),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__insert_at(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.insert_at),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_bdepth(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.n_bdepth),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_bdepth_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.n_bdepth_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.n_buffer),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_d(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.n_buffer_d),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_d_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.n_buffer_d_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_err(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.n_buffer_err),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_or_in(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.n_buffer_or_in),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_or_in_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.n_buffer_or_in_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_shf_out(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.n_buffer_shf_out),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_shf_out_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.n_buffer_shf_out_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_t0(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.n_buffer_t0),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_err_in(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.n_err_in),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_err_or_in(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.n_err_or_in),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_err_shf_out(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.n_err_shf_out),
.i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__update_buffer(
  i_pipeline.i_pipeline_s0_fetch.i_core_fetch_buffer.update_buffer),
.i_pipeline__i_pipeline_s1_decode__g_clk(
  i_pipeline.i_pipeline_s1_decode.g_clk),
.i_pipeline__i_pipeline_s1_decode__g_resetn(
  i_pipeline.i_pipeline_s1_decode.g_resetn),
.i_pipeline__i_pipeline_s1_decode__s1_valid(
  i_pipeline.i_pipeline_s1_decode.s1_valid),
.i_pipeline__i_pipeline_s1_decode__s1_busy(
  i_pipeline.i_pipeline_s1_decode.s1_busy),
.i_pipeline__i_pipeline_s1_decode__s1_data(
  i_pipeline.i_pipeline_s1_decode.s1_data),
.i_pipeline__i_pipeline_s1_decode__s1_error(
  i_pipeline.i_pipeline_s1_decode.s1_error),
.i_pipeline__i_pipeline_s1_decode__s1_flush(
  i_pipeline.i_pipeline_s1_decode.s1_flush),
.i_pipeline__i_pipeline_s1_decode__s1_bubble(
  i_pipeline.i_pipeline_s1_decode.s1_bubble),
.i_pipeline__i_pipeline_s1_decode__s1_rs1_addr(
  i_pipeline.i_pipeline_s1_decode.s1_rs1_addr),
.i_pipeline__i_pipeline_s1_decode__s1_rs2_addr(
  i_pipeline.i_pipeline_s1_decode.s1_rs2_addr),
.i_pipeline__i_pipeline_s1_decode__s1_rs3_addr(
  i_pipeline.i_pipeline_s1_decode.s1_rs3_addr),
.i_pipeline__i_pipeline_s1_decode__s1_rs1_rdata(
  i_pipeline.i_pipeline_s1_decode.s1_rs1_rdata),
.i_pipeline__i_pipeline_s1_decode__s1_rs2_rdata(
  i_pipeline.i_pipeline_s1_decode.s1_rs2_rdata),
.i_pipeline__i_pipeline_s1_decode__s1_rs3_rdata(
  i_pipeline.i_pipeline_s1_decode.s1_rs3_rdata),
.i_pipeline__i_pipeline_s1_decode__leak_prng(
  i_pipeline.i_pipeline_s1_decode.leak_prng),
.i_pipeline__i_pipeline_s1_decode__leak_lkgcfg(
  i_pipeline.i_pipeline_s1_decode.leak_lkgcfg),
.i_pipeline__i_pipeline_s1_decode__s1_leak_fence(
  i_pipeline.i_pipeline_s1_decode.s1_leak_fence),
.i_pipeline__i_pipeline_s1_decode__cf_req(
  i_pipeline.i_pipeline_s1_decode.cf_req),
.i_pipeline__i_pipeline_s1_decode__cf_target(
  i_pipeline.i_pipeline_s1_decode.cf_target),
.i_pipeline__i_pipeline_s1_decode__cf_ack(
  i_pipeline.i_pipeline_s1_decode.cf_ack),
.i_pipeline__i_pipeline_s1_decode__s2_valid(
  i_pipeline.i_pipeline_s1_decode.s2_valid),
.i_pipeline__i_pipeline_s1_decode__s2_busy(
  i_pipeline.i_pipeline_s1_decode.s2_busy),
.i_pipeline__i_pipeline_s1_decode__s2_rd(
  i_pipeline.i_pipeline_s1_decode.s2_rd),
.i_pipeline__i_pipeline_s1_decode__s2_opr_a(
  i_pipeline.i_pipeline_s1_decode.s2_opr_a),
.i_pipeline__i_pipeline_s1_decode__s2_opr_b(
  i_pipeline.i_pipeline_s1_decode.s2_opr_b),
.i_pipeline__i_pipeline_s1_decode__s2_opr_c(
  i_pipeline.i_pipeline_s1_decode.s2_opr_c),
.i_pipeline__i_pipeline_s1_decode__s2_uop(
  i_pipeline.i_pipeline_s1_decode.s2_uop),
.i_pipeline__i_pipeline_s1_decode__s2_fu(
  i_pipeline.i_pipeline_s1_decode.s2_fu),
.i_pipeline__i_pipeline_s1_decode__s2_pw(
  i_pipeline.i_pipeline_s1_decode.s2_pw),
.i_pipeline__i_pipeline_s1_decode__s2_trap(
  i_pipeline.i_pipeline_s1_decode.s2_trap),
.i_pipeline__i_pipeline_s1_decode__s2_size(
  i_pipeline.i_pipeline_s1_decode.s2_size),
.i_pipeline__i_pipeline_s1_decode__s2_instr(
  i_pipeline.i_pipeline_s1_decode.s2_instr),
.i_pipeline__i_pipeline_s1_decode__s2_valid_t0(
  i_pipeline.i_pipeline_s1_decode.s2_valid_t0),
.i_pipeline__i_pipeline_s1_decode__s2_uop_t0(
  i_pipeline.i_pipeline_s1_decode.s2_uop_t0),
.i_pipeline__i_pipeline_s1_decode__s2_trap_t0(
  i_pipeline.i_pipeline_s1_decode.s2_trap_t0),
.i_pipeline__i_pipeline_s1_decode__s2_size_t0(
  i_pipeline.i_pipeline_s1_decode.s2_size_t0),
.i_pipeline__i_pipeline_s1_decode__s2_rd_t0(
  i_pipeline.i_pipeline_s1_decode.s2_rd_t0),
.i_pipeline__i_pipeline_s1_decode__s2_pw_t0(
  i_pipeline.i_pipeline_s1_decode.s2_pw_t0),
.i_pipeline__i_pipeline_s1_decode__s2_opr_c_t0(
  i_pipeline.i_pipeline_s1_decode.s2_opr_c_t0),
.i_pipeline__i_pipeline_s1_decode__s2_opr_b_t0(
  i_pipeline.i_pipeline_s1_decode.s2_opr_b_t0),
.i_pipeline__i_pipeline_s1_decode__s2_opr_a_t0(
  i_pipeline.i_pipeline_s1_decode.s2_opr_a_t0),
.i_pipeline__i_pipeline_s1_decode__s2_instr_t0(
  i_pipeline.i_pipeline_s1_decode.s2_instr_t0),
.i_pipeline__i_pipeline_s1_decode__s2_fu_t0(
  i_pipeline.i_pipeline_s1_decode.s2_fu_t0),
.i_pipeline__i_pipeline_s1_decode__s2_busy_t0(
  i_pipeline.i_pipeline_s1_decode.s2_busy_t0),
.i_pipeline__i_pipeline_s1_decode__s1_rs3_rdata_t0(
  i_pipeline.i_pipeline_s1_decode.s1_rs3_rdata_t0),
.i_pipeline__i_pipeline_s1_decode__s1_rs3_addr_t0(
  i_pipeline.i_pipeline_s1_decode.s1_rs3_addr_t0),
.i_pipeline__i_pipeline_s1_decode__s1_rs2_rdata_t0(
  i_pipeline.i_pipeline_s1_decode.s1_rs2_rdata_t0),
.i_pipeline__i_pipeline_s1_decode__s1_rs2_addr_t0(
  i_pipeline.i_pipeline_s1_decode.s1_rs2_addr_t0),
.i_pipeline__i_pipeline_s1_decode__s1_rs1_rdata_t0(
  i_pipeline.i_pipeline_s1_decode.s1_rs1_rdata_t0),
.i_pipeline__i_pipeline_s1_decode__s1_rs1_addr_t0(
  i_pipeline.i_pipeline_s1_decode.s1_rs1_addr_t0),
.i_pipeline__i_pipeline_s1_decode__s1_leak_fence_t0(
  i_pipeline.i_pipeline_s1_decode.s1_leak_fence_t0),
.i_pipeline__i_pipeline_s1_decode__s1_flush_t0(
  i_pipeline.i_pipeline_s1_decode.s1_flush_t0),
.i_pipeline__i_pipeline_s1_decode__s1_bubble_t0(
  i_pipeline.i_pipeline_s1_decode.s1_bubble_t0),
.i_pipeline__i_pipeline_s1_decode__leak_lkgcfg_t0(
  i_pipeline.i_pipeline_s1_decode.leak_lkgcfg_t0),
.i_pipeline__i_pipeline_s1_decode__leak_prng_t0(
  i_pipeline.i_pipeline_s1_decode.leak_prng_t0),
.i_pipeline__i_pipeline_s1_decode__s1_valid_t0(
  i_pipeline.i_pipeline_s1_decode.s1_valid_t0),
.i_pipeline__i_pipeline_s1_decode__s1_error_t0(
  i_pipeline.i_pipeline_s1_decode.s1_error_t0),
.i_pipeline__i_pipeline_s1_decode__s1_data_t0(
  i_pipeline.i_pipeline_s1_decode.s1_data_t0),
.i_pipeline__i_pipeline_s1_decode__s1_busy_t0(
  i_pipeline.i_pipeline_s1_decode.s1_busy_t0),
.i_pipeline__i_pipeline_s1_decode__cf_target_t0(
  i_pipeline.i_pipeline_s1_decode.cf_target_t0),
.i_pipeline__i_pipeline_s1_decode__cf_req_t0(
  i_pipeline.i_pipeline_s1_decode.cf_req_t0),
.i_pipeline__i_pipeline_s1_decode__cf_ack_t0(
  i_pipeline.i_pipeline_s1_decode.cf_ack_t0),
.i_pipeline__i_pipeline_s1_decode__bubble_fu(
  i_pipeline.i_pipeline_s1_decode.bubble_fu),
.i_pipeline__i_pipeline_s1_decode__bubble_uop(
  i_pipeline.i_pipeline_s1_decode.bubble_uop),
.i_pipeline__i_pipeline_s1_decode__cfu_no_rd(
  i_pipeline.i_pipeline_s1_decode.cfu_no_rd),
.i_pipeline__i_pipeline_s1_decode__clr_rd_lsb(
  i_pipeline.i_pipeline_s1_decode.clr_rd_lsb),
.i_pipeline__i_pipeline_s1_decode__csr_no_read(
  i_pipeline.i_pipeline_s1_decode.csr_no_read),
.i_pipeline__i_pipeline_s1_decode__csr_no_write(
  i_pipeline.i_pipeline_s1_decode.csr_no_write),
.i_pipeline__i_pipeline_s1_decode__csr_op(
  i_pipeline.i_pipeline_s1_decode.csr_op),
.i_pipeline__i_pipeline_s1_decode__dec_add(
  i_pipeline.i_pipeline_s1_decode.dec_add),
.i_pipeline__i_pipeline_s1_decode__dec_addi(
  i_pipeline.i_pipeline_s1_decode.dec_addi),
.i_pipeline__i_pipeline_s1_decode__dec_and(
  i_pipeline.i_pipeline_s1_decode.dec_and),
.i_pipeline__i_pipeline_s1_decode__dec_andi(
  i_pipeline.i_pipeline_s1_decode.dec_andi),
.i_pipeline__i_pipeline_s1_decode__dec_auipc(
  i_pipeline.i_pipeline_s1_decode.dec_auipc),
.i_pipeline__i_pipeline_s1_decode__dec_b_bdep(
  i_pipeline.i_pipeline_s1_decode.dec_b_bdep),
.i_pipeline__i_pipeline_s1_decode__dec_b_bext(
  i_pipeline.i_pipeline_s1_decode.dec_b_bext),
.i_pipeline__i_pipeline_s1_decode__dec_b_clmul(
  i_pipeline.i_pipeline_s1_decode.dec_b_clmul),
.i_pipeline__i_pipeline_s1_decode__dec_b_clmulh(
  i_pipeline.i_pipeline_s1_decode.dec_b_clmulh),
.i_pipeline__i_pipeline_s1_decode__dec_b_clmulr(
  i_pipeline.i_pipeline_s1_decode.dec_b_clmulr),
.i_pipeline__i_pipeline_s1_decode__dec_b_cmov(
  i_pipeline.i_pipeline_s1_decode.dec_b_cmov),
.i_pipeline__i_pipeline_s1_decode__dec_b_fsl(
  i_pipeline.i_pipeline_s1_decode.dec_b_fsl),
.i_pipeline__i_pipeline_s1_decode__dec_b_fsr(
  i_pipeline.i_pipeline_s1_decode.dec_b_fsr),
.i_pipeline__i_pipeline_s1_decode__dec_b_fsri(
  i_pipeline.i_pipeline_s1_decode.dec_b_fsri),
.i_pipeline__i_pipeline_s1_decode__dec_b_grev(
  i_pipeline.i_pipeline_s1_decode.dec_b_grev),
.i_pipeline__i_pipeline_s1_decode__dec_b_grevi(
  i_pipeline.i_pipeline_s1_decode.dec_b_grevi),
.i_pipeline__i_pipeline_s1_decode__dec_b_ror(
  i_pipeline.i_pipeline_s1_decode.dec_b_ror),
.i_pipeline__i_pipeline_s1_decode__dec_b_rori(
  i_pipeline.i_pipeline_s1_decode.dec_b_rori),
.i_pipeline__i_pipeline_s1_decode__dec_beq(
  i_pipeline.i_pipeline_s1_decode.dec_beq),
.i_pipeline__i_pipeline_s1_decode__dec_bge(
  i_pipeline.i_pipeline_s1_decode.dec_bge),
.i_pipeline__i_pipeline_s1_decode__dec_bgeu(
  i_pipeline.i_pipeline_s1_decode.dec_bgeu),
.i_pipeline__i_pipeline_s1_decode__dec_blt(
  i_pipeline.i_pipeline_s1_decode.dec_blt),
.i_pipeline__i_pipeline_s1_decode__dec_bltu(
  i_pipeline.i_pipeline_s1_decode.dec_bltu),
.i_pipeline__i_pipeline_s1_decode__dec_bne(
  i_pipeline.i_pipeline_s1_decode.dec_bne),
.i_pipeline__i_pipeline_s1_decode__dec_c_add(
  i_pipeline.i_pipeline_s1_decode.dec_c_add),
.i_pipeline__i_pipeline_s1_decode__dec_c_addi(
  i_pipeline.i_pipeline_s1_decode.dec_c_addi),
.i_pipeline__i_pipeline_s1_decode__dec_c_addi16sp(
  i_pipeline.i_pipeline_s1_decode.dec_c_addi16sp),
.i_pipeline__i_pipeline_s1_decode__dec_c_addi4spn(
  i_pipeline.i_pipeline_s1_decode.dec_c_addi4spn),
.i_pipeline__i_pipeline_s1_decode__dec_c_and(
  i_pipeline.i_pipeline_s1_decode.dec_c_and),
.i_pipeline__i_pipeline_s1_decode__dec_c_andi(
  i_pipeline.i_pipeline_s1_decode.dec_c_andi),
.i_pipeline__i_pipeline_s1_decode__dec_c_beqz(
  i_pipeline.i_pipeline_s1_decode.dec_c_beqz),
.i_pipeline__i_pipeline_s1_decode__dec_c_bnez(
  i_pipeline.i_pipeline_s1_decode.dec_c_bnez),
.i_pipeline__i_pipeline_s1_decode__dec_c_ebreak(
  i_pipeline.i_pipeline_s1_decode.dec_c_ebreak),
.i_pipeline__i_pipeline_s1_decode__dec_c_j(
  i_pipeline.i_pipeline_s1_decode.dec_c_j),
.i_pipeline__i_pipeline_s1_decode__dec_c_jal(
  i_pipeline.i_pipeline_s1_decode.dec_c_jal),
.i_pipeline__i_pipeline_s1_decode__dec_c_jalr(
  i_pipeline.i_pipeline_s1_decode.dec_c_jalr),
.i_pipeline__i_pipeline_s1_decode__dec_c_jr(
  i_pipeline.i_pipeline_s1_decode.dec_c_jr),
.i_pipeline__i_pipeline_s1_decode__dec_c_li(
  i_pipeline.i_pipeline_s1_decode.dec_c_li),
.i_pipeline__i_pipeline_s1_decode__dec_c_lui(
  i_pipeline.i_pipeline_s1_decode.dec_c_lui),
.i_pipeline__i_pipeline_s1_decode__dec_c_lw(
  i_pipeline.i_pipeline_s1_decode.dec_c_lw),
.i_pipeline__i_pipeline_s1_decode__dec_c_lwsp(
  i_pipeline.i_pipeline_s1_decode.dec_c_lwsp),
.i_pipeline__i_pipeline_s1_decode__dec_c_mv(
  i_pipeline.i_pipeline_s1_decode.dec_c_mv),
.i_pipeline__i_pipeline_s1_decode__dec_c_nop(
  i_pipeline.i_pipeline_s1_decode.dec_c_nop),
.i_pipeline__i_pipeline_s1_decode__dec_c_or(
  i_pipeline.i_pipeline_s1_decode.dec_c_or),
.i_pipeline__i_pipeline_s1_decode__dec_c_slli(
  i_pipeline.i_pipeline_s1_decode.dec_c_slli),
.i_pipeline__i_pipeline_s1_decode__dec_c_srai(
  i_pipeline.i_pipeline_s1_decode.dec_c_srai),
.i_pipeline__i_pipeline_s1_decode__dec_c_srli(
  i_pipeline.i_pipeline_s1_decode.dec_c_srli),
.i_pipeline__i_pipeline_s1_decode__dec_c_sub(
  i_pipeline.i_pipeline_s1_decode.dec_c_sub),
.i_pipeline__i_pipeline_s1_decode__dec_c_sw(
  i_pipeline.i_pipeline_s1_decode.dec_c_sw),
.i_pipeline__i_pipeline_s1_decode__dec_c_swsp(
  i_pipeline.i_pipeline_s1_decode.dec_c_swsp),
.i_pipeline__i_pipeline_s1_decode__dec_c_xor(
  i_pipeline.i_pipeline_s1_decode.dec_c_xor),
.i_pipeline__i_pipeline_s1_decode__dec_csrrc(
  i_pipeline.i_pipeline_s1_decode.dec_csrrc),
.i_pipeline__i_pipeline_s1_decode__dec_csrrci(
  i_pipeline.i_pipeline_s1_decode.dec_csrrci),
.i_pipeline__i_pipeline_s1_decode__dec_csrrs(
  i_pipeline.i_pipeline_s1_decode.dec_csrrs),
.i_pipeline__i_pipeline_s1_decode__dec_csrrsi(
  i_pipeline.i_pipeline_s1_decode.dec_csrrsi),
.i_pipeline__i_pipeline_s1_decode__dec_csrrw(
  i_pipeline.i_pipeline_s1_decode.dec_csrrw),
.i_pipeline__i_pipeline_s1_decode__dec_csrrwi(
  i_pipeline.i_pipeline_s1_decode.dec_csrrwi),
.i_pipeline__i_pipeline_s1_decode__dec_div(
  i_pipeline.i_pipeline_s1_decode.dec_div),
.i_pipeline__i_pipeline_s1_decode__dec_divu(
  i_pipeline.i_pipeline_s1_decode.dec_divu),
.i_pipeline__i_pipeline_s1_decode__dec_ebreak(
  i_pipeline.i_pipeline_s1_decode.dec_ebreak),
.i_pipeline__i_pipeline_s1_decode__dec_ecall(
  i_pipeline.i_pipeline_s1_decode.dec_ecall),
.i_pipeline__i_pipeline_s1_decode__dec_fence(
  i_pipeline.i_pipeline_s1_decode.dec_fence),
.i_pipeline__i_pipeline_s1_decode__dec_fence_i(
  i_pipeline.i_pipeline_s1_decode.dec_fence_i),
.i_pipeline__i_pipeline_s1_decode__dec_jal(
  i_pipeline.i_pipeline_s1_decode.dec_jal),
.i_pipeline__i_pipeline_s1_decode__dec_jalr(
  i_pipeline.i_pipeline_s1_decode.dec_jalr),
.i_pipeline__i_pipeline_s1_decode__dec_lb(
  i_pipeline.i_pipeline_s1_decode.dec_lb),
.i_pipeline__i_pipeline_s1_decode__dec_lbu(
  i_pipeline.i_pipeline_s1_decode.dec_lbu),
.i_pipeline__i_pipeline_s1_decode__dec_lh(
  i_pipeline.i_pipeline_s1_decode.dec_lh),
.i_pipeline__i_pipeline_s1_decode__dec_lhu(
  i_pipeline.i_pipeline_s1_decode.dec_lhu),
.i_pipeline__i_pipeline_s1_decode__dec_lui(
  i_pipeline.i_pipeline_s1_decode.dec_lui),
.i_pipeline__i_pipeline_s1_decode__dec_lw(
  i_pipeline.i_pipeline_s1_decode.dec_lw),
.i_pipeline__i_pipeline_s1_decode__dec_mret(
  i_pipeline.i_pipeline_s1_decode.dec_mret),
.i_pipeline__i_pipeline_s1_decode__dec_mul(
  i_pipeline.i_pipeline_s1_decode.dec_mul),
.i_pipeline__i_pipeline_s1_decode__dec_mulh(
  i_pipeline.i_pipeline_s1_decode.dec_mulh),
.i_pipeline__i_pipeline_s1_decode__dec_mulhsu(
  i_pipeline.i_pipeline_s1_decode.dec_mulhsu),
.i_pipeline__i_pipeline_s1_decode__dec_mulhu(
  i_pipeline.i_pipeline_s1_decode.dec_mulhu),
.i_pipeline__i_pipeline_s1_decode__dec_or(
  i_pipeline.i_pipeline_s1_decode.dec_or),
.i_pipeline__i_pipeline_s1_decode__dec_ori(
  i_pipeline.i_pipeline_s1_decode.dec_ori),
.i_pipeline__i_pipeline_s1_decode__dec_rd_16(
  i_pipeline.i_pipeline_s1_decode.dec_rd_16),
.i_pipeline__i_pipeline_s1_decode__dec_rd_16_t0(
  i_pipeline.i_pipeline_s1_decode.dec_rd_16_t0),
.i_pipeline__i_pipeline_s1_decode__dec_rd_32(
  i_pipeline.i_pipeline_s1_decode.dec_rd_32),
.i_pipeline__i_pipeline_s1_decode__dec_rd_32_t0(
  i_pipeline.i_pipeline_s1_decode.dec_rd_32_t0),
.i_pipeline__i_pipeline_s1_decode__dec_rem(
  i_pipeline.i_pipeline_s1_decode.dec_rem),
.i_pipeline__i_pipeline_s1_decode__dec_remu(
  i_pipeline.i_pipeline_s1_decode.dec_remu),
.i_pipeline__i_pipeline_s1_decode__dec_rs1_16(
  i_pipeline.i_pipeline_s1_decode.dec_rs1_16),
.i_pipeline__i_pipeline_s1_decode__dec_rs1_16_t0(
  i_pipeline.i_pipeline_s1_decode.dec_rs1_16_t0),
.i_pipeline__i_pipeline_s1_decode__dec_rs2_16(
  i_pipeline.i_pipeline_s1_decode.dec_rs2_16),
.i_pipeline__i_pipeline_s1_decode__dec_rs2_16_t0(
  i_pipeline.i_pipeline_s1_decode.dec_rs2_16_t0),
.i_pipeline__i_pipeline_s1_decode__dec_sb(
  i_pipeline.i_pipeline_s1_decode.dec_sb),
.i_pipeline__i_pipeline_s1_decode__dec_sh(
  i_pipeline.i_pipeline_s1_decode.dec_sh),
.i_pipeline__i_pipeline_s1_decode__dec_sll(
  i_pipeline.i_pipeline_s1_decode.dec_sll),
.i_pipeline__i_pipeline_s1_decode__dec_slli(
  i_pipeline.i_pipeline_s1_decode.dec_slli),
.i_pipeline__i_pipeline_s1_decode__dec_slt(
  i_pipeline.i_pipeline_s1_decode.dec_slt),
.i_pipeline__i_pipeline_s1_decode__dec_slti(
  i_pipeline.i_pipeline_s1_decode.dec_slti),
.i_pipeline__i_pipeline_s1_decode__dec_sltiu(
  i_pipeline.i_pipeline_s1_decode.dec_sltiu),
.i_pipeline__i_pipeline_s1_decode__dec_sltu(
  i_pipeline.i_pipeline_s1_decode.dec_sltu),
.i_pipeline__i_pipeline_s1_decode__dec_sra(
  i_pipeline.i_pipeline_s1_decode.dec_sra),
.i_pipeline__i_pipeline_s1_decode__dec_srai(
  i_pipeline.i_pipeline_s1_decode.dec_srai),
.i_pipeline__i_pipeline_s1_decode__dec_srl(
  i_pipeline.i_pipeline_s1_decode.dec_srl),
.i_pipeline__i_pipeline_s1_decode__dec_srli(
  i_pipeline.i_pipeline_s1_decode.dec_srli),
.i_pipeline__i_pipeline_s1_decode__dec_sub(
  i_pipeline.i_pipeline_s1_decode.dec_sub),
.i_pipeline__i_pipeline_s1_decode__dec_sw(
  i_pipeline.i_pipeline_s1_decode.dec_sw),
.i_pipeline__i_pipeline_s1_decode__dec_wfi(
  i_pipeline.i_pipeline_s1_decode.dec_wfi),
.i_pipeline__i_pipeline_s1_decode__dec_xc_aesmix_dec(
  i_pipeline.i_pipeline_s1_decode.dec_xc_aesmix_dec),
.i_pipeline__i_pipeline_s1_decode__dec_xc_aesmix_enc(
  i_pipeline.i_pipeline_s1_decode.dec_xc_aesmix_enc),
.i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_dec(
  i_pipeline.i_pipeline_s1_decode.dec_xc_aessub_dec),
.i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_decrot(
  i_pipeline.i_pipeline_s1_decode.dec_xc_aessub_decrot),
.i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_enc(
  i_pipeline.i_pipeline_s1_decode.dec_xc_aessub_enc),
.i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_encrot(
  i_pipeline.i_pipeline_s1_decode.dec_xc_aessub_encrot),
.i_pipeline__i_pipeline_s1_decode__dec_xc_bop(
  i_pipeline.i_pipeline_s1_decode.dec_xc_bop),
.i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_b(
  i_pipeline.i_pipeline_s1_decode.dec_xc_ldr_b),
.i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_bu(
  i_pipeline.i_pipeline_s1_decode.dec_xc_ldr_bu),
.i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_h(
  i_pipeline.i_pipeline_s1_decode.dec_xc_ldr_h),
.i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_hu(
  i_pipeline.i_pipeline_s1_decode.dec_xc_ldr_hu),
.i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_w(
  i_pipeline.i_pipeline_s1_decode.dec_xc_ldr_w),
.i_pipeline__i_pipeline_s1_decode__dec_xc_lkgfence(
  i_pipeline.i_pipeline_s1_decode.dec_xc_lkgfence),
.i_pipeline__i_pipeline_s1_decode__dec_xc_lut(
  i_pipeline.i_pipeline_s1_decode.dec_xc_lut),
.i_pipeline__i_pipeline_s1_decode__dec_xc_macc_1(
  i_pipeline.i_pipeline_s1_decode.dec_xc_macc_1),
.i_pipeline__i_pipeline_s1_decode__dec_xc_madd_3(
  i_pipeline.i_pipeline_s1_decode.dec_xc_madd_3),
.i_pipeline__i_pipeline_s1_decode__dec_xc_mmul_3(
  i_pipeline.i_pipeline_s1_decode.dec_xc_mmul_3),
.i_pipeline__i_pipeline_s1_decode__dec_xc_mror(
  i_pipeline.i_pipeline_s1_decode.dec_xc_mror),
.i_pipeline__i_pipeline_s1_decode__dec_xc_msub_3(
  i_pipeline.i_pipeline_s1_decode.dec_xc_msub_3),
.i_pipeline__i_pipeline_s1_decode__dec_xc_padd(
  i_pipeline.i_pipeline_s1_decode.dec_xc_padd),
.i_pipeline__i_pipeline_s1_decode__dec_xc_pclmul_h(
  i_pipeline.i_pipeline_s1_decode.dec_xc_pclmul_h),
.i_pipeline__i_pipeline_s1_decode__dec_xc_pclmul_l(
  i_pipeline.i_pipeline_s1_decode.dec_xc_pclmul_l),
.i_pipeline__i_pipeline_s1_decode__dec_xc_pmul_h(
  i_pipeline.i_pipeline_s1_decode.dec_xc_pmul_h),
.i_pipeline__i_pipeline_s1_decode__dec_xc_pmul_l(
  i_pipeline.i_pipeline_s1_decode.dec_xc_pmul_l),
.i_pipeline__i_pipeline_s1_decode__dec_xc_pror(
  i_pipeline.i_pipeline_s1_decode.dec_xc_pror),
.i_pipeline__i_pipeline_s1_decode__dec_xc_pror_i(
  i_pipeline.i_pipeline_s1_decode.dec_xc_pror_i),
.i_pipeline__i_pipeline_s1_decode__dec_xc_psll(
  i_pipeline.i_pipeline_s1_decode.dec_xc_psll),
.i_pipeline__i_pipeline_s1_decode__dec_xc_psll_i(
  i_pipeline.i_pipeline_s1_decode.dec_xc_psll_i),
.i_pipeline__i_pipeline_s1_decode__dec_xc_psrl(
  i_pipeline.i_pipeline_s1_decode.dec_xc_psrl),
.i_pipeline__i_pipeline_s1_decode__dec_xc_psrl_i(
  i_pipeline.i_pipeline_s1_decode.dec_xc_psrl_i),
.i_pipeline__i_pipeline_s1_decode__dec_xc_psub(
  i_pipeline.i_pipeline_s1_decode.dec_xc_psub),
.i_pipeline__i_pipeline_s1_decode__dec_xc_rngsamp(
  i_pipeline.i_pipeline_s1_decode.dec_xc_rngsamp),
.i_pipeline__i_pipeline_s1_decode__dec_xc_rngseed(
  i_pipeline.i_pipeline_s1_decode.dec_xc_rngseed),
.i_pipeline__i_pipeline_s1_decode__dec_xc_rngtest(
  i_pipeline.i_pipeline_s1_decode.dec_xc_rngtest),
.i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s0(
  i_pipeline.i_pipeline_s1_decode.dec_xc_sha256_s0),
.i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s1(
  i_pipeline.i_pipeline_s1_decode.dec_xc_sha256_s1),
.i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s2(
  i_pipeline.i_pipeline_s1_decode.dec_xc_sha256_s2),
.i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s3(
  i_pipeline.i_pipeline_s1_decode.dec_xc_sha256_s3),
.i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_x1(
  i_pipeline.i_pipeline_s1_decode.dec_xc_sha3_x1),
.i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_x2(
  i_pipeline.i_pipeline_s1_decode.dec_xc_sha3_x2),
.i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_x4(
  i_pipeline.i_pipeline_s1_decode.dec_xc_sha3_x4),
.i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_xy(
  i_pipeline.i_pipeline_s1_decode.dec_xc_sha3_xy),
.i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_yx(
  i_pipeline.i_pipeline_s1_decode.dec_xc_sha3_yx),
.i_pipeline__i_pipeline_s1_decode__dec_xc_str_b(
  i_pipeline.i_pipeline_s1_decode.dec_xc_str_b),
.i_pipeline__i_pipeline_s1_decode__dec_xc_str_h(
  i_pipeline.i_pipeline_s1_decode.dec_xc_str_h),
.i_pipeline__i_pipeline_s1_decode__dec_xc_str_w(
  i_pipeline.i_pipeline_s1_decode.dec_xc_str_w),
.i_pipeline__i_pipeline_s1_decode__dec_xor(
  i_pipeline.i_pipeline_s1_decode.dec_xor),
.i_pipeline__i_pipeline_s1_decode__dec_xori(
  i_pipeline.i_pipeline_s1_decode.dec_xori),
.i_pipeline__i_pipeline_s1_decode__instr_16bit(
  i_pipeline.i_pipeline_s1_decode.instr_16bit),
.i_pipeline__i_pipeline_s1_decode__instr_32bit(
  i_pipeline.i_pipeline_s1_decode.instr_32bit),
.i_pipeline__i_pipeline_s1_decode__invalid_instr(
  i_pipeline.i_pipeline_s1_decode.invalid_instr),
.i_pipeline__i_pipeline_s1_decode__leak_stall(
  i_pipeline.i_pipeline_s1_decode.leak_stall),
.i_pipeline__i_pipeline_s1_decode__lf_count(
  i_pipeline.i_pipeline_s1_decode.lf_count),
.i_pipeline__i_pipeline_s1_decode__lf_count_ld(
  i_pipeline.i_pipeline_s1_decode.lf_count_ld),
.i_pipeline__i_pipeline_s1_decode__lsu_no_rd(
  i_pipeline.i_pipeline_s1_decode.lsu_no_rd),
.i_pipeline__i_pipeline_s1_decode__lsu_width(
  i_pipeline.i_pipeline_s1_decode.lsu_width),
.i_pipeline__i_pipeline_s1_decode__n_lf_count(
  i_pipeline.i_pipeline_s1_decode.n_lf_count),
.i_pipeline__i_pipeline_s1_decode__n_program_counter(
  i_pipeline.i_pipeline_s1_decode.n_program_counter),
.i_pipeline__i_pipeline_s1_decode__n_program_counter_t0(
  i_pipeline.i_pipeline_s1_decode.n_program_counter_t0),
.i_pipeline__i_pipeline_s1_decode__n_s2_fu(
  i_pipeline.i_pipeline_s1_decode.n_s2_fu),
.i_pipeline__i_pipeline_s1_decode__n_s2_imm(
  i_pipeline.i_pipeline_s1_decode.n_s2_imm),
.i_pipeline__i_pipeline_s1_decode__n_s2_imm_pc(
  i_pipeline.i_pipeline_s1_decode.n_s2_imm_pc),
.i_pipeline__i_pipeline_s1_decode__n_s2_imm_pc_t0(
  i_pipeline.i_pipeline_s1_decode.n_s2_imm_pc_t0),
.i_pipeline__i_pipeline_s1_decode__n_s2_imm_t0(
  i_pipeline.i_pipeline_s1_decode.n_s2_imm_t0),
.i_pipeline__i_pipeline_s1_decode__n_s2_instr(
  i_pipeline.i_pipeline_s1_decode.n_s2_instr),
.i_pipeline__i_pipeline_s1_decode__n_s2_instr_t0(
  i_pipeline.i_pipeline_s1_decode.n_s2_instr_t0),
.i_pipeline__i_pipeline_s1_decode__n_s2_opr_a(
  i_pipeline.i_pipeline_s1_decode.n_s2_opr_a),
.i_pipeline__i_pipeline_s1_decode__n_s2_opr_a_t0(
  i_pipeline.i_pipeline_s1_decode.n_s2_opr_a_t0),
.i_pipeline__i_pipeline_s1_decode__n_s2_opr_b(
  i_pipeline.i_pipeline_s1_decode.n_s2_opr_b),
.i_pipeline__i_pipeline_s1_decode__n_s2_opr_b_t0(
  i_pipeline.i_pipeline_s1_decode.n_s2_opr_b_t0),
.i_pipeline__i_pipeline_s1_decode__n_s2_opr_c(
  i_pipeline.i_pipeline_s1_decode.n_s2_opr_c),
.i_pipeline__i_pipeline_s1_decode__n_s2_opr_c_t0(
  i_pipeline.i_pipeline_s1_decode.n_s2_opr_c_t0),
.i_pipeline__i_pipeline_s1_decode__n_s2_pw(
  i_pipeline.i_pipeline_s1_decode.n_s2_pw),
.i_pipeline__i_pipeline_s1_decode__n_s2_pw_t0(
  i_pipeline.i_pipeline_s1_decode.n_s2_pw_t0),
.i_pipeline__i_pipeline_s1_decode__n_s2_rd(
  i_pipeline.i_pipeline_s1_decode.n_s2_rd),
.i_pipeline__i_pipeline_s1_decode__n_s2_rd_t0(
  i_pipeline.i_pipeline_s1_decode.n_s2_rd_t0),
.i_pipeline__i_pipeline_s1_decode__n_s2_trap(
  i_pipeline.i_pipeline_s1_decode.n_s2_trap),
.i_pipeline__i_pipeline_s1_decode__n_s2_uop(
  i_pipeline.i_pipeline_s1_decode.n_s2_uop),
.i_pipeline__i_pipeline_s1_decode__n_s2_valid(
  i_pipeline.i_pipeline_s1_decode.n_s2_valid),
.i_pipeline__i_pipeline_s1_decode__opra_flush(
  i_pipeline.i_pipeline_s1_decode.opra_flush),
.i_pipeline__i_pipeline_s1_decode__opra_ld_en(
  i_pipeline.i_pipeline_s1_decode.opra_ld_en),
.i_pipeline__i_pipeline_s1_decode__opra_src_csri(
  i_pipeline.i_pipeline_s1_decode.opra_src_csri),
.i_pipeline__i_pipeline_s1_decode__opra_src_rs1(
  i_pipeline.i_pipeline_s1_decode.opra_src_rs1),
.i_pipeline__i_pipeline_s1_decode__opra_src_zero(
  i_pipeline.i_pipeline_s1_decode.opra_src_zero),
.i_pipeline__i_pipeline_s1_decode__oprb_flush(
  i_pipeline.i_pipeline_s1_decode.oprb_flush),
.i_pipeline__i_pipeline_s1_decode__oprb_ld_en(
  i_pipeline.i_pipeline_s1_decode.oprb_ld_en),
.i_pipeline__i_pipeline_s1_decode__oprb_rs2_shf_1(
  i_pipeline.i_pipeline_s1_decode.oprb_rs2_shf_1),
.i_pipeline__i_pipeline_s1_decode__oprb_rs2_shf_2(
  i_pipeline.i_pipeline_s1_decode.oprb_rs2_shf_2),
.i_pipeline__i_pipeline_s1_decode__oprb_src_imm(
  i_pipeline.i_pipeline_s1_decode.oprb_src_imm),
.i_pipeline__i_pipeline_s1_decode__oprb_src_rs2(
  i_pipeline.i_pipeline_s1_decode.oprb_src_rs2),
.i_pipeline__i_pipeline_s1_decode__oprb_src_zero(
  i_pipeline.i_pipeline_s1_decode.oprb_src_zero),
.i_pipeline__i_pipeline_s1_decode__oprc_flush(
  i_pipeline.i_pipeline_s1_decode.oprc_flush),
.i_pipeline__i_pipeline_s1_decode__oprc_ld_en(
  i_pipeline.i_pipeline_s1_decode.oprc_ld_en),
.i_pipeline__i_pipeline_s1_decode__oprc_src_pcim(
  i_pipeline.i_pipeline_s1_decode.oprc_src_pcim),
.i_pipeline__i_pipeline_s1_decode__oprc_src_rs2(
  i_pipeline.i_pipeline_s1_decode.oprc_src_rs2),
.i_pipeline__i_pipeline_s1_decode__oprc_src_rs3(
  i_pipeline.i_pipeline_s1_decode.oprc_src_rs3),
.i_pipeline__i_pipeline_s1_decode__p_in(
  i_pipeline.i_pipeline_s1_decode.p_in),
.i_pipeline__i_pipeline_s1_decode__p_in_t0(
  i_pipeline.i_pipeline_s1_decode.p_in_t0),
.i_pipeline__i_pipeline_s1_decode__p_mr(
  i_pipeline.i_pipeline_s1_decode.p_mr),
.i_pipeline__i_pipeline_s1_decode__p_mr_t0(
  i_pipeline.i_pipeline_s1_decode.p_mr_t0),
.i_pipeline__i_pipeline_s1_decode__p_out(
  i_pipeline.i_pipeline_s1_decode.p_out),
.i_pipeline__i_pipeline_s1_decode__p_out_t0(
  i_pipeline.i_pipeline_s1_decode.p_out_t0),
.i_pipeline__i_pipeline_s1_decode__p_s2_busy(
  i_pipeline.i_pipeline_s1_decode.p_s2_busy),
.i_pipeline__i_pipeline_s1_decode__p_s2_busy_t0(
  i_pipeline.i_pipeline_s1_decode.p_s2_busy_t0),
.i_pipeline__i_pipeline_s1_decode__packed_instruction(
  i_pipeline.i_pipeline_s1_decode.packed_instruction),
.i_pipeline__i_pipeline_s1_decode__pc_plus_imm(
  i_pipeline.i_pipeline_s1_decode.pc_plus_imm),
.i_pipeline__i_pipeline_s1_decode__pc_plus_imm_t0(
  i_pipeline.i_pipeline_s1_decode.pc_plus_imm_t0),
.i_pipeline__i_pipeline_s1_decode__pipe_progress(
  i_pipeline.i_pipeline_s1_decode.pipe_progress),
.i_pipeline__i_pipeline_s1_decode__program_counter(
  i_pipeline.i_pipeline_s1_decode.program_counter),
.i_pipeline__i_pipeline_s1_decode__program_counter_t0(
  i_pipeline.i_pipeline_s1_decode.program_counter_t0),
.i_pipeline__i_pipeline_s1_decode__s1_rs2_shf(
  i_pipeline.i_pipeline_s1_decode.s1_rs2_shf),
.i_pipeline__i_pipeline_s1_decode__s1_rs2_shf_t0(
  i_pipeline.i_pipeline_s1_decode.s1_rs2_shf_t0),
.i_pipeline__i_pipeline_s1_decode__trap_cause(
  i_pipeline.i_pipeline_s1_decode.trap_cause),
.i_pipeline__i_pipeline_s1_decode__uop_alu(
  i_pipeline.i_pipeline_s1_decode.uop_alu),
.i_pipeline__i_pipeline_s1_decode__uop_asi(
  i_pipeline.i_pipeline_s1_decode.uop_asi),
.i_pipeline__i_pipeline_s1_decode__uop_bit(
  i_pipeline.i_pipeline_s1_decode.uop_bit),
.i_pipeline__i_pipeline_s1_decode__uop_cfu(
  i_pipeline.i_pipeline_s1_decode.uop_cfu),
.i_pipeline__i_pipeline_s1_decode__uop_csr(
  i_pipeline.i_pipeline_s1_decode.uop_csr),
.i_pipeline__i_pipeline_s1_decode__uop_lsu(
  i_pipeline.i_pipeline_s1_decode.uop_lsu),
.i_pipeline__i_pipeline_s1_decode__uop_mul(
  i_pipeline.i_pipeline_s1_decode.uop_mul),
.i_pipeline__i_pipeline_s1_decode__uop_rng(
  i_pipeline.i_pipeline_s1_decode.uop_rng),
.i_pipeline__i_pipeline_s1_decode__use_imm32_b(
  i_pipeline.i_pipeline_s1_decode.use_imm32_b),
.i_pipeline__i_pipeline_s1_decode__use_imm32_i(
  i_pipeline.i_pipeline_s1_decode.use_imm32_i),
.i_pipeline__i_pipeline_s1_decode__use_imm32_s(
  i_pipeline.i_pipeline_s1_decode.use_imm32_s),
.i_pipeline__i_pipeline_s1_decode__use_imm32_u(
  i_pipeline.i_pipeline_s1_decode.use_imm32_u),
.i_pipeline__i_pipeline_s1_decode__use_imm_csr(
  i_pipeline.i_pipeline_s1_decode.use_imm_csr),
.i_pipeline__i_pipeline_s1_decode__use_imm_sha3(
  i_pipeline.i_pipeline_s1_decode.use_imm_sha3),
.i_pipeline__i_pipeline_s1_decode__use_imm_shfi(
  i_pipeline.i_pipeline_s1_decode.use_imm_shfi),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__g_clk(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.g_clk),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__g_resetn(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.g_resetn),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_data(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.i_data),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_valid(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.i_valid),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_busy(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.o_busy),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__mr_data(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.mr_data),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__flush(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.flush),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__flush_dat(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.flush_dat),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_data(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.o_data),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_valid(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.o_valid),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_busy(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.i_busy),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__flush_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.flush_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_valid_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.o_valid_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_data_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.o_data_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_busy_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.o_busy_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__mr_data_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.mr_data_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_valid_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.i_valid_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_data_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.i_data_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_busy_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.i_busy_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__flush_dat_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.flush_dat_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__genblk1__progress(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg.\genblk1.progress ),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__g_clk(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.g_clk),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__g_resetn(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.g_resetn),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_data(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.i_data),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_valid(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.i_valid),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_busy(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.o_busy),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__mr_data(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.mr_data),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__flush(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.flush),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__flush_dat(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.flush_dat),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_data(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.o_data),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_valid(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.o_valid),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_busy(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.i_busy),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__flush_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.flush_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_valid_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.o_valid_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_data_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.o_data_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_busy_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.o_busy_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__mr_data_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.mr_data_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_valid_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.i_valid_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_data_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.i_data_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_busy_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.i_busy_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__flush_dat_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.flush_dat_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__genblk1__progress(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_a.\genblk1.progress ),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__g_clk(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.g_clk),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__g_resetn(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.g_resetn),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_data(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.i_data),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_valid(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.i_valid),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_busy(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.o_busy),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__mr_data(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.mr_data),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__flush(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.flush),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__flush_dat(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.flush_dat),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_data(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.o_data),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_valid(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.o_valid),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_busy(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.i_busy),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__flush_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.flush_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_valid_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.o_valid_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_data_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.o_data_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_busy_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.o_busy_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__mr_data_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.mr_data_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_valid_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.i_valid_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_data_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.i_data_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_busy_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.i_busy_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__flush_dat_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.flush_dat_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__genblk1__progress(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_b.\genblk1.progress ),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__g_clk(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.g_clk),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__g_resetn(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.g_resetn),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_data(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.i_data),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_valid(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.i_valid),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_busy(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.o_busy),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__mr_data(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.mr_data),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__flush(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.flush),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__flush_dat(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.flush_dat),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_data(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.o_data),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_valid(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.o_valid),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_busy(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.i_busy),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__flush_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.flush_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_valid_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.o_valid_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_data_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.o_data_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_busy_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.o_busy_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__mr_data_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.mr_data_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_valid_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.i_valid_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_data_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.i_data_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_busy_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.i_busy_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__flush_dat_t0(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.flush_dat_t0),
.i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__genblk1__progress(
  i_pipeline.i_pipeline_s1_decode.i_decode_pipereg_opr_c.\genblk1.progress ),
.i_pipeline__i_pipeline_s1_decode__i_frv_leak__g_clk(
  i_pipeline.i_pipeline_s1_decode.i_frv_leak.g_clk),
.i_pipeline__i_pipeline_s1_decode__i_frv_leak__g_resetn(
  i_pipeline.i_pipeline_s1_decode.i_frv_leak.g_resetn),
.i_pipeline__i_pipeline_s1_decode__i_frv_leak__leak_prng(
  i_pipeline.i_pipeline_s1_decode.i_frv_leak.leak_prng),
.i_pipeline__i_pipeline_s1_decode__i_frv_leak__leak_fence(
  i_pipeline.i_pipeline_s1_decode.i_frv_leak.leak_fence),
.i_pipeline__i_pipeline_s1_decode__i_frv_leak__leak_prng_t0(
  i_pipeline.i_pipeline_s1_decode.i_frv_leak.leak_prng_t0),
.i_pipeline__i_pipeline_s1_decode__i_frv_leak__leak_fence_t0(
  i_pipeline.i_pipeline_s1_decode.i_frv_leak.leak_fence_t0),
.i_pipeline__i_pipeline_s1_decode__i_frv_leak__genblk1__genblk1__n_prng_lsb(
  i_pipeline.i_pipeline_s1_decode.i_frv_leak.\genblk1.genblk1.n_prng_lsb ),
.i_pipeline__i_pipeline_s1_decode__i_frv_leak__genblk1__genblk1__n_prng_lsb_t0(
  i_pipeline.i_pipeline_s1_decode.i_frv_leak.\genblk1.genblk1.n_prng_lsb_t0 ),
.i_pipeline__i_pipeline_s2_execute__g_clk(
  i_pipeline.i_pipeline_s2_execute.g_clk),
.i_pipeline__i_pipeline_s2_execute__g_resetn(
  i_pipeline.i_pipeline_s2_execute.g_resetn),
.i_pipeline__i_pipeline_s2_execute__s2_rd(
  i_pipeline.i_pipeline_s2_execute.s2_rd),
.i_pipeline__i_pipeline_s2_execute__s2_opr_a(
  i_pipeline.i_pipeline_s2_execute.s2_opr_a),
.i_pipeline__i_pipeline_s2_execute__s2_opr_b(
  i_pipeline.i_pipeline_s2_execute.s2_opr_b),
.i_pipeline__i_pipeline_s2_execute__s2_opr_c(
  i_pipeline.i_pipeline_s2_execute.s2_opr_c),
.i_pipeline__i_pipeline_s2_execute__s2_uop(
  i_pipeline.i_pipeline_s2_execute.s2_uop),
.i_pipeline__i_pipeline_s2_execute__s2_fu(
  i_pipeline.i_pipeline_s2_execute.s2_fu),
.i_pipeline__i_pipeline_s2_execute__s2_pw(
  i_pipeline.i_pipeline_s2_execute.s2_pw),
.i_pipeline__i_pipeline_s2_execute__s2_trap(
  i_pipeline.i_pipeline_s2_execute.s2_trap),
.i_pipeline__i_pipeline_s2_execute__s2_size(
  i_pipeline.i_pipeline_s2_execute.s2_size),
.i_pipeline__i_pipeline_s2_execute__s2_instr(
  i_pipeline.i_pipeline_s2_execute.s2_instr),
.i_pipeline__i_pipeline_s2_execute__s2_busy(
  i_pipeline.i_pipeline_s2_execute.s2_busy),
.i_pipeline__i_pipeline_s2_execute__s2_valid(
  i_pipeline.i_pipeline_s2_execute.s2_valid),
.i_pipeline__i_pipeline_s2_execute__leak_prng(
  i_pipeline.i_pipeline_s2_execute.leak_prng),
.i_pipeline__i_pipeline_s2_execute__leak_lkgcfg(
  i_pipeline.i_pipeline_s2_execute.leak_lkgcfg),
.i_pipeline__i_pipeline_s2_execute__rng_req_valid(
  i_pipeline.i_pipeline_s2_execute.rng_req_valid),
.i_pipeline__i_pipeline_s2_execute__rng_req_op(
  i_pipeline.i_pipeline_s2_execute.rng_req_op),
.i_pipeline__i_pipeline_s2_execute__rng_req_data(
  i_pipeline.i_pipeline_s2_execute.rng_req_data),
.i_pipeline__i_pipeline_s2_execute__rng_req_ready(
  i_pipeline.i_pipeline_s2_execute.rng_req_ready),
.i_pipeline__i_pipeline_s2_execute__rng_rsp_valid(
  i_pipeline.i_pipeline_s2_execute.rng_rsp_valid),
.i_pipeline__i_pipeline_s2_execute__rng_rsp_status(
  i_pipeline.i_pipeline_s2_execute.rng_rsp_status),
.i_pipeline__i_pipeline_s2_execute__rng_rsp_data(
  i_pipeline.i_pipeline_s2_execute.rng_rsp_data),
.i_pipeline__i_pipeline_s2_execute__rng_rsp_ready(
  i_pipeline.i_pipeline_s2_execute.rng_rsp_ready),
.i_pipeline__i_pipeline_s2_execute__uxcrypto_ct(
  i_pipeline.i_pipeline_s2_execute.uxcrypto_ct),
.i_pipeline__i_pipeline_s2_execute__uxcrypto_b0(
  i_pipeline.i_pipeline_s2_execute.uxcrypto_b0),
.i_pipeline__i_pipeline_s2_execute__uxcrypto_b1(
  i_pipeline.i_pipeline_s2_execute.uxcrypto_b1),
.i_pipeline__i_pipeline_s2_execute__flush(
  i_pipeline.i_pipeline_s2_execute.flush),
.i_pipeline__i_pipeline_s2_execute__fwd_s2_rd(
  i_pipeline.i_pipeline_s2_execute.fwd_s2_rd),
.i_pipeline__i_pipeline_s2_execute__fwd_s2_wide(
  i_pipeline.i_pipeline_s2_execute.fwd_s2_wide),
.i_pipeline__i_pipeline_s2_execute__fwd_s2_wdata(
  i_pipeline.i_pipeline_s2_execute.fwd_s2_wdata),
.i_pipeline__i_pipeline_s2_execute__fwd_s2_wdata_hi(
  i_pipeline.i_pipeline_s2_execute.fwd_s2_wdata_hi),
.i_pipeline__i_pipeline_s2_execute__fwd_s2_load(
  i_pipeline.i_pipeline_s2_execute.fwd_s2_load),
.i_pipeline__i_pipeline_s2_execute__fwd_s2_csr(
  i_pipeline.i_pipeline_s2_execute.fwd_s2_csr),
.i_pipeline__i_pipeline_s2_execute__s3_rd(
  i_pipeline.i_pipeline_s2_execute.s3_rd),
.i_pipeline__i_pipeline_s2_execute__s3_opr_a(
  i_pipeline.i_pipeline_s2_execute.s3_opr_a),
.i_pipeline__i_pipeline_s2_execute__s3_opr_b(
  i_pipeline.i_pipeline_s2_execute.s3_opr_b),
.i_pipeline__i_pipeline_s2_execute__s3_uop(
  i_pipeline.i_pipeline_s2_execute.s3_uop),
.i_pipeline__i_pipeline_s2_execute__s3_fu(
  i_pipeline.i_pipeline_s2_execute.s3_fu),
.i_pipeline__i_pipeline_s2_execute__s3_trap(
  i_pipeline.i_pipeline_s2_execute.s3_trap),
.i_pipeline__i_pipeline_s2_execute__s3_size(
  i_pipeline.i_pipeline_s2_execute.s3_size),
.i_pipeline__i_pipeline_s2_execute__s3_instr(
  i_pipeline.i_pipeline_s2_execute.s3_instr),
.i_pipeline__i_pipeline_s2_execute__s3_busy(
  i_pipeline.i_pipeline_s2_execute.s3_busy),
.i_pipeline__i_pipeline_s2_execute__s3_valid(
  i_pipeline.i_pipeline_s2_execute.s3_valid),
.i_pipeline__i_pipeline_s2_execute__flush_t0(
  i_pipeline.i_pipeline_s2_execute.flush_t0),
.i_pipeline__i_pipeline_s2_execute__s2_valid_t0(
  i_pipeline.i_pipeline_s2_execute.s2_valid_t0),
.i_pipeline__i_pipeline_s2_execute__s2_uop_t0(
  i_pipeline.i_pipeline_s2_execute.s2_uop_t0),
.i_pipeline__i_pipeline_s2_execute__s2_trap_t0(
  i_pipeline.i_pipeline_s2_execute.s2_trap_t0),
.i_pipeline__i_pipeline_s2_execute__s2_size_t0(
  i_pipeline.i_pipeline_s2_execute.s2_size_t0),
.i_pipeline__i_pipeline_s2_execute__s2_rd_t0(
  i_pipeline.i_pipeline_s2_execute.s2_rd_t0),
.i_pipeline__i_pipeline_s2_execute__s2_pw_t0(
  i_pipeline.i_pipeline_s2_execute.s2_pw_t0),
.i_pipeline__i_pipeline_s2_execute__s2_opr_c_t0(
  i_pipeline.i_pipeline_s2_execute.s2_opr_c_t0),
.i_pipeline__i_pipeline_s2_execute__s2_opr_b_t0(
  i_pipeline.i_pipeline_s2_execute.s2_opr_b_t0),
.i_pipeline__i_pipeline_s2_execute__s2_opr_a_t0(
  i_pipeline.i_pipeline_s2_execute.s2_opr_a_t0),
.i_pipeline__i_pipeline_s2_execute__s2_instr_t0(
  i_pipeline.i_pipeline_s2_execute.s2_instr_t0),
.i_pipeline__i_pipeline_s2_execute__s2_fu_t0(
  i_pipeline.i_pipeline_s2_execute.s2_fu_t0),
.i_pipeline__i_pipeline_s2_execute__s2_busy_t0(
  i_pipeline.i_pipeline_s2_execute.s2_busy_t0),
.i_pipeline__i_pipeline_s2_execute__leak_lkgcfg_t0(
  i_pipeline.i_pipeline_s2_execute.leak_lkgcfg_t0),
.i_pipeline__i_pipeline_s2_execute__leak_prng_t0(
  i_pipeline.i_pipeline_s2_execute.leak_prng_t0),
.i_pipeline__i_pipeline_s2_execute__rng_req_data_t0(
  i_pipeline.i_pipeline_s2_execute.rng_req_data_t0),
.i_pipeline__i_pipeline_s2_execute__rng_req_op_t0(
  i_pipeline.i_pipeline_s2_execute.rng_req_op_t0),
.i_pipeline__i_pipeline_s2_execute__rng_req_ready_t0(
  i_pipeline.i_pipeline_s2_execute.rng_req_ready_t0),
.i_pipeline__i_pipeline_s2_execute__rng_req_valid_t0(
  i_pipeline.i_pipeline_s2_execute.rng_req_valid_t0),
.i_pipeline__i_pipeline_s2_execute__rng_rsp_data_t0(
  i_pipeline.i_pipeline_s2_execute.rng_rsp_data_t0),
.i_pipeline__i_pipeline_s2_execute__rng_rsp_ready_t0(
  i_pipeline.i_pipeline_s2_execute.rng_rsp_ready_t0),
.i_pipeline__i_pipeline_s2_execute__rng_rsp_status_t0(
  i_pipeline.i_pipeline_s2_execute.rng_rsp_status_t0),
.i_pipeline__i_pipeline_s2_execute__rng_rsp_valid_t0(
  i_pipeline.i_pipeline_s2_execute.rng_rsp_valid_t0),
.i_pipeline__i_pipeline_s2_execute__fwd_s2_csr_t0(
  i_pipeline.i_pipeline_s2_execute.fwd_s2_csr_t0),
.i_pipeline__i_pipeline_s2_execute__fwd_s2_load_t0(
  i_pipeline.i_pipeline_s2_execute.fwd_s2_load_t0),
.i_pipeline__i_pipeline_s2_execute__fwd_s2_rd_t0(
  i_pipeline.i_pipeline_s2_execute.fwd_s2_rd_t0),
.i_pipeline__i_pipeline_s2_execute__fwd_s2_wdata_t0(
  i_pipeline.i_pipeline_s2_execute.fwd_s2_wdata_t0),
.i_pipeline__i_pipeline_s2_execute__fwd_s2_wdata_hi_t0(
  i_pipeline.i_pipeline_s2_execute.fwd_s2_wdata_hi_t0),
.i_pipeline__i_pipeline_s2_execute__fwd_s2_wide_t0(
  i_pipeline.i_pipeline_s2_execute.fwd_s2_wide_t0),
.i_pipeline__i_pipeline_s2_execute__s3_busy_t0(
  i_pipeline.i_pipeline_s2_execute.s3_busy_t0),
.i_pipeline__i_pipeline_s2_execute__s3_fu_t0(
  i_pipeline.i_pipeline_s2_execute.s3_fu_t0),
.i_pipeline__i_pipeline_s2_execute__s3_instr_t0(
  i_pipeline.i_pipeline_s2_execute.s3_instr_t0),
.i_pipeline__i_pipeline_s2_execute__s3_opr_a_t0(
  i_pipeline.i_pipeline_s2_execute.s3_opr_a_t0),
.i_pipeline__i_pipeline_s2_execute__s3_opr_b_t0(
  i_pipeline.i_pipeline_s2_execute.s3_opr_b_t0),
.i_pipeline__i_pipeline_s2_execute__s3_rd_t0(
  i_pipeline.i_pipeline_s2_execute.s3_rd_t0),
.i_pipeline__i_pipeline_s2_execute__s3_size_t0(
  i_pipeline.i_pipeline_s2_execute.s3_size_t0),
.i_pipeline__i_pipeline_s2_execute__s3_trap_t0(
  i_pipeline.i_pipeline_s2_execute.s3_trap_t0),
.i_pipeline__i_pipeline_s2_execute__s3_uop_t0(
  i_pipeline.i_pipeline_s2_execute.s3_uop_t0),
.i_pipeline__i_pipeline_s2_execute__s3_valid_t0(
  i_pipeline.i_pipeline_s2_execute.s3_valid_t0),
.i_pipeline__i_pipeline_s2_execute__uxcrypto_b0_t0(
  i_pipeline.i_pipeline_s2_execute.uxcrypto_b0_t0),
.i_pipeline__i_pipeline_s2_execute__uxcrypto_b1_t0(
  i_pipeline.i_pipeline_s2_execute.uxcrypto_b1_t0),
.i_pipeline__i_pipeline_s2_execute__uxcrypto_ct_t0(
  i_pipeline.i_pipeline_s2_execute.uxcrypto_ct_t0),
.i_pipeline__i_pipeline_s2_execute__alu_add_result(
  i_pipeline.i_pipeline_s2_execute.alu_add_result),
.i_pipeline__i_pipeline_s2_execute__alu_add_result_t0(
  i_pipeline.i_pipeline_s2_execute.alu_add_result_t0),
.i_pipeline__i_pipeline_s2_execute__alu_eq(
  i_pipeline.i_pipeline_s2_execute.alu_eq),
.i_pipeline__i_pipeline_s2_execute__alu_eq_t0(
  i_pipeline.i_pipeline_s2_execute.alu_eq_t0),
.i_pipeline__i_pipeline_s2_execute__alu_lt(
  i_pipeline.i_pipeline_s2_execute.alu_lt),
.i_pipeline__i_pipeline_s2_execute__alu_lt_t0(
  i_pipeline.i_pipeline_s2_execute.alu_lt_t0),
.i_pipeline__i_pipeline_s2_execute__alu_op_add(
  i_pipeline.i_pipeline_s2_execute.alu_op_add),
.i_pipeline__i_pipeline_s2_execute__alu_op_and(
  i_pipeline.i_pipeline_s2_execute.alu_op_and),
.i_pipeline__i_pipeline_s2_execute__alu_op_cmp(
  i_pipeline.i_pipeline_s2_execute.alu_op_cmp),
.i_pipeline__i_pipeline_s2_execute__alu_op_or(
  i_pipeline.i_pipeline_s2_execute.alu_op_or),
.i_pipeline__i_pipeline_s2_execute__alu_op_rot(
  i_pipeline.i_pipeline_s2_execute.alu_op_rot),
.i_pipeline__i_pipeline_s2_execute__alu_op_shf(
  i_pipeline.i_pipeline_s2_execute.alu_op_shf),
.i_pipeline__i_pipeline_s2_execute__alu_op_shf_arith(
  i_pipeline.i_pipeline_s2_execute.alu_op_shf_arith),
.i_pipeline__i_pipeline_s2_execute__alu_op_shf_left(
  i_pipeline.i_pipeline_s2_execute.alu_op_shf_left),
.i_pipeline__i_pipeline_s2_execute__alu_op_sub(
  i_pipeline.i_pipeline_s2_execute.alu_op_sub),
.i_pipeline__i_pipeline_s2_execute__alu_op_unsigned(
  i_pipeline.i_pipeline_s2_execute.alu_op_unsigned),
.i_pipeline__i_pipeline_s2_execute__alu_op_xor(
  i_pipeline.i_pipeline_s2_execute.alu_op_xor),
.i_pipeline__i_pipeline_s2_execute__alu_ready(
  i_pipeline.i_pipeline_s2_execute.alu_ready),
.i_pipeline__i_pipeline_s2_execute__alu_ready_t0(
  i_pipeline.i_pipeline_s2_execute.alu_ready_t0),
.i_pipeline__i_pipeline_s2_execute__alu_result(
  i_pipeline.i_pipeline_s2_execute.alu_result),
.i_pipeline__i_pipeline_s2_execute__alu_result_t0(
  i_pipeline.i_pipeline_s2_execute.alu_result_t0),
.i_pipeline__i_pipeline_s2_execute__asi_done(
  i_pipeline.i_pipeline_s2_execute.asi_done),
.i_pipeline__i_pipeline_s2_execute__asi_finished(
  i_pipeline.i_pipeline_s2_execute.asi_finished),
.i_pipeline__i_pipeline_s2_execute__asi_flush_aesmix(
  i_pipeline.i_pipeline_s2_execute.asi_flush_aesmix),
.i_pipeline__i_pipeline_s2_execute__asi_flush_aessub(
  i_pipeline.i_pipeline_s2_execute.asi_flush_aessub),
.i_pipeline__i_pipeline_s2_execute__asi_ready(
  i_pipeline.i_pipeline_s2_execute.asi_ready),
.i_pipeline__i_pipeline_s2_execute__asi_ready_t0(
  i_pipeline.i_pipeline_s2_execute.asi_ready_t0),
.i_pipeline__i_pipeline_s2_execute__asi_result(
  i_pipeline.i_pipeline_s2_execute.asi_result),
.i_pipeline__i_pipeline_s2_execute__asi_result_t0(
  i_pipeline.i_pipeline_s2_execute.asi_result_t0),
.i_pipeline__i_pipeline_s2_execute__bitw_bop(
  i_pipeline.i_pipeline_s2_execute.bitw_bop),
.i_pipeline__i_pipeline_s2_execute__bitw_bop_lut(
  i_pipeline.i_pipeline_s2_execute.bitw_bop_lut),
.i_pipeline__i_pipeline_s2_execute__bitw_bop_lut_t0(
  i_pipeline.i_pipeline_s2_execute.bitw_bop_lut_t0),
.i_pipeline__i_pipeline_s2_execute__bitw_cmov(
  i_pipeline.i_pipeline_s2_execute.bitw_cmov),
.i_pipeline__i_pipeline_s2_execute__bitw_flush(
  i_pipeline.i_pipeline_s2_execute.bitw_flush),
.i_pipeline__i_pipeline_s2_execute__bitw_fsl(
  i_pipeline.i_pipeline_s2_execute.bitw_fsl),
.i_pipeline__i_pipeline_s2_execute__bitw_fsr(
  i_pipeline.i_pipeline_s2_execute.bitw_fsr),
.i_pipeline__i_pipeline_s2_execute__bitw_gpr_wide(
  i_pipeline.i_pipeline_s2_execute.bitw_gpr_wide),
.i_pipeline__i_pipeline_s2_execute__bitw_lut(
  i_pipeline.i_pipeline_s2_execute.bitw_lut),
.i_pipeline__i_pipeline_s2_execute__bitw_ready(
  i_pipeline.i_pipeline_s2_execute.bitw_ready),
.i_pipeline__i_pipeline_s2_execute__bitw_ready_t0(
  i_pipeline.i_pipeline_s2_execute.bitw_ready_t0),
.i_pipeline__i_pipeline_s2_execute__bitw_result_wide(
  i_pipeline.i_pipeline_s2_execute.bitw_result_wide),
.i_pipeline__i_pipeline_s2_execute__bitw_result_wide_t0(
  i_pipeline.i_pipeline_s2_execute.bitw_result_wide_t0),
.i_pipeline__i_pipeline_s2_execute__cfu_cond(
  i_pipeline.i_pipeline_s2_execute.cfu_cond),
.i_pipeline__i_pipeline_s2_execute__cfu_cond_taken(
  i_pipeline.i_pipeline_s2_execute.cfu_cond_taken),
.i_pipeline__i_pipeline_s2_execute__cfu_jalr(
  i_pipeline.i_pipeline_s2_execute.cfu_jalr),
.i_pipeline__i_pipeline_s2_execute__cond_beq(
  i_pipeline.i_pipeline_s2_execute.cond_beq),
.i_pipeline__i_pipeline_s2_execute__cond_bge(
  i_pipeline.i_pipeline_s2_execute.cond_bge),
.i_pipeline__i_pipeline_s2_execute__cond_bgeu(
  i_pipeline.i_pipeline_s2_execute.cond_bgeu),
.i_pipeline__i_pipeline_s2_execute__cond_blt(
  i_pipeline.i_pipeline_s2_execute.cond_blt),
.i_pipeline__i_pipeline_s2_execute__cond_bltu(
  i_pipeline.i_pipeline_s2_execute.cond_bltu),
.i_pipeline__i_pipeline_s2_execute__cond_bne(
  i_pipeline.i_pipeline_s2_execute.cond_bne),
.i_pipeline__i_pipeline_s2_execute__imul_clmul(
  i_pipeline.i_pipeline_s2_execute.imul_clmul),
.i_pipeline__i_pipeline_s2_execute__imul_clmul_r(
  i_pipeline.i_pipeline_s2_execute.imul_clmul_r),
.i_pipeline__i_pipeline_s2_execute__imul_div(
  i_pipeline.i_pipeline_s2_execute.imul_div),
.i_pipeline__i_pipeline_s2_execute__imul_divu(
  i_pipeline.i_pipeline_s2_execute.imul_divu),
.i_pipeline__i_pipeline_s2_execute__imul_flush(
  i_pipeline.i_pipeline_s2_execute.imul_flush),
.i_pipeline__i_pipeline_s2_execute__imul_gpr_wide(
  i_pipeline.i_pipeline_s2_execute.imul_gpr_wide),
.i_pipeline__i_pipeline_s2_execute__imul_macc(
  i_pipeline.i_pipeline_s2_execute.imul_macc),
.i_pipeline__i_pipeline_s2_execute__imul_madd(
  i_pipeline.i_pipeline_s2_execute.imul_madd),
.i_pipeline__i_pipeline_s2_execute__imul_mmul(
  i_pipeline.i_pipeline_s2_execute.imul_mmul),
.i_pipeline__i_pipeline_s2_execute__imul_msub(
  i_pipeline.i_pipeline_s2_execute.imul_msub),
.i_pipeline__i_pipeline_s2_execute__imul_mul(
  i_pipeline.i_pipeline_s2_execute.imul_mul),
.i_pipeline__i_pipeline_s2_execute__imul_mulhsu(
  i_pipeline.i_pipeline_s2_execute.imul_mulhsu),
.i_pipeline__i_pipeline_s2_execute__imul_mulhu(
  i_pipeline.i_pipeline_s2_execute.imul_mulhu),
.i_pipeline__i_pipeline_s2_execute__imul_pclmul(
  i_pipeline.i_pipeline_s2_execute.imul_pclmul),
.i_pipeline__i_pipeline_s2_execute__imul_pmul(
  i_pipeline.i_pipeline_s2_execute.imul_pmul),
.i_pipeline__i_pipeline_s2_execute__imul_pw_16(
  i_pipeline.i_pipeline_s2_execute.imul_pw_16),
.i_pipeline__i_pipeline_s2_execute__imul_pw_2(
  i_pipeline.i_pipeline_s2_execute.imul_pw_2),
.i_pipeline__i_pipeline_s2_execute__imul_pw_32(
  i_pipeline.i_pipeline_s2_execute.imul_pw_32),
.i_pipeline__i_pipeline_s2_execute__imul_pw_4(
  i_pipeline.i_pipeline_s2_execute.imul_pw_4),
.i_pipeline__i_pipeline_s2_execute__imul_pw_8(
  i_pipeline.i_pipeline_s2_execute.imul_pw_8),
.i_pipeline__i_pipeline_s2_execute__imul_ready(
  i_pipeline.i_pipeline_s2_execute.imul_ready),
.i_pipeline__i_pipeline_s2_execute__imul_ready_t0(
  i_pipeline.i_pipeline_s2_execute.imul_ready_t0),
.i_pipeline__i_pipeline_s2_execute__imul_rem(
  i_pipeline.i_pipeline_s2_execute.imul_rem),
.i_pipeline__i_pipeline_s2_execute__imul_remu(
  i_pipeline.i_pipeline_s2_execute.imul_remu),
.i_pipeline__i_pipeline_s2_execute__imul_result(
  i_pipeline.i_pipeline_s2_execute.imul_result),
.i_pipeline__i_pipeline_s2_execute__imul_result_hi(
  i_pipeline.i_pipeline_s2_execute.imul_result_hi),
.i_pipeline__i_pipeline_s2_execute__imul_result_t0(
  i_pipeline.i_pipeline_s2_execute.imul_result_t0),
.i_pipeline__i_pipeline_s2_execute__imul_result_wide(
  i_pipeline.i_pipeline_s2_execute.imul_result_wide),
.i_pipeline__i_pipeline_s2_execute__imul_result_wide_t0(
  i_pipeline.i_pipeline_s2_execute.imul_result_wide_t0),
.i_pipeline__i_pipeline_s2_execute__leak_fence(
  i_pipeline.i_pipeline_s2_execute.leak_fence),
.i_pipeline__i_pipeline_s2_execute__lsu_load(
  i_pipeline.i_pipeline_s2_execute.lsu_load),
.i_pipeline__i_pipeline_s2_execute__lsu_store(
  i_pipeline.i_pipeline_s2_execute.lsu_store),
.i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_cfu(
  i_pipeline.i_pipeline_s2_execute.n_s3_opr_a_cfu),
.i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_cfu_t0(
  i_pipeline.i_pipeline_s2_execute.n_s3_opr_a_cfu_t0),
.i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_mul(
  i_pipeline.i_pipeline_s2_execute.n_s3_opr_a_mul),
.i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_mul_t0(
  i_pipeline.i_pipeline_s2_execute.n_s3_opr_a_mul_t0),
.i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_rng(
  i_pipeline.i_pipeline_s2_execute.n_s3_opr_a_rng),
.i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_rng_t0(
  i_pipeline.i_pipeline_s2_execute.n_s3_opr_a_rng_t0),
.i_pipeline__i_pipeline_s2_execute__n_s3_opr_b(
  i_pipeline.i_pipeline_s2_execute.n_s3_opr_b),
.i_pipeline__i_pipeline_s2_execute__n_s3_opr_b_t0(
  i_pipeline.i_pipeline_s2_execute.n_s3_opr_b_t0),
.i_pipeline__i_pipeline_s2_execute__n_s3_uop(
  i_pipeline.i_pipeline_s2_execute.n_s3_uop),
.i_pipeline__i_pipeline_s2_execute__n_s3_uop_cfu(
  i_pipeline.i_pipeline_s2_execute.n_s3_uop_cfu),
.i_pipeline__i_pipeline_s2_execute__n_s3_uop_cfu_t0(
  i_pipeline.i_pipeline_s2_execute.n_s3_uop_cfu_t0),
.i_pipeline__i_pipeline_s2_execute__n_s3_uop_t0(
  i_pipeline.i_pipeline_s2_execute.n_s3_uop_t0),
.i_pipeline__i_pipeline_s2_execute__opra_flush(
  i_pipeline.i_pipeline_s2_execute.opra_flush),
.i_pipeline__i_pipeline_s2_execute__opra_ld_en(
  i_pipeline.i_pipeline_s2_execute.opra_ld_en),
.i_pipeline__i_pipeline_s2_execute__oprb_flush(
  i_pipeline.i_pipeline_s2_execute.oprb_flush),
.i_pipeline__i_pipeline_s2_execute__oprb_ld_en(
  i_pipeline.i_pipeline_s2_execute.oprb_ld_en),
.i_pipeline__i_pipeline_s2_execute__p_busy(
  i_pipeline.i_pipeline_s2_execute.p_busy),
.i_pipeline__i_pipeline_s2_execute__p_busy_t0(
  i_pipeline.i_pipeline_s2_execute.p_busy_t0),
.i_pipeline__i_pipeline_s2_execute__p_valid(
  i_pipeline.i_pipeline_s2_execute.p_valid),
.i_pipeline__i_pipeline_s2_execute__pipe_reg_out(
  i_pipeline.i_pipeline_s2_execute.pipe_reg_out),
.i_pipeline__i_pipeline_s2_execute__pipe_reg_out_t0(
  i_pipeline.i_pipeline_s2_execute.pipe_reg_out_t0),
.i_pipeline__i_pipeline_s2_execute__rng_if_ready(
  i_pipeline.i_pipeline_s2_execute.rng_if_ready),
.i_pipeline__i_pipeline_s2_execute__rng_if_ready_t0(
  i_pipeline.i_pipeline_s2_execute.rng_if_ready_t0),
.i_pipeline__i_pipeline_s2_execute__rng_ready(
  i_pipeline.i_pipeline_s2_execute.rng_ready),
.i_pipeline__i_pipeline_s2_execute__rng_uop_samp(
  i_pipeline.i_pipeline_s2_execute.rng_uop_samp),
.i_pipeline__i_pipeline_s2_execute__rng_uop_seed(
  i_pipeline.i_pipeline_s2_execute.rng_uop_seed),
.i_pipeline__i_pipeline_s2_execute__rng_uop_test(
  i_pipeline.i_pipeline_s2_execute.rng_uop_test),
.i_pipeline__i_pipeline_s2_execute__rng_valid(
  i_pipeline.i_pipeline_s2_execute.rng_valid),
.i_pipeline__i_pipeline_s2_execute__i_alu__g_clk(
  i_pipeline.i_pipeline_s2_execute.i_alu.g_clk),
.i_pipeline__i_pipeline_s2_execute__i_alu__g_resetn(
  i_pipeline.i_pipeline_s2_execute.i_alu.g_resetn),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_valid(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_valid),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_flush(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_flush),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_ready(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_ready),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_pw(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_pw),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_add(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_add),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_sub(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_sub),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_xor(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_xor),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_or(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_or),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_and(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_and),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_shf),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_rot(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_rot),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf_left(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_shf_left),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf_arith(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_shf_arith),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_cmp(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_cmp),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_unsigned(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_unsigned),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_lt(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_lt),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_eq(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_eq),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_add_result(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_add_result),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_lhs(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_lhs),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_rhs(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_rhs),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_result(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_result),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_add_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_add_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_eq_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_eq_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_flush_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_flush_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_lhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_lhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_lt_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_lt_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_add_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_add_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_and_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_and_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_cmp_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_cmp_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_or_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_or_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_rot_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_rot_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_shf_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf_arith_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_shf_arith_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf_left_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_shf_left_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_sub_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_sub_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_unsigned_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_unsigned_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_xor_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_op_xor_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_pw_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_pw_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_lt_signed(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_lt_signed),
.i_pipeline__i_pipeline_s2_execute__i_alu__alu_lt_unsigned(
  i_pipeline.i_pipeline_s2_execute.i_alu.alu_lt_unsigned),
.i_pipeline__i_pipeline_s2_execute__i_alu__bw_result(
  i_pipeline.i_pipeline_s2_execute.i_alu.bw_result),
.i_pipeline__i_pipeline_s2_execute__i_alu__bw_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.bw_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__out_adder(
  i_pipeline.i_pipeline_s2_execute.i_alu.out_adder),
.i_pipeline__i_pipeline_s2_execute__i_alu__out_bw(
  i_pipeline.i_pipeline_s2_execute.i_alu.out_bw),
.i_pipeline__i_pipeline_s2_execute__i_alu__out_shift(
  i_pipeline.i_pipeline_s2_execute.i_alu.out_shift),
.i_pipeline__i_pipeline_s2_execute__i_alu__pw_d(
  i_pipeline.i_pipeline_s2_execute.i_alu.pw_d),
.i_pipeline__i_pipeline_s2_execute__i_alu__shift_arith(
  i_pipeline.i_pipeline_s2_execute.i_alu.shift_arith),
.i_pipeline__i_pipeline_s2_execute__i_alu__shift_arith_mask(
  i_pipeline.i_pipeline_s2_execute.i_alu.shift_arith_mask),
.i_pipeline__i_pipeline_s2_execute__i_alu__shift_arith_mask_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.shift_arith_mask_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__shift_out(
  i_pipeline.i_pipeline_s2_execute.i_alu.shift_out),
.i_pipeline__i_pipeline_s2_execute__i_alu__shift_out_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.shift_out_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__shift_result(
  i_pipeline.i_pipeline_s2_execute.i_alu.shift_result),
.i_pipeline__i_pipeline_s2_execute__i_alu__shift_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.shift_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__lhs(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.lhs),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__rhs(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.rhs),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__pw(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.pw),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__cin(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.cin),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__sub(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.sub),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__c_en(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.c_en),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__c_out(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.c_out),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__result(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.result),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__sub_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.sub_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__result_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.result_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__pw_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.pw_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__lhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.lhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__cin_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.cin_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__c_out_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.c_out_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__c_en_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.c_en_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__carry_mask(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.carry_mask),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__carry_mask_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.carry_mask_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_0___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[0].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_0___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[0].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_10___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[10].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_10___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[10].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_11___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[11].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_11___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[11].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_11___force_carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[11].force_carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_12___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[12].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_12___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[12].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_13___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[13].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_13___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[13].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_13___force_carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[13].force_carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_14___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[14].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_14___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[14].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_15___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[15].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_15___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[15].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_15___force_carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[15].force_carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_16___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[16].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_16___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[16].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_17___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[17].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_17___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[17].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_18___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[18].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_18___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[18].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_19___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[19].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_19___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[19].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_1___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[1].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_1___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[1].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_20___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[20].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_20___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[20].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_21___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[21].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_21___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[21].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_22___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[22].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_22___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[22].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_23___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[23].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_23___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[23].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_23___force_carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[23].force_carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_24___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[24].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_24___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[24].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_25___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[25].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_25___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[25].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_26___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[26].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_26___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[26].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_27___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[27].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_27___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[27].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_28___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[28].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_28___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[28].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_29___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[29].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_29___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[29].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_2___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[2].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_2___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[2].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_30___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[30].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_30___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[30].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_31___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[31].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_31___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[31].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_3___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[3].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_3___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[3].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_4___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[4].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_4___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[4].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_5___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[5].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_5___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[5].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_6___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[6].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_6___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[6].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_7___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[7].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_7___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[7].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_8___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[8].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_8___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[8].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_9___c_in(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[9].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_9___carry(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.\genblk1[9].carry ),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__rhs_m(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.rhs_m),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__rhs_m_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_addsub.rhs_m_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__crs1(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.crs1),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__shamt(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.shamt),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__pw(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.pw),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__shift(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.shift),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__rotate(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.rotate),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__left(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.left),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__right(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.right),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__result(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.result),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__shift_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.shift_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__shamt_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.shamt_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__rotate_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.rotate_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__right_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.right_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__left_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.left_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__crs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.crs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__result_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.result_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__pw_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.pw_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l1),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_16(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l16_16),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_16_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l16_16_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_32_left(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l16_32_left),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_32_left_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l16_32_left_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_32_right(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l16_32_right),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_32_right_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l16_32_right_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_16_left(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l1_16_left),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_16_right(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l1_16_right),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_2_left(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l1_2_left),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_2_right(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l1_2_right),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l1_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l2),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_16_left(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l2_16_left),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_16_left_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l2_16_left_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_16_right(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l2_16_right),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_16_right_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l2_16_right_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_2(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l2_2),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_2_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l2_2_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_4_left(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l2_4_left),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_4_left_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l2_4_left_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_4_right(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l2_4_right),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_4_right_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l2_4_right_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l2_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l4),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_16_left(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l4_16_left),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_16_left_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l4_16_left_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_16_right(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l4_16_right),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_16_right_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l4_16_right_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_2(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l4_2),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_2_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l4_2_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_8_left(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l4_8_left),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_8_left_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l4_8_left_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_8_right(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l4_8_right),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_8_right_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l4_8_right_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l4_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l8),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_16_left(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l8_16_left),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_16_left_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l8_16_left_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_16_right(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l8_16_right),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_16_right_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l8_16_right_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_2(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l8_2),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_2_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l8_2_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_t0(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.l8_t0),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_16(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l16_l_16),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_2(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l16_l_2),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_32(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l16_l_32),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_4(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l16_l_4),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_8(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l16_l_8),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_n_n(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l16_n_n),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_16(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l16_r_16),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_2(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l16_r_2),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_32(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l16_r_32),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_4(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l16_r_4),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_8(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l16_r_8),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_16(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l1_l_16),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_2(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l1_l_2),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_32(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l1_l_32),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_4(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l1_l_4),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_8(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l1_l_8),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_n_n(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l1_n_n),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_16(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l1_r_16),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_2(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l1_r_2),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_32(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l1_r_32),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_4(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l1_r_4),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_8(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l1_r_8),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_2(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l2_2),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_16(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l2_l_16),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_32(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l2_l_32),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_4(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l2_l_4),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_8(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l2_l_8),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_n_n(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l2_n_n),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_16(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l2_r_16),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_32(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l2_r_32),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_4(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l2_r_4),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_8(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l2_r_8),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_16(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l4_l_16),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_2(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l4_l_2),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_32(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l4_l_32),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_4(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l4_l_4),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_8(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l4_l_8),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_n_n(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l4_n_n),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_16(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l4_r_16),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_2(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l4_r_2),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_32(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l4_r_32),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_4(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l4_r_4),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_8(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l4_r_8),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_16(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l8_l_16),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_2(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l8_l_2),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_32(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l8_l_32),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_4(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l8_l_4),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_8(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l8_l_8),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_n_n(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l8_n_n),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_16(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l8_r_16),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_2(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l8_r_2),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_32(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l8_r_32),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_4(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l8_r_4),
.i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_8(
  i_pipeline.i_pipeline_s2_execute.i_alu.i_p_shfrot.ld_l8_r_8),
.i_pipeline__i_pipeline_s2_execute__i_asi__g_clk(
  i_pipeline.i_pipeline_s2_execute.i_asi.g_clk),
.i_pipeline__i_pipeline_s2_execute__i_asi__g_resetn(
  i_pipeline.i_pipeline_s2_execute.i_asi.g_resetn),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_valid(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_valid),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_ready(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_ready),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_aessub(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_flush_aessub),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_aesmix(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_flush_aesmix),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_data(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_flush_data),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_uop(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_uop),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_rs1(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_rs1),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_rs2(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_rs2),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_shamt(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_shamt),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_result(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_result),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_aesmix_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_flush_aesmix_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_aessub_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_flush_aessub_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_data_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_flush_data_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_rs2_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_rs2_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_shamt_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_shamt_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_uop_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_uop_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__asi_valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.asi_valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_enc(
  i_pipeline.i_pipeline_s2_execute.i_asi.aes_mix_enc),
.i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_ready(
  i_pipeline.i_pipeline_s2_execute.i_asi.aes_mix_ready),
.i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.aes_mix_ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_rs1(
  i_pipeline.i_pipeline_s2_execute.i_asi.aes_mix_rs1),
.i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.aes_mix_rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_rs2(
  i_pipeline.i_pipeline_s2_execute.i_asi.aes_mix_rs2),
.i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_rs2_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.aes_mix_rs2_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_ready(
  i_pipeline.i_pipeline_s2_execute.i_asi.aes_sub_ready),
.i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.aes_sub_ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_rs1(
  i_pipeline.i_pipeline_s2_execute.i_asi.aes_sub_rs1),
.i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.aes_sub_rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_rs2(
  i_pipeline.i_pipeline_s2_execute.i_asi.aes_sub_rs2),
.i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_rs2_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.aes_sub_rs2_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__insn_aes(
  i_pipeline.i_pipeline_s2_execute.i_asi.insn_aes),
.i_pipeline__i_pipeline_s2_execute__i_asi__insn_aes_mix(
  i_pipeline.i_pipeline_s2_execute.i_asi.insn_aes_mix),
.i_pipeline__i_pipeline_s2_execute__i_asi__insn_aes_sub(
  i_pipeline.i_pipeline_s2_execute.i_asi.insn_aes_sub),
.i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha2(
  i_pipeline.i_pipeline_s2_execute.i_asi.insn_sha2),
.i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3(
  i_pipeline.i_pipeline_s2_execute.i_asi.insn_sha3),
.i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_x1(
  i_pipeline.i_pipeline_s2_execute.i_asi.insn_sha3_x1),
.i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_x2(
  i_pipeline.i_pipeline_s2_execute.i_asi.insn_sha3_x2),
.i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_x4(
  i_pipeline.i_pipeline_s2_execute.i_asi.insn_sha3_x4),
.i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_xy(
  i_pipeline.i_pipeline_s2_execute.i_asi.insn_sha3_xy),
.i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_yx(
  i_pipeline.i_pipeline_s2_execute.i_asi.insn_sha3_yx),
.i_pipeline__i_pipeline_s2_execute__i_asi__result_aesmix(
  i_pipeline.i_pipeline_s2_execute.i_asi.result_aesmix),
.i_pipeline__i_pipeline_s2_execute__i_asi__result_aesmix_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.result_aesmix_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__result_aessub(
  i_pipeline.i_pipeline_s2_execute.i_asi.result_aessub),
.i_pipeline__i_pipeline_s2_execute__i_asi__result_aessub_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.result_aessub_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__result_sha2(
  i_pipeline.i_pipeline_s2_execute.i_asi.result_sha2),
.i_pipeline__i_pipeline_s2_execute__i_asi__result_sha2_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.result_sha2_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__result_sha3(
  i_pipeline.i_pipeline_s2_execute.i_asi.result_sha3),
.i_pipeline__i_pipeline_s2_execute__i_asi__result_sha3_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.result_sha3_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__sha2_rs1(
  i_pipeline.i_pipeline_s2_execute.i_asi.sha2_rs1),
.i_pipeline__i_pipeline_s2_execute__i_asi__sha2_rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.sha2_rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__clock(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.clock),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__reset(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.reset),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__flush(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.flush),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__flush_data(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.flush_data),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__valid(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.valid),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__rs1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.rs1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__rs2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.rs2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__enc(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.enc),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__ready(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.ready),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.result),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__flush_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.flush_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.result_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__rs2_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.rs2_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__flush_data_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.flush_data_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__enc_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.enc_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.d0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d0_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.d0_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.d1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d1_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.d1_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.d2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d2_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.d2_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.d3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d3_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.d3_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.e0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e0_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.e0_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.e1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e1_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.e1_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.e2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e2_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.e2_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.e3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e3_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.e3_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__mix_dec_0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\genblk1.mix_dec_0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__mix_dec_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\genblk1.mix_dec_0_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__mix_dec_1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\genblk1.mix_dec_1 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__mix_dec_1_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\genblk1.mix_dec_1_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__mix_dec_2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\genblk1.mix_dec_2 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__mix_dec_2_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\genblk1.mix_dec_2_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__mix_dec_3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\genblk1.mix_dec_3 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__mix_dec_3_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\genblk1.mix_dec_3_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__mix_enc_0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\genblk1.mix_enc_0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__mix_enc_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\genblk1.mix_enc_0_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__mix_enc_1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\genblk1.mix_enc_1 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__mix_enc_1_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\genblk1.mix_enc_1_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__mix_enc_2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\genblk1.mix_enc_2 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__mix_enc_2_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\genblk1.mix_enc_2_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__mix_enc_3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\genblk1.mix_enc_3 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__mix_enc_3_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\genblk1.mix_enc_3_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtime2_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_506_5988___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtime2$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:506$5988.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtime2_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_506_5988___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtime2$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:506$5988.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtime2_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_507_5990___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtime2$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:507$5990.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtime2_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_507_5990___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtime2$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:507$5990.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtime2_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_508_5992___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtime2$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:508$5992.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtime2_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_508_5992___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtime2$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:508$5992.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtime2_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_509_5994___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtime2$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:509$5994.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtime2_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_509_5994___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtime2$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:509$5994.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtime3_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_506_5989___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtime3$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:506$5989.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtime3_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_506_5989___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtime3$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:506$5989.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtime3_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_507_5991___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtime3$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:507$5991.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtime3_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_507_5991___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtime3$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:507$5991.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtime3_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_508_5993___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtime3$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:508$5993.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtime3_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_508_5993___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtime3$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:508$5993.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtime3_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_509_5995___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtime3$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:509$5995.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtime3_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_509_5995___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtime3$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:509$5995.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_511_5996___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:511$5996.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_511_5996___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:511$5996.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_511_5997___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:511$5997.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_511_5997___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:511$5997.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_511_5998___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:511$5998.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_511_5998___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:511$5998.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_511_5999___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:511$5999.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_511_5999___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:511$5999.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_512_6000___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:512$6000.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_512_6000___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:512$6000.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_512_6001___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:512$6001.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_512_6001___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:512$6001.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_512_6002___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:512$6002.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_512_6002___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:512$6002.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_512_6003___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:512$6003.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_512_6003___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:512$6003.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_513_6004___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:513$6004.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_513_6004___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:513$6004.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_513_6005___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:513$6005.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_513_6005___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:513$6005.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_513_6006___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:513$6006.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_513_6006___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:513$6006.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_513_6007___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:513$6007.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_513_6007___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:513$6007.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_514_6008___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:514$6008.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_514_6008___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:514$6008.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_514_6009___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:514$6009.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_514_6009___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:514$6009.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_514_6010___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:514$6010.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_514_6010___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:514$6010.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_514_6011___result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:514$6011.$result ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__xtimeN_func__data_kceesay_workspace_mucfi_cpus_scarv_scarv_unclocked_cellift_generated_sv2v_out__v_514_6011___result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aesmix.\xtimeN$func$/data/kceesay/workspace/mucfi/cpus/scarv/scarv_unclocked/cellift/generated/sv2v_out.v:514$6011.$result_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__clock(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.clock),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__reset(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.reset),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__flush(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.flush),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__flush_data(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.flush_data),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__valid(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.valid),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rs1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.rs1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rs2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.rs2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__enc(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.enc),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rot(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.rot),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__ready(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.ready),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.result),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__flush_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.flush_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.result_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rs2_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.rs2_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__flush_data_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.flush_data_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__enc_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.enc_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rot_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.rot_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sb_in_0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sb_in_0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sb_in_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sb_in_0_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sb_in_1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sb_in_1 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sb_in_1_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sb_in_1_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sb_in_2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sb_in_2 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sb_in_2_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sb_in_2_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sb_in_3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sb_in_3 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sb_in_3_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sb_in_3_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sb_out_0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sb_out_0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sb_out_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sb_out_0_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sb_out_1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sb_out_1 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sb_out_1_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sb_out_1_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sb_out_2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sb_out_2 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sb_out_2_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sb_out_2_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sb_out_3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sb_out_3 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sb_out_3_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sb_out_3_t0 ),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__in(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .in),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__inv(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .inv),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .out),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__in_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .in_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .out_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__inv_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .inv_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out_fwd(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .out_fwd),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out_fwd_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .out_fwd_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out_inv(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .out_inv),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out_inv_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .out_inv_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__in(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.in),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__out(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.out),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__in_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.in_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__out_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.out_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.s0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.s1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.s2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.s3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.s4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.s5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.s6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.s7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t15(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t15),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t17(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t17),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t18(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t18),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t19(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t19),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t20(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t20),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t21(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t21),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t22(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t22),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t23(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t23),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t24(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t24),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t25(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t25),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t26(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t26),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t27(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t27),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t28(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t28),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t29(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t29),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t30(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t30),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t31(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t31),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t32(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t32),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t33(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t33),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t34(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t34),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t35(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t35),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t36(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t36),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t37(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t37),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t38(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t38),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t39(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t39),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t40(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t40),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t41(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t41),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t42(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t42),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t43(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t43),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t44(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t44),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t45(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t45),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.t9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc17(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc17),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc18(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc18),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc20(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc20),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc21(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc21),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc26(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc26),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.tc9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y15(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y15),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y17(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y17),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y18(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y18),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y19(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y19),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y20(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y20),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y21(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y21),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.y9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z15(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z15),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z17(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z17),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_fwd.z9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__in(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.in),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__out(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.out),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__in_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.in_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__out_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.out_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__aa(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.aa),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.ab0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.ab1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.ab2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab20(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.ab20),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab21(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.ab21),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab22(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.ab22),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab23(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.ab23),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.ab3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.abcd1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.abcd2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.abcd3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.abcd4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.abcd5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.abcd6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ah(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.ah),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__al(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.al),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__bb(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.bb),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__bh(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.bh),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__bl(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.bl),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.cp1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.cp2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.cp3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.cp4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.d0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.d1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.d2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.d3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__dd(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.dd),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__dh(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.dh),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__dl(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.dl),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.p0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.p1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.p2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.p3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.p4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.p6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.p7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph01(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.ph01),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph02(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.ph02),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph03(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.ph03),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.ph11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.ph12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.ph13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl01(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.pl01),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl02(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.pl02),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl03(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.pl03),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.pl11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.pl12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.pl13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.pr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.pr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pr3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.pr3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__qr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.qr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__qr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.qr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__qr3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.qr3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.r1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.r10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.r11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.r2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.r3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.r4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.r5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.r6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.r7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.r8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.r9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.rr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.rr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rtl0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.rtl0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rtl1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.rtl1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rtl2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.rtl2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.s0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.s1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.s2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.s3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.s4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.s5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.s6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.s7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sa0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.sa0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sa1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.sa1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sb0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.sb0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sb1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.sb1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sd0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.sd0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sd1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.sd1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__t01(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.t01),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__t02(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.t02),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.tinv1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.tinv10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.tinv11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.tinv12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.tinv13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.tinv2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.tinv3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.tinv4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.tinv5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.tinv6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.tinv7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.tinv8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.tinv9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__vr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.vr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__vr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.vr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__vr3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.vr3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__wr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.wr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__wr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.wr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__wr3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.wr3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.x11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.x13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.x14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.x16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x18(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.x18),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x19(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.x19),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.y0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.y1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.y2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.y3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.y4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.y5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.y6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_0 .i_sbox_inv.y7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__in(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .in),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__inv(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .inv),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__out(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .out),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__in_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .in_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__out_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .out_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__inv_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .inv_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__out_fwd(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .out_fwd),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__out_fwd_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .out_fwd_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__out_inv(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .out_inv),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__out_inv_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .out_inv_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__in(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.in),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__out(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.out),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__in_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.in_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__out_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.out_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__s0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.s0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__s1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.s1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__s2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.s2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__s3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.s3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__s4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.s4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__s5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.s5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__s6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.s6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__s7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.s7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t15(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t15),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t17(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t17),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t18(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t18),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t19(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t19),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t20(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t20),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t21(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t21),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t22(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t22),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t23(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t23),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t24(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t24),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t25(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t25),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t26(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t26),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t27(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t27),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t28(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t28),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t29(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t29),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t30(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t30),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t31(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t31),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t32(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t32),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t33(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t33),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t34(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t34),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t35(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t35),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t36(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t36),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t37(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t37),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t38(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t38),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t39(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t39),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t40(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t40),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t41(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t41),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t42(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t42),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t43(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t43),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t44(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t44),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t45(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t45),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__t9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.t9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc17(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc17),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc18(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc18),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc20(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc20),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc21(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc21),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc26(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc26),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__tc9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.tc9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y15(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y15),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y17(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y17),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y18(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y18),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y19(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y19),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y20(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y20),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y21(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y21),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__y9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.y9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z15(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z15),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z17(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z17),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_fwd__z9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_fwd.z9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__in(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.in),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__out(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.out),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__in_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.in_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__out_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.out_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__aa(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.aa),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__ab0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.ab0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__ab1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.ab1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__ab2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.ab2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__ab20(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.ab20),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__ab21(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.ab21),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__ab22(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.ab22),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__ab23(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.ab23),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__ab3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.ab3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__abcd1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.abcd1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__abcd2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.abcd2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__abcd3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.abcd3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__abcd4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.abcd4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__abcd5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.abcd5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__abcd6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.abcd6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__ah(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.ah),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__al(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.al),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__bb(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.bb),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__bh(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.bh),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__bl(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.bl),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__cp1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.cp1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__cp2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.cp2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__cp3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.cp3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__cp4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.cp4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__d0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.d0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__d1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.d1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__d2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.d2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__d3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.d3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__dd(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.dd),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__dh(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.dh),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__dl(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.dl),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__p0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.p0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__p1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.p1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__p2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.p2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__p3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.p3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__p4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.p4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__p6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.p6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__p7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.p7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__ph01(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.ph01),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__ph02(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.ph02),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__ph03(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.ph03),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__ph11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.ph11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__ph12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.ph12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__ph13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.ph13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__pl01(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.pl01),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__pl02(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.pl02),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__pl03(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.pl03),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__pl11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.pl11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__pl12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.pl12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__pl13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.pl13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__pr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.pr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__pr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.pr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__pr3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.pr3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__qr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.qr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__qr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.qr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__qr3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.qr3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__r1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.r1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__r10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.r10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__r11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.r11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__r2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.r2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__r3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.r3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__r4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.r4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__r5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.r5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__r6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.r6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__r7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.r7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__r8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.r8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__r9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.r9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__rr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.rr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__rr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.rr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__rtl0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.rtl0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__rtl1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.rtl1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__rtl2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.rtl2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__s0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.s0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__s1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.s1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__s2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.s2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__s3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.s3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__s4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.s4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__s5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.s5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__s6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.s6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__s7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.s7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__sa0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.sa0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__sa1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.sa1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__sb0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.sb0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__sb1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.sb1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__sd0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.sd0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__sd1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.sd1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__t01(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.t01),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__t02(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.t02),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__tinv1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.tinv1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__tinv10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.tinv10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__tinv11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.tinv11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__tinv12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.tinv12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__tinv13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.tinv13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__tinv2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.tinv2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__tinv3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.tinv3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__tinv4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.tinv4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__tinv5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.tinv5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__tinv6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.tinv6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__tinv7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.tinv7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__tinv8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.tinv8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__tinv9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.tinv9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__vr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.vr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__vr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.vr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__vr3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.vr3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__wr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.wr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__wr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.wr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__wr3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.wr3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__x11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.x11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__x13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.x13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__x14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.x14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__x16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.x16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__x18(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.x18),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__x19(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.x19),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__y0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.y0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__y1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.y1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__y2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.y2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__y3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.y3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__y4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.y4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__y5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.y5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__y6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.y6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_1__i_sbox_inv__y7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_1 .i_sbox_inv.y7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__in(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .in),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__inv(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .inv),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__out(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .out),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__in_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .in_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__out_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .out_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__inv_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .inv_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__out_fwd(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .out_fwd),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__out_fwd_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .out_fwd_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__out_inv(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .out_inv),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__out_inv_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .out_inv_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__in(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.in),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__out(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.out),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__in_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.in_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__out_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.out_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__s0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.s0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__s1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.s1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__s2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.s2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__s3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.s3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__s4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.s4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__s5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.s5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__s6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.s6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__s7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.s7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t15(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t15),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t17(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t17),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t18(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t18),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t19(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t19),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t20(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t20),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t21(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t21),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t22(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t22),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t23(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t23),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t24(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t24),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t25(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t25),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t26(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t26),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t27(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t27),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t28(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t28),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t29(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t29),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t30(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t30),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t31(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t31),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t32(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t32),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t33(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t33),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t34(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t34),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t35(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t35),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t36(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t36),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t37(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t37),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t38(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t38),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t39(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t39),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t40(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t40),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t41(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t41),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t42(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t42),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t43(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t43),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t44(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t44),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t45(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t45),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__t9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.t9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc17(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc17),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc18(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc18),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc20(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc20),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc21(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc21),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc26(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc26),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__tc9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.tc9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y15(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y15),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y17(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y17),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y18(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y18),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y19(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y19),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y20(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y20),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y21(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y21),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__y9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.y9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z15(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z15),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z17(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z17),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_fwd__z9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_fwd.z9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__in(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.in),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__out(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.out),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__in_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.in_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__out_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.out_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__aa(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.aa),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__ab0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.ab0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__ab1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.ab1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__ab2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.ab2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__ab20(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.ab20),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__ab21(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.ab21),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__ab22(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.ab22),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__ab23(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.ab23),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__ab3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.ab3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__abcd1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.abcd1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__abcd2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.abcd2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__abcd3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.abcd3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__abcd4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.abcd4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__abcd5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.abcd5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__abcd6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.abcd6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__ah(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.ah),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__al(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.al),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__bb(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.bb),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__bh(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.bh),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__bl(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.bl),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__cp1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.cp1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__cp2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.cp2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__cp3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.cp3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__cp4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.cp4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__d0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.d0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__d1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.d1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__d2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.d2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__d3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.d3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__dd(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.dd),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__dh(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.dh),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__dl(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.dl),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__p0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.p0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__p1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.p1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__p2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.p2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__p3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.p3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__p4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.p4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__p6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.p6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__p7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.p7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__ph01(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.ph01),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__ph02(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.ph02),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__ph03(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.ph03),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__ph11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.ph11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__ph12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.ph12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__ph13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.ph13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__pl01(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.pl01),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__pl02(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.pl02),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__pl03(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.pl03),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__pl11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.pl11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__pl12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.pl12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__pl13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.pl13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__pr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.pr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__pr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.pr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__pr3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.pr3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__qr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.qr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__qr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.qr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__qr3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.qr3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__r1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.r1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__r10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.r10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__r11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.r11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__r2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.r2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__r3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.r3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__r4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.r4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__r5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.r5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__r6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.r6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__r7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.r7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__r8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.r8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__r9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.r9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__rr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.rr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__rr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.rr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__rtl0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.rtl0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__rtl1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.rtl1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__rtl2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.rtl2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__s0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.s0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__s1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.s1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__s2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.s2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__s3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.s3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__s4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.s4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__s5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.s5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__s6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.s6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__s7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.s7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__sa0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.sa0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__sa1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.sa1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__sb0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.sb0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__sb1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.sb1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__sd0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.sd0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__sd1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.sd1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__t01(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.t01),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__t02(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.t02),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__tinv1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.tinv1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__tinv10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.tinv10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__tinv11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.tinv11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__tinv12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.tinv12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__tinv13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.tinv13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__tinv2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.tinv2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__tinv3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.tinv3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__tinv4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.tinv4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__tinv5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.tinv5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__tinv6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.tinv6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__tinv7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.tinv7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__tinv8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.tinv8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__tinv9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.tinv9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__vr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.vr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__vr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.vr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__vr3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.vr3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__wr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.wr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__wr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.wr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__wr3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.wr3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__x11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.x11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__x13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.x13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__x14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.x14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__x16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.x16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__x18(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.x18),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__x19(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.x19),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__y0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.y0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__y1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.y1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__y2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.y2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__y3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.y3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__y4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.y4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__y5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.y5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__y6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.y6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_2__i_sbox_inv__y7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_2 .i_sbox_inv.y7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__in(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .in),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__inv(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .inv),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__out(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .out),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__in_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .in_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__out_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .out_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__inv_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .inv_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__out_fwd(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .out_fwd),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__out_fwd_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .out_fwd_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__out_inv(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .out_inv),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__out_inv_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .out_inv_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__in(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.in),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__out(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.out),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__in_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.in_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__out_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.out_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__s0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.s0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__s1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.s1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__s2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.s2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__s3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.s3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__s4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.s4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__s5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.s5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__s6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.s6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__s7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.s7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t15(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t15),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t17(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t17),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t18(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t18),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t19(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t19),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t20(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t20),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t21(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t21),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t22(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t22),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t23(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t23),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t24(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t24),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t25(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t25),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t26(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t26),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t27(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t27),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t28(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t28),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t29(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t29),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t30(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t30),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t31(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t31),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t32(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t32),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t33(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t33),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t34(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t34),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t35(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t35),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t36(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t36),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t37(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t37),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t38(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t38),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t39(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t39),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t40(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t40),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t41(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t41),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t42(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t42),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t43(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t43),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t44(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t44),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t45(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t45),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__t9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.t9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc17(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc17),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc18(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc18),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc20(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc20),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc21(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc21),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc26(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc26),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__tc9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.tc9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y15(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y15),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y17(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y17),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y18(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y18),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y19(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y19),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y20(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y20),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y21(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y21),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__y9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.y9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z15(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z15),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z17(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z17),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_fwd__z9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_fwd.z9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__in(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.in),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__out(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.out),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__in_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.in_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__out_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.out_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__aa(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.aa),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__ab0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.ab0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__ab1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.ab1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__ab2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.ab2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__ab20(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.ab20),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__ab21(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.ab21),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__ab22(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.ab22),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__ab23(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.ab23),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__ab3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.ab3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__abcd1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.abcd1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__abcd2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.abcd2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__abcd3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.abcd3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__abcd4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.abcd4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__abcd5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.abcd5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__abcd6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.abcd6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__ah(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.ah),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__al(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.al),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__bb(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.bb),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__bh(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.bh),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__bl(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.bl),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__cp1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.cp1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__cp2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.cp2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__cp3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.cp3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__cp4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.cp4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__d0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.d0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__d1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.d1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__d2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.d2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__d3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.d3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__dd(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.dd),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__dh(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.dh),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__dl(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.dl),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__p0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.p0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__p1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.p1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__p2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.p2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__p3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.p3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__p4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.p4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__p6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.p6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__p7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.p7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__ph01(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.ph01),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__ph02(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.ph02),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__ph03(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.ph03),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__ph11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.ph11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__ph12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.ph12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__ph13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.ph13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__pl01(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.pl01),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__pl02(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.pl02),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__pl03(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.pl03),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__pl11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.pl11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__pl12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.pl12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__pl13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.pl13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__pr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.pr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__pr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.pr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__pr3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.pr3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__qr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.qr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__qr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.qr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__qr3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.qr3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__r1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.r1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__r10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.r10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__r11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.r11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__r2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.r2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__r3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.r3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__r4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.r4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__r5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.r5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__r6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.r6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__r7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.r7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__r8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.r8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__r9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.r9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__rr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.rr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__rr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.rr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__rtl0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.rtl0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__rtl1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.rtl1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__rtl2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.rtl2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__s0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.s0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__s1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.s1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__s2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.s2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__s3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.s3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__s4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.s4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__s5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.s5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__s6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.s6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__s7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.s7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__sa0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.sa0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__sa1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.sa1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__sb0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.sb0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__sb1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.sb1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__sd0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.sd0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__sd1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.sd1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__t01(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.t01),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__t02(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.t02),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__tinv1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.tinv1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__tinv10(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.tinv10),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__tinv11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.tinv11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__tinv12(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.tinv12),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__tinv13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.tinv13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__tinv2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.tinv2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__tinv3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.tinv3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__tinv4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.tinv4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__tinv5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.tinv5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__tinv6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.tinv6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__tinv7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.tinv7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__tinv8(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.tinv8),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__tinv9(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.tinv9),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__vr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.vr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__vr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.vr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__vr3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.vr3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__wr1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.wr1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__wr2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.wr2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__wr3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.wr3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__x11(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.x11),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__x13(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.x13),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__x14(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.x14),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__x16(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.x16),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__x18(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.x18),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__x19(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.x19),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__y0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.y0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__y1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.y1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__y2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.y2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__y3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.y3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__y4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.y4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__y5(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.y5),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__y6(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.y6),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_3__i_sbox_inv__y7(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_aessub.\genblk1.sbox_3 .i_sbox_inv.y7),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__rs1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.rs1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__ss(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.ss),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.result),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.result_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__ss_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.ss_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.s0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s0_result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.s0_result),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s0_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.s0_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.s1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s1_result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.s1_result),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s1_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.s1_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.s2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s2_result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.s2_result),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s2_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.s2_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s3(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.s3),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s3_result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.s3_result),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s3_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha256.s3_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__rs1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.rs1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__rs2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.rs2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shamt(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.shamt),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_xy(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.f_xy),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.f_x1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.f_x2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x4(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.f_x4),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_yx(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.f_yx),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__result(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.result),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shamt_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.shamt_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__result_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.result_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__rs2_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.rs2_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x1_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.f_x1_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x2_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.f_x2_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x4_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.f_x4_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_xy_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.f_xy_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_yx_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.f_yx_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__in_x_plus(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.in_x_plus),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__in_y_plus(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.in_y_plus),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_in_lhs(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.lut_in_lhs),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_in_rhs(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.lut_in_rhs),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_out_lhs(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.lut_out_lhs),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_out_rhs(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.lut_out_rhs),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__result_sum(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.result_sum),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__result_sum_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.result_sum_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shf_1(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.shf_1),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shf_1_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.shf_1_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shf_2(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.shf_2),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shf_2_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.shf_2_t0),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__sum_rhs(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.sum_rhs),
.i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__sum_rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_asi.i_xc_sha3.sum_rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__g_clk(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.g_clk),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__g_resetn(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.g_resetn),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_data(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.i_data),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_valid(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.i_valid),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_busy(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.o_busy),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__mr_data(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.mr_data),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__flush(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.flush),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__flush_dat(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.flush_dat),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_data(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.o_data),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_valid(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.o_valid),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_busy(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.i_busy),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__flush_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.flush_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.o_valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_data_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.o_data_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_busy_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.o_busy_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__mr_data_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.mr_data_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.i_valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_data_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.i_data_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_busy_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.i_busy_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__flush_dat_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.flush_dat_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__genblk1__progress(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg.\genblk1.progress ),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__g_clk(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.g_clk),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__g_resetn(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.g_resetn),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_data(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.i_data),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_valid(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.i_valid),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_busy(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.o_busy),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__mr_data(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.mr_data),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__flush(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.flush),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__flush_dat(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.flush_dat),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_data(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.o_data),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_valid(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.o_valid),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_busy(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.i_busy),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__flush_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.flush_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.o_valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_data_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.o_data_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_busy_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.o_busy_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__mr_data_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.mr_data_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.i_valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_data_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.i_data_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_busy_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.i_busy_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__flush_dat_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.flush_dat_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__genblk1__progress(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_a.\genblk1.progress ),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__g_clk(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.g_clk),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__g_resetn(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.g_resetn),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_data(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.i_data),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_valid(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.i_valid),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_busy(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.o_busy),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__mr_data(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.mr_data),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__flush(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.flush),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__flush_dat(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.flush_dat),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_data(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.o_data),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_valid(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.o_valid),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_busy(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.i_busy),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__flush_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.flush_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.o_valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_data_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.o_data_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_busy_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.o_busy_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__mr_data_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.mr_data_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.i_valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_data_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.i_data_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_busy_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.i_busy_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__flush_dat_t0(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.flush_dat_t0),
.i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__genblk1__progress(
  i_pipeline.i_pipeline_s2_execute.i_execute_pipe_reg_opr_b.\genblk1.progress ),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs1(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rs1),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs2(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rs2),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs3(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rs3),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__bop_lut(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.bop_lut),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__flush(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.flush),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__valid(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.valid),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_fsl(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.uop_fsl),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_fsr(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.uop_fsr),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_mror(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.uop_mror),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_cmov(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.uop_cmov),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_lut(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.uop_lut),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_bop(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.uop_bop),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.result),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__ready(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.ready),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__flush_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.flush_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.result_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs2_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rs2_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs3_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rs3_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__bop_lut_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.bop_lut_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_bop_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.uop_bop_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_cmov_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.uop_cmov_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_fsl_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.uop_fsl_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_fsr_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.uop_fsr_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_lut_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.uop_lut_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_mror_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.uop_mror_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__r_in(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.r_in),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__r_in_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.r_in_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__r_out(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.r_out),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__r_out_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.r_out_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__ramt(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.ramt),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_bop(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.result_bop),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_bop_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.result_bop_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_cmov(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.result_cmov),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_cmov_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.result_cmov_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_fsl(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.result_fsl),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_lut(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.result_lut),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_lut_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.result_lut_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rt_0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rt_0_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_1(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rt_1),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_1_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rt_1_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_2(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rt_2),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_2_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rt_2_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_3(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rt_3),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_3_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rt_3_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_4(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rt_4),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_4_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rt_4_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_5(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rt_5),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_5_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rt_5_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rword_l(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rword_l),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rword_l_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.rword_l_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs1(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk2.i_b_lut .crs1),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs2(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk2.i_b_lut .crs2),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs3(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk2.i_b_lut .crs3),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__result(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk2.i_b_lut .result),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk2.i_b_lut .crs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__result_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk2.i_b_lut .result_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs2_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk2.i_b_lut .crs2_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs3_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk2.i_b_lut .crs3_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rd(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk3.i_b_bop .rd),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rs1(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk3.i_b_bop .rs1),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rs2(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk3.i_b_bop .rs2),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__lut(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk3.i_b_bop .lut),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__result(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk3.i_b_bop .result),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__result_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk3.i_b_bop .result_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk3.i_b_bop .rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rs2_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk3.i_b_bop .rs2_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__lut_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk3.i_b_bop .lut_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rd_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_bitwise.\genblk3.i_b_bop .rd_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__g_clk(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.g_clk),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__g_resetn(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.g_resetn),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__flush(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.flush),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__pipeline_progress(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.pipeline_progress),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__valid(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.valid),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rs1(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rs1),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_valid(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rng_req_valid),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_op(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rng_req_op),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_data(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rng_req_data),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_ready(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rng_req_ready),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_valid(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rng_rsp_valid),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_status(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rng_rsp_status),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_data(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rng_rsp_data),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_ready(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rng_rsp_ready),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_test(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.uop_test),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_seed(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.uop_seed),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_samp(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.uop_samp),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__result(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.result),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__ready(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.ready),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__flush_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.flush_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__result_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.result_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__pipeline_progress_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.pipeline_progress_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_data_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rng_req_data_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_op_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rng_req_op_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rng_req_ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rng_req_valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_data_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rng_rsp_data_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rng_rsp_ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_status_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rng_rsp_status_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.rng_rsp_valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_samp_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.uop_samp_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_seed_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.uop_seed_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_test_t0(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.uop_test_t0),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__n_req_done(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.n_req_done),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__req_done(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.req_done),
.i_pipeline__i_pipeline_s2_execute__i_frv_rngif__status_healthy(
  i_pipeline.i_pipeline_s2_execute.i_frv_rngif.status_healthy),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__clock(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.clock),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__resetn(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.resetn),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs1(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.rs1),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs2(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.rs2),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs3(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.rs3),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__flush(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.flush),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__flush_data(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.flush_data),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__valid(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.valid),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_div(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_div),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_divu(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_divu),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_rem(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_rem),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_remu(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_remu),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mul(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_mul),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mulu(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_mulu),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mulsu(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_mulsu),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_clmul(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_clmul),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_pmul(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_pmul),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_pclmul(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_pclmul),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_madd(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_madd),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_msub(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_msub),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_macc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_macc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mmul(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_mmul),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_32(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.pw_32),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_16(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.pw_16),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_8(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.pw_8),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_4(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.pw_4),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_2(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.pw_2),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__result(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.result),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__ready(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.ready),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__flush_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.flush_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__result_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.result_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mul_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_mul_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_16_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.pw_16_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_2_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.pw_2_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_32_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.pw_32_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_4_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.pw_4_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_8_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.pw_8_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs2_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.rs2_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs3_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.rs3_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_macc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_macc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_madd_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_madd_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mmul_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_mmul_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_msub_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_msub_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__flush_data_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.flush_data_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_clmul_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_clmul_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_div_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_div_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_divu_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_divu_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mulsu_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_mulsu_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mulu_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_mulu_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_pclmul_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_pclmul_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_pmul_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_pmul_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_rem_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_rem_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_remu_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.uop_remu_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__arg_0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.arg_0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__arg_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.arg_0_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__arg_1(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.arg_1),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__arg_1_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.arg_1_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.carry),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__carry_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.carry_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__count(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.count),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__count_en(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.count_en),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__count_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.count_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__do_mulu(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.do_mulu),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__fsm(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.fsm),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__insn_divrem(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.insn_divrem),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__insn_long(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.insn_long),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__insn_mdr(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.insn_mdr),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__ld_long(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.ld_long),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__ld_mdr(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.ld_mdr),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__ld_on_init(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.ld_on_init),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_n_acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.long_n_acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_n_acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.long_n_acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_n_carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.long_n_carry),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_n_carry_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.long_n_carry_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_cin(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.long_padd_cin),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_cin_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.long_padd_cin_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_lhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.long_padd_lhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_lhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.long_padd_lhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_rhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.long_padd_rhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.long_padd_rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_sub(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.long_padd_sub),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_sub_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.long_padd_sub_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_ready(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.long_ready),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.long_ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_result(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.long_result),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.long_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_n_acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_n_acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_arg_0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_n_arg_0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_arg_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_n_arg_0_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_arg_1(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_n_arg_1),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_arg_1_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_n_arg_1_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_cen(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_padd_cen),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_cen_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_padd_cen_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_cin(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_padd_cin),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_cin_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_padd_cin_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_lhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_padd_lhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_lhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_padd_lhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_rhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_padd_rhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_padd_rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_sub(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_padd_sub),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_sub_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_padd_sub_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_ready(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_ready),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_result(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_result),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.mdr_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.n_acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.n_acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_arg_0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.n_arg_0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_arg_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.n_arg_0_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.n_carry),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_count(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.n_count),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_count_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.n_count_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_fsm(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.n_fsm),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_cen(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.padd_cen),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_cin(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.padd_cin),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_cout(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.padd_cout),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_cout_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.padd_cout_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_lhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.padd_lhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_lhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.padd_lhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_result(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.padd_result),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.padd_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_rhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.padd_rhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.padd_rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_sub(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.padd_sub),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__reg_ld_en(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.reg_ld_en),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__clock(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.clock),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__resetn(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.resetn),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs1(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.rs1),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs2(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.rs2),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs3(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.rs3),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__flush(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.flush),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__valid(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.valid),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_div(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_div),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_divu(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_divu),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_rem(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_rem),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_remu(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_remu),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mul(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_mul),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mulu(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_mulu),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mulsu(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_mulsu),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_clmul(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_clmul),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_pmul(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_pmul),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_pclmul(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_pclmul),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_32(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pw_32),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_16(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pw_16),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_8(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pw_8),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_4(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pw_4),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_2(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pw_2),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__count(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.count),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.arg_0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_1(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.arg_1),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.n_acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_arg_0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.n_arg_0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_arg_1(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.n_arg_1),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_lhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.padd_lhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_rhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.padd_rhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_sub(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.padd_sub),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cin(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.padd_cin),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cen(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.padd_cen),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cout(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.padd_cout),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_result(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.padd_result),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__result(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.result),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__ready(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.ready),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__flush_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.flush_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__result_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.result_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.arg_0_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__count_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.count_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.n_acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_arg_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.n_arg_0_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cen_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.padd_cen_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cin_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.padd_cin_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cout_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.padd_cout_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_lhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.padd_lhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.padd_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.padd_rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_sub_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.padd_sub_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_16_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pw_16_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_2_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pw_2_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_32_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pw_32_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_4_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pw_4_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_8_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pw_8_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs2_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.rs2_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_1_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.arg_1_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_arg_1_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.n_arg_1_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_clmul_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_clmul_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_div_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_div_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_divu_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_divu_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mul_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_mul_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mulsu_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_mulsu_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mulu_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_mulu_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_pclmul_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_pclmul_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_pmul_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_pmul_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_rem_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_rem_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_remu_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.do_remu_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs3_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.rs3_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_sel(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.arg_sel),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_sel_neg(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.arg_sel_neg),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_sel_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.arg_sel_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_n_acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.div_n_acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_n_acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.div_n_acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_n_arg_0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.div_n_arg_0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_n_arg_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.div_n_arg_0_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_outsign(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.div_outsign),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_ready(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.div_ready),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.div_ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_signed(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.div_signed),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__divrem_result(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.divrem_result),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__divrem_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.divrem_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_carryless(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_carryless),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_lhs_sign(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_lhs_sign),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_n_acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_n_acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_n_acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_n_acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_n_arg_0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_n_arg_0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_n_arg_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_n_arg_0_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_cen(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_padd_cen),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_cen_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_padd_cen_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_cin(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_padd_cin),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_cin_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_padd_cin_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_lhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_padd_lhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_lhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_padd_lhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_rhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_padd_rhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_padd_rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_sub(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_padd_sub),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_sub_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_padd_sub_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_ready(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_ready),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.mul_ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_n_acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pmul_n_acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_n_acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pmul_n_acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_n_arg_0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pmul_n_arg_0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_n_arg_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pmul_n_arg_0_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_cen(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pmul_padd_cen),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_cen_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pmul_padd_cen_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_lhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pmul_padd_lhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_lhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pmul_padd_lhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_rhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pmul_padd_rhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pmul_padd_rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_sub(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pmul_padd_sub),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_sub_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pmul_padd_sub_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_ready(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pmul_ready),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pmul_ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_result(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pmul_result),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.pmul_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rem_outsign(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.rem_outsign),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__result_div(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.result_div),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__result_rem(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.result_rem),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__route_div(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.route_div),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__route_mul(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.route_mul),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__route_pmul(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.route_pmul),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__rs1(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.rs1),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__rs2(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.rs2),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__count(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.count),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__arg_0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.arg_0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__carryless(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.carryless),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_16(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.pw_16),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_8(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.pw_8),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_4(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.pw_4),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_2(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.pw_2),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_lhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.padd_lhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_rhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.padd_rhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_sub(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.padd_sub),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_cen(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.padd_cen),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_cout(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.padd_cout),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_result(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.padd_result),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__n_acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.n_acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__n_arg_0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.n_arg_0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__result(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.result),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__ready(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.ready),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__result_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.result_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__arg_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.arg_0_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__carryless_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.carryless_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__count_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.count_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__n_acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.n_acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__n_arg_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.n_arg_0_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_cen_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.padd_cen_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_cout_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.padd_cout_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_lhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.padd_lhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.padd_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.padd_rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_sub_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.padd_sub_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_16_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.pw_16_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_2_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.pw_2_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_4_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.pw_4_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_8_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.pw_8_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__rs2_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.rs2_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_mask(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.padd_mask),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_mask_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.padd_mask_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pmul_result_0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.pmul_result_0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pmul_result_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_malu_pmul.pmul_result_0_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__clock(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.clock),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__resetn(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.resetn),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__rs1(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.rs1),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__rs2(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.rs2),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__valid(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.valid),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__op_signed(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.op_signed),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__flush(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.flush),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__count(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.count),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__arg_0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.arg_0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__arg_1(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.arg_1),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.n_acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_arg_0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.n_arg_0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_arg_1(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.n_arg_1),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__ready(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.ready),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__flush_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.flush_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__arg_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.arg_0_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__count_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.count_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.n_acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_arg_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.n_arg_0_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__rs2_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.rs2_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__arg_1_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.arg_1_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_arg_1_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.n_arg_1_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__op_signed_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.op_signed_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__valid_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.valid_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__div_less(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.div_less),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__div_run(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.div_run),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__div_start(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.div_start),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__divisor_start(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.divisor_start),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__divisor_start_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.divisor_start_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__qmask(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.qmask),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__qmask_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.qmask_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__signed_lhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.signed_lhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__signed_rhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.signed_rhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__sub_result(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.sub_result),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__sub_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_divrem.sub_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rs1(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.rs1),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rs2(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.rs2),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__count(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.count),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__arg_0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.arg_0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__carryless(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.carryless),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_32(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.pw_32),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_16(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.pw_16),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_8(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.pw_8),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_4(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.pw_4),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_2(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.pw_2),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__lhs_sign(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.lhs_sign),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rhs_sign(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.rhs_sign),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_lhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.padd_lhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_rhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.padd_rhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_sub(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.padd_sub),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cin(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.padd_cin),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cen(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.padd_cen),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cout(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.padd_cout),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_result(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.padd_result),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__n_acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.n_acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__n_arg_0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.n_arg_0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__ready(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.ready),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__arg_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.arg_0_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__carryless_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.carryless_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__count_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.count_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__lhs_sign_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.lhs_sign_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__n_acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.n_acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__n_arg_0_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.n_arg_0_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cen_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.padd_cen_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cin_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.padd_cin_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cout_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.padd_cout_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_lhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.padd_lhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.padd_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.padd_rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_sub_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.padd_sub_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_16_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.pw_16_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_2_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.pw_2_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_32_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.pw_32_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_4_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.pw_4_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_8_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.pw_8_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rhs_sign_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.rhs_sign_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rs2_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.rs2_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_32(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.add_32),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_32_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.add_32_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_lhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.add_lhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_rhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.add_rhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_malu_muldivrem.i_xc_malu_mul.add_rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__lhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.lhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__rhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.rhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__pw(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.pw),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__cin(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.cin),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__sub(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.sub),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__c_en(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.c_en),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__c_out(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.c_out),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__result(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.result),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__sub_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.sub_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__result_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.result_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__pw_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.pw_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__lhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.lhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__cin_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.cin_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__c_out_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.c_out_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__c_en_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.c_en_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__carry_mask(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.carry_mask),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__carry_mask_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.carry_mask_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_0___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[0].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_0___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[0].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_10___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[10].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_10___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[10].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_11___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[11].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_11___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[11].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_11___force_carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[11].force_carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_12___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[12].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_12___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[12].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_13___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[13].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_13___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[13].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_13___force_carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[13].force_carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_14___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[14].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_14___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[14].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_15___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[15].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_15___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[15].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_15___force_carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[15].force_carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_16___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[16].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_16___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[16].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_17___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[17].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_17___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[17].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_18___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[18].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_18___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[18].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_19___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[19].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_19___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[19].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_1___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[1].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_1___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[1].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_20___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[20].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_20___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[20].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_21___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[21].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_21___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[21].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_22___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[22].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_22___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[22].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_23___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[23].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_23___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[23].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_23___force_carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[23].force_carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_24___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[24].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_24___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[24].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_25___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[25].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_25___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[25].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_26___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[26].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_26___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[26].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_27___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[27].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_27___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[27].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_28___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[28].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_28___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[28].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_29___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[29].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_29___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[29].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_2___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[2].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_2___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[2].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_30___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[30].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_30___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[30].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_31___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[31].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_31___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[31].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_3___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[3].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_3___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[3].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_4___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[4].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_4___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[4].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_5___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[5].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_5___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[5].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_6___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[6].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_6___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[6].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_7___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[7].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_7___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[7].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_8___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[8].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_8___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[8].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_9___c_in(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[9].c_in ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_9___carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.\genblk1[9].carry ),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__rhs_m(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.rhs_m),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__rhs_m_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_p_addsub.rhs_m_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs1(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.rs1),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs2(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.rs2),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs3(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.rs3),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_init(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.fsm_init),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mdr(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.fsm_mdr),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_msub_1(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.fsm_msub_1),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_macc_1(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.fsm_macc_1),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mmul_1(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.fsm_mmul_1),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mmul_2(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.fsm_mmul_2),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_done(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.fsm_done),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.carry),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__count(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.count),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_lhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.padd_lhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_rhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.padd_rhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_cin(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.padd_cin),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_sub(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.padd_sub),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_cout(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.padd_cout),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_result(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.padd_result),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_madd(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.uop_madd),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_msub(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.uop_msub),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_macc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.uop_macc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_mmul(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.uop_mmul),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__n_carry(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.n_carry),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__n_acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.n_acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__result(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.result),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__ready(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.ready),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__result_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.result_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__count_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.count_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__n_acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.n_acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_cin_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.padd_cin_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_cout_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.padd_cout_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_lhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.padd_lhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.padd_result_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.padd_rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_sub_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.padd_sub_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__ready_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.ready_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs1_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.rs1_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs2_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.rs2_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs3_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.rs3_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__carry_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.carry_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_done_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.fsm_done_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_init_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.fsm_init_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_macc_1_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.fsm_macc_1_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mdr_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.fsm_mdr_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mmul_1_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.fsm_mmul_1_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mmul_2_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.fsm_mmul_2_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_msub_1_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.fsm_msub_1_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__n_carry_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.n_carry_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_macc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.uop_macc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_madd_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.uop_madd_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_mmul_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.uop_mmul_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_msub_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.uop_msub_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_lhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.macc_lhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_lhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.macc_lhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_n_acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.macc_n_acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_n_acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.macc_n_acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_rhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.macc_rhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.macc_rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_lhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.mmul_lhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_lhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.mmul_lhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_n_acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.mmul_n_acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_n_acc_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.mmul_n_acc_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_rhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.mmul_rhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.mmul_rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__msub_lhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.msub_lhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__msub_lhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.msub_lhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__msub_rhs(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.msub_rhs),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__msub_rhs_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.msub_rhs_t0),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__result_acc(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.result_acc),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__sub_result(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.sub_result),
.i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__sub_result_t0(
  i_pipeline.i_pipeline_s2_execute.i_xc_malu.i_xc_malu_long.sub_result_t0),
.i_pipeline__i_pipeline_s3_memory__g_clk(
  i_pipeline.i_pipeline_s3_memory.g_clk),
.i_pipeline__i_pipeline_s3_memory__g_resetn(
  i_pipeline.i_pipeline_s3_memory.g_resetn),
.i_pipeline__i_pipeline_s3_memory__flush(
  i_pipeline.i_pipeline_s3_memory.flush),
.i_pipeline__i_pipeline_s3_memory__s3_rd(
  i_pipeline.i_pipeline_s3_memory.s3_rd),
.i_pipeline__i_pipeline_s3_memory__s3_opr_a(
  i_pipeline.i_pipeline_s3_memory.s3_opr_a),
.i_pipeline__i_pipeline_s3_memory__s3_opr_b(
  i_pipeline.i_pipeline_s3_memory.s3_opr_b),
.i_pipeline__i_pipeline_s3_memory__s3_uop(
  i_pipeline.i_pipeline_s3_memory.s3_uop),
.i_pipeline__i_pipeline_s3_memory__s3_fu(
  i_pipeline.i_pipeline_s3_memory.s3_fu),
.i_pipeline__i_pipeline_s3_memory__s3_trap(
  i_pipeline.i_pipeline_s3_memory.s3_trap),
.i_pipeline__i_pipeline_s3_memory__s3_size(
  i_pipeline.i_pipeline_s3_memory.s3_size),
.i_pipeline__i_pipeline_s3_memory__s3_instr(
  i_pipeline.i_pipeline_s3_memory.s3_instr),
.i_pipeline__i_pipeline_s3_memory__s3_busy(
  i_pipeline.i_pipeline_s3_memory.s3_busy),
.i_pipeline__i_pipeline_s3_memory__s3_valid(
  i_pipeline.i_pipeline_s3_memory.s3_valid),
.i_pipeline__i_pipeline_s3_memory__leak_prng(
  i_pipeline.i_pipeline_s3_memory.leak_prng),
.i_pipeline__i_pipeline_s3_memory__leak_lkgcfg(
  i_pipeline.i_pipeline_s3_memory.leak_lkgcfg),
.i_pipeline__i_pipeline_s3_memory__leak_fence_unc0(
  i_pipeline.i_pipeline_s3_memory.leak_fence_unc0),
.i_pipeline__i_pipeline_s3_memory__leak_fence_unc1(
  i_pipeline.i_pipeline_s3_memory.leak_fence_unc1),
.i_pipeline__i_pipeline_s3_memory__leak_fence_unc2(
  i_pipeline.i_pipeline_s3_memory.leak_fence_unc2),
.i_pipeline__i_pipeline_s3_memory__fwd_s3_rd(
  i_pipeline.i_pipeline_s3_memory.fwd_s3_rd),
.i_pipeline__i_pipeline_s3_memory__fwd_s3_wide(
  i_pipeline.i_pipeline_s3_memory.fwd_s3_wide),
.i_pipeline__i_pipeline_s3_memory__fwd_s3_wdata(
  i_pipeline.i_pipeline_s3_memory.fwd_s3_wdata),
.i_pipeline__i_pipeline_s3_memory__fwd_s3_wdata_hi(
  i_pipeline.i_pipeline_s3_memory.fwd_s3_wdata_hi),
.i_pipeline__i_pipeline_s3_memory__fwd_s3_load(
  i_pipeline.i_pipeline_s3_memory.fwd_s3_load),
.i_pipeline__i_pipeline_s3_memory__fwd_s3_csr(
  i_pipeline.i_pipeline_s3_memory.fwd_s3_csr),
.i_pipeline__i_pipeline_s3_memory__hold_lsu_req(
  i_pipeline.i_pipeline_s3_memory.hold_lsu_req),
.i_pipeline__i_pipeline_s3_memory__mmio_en(
  i_pipeline.i_pipeline_s3_memory.mmio_en),
.i_pipeline__i_pipeline_s3_memory__mmio_wen(
  i_pipeline.i_pipeline_s3_memory.mmio_wen),
.i_pipeline__i_pipeline_s3_memory__mmio_addr(
  i_pipeline.i_pipeline_s3_memory.mmio_addr),
.i_pipeline__i_pipeline_s3_memory__mmio_wdata(
  i_pipeline.i_pipeline_s3_memory.mmio_wdata),
.i_pipeline__i_pipeline_s3_memory__dmem_req(
  i_pipeline.i_pipeline_s3_memory.dmem_req),
.i_pipeline__i_pipeline_s3_memory__dmem_wen(
  i_pipeline.i_pipeline_s3_memory.dmem_wen),
.i_pipeline__i_pipeline_s3_memory__dmem_strb(
  i_pipeline.i_pipeline_s3_memory.dmem_strb),
.i_pipeline__i_pipeline_s3_memory__dmem_wdata(
  i_pipeline.i_pipeline_s3_memory.dmem_wdata),
.i_pipeline__i_pipeline_s3_memory__dmem_addr(
  i_pipeline.i_pipeline_s3_memory.dmem_addr),
.i_pipeline__i_pipeline_s3_memory__dmem_gnt(
  i_pipeline.i_pipeline_s3_memory.dmem_gnt),
.i_pipeline__i_pipeline_s3_memory__s4_rd(
  i_pipeline.i_pipeline_s3_memory.s4_rd),
.i_pipeline__i_pipeline_s3_memory__s4_opr_a(
  i_pipeline.i_pipeline_s3_memory.s4_opr_a),
.i_pipeline__i_pipeline_s3_memory__s4_opr_b(
  i_pipeline.i_pipeline_s3_memory.s4_opr_b),
.i_pipeline__i_pipeline_s3_memory__s4_uop(
  i_pipeline.i_pipeline_s3_memory.s4_uop),
.i_pipeline__i_pipeline_s3_memory__s4_fu(
  i_pipeline.i_pipeline_s3_memory.s4_fu),
.i_pipeline__i_pipeline_s3_memory__s4_trap(
  i_pipeline.i_pipeline_s3_memory.s4_trap),
.i_pipeline__i_pipeline_s3_memory__s4_size(
  i_pipeline.i_pipeline_s3_memory.s4_size),
.i_pipeline__i_pipeline_s3_memory__s4_instr(
  i_pipeline.i_pipeline_s3_memory.s4_instr),
.i_pipeline__i_pipeline_s3_memory__s4_busy(
  i_pipeline.i_pipeline_s3_memory.s4_busy),
.i_pipeline__i_pipeline_s3_memory__s4_valid(
  i_pipeline.i_pipeline_s3_memory.s4_valid),
.i_pipeline__i_pipeline_s3_memory__flush_t0(
  i_pipeline.i_pipeline_s3_memory.flush_t0),
.i_pipeline__i_pipeline_s3_memory__leak_lkgcfg_t0(
  i_pipeline.i_pipeline_s3_memory.leak_lkgcfg_t0),
.i_pipeline__i_pipeline_s3_memory__leak_prng_t0(
  i_pipeline.i_pipeline_s3_memory.leak_prng_t0),
.i_pipeline__i_pipeline_s3_memory__mmio_wen_t0(
  i_pipeline.i_pipeline_s3_memory.mmio_wen_t0),
.i_pipeline__i_pipeline_s3_memory__mmio_wdata_t0(
  i_pipeline.i_pipeline_s3_memory.mmio_wdata_t0),
.i_pipeline__i_pipeline_s3_memory__mmio_en_t0(
  i_pipeline.i_pipeline_s3_memory.mmio_en_t0),
.i_pipeline__i_pipeline_s3_memory__mmio_addr_t0(
  i_pipeline.i_pipeline_s3_memory.mmio_addr_t0),
.i_pipeline__i_pipeline_s3_memory__s3_busy_t0(
  i_pipeline.i_pipeline_s3_memory.s3_busy_t0),
.i_pipeline__i_pipeline_s3_memory__s3_fu_t0(
  i_pipeline.i_pipeline_s3_memory.s3_fu_t0),
.i_pipeline__i_pipeline_s3_memory__s3_instr_t0(
  i_pipeline.i_pipeline_s3_memory.s3_instr_t0),
.i_pipeline__i_pipeline_s3_memory__s3_opr_a_t0(
  i_pipeline.i_pipeline_s3_memory.s3_opr_a_t0),
.i_pipeline__i_pipeline_s3_memory__s3_opr_b_t0(
  i_pipeline.i_pipeline_s3_memory.s3_opr_b_t0),
.i_pipeline__i_pipeline_s3_memory__s3_rd_t0(
  i_pipeline.i_pipeline_s3_memory.s3_rd_t0),
.i_pipeline__i_pipeline_s3_memory__s3_size_t0(
  i_pipeline.i_pipeline_s3_memory.s3_size_t0),
.i_pipeline__i_pipeline_s3_memory__s3_trap_t0(
  i_pipeline.i_pipeline_s3_memory.s3_trap_t0),
.i_pipeline__i_pipeline_s3_memory__s3_uop_t0(
  i_pipeline.i_pipeline_s3_memory.s3_uop_t0),
.i_pipeline__i_pipeline_s3_memory__s3_valid_t0(
  i_pipeline.i_pipeline_s3_memory.s3_valid_t0),
.i_pipeline__i_pipeline_s3_memory__dmem_addr_t0(
  i_pipeline.i_pipeline_s3_memory.dmem_addr_t0),
.i_pipeline__i_pipeline_s3_memory__dmem_gnt_t0(
  i_pipeline.i_pipeline_s3_memory.dmem_gnt_t0),
.i_pipeline__i_pipeline_s3_memory__dmem_req_t0(
  i_pipeline.i_pipeline_s3_memory.dmem_req_t0),
.i_pipeline__i_pipeline_s3_memory__dmem_strb_t0(
  i_pipeline.i_pipeline_s3_memory.dmem_strb_t0),
.i_pipeline__i_pipeline_s3_memory__dmem_wdata_t0(
  i_pipeline.i_pipeline_s3_memory.dmem_wdata_t0),
.i_pipeline__i_pipeline_s3_memory__dmem_wen_t0(
  i_pipeline.i_pipeline_s3_memory.dmem_wen_t0),
.i_pipeline__i_pipeline_s3_memory__hold_lsu_req_t0(
  i_pipeline.i_pipeline_s3_memory.hold_lsu_req_t0),
.i_pipeline__i_pipeline_s3_memory__fwd_s3_csr_t0(
  i_pipeline.i_pipeline_s3_memory.fwd_s3_csr_t0),
.i_pipeline__i_pipeline_s3_memory__fwd_s3_load_t0(
  i_pipeline.i_pipeline_s3_memory.fwd_s3_load_t0),
.i_pipeline__i_pipeline_s3_memory__fwd_s3_rd_t0(
  i_pipeline.i_pipeline_s3_memory.fwd_s3_rd_t0),
.i_pipeline__i_pipeline_s3_memory__fwd_s3_wdata_t0(
  i_pipeline.i_pipeline_s3_memory.fwd_s3_wdata_t0),
.i_pipeline__i_pipeline_s3_memory__fwd_s3_wdata_hi_t0(
  i_pipeline.i_pipeline_s3_memory.fwd_s3_wdata_hi_t0),
.i_pipeline__i_pipeline_s3_memory__fwd_s3_wide_t0(
  i_pipeline.i_pipeline_s3_memory.fwd_s3_wide_t0),
.i_pipeline__i_pipeline_s3_memory__leak_fence_unc0_t0(
  i_pipeline.i_pipeline_s3_memory.leak_fence_unc0_t0),
.i_pipeline__i_pipeline_s3_memory__leak_fence_unc1_t0(
  i_pipeline.i_pipeline_s3_memory.leak_fence_unc1_t0),
.i_pipeline__i_pipeline_s3_memory__leak_fence_unc2_t0(
  i_pipeline.i_pipeline_s3_memory.leak_fence_unc2_t0),
.i_pipeline__i_pipeline_s3_memory__s4_busy_t0(
  i_pipeline.i_pipeline_s3_memory.s4_busy_t0),
.i_pipeline__i_pipeline_s3_memory__s4_fu_t0(
  i_pipeline.i_pipeline_s3_memory.s4_fu_t0),
.i_pipeline__i_pipeline_s3_memory__s4_instr_t0(
  i_pipeline.i_pipeline_s3_memory.s4_instr_t0),
.i_pipeline__i_pipeline_s3_memory__s4_opr_a_t0(
  i_pipeline.i_pipeline_s3_memory.s4_opr_a_t0),
.i_pipeline__i_pipeline_s3_memory__s4_opr_b_t0(
  i_pipeline.i_pipeline_s3_memory.s4_opr_b_t0),
.i_pipeline__i_pipeline_s3_memory__s4_rd_t0(
  i_pipeline.i_pipeline_s3_memory.s4_rd_t0),
.i_pipeline__i_pipeline_s3_memory__s4_size_t0(
  i_pipeline.i_pipeline_s3_memory.s4_size_t0),
.i_pipeline__i_pipeline_s3_memory__s4_trap_t0(
  i_pipeline.i_pipeline_s3_memory.s4_trap_t0),
.i_pipeline__i_pipeline_s3_memory__s4_uop_t0(
  i_pipeline.i_pipeline_s3_memory.s4_uop_t0),
.i_pipeline__i_pipeline_s3_memory__s4_valid_t0(
  i_pipeline.i_pipeline_s3_memory.s4_valid_t0),
.i_pipeline__i_pipeline_s3_memory__bitw_gpr_wide(
  i_pipeline.i_pipeline_s3_memory.bitw_gpr_wide),
.i_pipeline__i_pipeline_s3_memory__imul_gpr_wide(
  i_pipeline.i_pipeline_s3_memory.imul_gpr_wide),
.i_pipeline__i_pipeline_s3_memory__leak_fence(
  i_pipeline.i_pipeline_s3_memory.leak_fence),
.i_pipeline__i_pipeline_s3_memory__lsu_a_error(
  i_pipeline.i_pipeline_s3_memory.lsu_a_error),
.i_pipeline__i_pipeline_s3_memory__lsu_a_error_t0(
  i_pipeline.i_pipeline_s3_memory.lsu_a_error_t0),
.i_pipeline__i_pipeline_s3_memory__lsu_byte(
  i_pipeline.i_pipeline_s3_memory.lsu_byte),
.i_pipeline__i_pipeline_s3_memory__lsu_cause(
  i_pipeline.i_pipeline_s3_memory.lsu_cause),
.i_pipeline__i_pipeline_s3_memory__lsu_half(
  i_pipeline.i_pipeline_s3_memory.lsu_half),
.i_pipeline__i_pipeline_s3_memory__lsu_mmio(
  i_pipeline.i_pipeline_s3_memory.lsu_mmio),
.i_pipeline__i_pipeline_s3_memory__lsu_mmio_t0(
  i_pipeline.i_pipeline_s3_memory.lsu_mmio_t0),
.i_pipeline__i_pipeline_s3_memory__lsu_ready(
  i_pipeline.i_pipeline_s3_memory.lsu_ready),
.i_pipeline__i_pipeline_s3_memory__lsu_ready_t0(
  i_pipeline.i_pipeline_s3_memory.lsu_ready_t0),
.i_pipeline__i_pipeline_s3_memory__lsu_word(
  i_pipeline.i_pipeline_s3_memory.lsu_word),
.i_pipeline__i_pipeline_s3_memory__n_s4_opr_a(
  i_pipeline.i_pipeline_s3_memory.n_s4_opr_a),
.i_pipeline__i_pipeline_s3_memory__n_s4_opr_a_t0(
  i_pipeline.i_pipeline_s3_memory.n_s4_opr_a_t0),
.i_pipeline__i_pipeline_s3_memory__n_s4_opr_b(
  i_pipeline.i_pipeline_s3_memory.n_s4_opr_b),
.i_pipeline__i_pipeline_s3_memory__n_s4_opr_b_t0(
  i_pipeline.i_pipeline_s3_memory.n_s4_opr_b_t0),
.i_pipeline__i_pipeline_s3_memory__n_s4_rd(
  i_pipeline.i_pipeline_s3_memory.n_s4_rd),
.i_pipeline__i_pipeline_s3_memory__n_s4_rd_t0(
  i_pipeline.i_pipeline_s3_memory.n_s4_rd_t0),
.i_pipeline__i_pipeline_s3_memory__n_s4_trap(
  i_pipeline.i_pipeline_s3_memory.n_s4_trap),
.i_pipeline__i_pipeline_s3_memory__opra_flush(
  i_pipeline.i_pipeline_s3_memory.opra_flush),
.i_pipeline__i_pipeline_s3_memory__opra_ld_en(
  i_pipeline.i_pipeline_s3_memory.opra_ld_en),
.i_pipeline__i_pipeline_s3_memory__oprb_flush(
  i_pipeline.i_pipeline_s3_memory.oprb_flush),
.i_pipeline__i_pipeline_s3_memory__oprb_ld_en(
  i_pipeline.i_pipeline_s3_memory.oprb_ld_en),
.i_pipeline__i_pipeline_s3_memory__p_busy(
  i_pipeline.i_pipeline_s3_memory.p_busy),
.i_pipeline__i_pipeline_s3_memory__p_busy_t0(
  i_pipeline.i_pipeline_s3_memory.p_busy_t0),
.i_pipeline__i_pipeline_s3_memory__p_valid(
  i_pipeline.i_pipeline_s3_memory.p_valid),
.i_pipeline__i_pipeline_s3_memory__pipe_reg_out(
  i_pipeline.i_pipeline_s3_memory.pipe_reg_out),
.i_pipeline__i_pipeline_s3_memory__pipe_reg_out_t0(
  i_pipeline.i_pipeline_s3_memory.pipe_reg_out_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__g_clk(
  i_pipeline.i_pipeline_s3_memory.i_lsu.g_clk),
.i_pipeline__i_pipeline_s3_memory__i_lsu__g_resetn(
  i_pipeline.i_pipeline_s3_memory.i_lsu.g_resetn),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_valid(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_valid),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_a_error(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_a_error),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_ready(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_ready),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_mmio(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_mmio),
.i_pipeline__i_pipeline_s3_memory__i_lsu__pipe_prog(
  i_pipeline.i_pipeline_s3_memory.i_lsu.pipe_prog),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_addr(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_addr),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_wdata(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_wdata),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_load(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_load),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_store(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_store),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_byte(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_byte),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_half(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_half),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_word(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_word),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_signed(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_signed),
.i_pipeline__i_pipeline_s3_memory__i_lsu__hold_lsu_req(
  i_pipeline.i_pipeline_s3_memory.i_lsu.hold_lsu_req),
.i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_en(
  i_pipeline.i_pipeline_s3_memory.i_lsu.mmio_en),
.i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_wen(
  i_pipeline.i_pipeline_s3_memory.i_lsu.mmio_wen),
.i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_addr(
  i_pipeline.i_pipeline_s3_memory.i_lsu.mmio_addr),
.i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_wdata(
  i_pipeline.i_pipeline_s3_memory.i_lsu.mmio_wdata),
.i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_req(
  i_pipeline.i_pipeline_s3_memory.i_lsu.dmem_req),
.i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_wen(
  i_pipeline.i_pipeline_s3_memory.i_lsu.dmem_wen),
.i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_strb(
  i_pipeline.i_pipeline_s3_memory.i_lsu.dmem_strb),
.i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_wdata(
  i_pipeline.i_pipeline_s3_memory.i_lsu.dmem_wdata),
.i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_addr(
  i_pipeline.i_pipeline_s3_memory.i_lsu.dmem_addr),
.i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_gnt(
  i_pipeline.i_pipeline_s3_memory.i_lsu.dmem_gnt),
.i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_wen_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.mmio_wen_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_wdata_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.mmio_wdata_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_en_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.mmio_en_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_addr_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.mmio_addr_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_load_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_load_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_store_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_store_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_addr_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.dmem_addr_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_gnt_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.dmem_gnt_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_req_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.dmem_req_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_strb_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.dmem_strb_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_wdata_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.dmem_wdata_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_wen_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.dmem_wen_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__hold_lsu_req_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.hold_lsu_req_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_a_error_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_a_error_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_addr_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_addr_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_byte_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_byte_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_half_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_half_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_mmio_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_mmio_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_ready_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_ready_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_signed_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_signed_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_valid_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_valid_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_wdata_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_wdata_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_word_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_word_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__pipe_prog_t0(
  i_pipeline.i_pipeline_s3_memory.i_lsu.pipe_prog_t0),
.i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_txn_done(
  i_pipeline.i_pipeline_s3_memory.i_lsu.dmem_txn_done),
.i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_finished(
  i_pipeline.i_pipeline_s3_memory.i_lsu.lsu_finished),
.i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_done(
  i_pipeline.i_pipeline_s3_memory.i_lsu.mmio_done),
.i_pipeline__i_pipeline_s3_memory__i_lsu__n_lsu_finished(
  i_pipeline.i_pipeline_s3_memory.i_lsu.n_lsu_finished),
.i_pipeline__i_pipeline_s3_memory__i_lsu__n_mmio_done(
  i_pipeline.i_pipeline_s3_memory.i_lsu.n_mmio_done),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__g_clk(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.g_clk),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__g_resetn(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.g_resetn),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_data(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.i_data),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_valid(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.i_valid),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_busy(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.o_busy),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__mr_data(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.mr_data),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__flush(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.flush),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__flush_dat(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.flush_dat),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_data(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.o_data),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_valid(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.o_valid),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_busy(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.i_busy),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__flush_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.flush_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_valid_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.o_valid_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_data_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.o_data_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_busy_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.o_busy_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__mr_data_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.mr_data_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_valid_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.i_valid_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_data_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.i_data_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_busy_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.i_busy_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__flush_dat_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.flush_dat_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__genblk1__progress(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg.\genblk1.progress ),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__g_clk(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.g_clk),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__g_resetn(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.g_resetn),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_data(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.i_data),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_valid(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.i_valid),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_busy(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.o_busy),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__mr_data(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.mr_data),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__flush(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.flush),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__flush_dat(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.flush_dat),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_data(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.o_data),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_valid(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.o_valid),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_busy(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.i_busy),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__flush_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.flush_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_valid_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.o_valid_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_data_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.o_data_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_busy_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.o_busy_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__mr_data_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.mr_data_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_valid_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.i_valid_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_data_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.i_data_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_busy_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.i_busy_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__flush_dat_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.flush_dat_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__genblk1__progress(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_a.\genblk1.progress ),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__g_clk(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.g_clk),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__g_resetn(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.g_resetn),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_data(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.i_data),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_valid(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.i_valid),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_busy(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.o_busy),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__mr_data(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.mr_data),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__flush(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.flush),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__flush_dat(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.flush_dat),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_data(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.o_data),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_valid(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.o_valid),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_busy(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.i_busy),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__flush_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.flush_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_valid_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.o_valid_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_data_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.o_data_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_busy_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.o_busy_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__mr_data_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.mr_data_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_valid_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.i_valid_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_data_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.i_data_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_busy_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.i_busy_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__flush_dat_t0(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.flush_dat_t0),
.i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__genblk1__progress(
  i_pipeline.i_pipeline_s3_memory.i_mem_pipereg_opr_b.\genblk1.progress ),
.i_pipeline__i_pipeline_s4_writeback__g_clk(
  i_pipeline.i_pipeline_s4_writeback.g_clk),
.i_pipeline__i_pipeline_s4_writeback__g_resetn(
  i_pipeline.i_pipeline_s4_writeback.g_resetn),
.i_pipeline__i_pipeline_s4_writeback__s4_rd(
  i_pipeline.i_pipeline_s4_writeback.s4_rd),
.i_pipeline__i_pipeline_s4_writeback__s4_opr_a(
  i_pipeline.i_pipeline_s4_writeback.s4_opr_a),
.i_pipeline__i_pipeline_s4_writeback__s4_opr_b(
  i_pipeline.i_pipeline_s4_writeback.s4_opr_b),
.i_pipeline__i_pipeline_s4_writeback__s4_uop(
  i_pipeline.i_pipeline_s4_writeback.s4_uop),
.i_pipeline__i_pipeline_s4_writeback__s4_fu(
  i_pipeline.i_pipeline_s4_writeback.s4_fu),
.i_pipeline__i_pipeline_s4_writeback__s4_trap(
  i_pipeline.i_pipeline_s4_writeback.s4_trap),
.i_pipeline__i_pipeline_s4_writeback__s4_size(
  i_pipeline.i_pipeline_s4_writeback.s4_size),
.i_pipeline__i_pipeline_s4_writeback__s4_instr(
  i_pipeline.i_pipeline_s4_writeback.s4_instr),
.i_pipeline__i_pipeline_s4_writeback__s4_busy(
  i_pipeline.i_pipeline_s4_writeback.s4_busy),
.i_pipeline__i_pipeline_s4_writeback__s4_valid(
  i_pipeline.i_pipeline_s4_writeback.s4_valid),
.i_pipeline__i_pipeline_s4_writeback__fwd_s4_rd(
  i_pipeline.i_pipeline_s4_writeback.fwd_s4_rd),
.i_pipeline__i_pipeline_s4_writeback__fwd_s4_wdata(
  i_pipeline.i_pipeline_s4_writeback.fwd_s4_wdata),
.i_pipeline__i_pipeline_s4_writeback__fwd_s4_load(
  i_pipeline.i_pipeline_s4_writeback.fwd_s4_load),
.i_pipeline__i_pipeline_s4_writeback__fwd_s4_csr(
  i_pipeline.i_pipeline_s4_writeback.fwd_s4_csr),
.i_pipeline__i_pipeline_s4_writeback__gpr_wen(
  i_pipeline.i_pipeline_s4_writeback.gpr_wen),
.i_pipeline__i_pipeline_s4_writeback__gpr_wide(
  i_pipeline.i_pipeline_s4_writeback.gpr_wide),
.i_pipeline__i_pipeline_s4_writeback__gpr_rd(
  i_pipeline.i_pipeline_s4_writeback.gpr_rd),
.i_pipeline__i_pipeline_s4_writeback__gpr_wdata(
  i_pipeline.i_pipeline_s4_writeback.gpr_wdata),
.i_pipeline__i_pipeline_s4_writeback__gpr_wdata_hi(
  i_pipeline.i_pipeline_s4_writeback.gpr_wdata_hi),
.i_pipeline__i_pipeline_s4_writeback__int_trap_req(
  i_pipeline.i_pipeline_s4_writeback.int_trap_req),
.i_pipeline__i_pipeline_s4_writeback__int_trap_cause(
  i_pipeline.i_pipeline_s4_writeback.int_trap_cause),
.i_pipeline__i_pipeline_s4_writeback__int_trap_ack(
  i_pipeline.i_pipeline_s4_writeback.int_trap_ack),
.i_pipeline__i_pipeline_s4_writeback__trap_cpu(
  i_pipeline.i_pipeline_s4_writeback.trap_cpu),
.i_pipeline__i_pipeline_s4_writeback__trap_int(
  i_pipeline.i_pipeline_s4_writeback.trap_int),
.i_pipeline__i_pipeline_s4_writeback__trap_cause(
  i_pipeline.i_pipeline_s4_writeback.trap_cause),
.i_pipeline__i_pipeline_s4_writeback__trap_mtval(
  i_pipeline.i_pipeline_s4_writeback.trap_mtval),
.i_pipeline__i_pipeline_s4_writeback__trap_pc(
  i_pipeline.i_pipeline_s4_writeback.trap_pc),
.i_pipeline__i_pipeline_s4_writeback__exec_mret(
  i_pipeline.i_pipeline_s4_writeback.exec_mret),
.i_pipeline__i_pipeline_s4_writeback__csr_mepc(
  i_pipeline.i_pipeline_s4_writeback.csr_mepc),
.i_pipeline__i_pipeline_s4_writeback__csr_mtvec(
  i_pipeline.i_pipeline_s4_writeback.csr_mtvec),
.i_pipeline__i_pipeline_s4_writeback__vector_intrs(
  i_pipeline.i_pipeline_s4_writeback.vector_intrs),
.i_pipeline__i_pipeline_s4_writeback__trs_pc(
  i_pipeline.i_pipeline_s4_writeback.trs_pc),
.i_pipeline__i_pipeline_s4_writeback__trs_instr(
  i_pipeline.i_pipeline_s4_writeback.trs_instr),
.i_pipeline__i_pipeline_s4_writeback__trs_valid(
  i_pipeline.i_pipeline_s4_writeback.trs_valid),
.i_pipeline__i_pipeline_s4_writeback__csr_en(
  i_pipeline.i_pipeline_s4_writeback.csr_en),
.i_pipeline__i_pipeline_s4_writeback__csr_wr(
  i_pipeline.i_pipeline_s4_writeback.csr_wr),
.i_pipeline__i_pipeline_s4_writeback__csr_wr_set(
  i_pipeline.i_pipeline_s4_writeback.csr_wr_set),
.i_pipeline__i_pipeline_s4_writeback__csr_wr_clr(
  i_pipeline.i_pipeline_s4_writeback.csr_wr_clr),
.i_pipeline__i_pipeline_s4_writeback__csr_addr(
  i_pipeline.i_pipeline_s4_writeback.csr_addr),
.i_pipeline__i_pipeline_s4_writeback__csr_wdata(
  i_pipeline.i_pipeline_s4_writeback.csr_wdata),
.i_pipeline__i_pipeline_s4_writeback__csr_rdata(
  i_pipeline.i_pipeline_s4_writeback.csr_rdata),
.i_pipeline__i_pipeline_s4_writeback__csr_error(
  i_pipeline.i_pipeline_s4_writeback.csr_error),
.i_pipeline__i_pipeline_s4_writeback__cf_req(
  i_pipeline.i_pipeline_s4_writeback.cf_req),
.i_pipeline__i_pipeline_s4_writeback__cf_target(
  i_pipeline.i_pipeline_s4_writeback.cf_target),
.i_pipeline__i_pipeline_s4_writeback__cf_ack(
  i_pipeline.i_pipeline_s4_writeback.cf_ack),
.i_pipeline__i_pipeline_s4_writeback__hold_lsu_req(
  i_pipeline.i_pipeline_s4_writeback.hold_lsu_req),
.i_pipeline__i_pipeline_s4_writeback__mmio_rdata(
  i_pipeline.i_pipeline_s4_writeback.mmio_rdata),
.i_pipeline__i_pipeline_s4_writeback__mmio_error(
  i_pipeline.i_pipeline_s4_writeback.mmio_error),
.i_pipeline__i_pipeline_s4_writeback__dmem_recv(
  i_pipeline.i_pipeline_s4_writeback.dmem_recv),
.i_pipeline__i_pipeline_s4_writeback__dmem_ack(
  i_pipeline.i_pipeline_s4_writeback.dmem_ack),
.i_pipeline__i_pipeline_s4_writeback__dmem_error(
  i_pipeline.i_pipeline_s4_writeback.dmem_error),
.i_pipeline__i_pipeline_s4_writeback__dmem_rdata(
  i_pipeline.i_pipeline_s4_writeback.dmem_rdata),
.i_pipeline__i_pipeline_s4_writeback__trap_cause_t0(
  i_pipeline.i_pipeline_s4_writeback.trap_cause_t0),
.i_pipeline__i_pipeline_s4_writeback__cf_target_t0(
  i_pipeline.i_pipeline_s4_writeback.cf_target_t0),
.i_pipeline__i_pipeline_s4_writeback__cf_req_t0(
  i_pipeline.i_pipeline_s4_writeback.cf_req_t0),
.i_pipeline__i_pipeline_s4_writeback__cf_ack_t0(
  i_pipeline.i_pipeline_s4_writeback.cf_ack_t0),
.i_pipeline__i_pipeline_s4_writeback__int_trap_req_t0(
  i_pipeline.i_pipeline_s4_writeback.int_trap_req_t0),
.i_pipeline__i_pipeline_s4_writeback__mmio_rdata_t0(
  i_pipeline.i_pipeline_s4_writeback.mmio_rdata_t0),
.i_pipeline__i_pipeline_s4_writeback__mmio_error_t0(
  i_pipeline.i_pipeline_s4_writeback.mmio_error_t0),
.i_pipeline__i_pipeline_s4_writeback__int_trap_cause_t0(
  i_pipeline.i_pipeline_s4_writeback.int_trap_cause_t0),
.i_pipeline__i_pipeline_s4_writeback__int_trap_ack_t0(
  i_pipeline.i_pipeline_s4_writeback.int_trap_ack_t0),
.i_pipeline__i_pipeline_s4_writeback__hold_lsu_req_t0(
  i_pipeline.i_pipeline_s4_writeback.hold_lsu_req_t0),
.i_pipeline__i_pipeline_s4_writeback__s4_busy_t0(
  i_pipeline.i_pipeline_s4_writeback.s4_busy_t0),
.i_pipeline__i_pipeline_s4_writeback__s4_fu_t0(
  i_pipeline.i_pipeline_s4_writeback.s4_fu_t0),
.i_pipeline__i_pipeline_s4_writeback__s4_instr_t0(
  i_pipeline.i_pipeline_s4_writeback.s4_instr_t0),
.i_pipeline__i_pipeline_s4_writeback__s4_opr_a_t0(
  i_pipeline.i_pipeline_s4_writeback.s4_opr_a_t0),
.i_pipeline__i_pipeline_s4_writeback__s4_opr_b_t0(
  i_pipeline.i_pipeline_s4_writeback.s4_opr_b_t0),
.i_pipeline__i_pipeline_s4_writeback__s4_rd_t0(
  i_pipeline.i_pipeline_s4_writeback.s4_rd_t0),
.i_pipeline__i_pipeline_s4_writeback__s4_size_t0(
  i_pipeline.i_pipeline_s4_writeback.s4_size_t0),
.i_pipeline__i_pipeline_s4_writeback__s4_trap_t0(
  i_pipeline.i_pipeline_s4_writeback.s4_trap_t0),
.i_pipeline__i_pipeline_s4_writeback__s4_uop_t0(
  i_pipeline.i_pipeline_s4_writeback.s4_uop_t0),
.i_pipeline__i_pipeline_s4_writeback__s4_valid_t0(
  i_pipeline.i_pipeline_s4_writeback.s4_valid_t0),
.i_pipeline__i_pipeline_s4_writeback__csr_addr_t0(
  i_pipeline.i_pipeline_s4_writeback.csr_addr_t0),
.i_pipeline__i_pipeline_s4_writeback__csr_en_t0(
  i_pipeline.i_pipeline_s4_writeback.csr_en_t0),
.i_pipeline__i_pipeline_s4_writeback__csr_error_t0(
  i_pipeline.i_pipeline_s4_writeback.csr_error_t0),
.i_pipeline__i_pipeline_s4_writeback__csr_mepc_t0(
  i_pipeline.i_pipeline_s4_writeback.csr_mepc_t0),
.i_pipeline__i_pipeline_s4_writeback__csr_mtvec_t0(
  i_pipeline.i_pipeline_s4_writeback.csr_mtvec_t0),
.i_pipeline__i_pipeline_s4_writeback__csr_rdata_t0(
  i_pipeline.i_pipeline_s4_writeback.csr_rdata_t0),
.i_pipeline__i_pipeline_s4_writeback__csr_wdata_t0(
  i_pipeline.i_pipeline_s4_writeback.csr_wdata_t0),
.i_pipeline__i_pipeline_s4_writeback__csr_wr_t0(
  i_pipeline.i_pipeline_s4_writeback.csr_wr_t0),
.i_pipeline__i_pipeline_s4_writeback__csr_wr_clr_t0(
  i_pipeline.i_pipeline_s4_writeback.csr_wr_clr_t0),
.i_pipeline__i_pipeline_s4_writeback__csr_wr_set_t0(
  i_pipeline.i_pipeline_s4_writeback.csr_wr_set_t0),
.i_pipeline__i_pipeline_s4_writeback__dmem_ack_t0(
  i_pipeline.i_pipeline_s4_writeback.dmem_ack_t0),
.i_pipeline__i_pipeline_s4_writeback__dmem_error_t0(
  i_pipeline.i_pipeline_s4_writeback.dmem_error_t0),
.i_pipeline__i_pipeline_s4_writeback__dmem_rdata_t0(
  i_pipeline.i_pipeline_s4_writeback.dmem_rdata_t0),
.i_pipeline__i_pipeline_s4_writeback__dmem_recv_t0(
  i_pipeline.i_pipeline_s4_writeback.dmem_recv_t0),
.i_pipeline__i_pipeline_s4_writeback__exec_mret_t0(
  i_pipeline.i_pipeline_s4_writeback.exec_mret_t0),
.i_pipeline__i_pipeline_s4_writeback__fwd_s4_csr_t0(
  i_pipeline.i_pipeline_s4_writeback.fwd_s4_csr_t0),
.i_pipeline__i_pipeline_s4_writeback__fwd_s4_load_t0(
  i_pipeline.i_pipeline_s4_writeback.fwd_s4_load_t0),
.i_pipeline__i_pipeline_s4_writeback__fwd_s4_rd_t0(
  i_pipeline.i_pipeline_s4_writeback.fwd_s4_rd_t0),
.i_pipeline__i_pipeline_s4_writeback__fwd_s4_wdata_t0(
  i_pipeline.i_pipeline_s4_writeback.fwd_s4_wdata_t0),
.i_pipeline__i_pipeline_s4_writeback__gpr_rd_t0(
  i_pipeline.i_pipeline_s4_writeback.gpr_rd_t0),
.i_pipeline__i_pipeline_s4_writeback__gpr_wdata_t0(
  i_pipeline.i_pipeline_s4_writeback.gpr_wdata_t0),
.i_pipeline__i_pipeline_s4_writeback__gpr_wdata_hi_t0(
  i_pipeline.i_pipeline_s4_writeback.gpr_wdata_hi_t0),
.i_pipeline__i_pipeline_s4_writeback__gpr_wen_t0(
  i_pipeline.i_pipeline_s4_writeback.gpr_wen_t0),
.i_pipeline__i_pipeline_s4_writeback__gpr_wide_t0(
  i_pipeline.i_pipeline_s4_writeback.gpr_wide_t0),
.i_pipeline__i_pipeline_s4_writeback__trap_cpu_t0(
  i_pipeline.i_pipeline_s4_writeback.trap_cpu_t0),
.i_pipeline__i_pipeline_s4_writeback__trap_int_t0(
  i_pipeline.i_pipeline_s4_writeback.trap_int_t0),
.i_pipeline__i_pipeline_s4_writeback__trap_mtval_t0(
  i_pipeline.i_pipeline_s4_writeback.trap_mtval_t0),
.i_pipeline__i_pipeline_s4_writeback__trap_pc_t0(
  i_pipeline.i_pipeline_s4_writeback.trap_pc_t0),
.i_pipeline__i_pipeline_s4_writeback__trs_instr_t0(
  i_pipeline.i_pipeline_s4_writeback.trs_instr_t0),
.i_pipeline__i_pipeline_s4_writeback__trs_pc_t0(
  i_pipeline.i_pipeline_s4_writeback.trs_pc_t0),
.i_pipeline__i_pipeline_s4_writeback__trs_valid_t0(
  i_pipeline.i_pipeline_s4_writeback.trs_valid_t0),
.i_pipeline__i_pipeline_s4_writeback__vector_intrs_t0(
  i_pipeline.i_pipeline_s4_writeback.vector_intrs_t0),
.i_pipeline__i_pipeline_s4_writeback__cf_req_noint(
  i_pipeline.i_pipeline_s4_writeback.cf_req_noint),
.i_pipeline__i_pipeline_s4_writeback__cf_target_noint(
  i_pipeline.i_pipeline_s4_writeback.cf_target_noint),
.i_pipeline__i_pipeline_s4_writeback__cf_target_noint_t0(
  i_pipeline.i_pipeline_s4_writeback.cf_target_noint_t0),
.i_pipeline__i_pipeline_s4_writeback__cfu_busy(
  i_pipeline.i_pipeline_s4_writeback.cfu_busy),
.i_pipeline__i_pipeline_s4_writeback__cfu_cf_taken(
  i_pipeline.i_pipeline_s4_writeback.cfu_cf_taken),
.i_pipeline__i_pipeline_s4_writeback__cfu_done(
  i_pipeline.i_pipeline_s4_writeback.cfu_done),
.i_pipeline__i_pipeline_s4_writeback__cfu_ebreak(
  i_pipeline.i_pipeline_s4_writeback.cfu_ebreak),
.i_pipeline__i_pipeline_s4_writeback__cfu_ecall(
  i_pipeline.i_pipeline_s4_writeback.cfu_ecall),
.i_pipeline__i_pipeline_s4_writeback__cfu_finish_now(
  i_pipeline.i_pipeline_s4_writeback.cfu_finish_now),
.i_pipeline__i_pipeline_s4_writeback__cfu_gpr_wdata(
  i_pipeline.i_pipeline_s4_writeback.cfu_gpr_wdata),
.i_pipeline__i_pipeline_s4_writeback__cfu_gpr_wdata_t0(
  i_pipeline.i_pipeline_s4_writeback.cfu_gpr_wdata_t0),
.i_pipeline__i_pipeline_s4_writeback__cfu_gpr_wen(
  i_pipeline.i_pipeline_s4_writeback.cfu_gpr_wen),
.i_pipeline__i_pipeline_s4_writeback__cfu_mret(
  i_pipeline.i_pipeline_s4_writeback.cfu_mret),
.i_pipeline__i_pipeline_s4_writeback__cfu_tgt_trap(
  i_pipeline.i_pipeline_s4_writeback.cfu_tgt_trap),
.i_pipeline__i_pipeline_s4_writeback__cfu_trap(
  i_pipeline.i_pipeline_s4_writeback.cfu_trap),
.i_pipeline__i_pipeline_s4_writeback__csr_done(
  i_pipeline.i_pipeline_s4_writeback.csr_done),
.i_pipeline__i_pipeline_s4_writeback__csr_gpr_wen(
  i_pipeline.i_pipeline_s4_writeback.csr_gpr_wen),
.i_pipeline__i_pipeline_s4_writeback__csr_read(
  i_pipeline.i_pipeline_s4_writeback.csr_read),
.i_pipeline__i_pipeline_s4_writeback__dmem_error_seen(
  i_pipeline.i_pipeline_s4_writeback.dmem_error_seen),
.i_pipeline__i_pipeline_s4_writeback__lsu_b_error(
  i_pipeline.i_pipeline_s4_writeback.lsu_b_error),
.i_pipeline__i_pipeline_s4_writeback__lsu_busy(
  i_pipeline.i_pipeline_s4_writeback.lsu_busy),
.i_pipeline__i_pipeline_s4_writeback__lsu_byte(
  i_pipeline.i_pipeline_s4_writeback.lsu_byte),
.i_pipeline__i_pipeline_s4_writeback__lsu_gpr_wen(
  i_pipeline.i_pipeline_s4_writeback.lsu_gpr_wen),
.i_pipeline__i_pipeline_s4_writeback__lsu_half(
  i_pipeline.i_pipeline_s4_writeback.lsu_half),
.i_pipeline__i_pipeline_s4_writeback__lsu_load(
  i_pipeline.i_pipeline_s4_writeback.lsu_load),
.i_pipeline__i_pipeline_s4_writeback__lsu_mmio(
  i_pipeline.i_pipeline_s4_writeback.lsu_mmio),
.i_pipeline__i_pipeline_s4_writeback__lsu_rsp_seen(
  i_pipeline.i_pipeline_s4_writeback.lsu_rsp_seen),
.i_pipeline__i_pipeline_s4_writeback__lsu_store(
  i_pipeline.i_pipeline_s4_writeback.lsu_store),
.i_pipeline__i_pipeline_s4_writeback__lsu_txn_recv(
  i_pipeline.i_pipeline_s4_writeback.lsu_txn_recv),
.i_pipeline__i_pipeline_s4_writeback__lsu_word(
  i_pipeline.i_pipeline_s4_writeback.lsu_word),
.i_pipeline__i_pipeline_s4_writeback__mem_rdata(
  i_pipeline.i_pipeline_s4_writeback.mem_rdata),
.i_pipeline__i_pipeline_s4_writeback__mem_rdata_t0(
  i_pipeline.i_pipeline_s4_writeback.mem_rdata_t0),
.i_pipeline__i_pipeline_s4_writeback__n_cfu_done(
  i_pipeline.i_pipeline_s4_writeback.n_cfu_done),
.i_pipeline__i_pipeline_s4_writeback__n_csr_done(
  i_pipeline.i_pipeline_s4_writeback.n_csr_done),
.i_pipeline__i_pipeline_s4_writeback__n_dmem_error_seen(
  i_pipeline.i_pipeline_s4_writeback.n_dmem_error_seen),
.i_pipeline__i_pipeline_s4_writeback__n_lsu_rsp_seen(
  i_pipeline.i_pipeline_s4_writeback.n_lsu_rsp_seen),
.i_pipeline__i_pipeline_s4_writeback__pipe_progress(
  i_pipeline.i_pipeline_s4_writeback.pipe_progress),
.i_pipeline__i_pipeline_s4_writeback__rdata_b0(
  i_pipeline.i_pipeline_s4_writeback.rdata_b0),
.i_pipeline__i_pipeline_s4_writeback__rdata_b0_t0(
  i_pipeline.i_pipeline_s4_writeback.rdata_b0_t0),
.i_pipeline__i_pipeline_s4_writeback__rdata_b1(
  i_pipeline.i_pipeline_s4_writeback.rdata_b1),
.i_pipeline__i_pipeline_s4_writeback__rdata_b1_t0(
  i_pipeline.i_pipeline_s4_writeback.rdata_b1_t0),
.i_pipeline__i_pipeline_s4_writeback__rdata_h1(
  i_pipeline.i_pipeline_s4_writeback.rdata_h1),
.i_pipeline__i_pipeline_s4_writeback__rdata_h1_t0(
  i_pipeline.i_pipeline_s4_writeback.rdata_h1_t0),
.i_pipeline__i_pipeline_s4_writeback__rng_gpr_wen(
  i_pipeline.i_pipeline_s4_writeback.rng_gpr_wen),
.i_pipeline__i_pipeline_s4_writeback__trap_int_pending(
  i_pipeline.i_pipeline_s4_writeback.trap_int_pending),
.i_pipeline__i_pipeline_s4_writeback__trap_target_addr(
  i_pipeline.i_pipeline_s4_writeback.trap_target_addr),
.i_pipeline__i_pipeline_s4_writeback__trap_target_addr_t0(
  i_pipeline.i_pipeline_s4_writeback.trap_target_addr_t0),
.i_pipeline__i_pipeline_s4_writeback__trap_vector_offset(
  i_pipeline.i_pipeline_s4_writeback.trap_vector_offset),
.i_pipeline__i_pipeline_s4_writeback__trap_vector_offset_t0(
  i_pipeline.i_pipeline_s4_writeback.trap_vector_offset_t0)
);
