    asm_no_taint_top_boot_addr_i_t0: assume property(boot_addr_i_t0 == 0);
    asm_no_taint_top_data_err_i_t0: assume property(data_err_i_t0 == 0);
    asm_no_taint_top_data_gnt_i_t0: assume property(data_gnt_i_t0 == 0);
    asm_no_taint_top_data_rdata_i_t0: assume property(data_rdata_i_t0 == 0);
    asm_no_taint_top_data_rdata_intg_i_t0: assume property(data_rdata_intg_i_t0 == 0);
    asm_no_taint_top_data_rvalid_i_t0: assume property(data_rvalid_i_t0 == 0);
    asm_no_taint_top_debug_req_i_t0: assume property(debug_req_i_t0 == 0);
    asm_no_taint_top_fetch_enable_i_t0: assume property(fetch_enable_i_t0 == 0);
    asm_no_taint_top_hart_id_i_t0: assume property(hart_id_i_t0 == 0);
    asm_no_taint_top_instr_err_i_t0: assume property(instr_err_i_t0 == 0);
    asm_no_taint_top_instr_gnt_i_t0: assume property(instr_gnt_i_t0 == 0);
    asm_no_taint_top_instr_rdata_i_t0: assume property(instr_rdata_i_t0 == 0);
    asm_no_taint_top_instr_rdata_intg_i_t0: assume property(instr_rdata_intg_i_t0 == 0);
    asm_no_taint_top_instr_rvalid_i_t0: assume property(instr_rvalid_i_t0 == 0);
    asm_no_taint_top_irq_external_i_t0: assume property(irq_external_i_t0 == 0);
    asm_no_taint_top_irq_fast_i_t0: assume property(irq_fast_i_t0 == 0);
    asm_no_taint_top_irq_nm_i_t0: assume property(irq_nm_i_t0 == 0);
    asm_no_taint_top_irq_software_i_t0: assume property(irq_software_i_t0 == 0);
    asm_no_taint_top_irq_timer_i_t0: assume property(irq_timer_i_t0 == 0);
    asm_no_taint_top_ram_cfg_i_t0: assume property(ram_cfg_i_t0 == 0);
    asm_no_taint_top_scan_rst_ni_t0: assume property(scan_rst_ni_t0 == 0);
    asm_no_taint_top_scramble_key_i_t0: assume property(scramble_key_i_t0 == 0);
    asm_no_taint_top_scramble_key_valid_i_t0: assume property(scramble_key_valid_i_t0 == 0);
    asm_no_taint_top_scramble_nonce_i_t0: assume property(scramble_nonce_i_t0 == 0);
    asm_no_taint_top_test_en_i_t0: assume property(test_en_i_t0 == 0);