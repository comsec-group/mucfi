bit gen_uc_rs2;
assign gen_uc_rs2 =  ((1'h1));
