bit gen_regrd_rs1;
assign gen_regrd_rs1 = 
 (((~ (| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h10), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h11), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h14), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h15), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h18), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h19), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1c), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1d), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h12) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h13)), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h16) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h17)), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1a) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1b)), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1e) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1f)) })) &
((~ (| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h08), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h09), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0c), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0d), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0a) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0b)), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0e) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0f)) })) &
((~ (| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h04), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h05), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h06) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h07)) })) &
((~ ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h02) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h03))) &
(~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h01)))))));
;