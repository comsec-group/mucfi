    asm_no_taint_top_irq_t0: assume property(irq_t0 == 0);
    asm_no_taint_top_mem_rdata_t0: assume property(mem_rdata_t0 == 0);
    asm_no_taint_top_mem_ready_t0: assume property(mem_ready_t0 == 0);
    asm_no_taint_top_pcpi_rd_t0: assume property(pcpi_rd_t0 == 0);
    asm_no_taint_top_pcpi_ready_t0: assume property(pcpi_ready_t0 == 0);
    asm_no_taint_top_pcpi_wait_t0: assume property(pcpi_wait_t0 == 0);
    asm_no_taint_top_pcpi_wr_t0: assume property(pcpi_wr_t0 == 0);