`include "formal/properties/taint_conditions/uc_iw.sv"
`include "formal/properties/taint_conditions/uc_regrd_rs1.sv"
`include "formal/properties/taint_conditions/uc_regrd_rs2.sv"
`include "formal/properties/taint_conditions/uc_rs1.sv"
`include "formal/properties/taint_conditions/uc_rs2.sv"
