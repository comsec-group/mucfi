


bit gen_rs1_uc;

reg [4:0] tmp0046;
always_ff @(posedge clk)
tmp0046 <= ((mem_do_rinst &&  mem_done) ? mem_rdata_latched[19:15] : decoded_rs1);

assign gen_rs1_uc =
$past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'hxx) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'hxx) >> 1) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'hxx) >> 2) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'hxx) >> 3) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'hxx) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1))));


bit gen_rs1_uc_cpuregs_rs1;
assign gen_rs1_uc_cpuregs_rs1 = (((1'h1 | (tmp0046[4] & ((1'h1 | (tmp0046[3] & ((1'h1 | (tmp0046[2] & ((1'h1 | (tmp0046[1] & ((1'h1 | (tmp0046[0] & $past((((((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1 & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1 & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1 & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))) | ((~ tmp0046[0]) & $past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1 & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1 & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))))) | ((~ tmp0046[1]) & ((1'h1 | (tmp0046[0] & $past((((((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1 & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1)) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1 & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1 & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))) | ((~ tmp0046[0]) & $past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1)) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1 & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1 & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))))))) | ((~ tmp0046[2]) & ((1'h1 | (tmp0046[1] & ((1'h1 | (tmp0046[0] & $past((((((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1 & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1 & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))) | ((~ tmp0046[0]) & $past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1 & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))))) | ((~ tmp0046[1]) & ((1'h1 | (tmp0046[0] & $past((((((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1 & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1)) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1 & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))) | ((~ tmp0046[0]) & $past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1)) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1 & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))))))))) | ((~ tmp0046[3]) & ((1'h1 | (tmp0046[2] & ((1'h1 | (tmp0046[1] & ((1'h1 | (tmp0046[0] & $past((((((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1 & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1 & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))) | ((~ tmp0046[0]) & $past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1 & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))))) | ((~ tmp0046[1]) & ((1'h1 | (tmp0046[0] & $past((((((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1 & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1)) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1 & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))) | ((~ tmp0046[0]) & $past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1)) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1 & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))))))) | ((~ tmp0046[2]) & ((1'h1 | (tmp0046[1] & ((1'h1 | (tmp0046[0] & $past((((((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1 & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))) | ((~ tmp0046[0]) & $past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))))) | ((~ tmp0046[1]) & ((1'h1 | (tmp0046[0] & $past((((((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1 & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1)) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))) | ((~ tmp0046[0]) & $past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1)) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))))))))))) | ((~ tmp0046[4]) & ((1'h1 | (tmp0046[3] & ((1'h1 | (tmp0046[2] & ((1'h1 | (tmp0046[1] & ((1'h1 | (tmp0046[0] & $past((((((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1 & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1 & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1 & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))) | ((~ tmp0046[0]) & $past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1 & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1 & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))))) | ((~ tmp0046[1]) & ((1'h1 | (tmp0046[0] & $past((((((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1 & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1)) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1 & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1 & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))) | ((~ tmp0046[0]) & $past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1)) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1 & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1 & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))))))) | ((~ tmp0046[2]) & ((1'h1 | (tmp0046[1] & ((1'h1 | (tmp0046[0] & $past((((((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1 & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1 & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))) | ((~ tmp0046[0]) & $past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1 & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))))) | ((~ tmp0046[1]) & ((1'h1 | (tmp0046[0] & $past((((((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1 & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1)) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1 & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))) | ((~ tmp0046[0]) & $past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1)) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1 & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))))))))) | ((~ tmp0046[3]) & ((1'h1 | (tmp0046[2] & ((1'h1 | (tmp0046[1] & ((1'h1 | (tmp0046[0] & $past((((((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1 & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1 & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))) | ((~ tmp0046[0]) & $past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1 & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))))) | ((~ tmp0046[1]) & ((1'h1 | (tmp0046[0] & $past((((((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1 & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1)) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1 & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))) | ((~ tmp0046[0]) & $past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1)) & (((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1 & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))))))) | ((~ tmp0046[2]) & ((1'h1 | (tmp0046[1] & ((1'h1 | (tmp0046[0] & $past((((((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1 & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))) | ((~ tmp0046[0]) & $past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))))) | ((~ tmp0046[1]) & ((1'h1 | (tmp0046[0] & $past((((((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1 & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1)) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))) | ((~ tmp0046[0]) & $past((((((~ (((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 1) & 1'b1)) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 2) & 1'b1) & ((~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 3) & 1'b1) & (~ ((((resetn &&  cpuregs_write) &&  latched_rd) ?  latched_rd : 5'h0) >> 4) & 1'b1)))) & ((((resetn &&  cpuregs_write) &&  latched_rd) ?  1'h1 : 1'h0) & 1'b1)) == 32'd1)))))))))))));