module alert_handler_reg_top (
	clk_i,
	rst_ni,
	rst_shadowed_ni,
	tl_i,
	tl_o,
	reg2hw,
	hw2reg,
	shadowed_storage_err_o,
	shadowed_update_err_o,
	intg_err_o,
	devmode_i
);
	input clk_i;
	input rst_ni;
	input rst_shadowed_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_i;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	output wire [1161:0] reg2hw;
	input wire [363:0] hw2reg;
	output wire shadowed_storage_err_o;
	output wire shadowed_update_err_o;
	output wire intg_err_o;
	input devmode_i;
	localparam signed [31:0] AW = 11;
	localparam signed [31:0] DW = 32;
	localparam signed [31:0] DBW = 4;
	wire reg_we;
	wire reg_re;
	wire [10:0] reg_addr;
	wire [31:0] reg_wdata;
	wire [3:0] reg_be;
	wire [31:0] reg_rdata;
	wire reg_error;
	wire addrmiss;
	reg wr_err;
	reg [31:0] reg_rdata_next;
	wire reg_busy;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_reg_h2d;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_reg_d2h;
	wire intg_err;
	tlul_cmd_intg_chk u_chk(
		.tl_i(tl_i),
		.err_o(intg_err)
	);
	wire reg_we_err;
	reg [349:0] reg_we_check;
	prim_reg_we_check #(.OneHotWidth(350)) u_prim_reg_we_check(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.oh_i(reg_we_check),
		.en_i(reg_we && !addrmiss),
		.err_o(reg_we_err)
	);
	reg err_q;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			err_q <= 1'sb0;
		else if (intg_err || reg_we_err)
			err_q <= 1'b1;
	assign intg_err_o = (err_q | intg_err) | reg_we_err;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o_pre;
	tlul_rsp_intg_gen #(
		.EnableRspIntgGen(1),
		.EnableDataIntgGen(1)
	) u_rsp_intg_gen(
		.tl_i(tl_o_pre),
		.tl_o(tl_o)
	);
	assign tl_reg_h2d = tl_i;
	assign tl_o_pre = tl_reg_d2h;
	function automatic [3:0] sv2v_cast_E4F5B;
		input reg [3:0] inp;
		sv2v_cast_E4F5B = inp;
	endfunction
	tlul_adapter_reg #(
		.RegAw(AW),
		.RegDw(DW),
		.EnableDataIntgGen(0)
	) u_reg_if(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_reg_h2d),
		.tl_o(tl_reg_d2h),
		.en_ifetch_i(sv2v_cast_E4F5B(4'h9)),
		.we_o(reg_we),
		.re_o(reg_re),
		.addr_o(reg_addr),
		.wdata_o(reg_wdata),
		.be_o(reg_be),
		.busy_i(reg_busy),
		.rdata_i(reg_rdata),
		.error_i(reg_error)
	);
	assign reg_rdata = reg_rdata_next;
	assign reg_error = ((devmode_i & addrmiss) | wr_err) | intg_err;
	wire intr_state_we;
	wire intr_state_classa_qs;
	wire intr_state_classa_wd;
	wire intr_state_classb_qs;
	wire intr_state_classb_wd;
	wire intr_state_classc_qs;
	wire intr_state_classc_wd;
	wire intr_state_classd_qs;
	wire intr_state_classd_wd;
	wire intr_enable_we;
	wire intr_enable_classa_qs;
	wire intr_enable_classa_wd;
	wire intr_enable_classb_qs;
	wire intr_enable_classb_wd;
	wire intr_enable_classc_qs;
	wire intr_enable_classc_wd;
	wire intr_enable_classd_qs;
	wire intr_enable_classd_wd;
	wire intr_test_we;
	wire intr_test_classa_wd;
	wire intr_test_classb_wd;
	wire intr_test_classc_wd;
	wire intr_test_classd_wd;
	wire ping_timer_regwen_we;
	wire ping_timer_regwen_qs;
	wire ping_timer_regwen_wd;
	wire ping_timeout_cyc_shadowed_re;
	wire ping_timeout_cyc_shadowed_we;
	wire [15:0] ping_timeout_cyc_shadowed_qs;
	wire [15:0] ping_timeout_cyc_shadowed_wd;
	wire ping_timeout_cyc_shadowed_storage_err;
	wire ping_timeout_cyc_shadowed_update_err;
	wire ping_timer_en_shadowed_re;
	wire ping_timer_en_shadowed_we;
	wire ping_timer_en_shadowed_qs;
	wire ping_timer_en_shadowed_wd;
	wire ping_timer_en_shadowed_storage_err;
	wire ping_timer_en_shadowed_update_err;
	wire alert_regwen_0_we;
	wire alert_regwen_0_qs;
	wire alert_regwen_0_wd;
	wire alert_regwen_1_we;
	wire alert_regwen_1_qs;
	wire alert_regwen_1_wd;
	wire alert_regwen_2_we;
	wire alert_regwen_2_qs;
	wire alert_regwen_2_wd;
	wire alert_regwen_3_we;
	wire alert_regwen_3_qs;
	wire alert_regwen_3_wd;
	wire alert_regwen_4_we;
	wire alert_regwen_4_qs;
	wire alert_regwen_4_wd;
	wire alert_regwen_5_we;
	wire alert_regwen_5_qs;
	wire alert_regwen_5_wd;
	wire alert_regwen_6_we;
	wire alert_regwen_6_qs;
	wire alert_regwen_6_wd;
	wire alert_regwen_7_we;
	wire alert_regwen_7_qs;
	wire alert_regwen_7_wd;
	wire alert_regwen_8_we;
	wire alert_regwen_8_qs;
	wire alert_regwen_8_wd;
	wire alert_regwen_9_we;
	wire alert_regwen_9_qs;
	wire alert_regwen_9_wd;
	wire alert_regwen_10_we;
	wire alert_regwen_10_qs;
	wire alert_regwen_10_wd;
	wire alert_regwen_11_we;
	wire alert_regwen_11_qs;
	wire alert_regwen_11_wd;
	wire alert_regwen_12_we;
	wire alert_regwen_12_qs;
	wire alert_regwen_12_wd;
	wire alert_regwen_13_we;
	wire alert_regwen_13_qs;
	wire alert_regwen_13_wd;
	wire alert_regwen_14_we;
	wire alert_regwen_14_qs;
	wire alert_regwen_14_wd;
	wire alert_regwen_15_we;
	wire alert_regwen_15_qs;
	wire alert_regwen_15_wd;
	wire alert_regwen_16_we;
	wire alert_regwen_16_qs;
	wire alert_regwen_16_wd;
	wire alert_regwen_17_we;
	wire alert_regwen_17_qs;
	wire alert_regwen_17_wd;
	wire alert_regwen_18_we;
	wire alert_regwen_18_qs;
	wire alert_regwen_18_wd;
	wire alert_regwen_19_we;
	wire alert_regwen_19_qs;
	wire alert_regwen_19_wd;
	wire alert_regwen_20_we;
	wire alert_regwen_20_qs;
	wire alert_regwen_20_wd;
	wire alert_regwen_21_we;
	wire alert_regwen_21_qs;
	wire alert_regwen_21_wd;
	wire alert_regwen_22_we;
	wire alert_regwen_22_qs;
	wire alert_regwen_22_wd;
	wire alert_regwen_23_we;
	wire alert_regwen_23_qs;
	wire alert_regwen_23_wd;
	wire alert_regwen_24_we;
	wire alert_regwen_24_qs;
	wire alert_regwen_24_wd;
	wire alert_regwen_25_we;
	wire alert_regwen_25_qs;
	wire alert_regwen_25_wd;
	wire alert_regwen_26_we;
	wire alert_regwen_26_qs;
	wire alert_regwen_26_wd;
	wire alert_regwen_27_we;
	wire alert_regwen_27_qs;
	wire alert_regwen_27_wd;
	wire alert_regwen_28_we;
	wire alert_regwen_28_qs;
	wire alert_regwen_28_wd;
	wire alert_regwen_29_we;
	wire alert_regwen_29_qs;
	wire alert_regwen_29_wd;
	wire alert_regwen_30_we;
	wire alert_regwen_30_qs;
	wire alert_regwen_30_wd;
	wire alert_regwen_31_we;
	wire alert_regwen_31_qs;
	wire alert_regwen_31_wd;
	wire alert_regwen_32_we;
	wire alert_regwen_32_qs;
	wire alert_regwen_32_wd;
	wire alert_regwen_33_we;
	wire alert_regwen_33_qs;
	wire alert_regwen_33_wd;
	wire alert_regwen_34_we;
	wire alert_regwen_34_qs;
	wire alert_regwen_34_wd;
	wire alert_regwen_35_we;
	wire alert_regwen_35_qs;
	wire alert_regwen_35_wd;
	wire alert_regwen_36_we;
	wire alert_regwen_36_qs;
	wire alert_regwen_36_wd;
	wire alert_regwen_37_we;
	wire alert_regwen_37_qs;
	wire alert_regwen_37_wd;
	wire alert_regwen_38_we;
	wire alert_regwen_38_qs;
	wire alert_regwen_38_wd;
	wire alert_regwen_39_we;
	wire alert_regwen_39_qs;
	wire alert_regwen_39_wd;
	wire alert_regwen_40_we;
	wire alert_regwen_40_qs;
	wire alert_regwen_40_wd;
	wire alert_regwen_41_we;
	wire alert_regwen_41_qs;
	wire alert_regwen_41_wd;
	wire alert_regwen_42_we;
	wire alert_regwen_42_qs;
	wire alert_regwen_42_wd;
	wire alert_regwen_43_we;
	wire alert_regwen_43_qs;
	wire alert_regwen_43_wd;
	wire alert_regwen_44_we;
	wire alert_regwen_44_qs;
	wire alert_regwen_44_wd;
	wire alert_regwen_45_we;
	wire alert_regwen_45_qs;
	wire alert_regwen_45_wd;
	wire alert_regwen_46_we;
	wire alert_regwen_46_qs;
	wire alert_regwen_46_wd;
	wire alert_regwen_47_we;
	wire alert_regwen_47_qs;
	wire alert_regwen_47_wd;
	wire alert_regwen_48_we;
	wire alert_regwen_48_qs;
	wire alert_regwen_48_wd;
	wire alert_regwen_49_we;
	wire alert_regwen_49_qs;
	wire alert_regwen_49_wd;
	wire alert_regwen_50_we;
	wire alert_regwen_50_qs;
	wire alert_regwen_50_wd;
	wire alert_regwen_51_we;
	wire alert_regwen_51_qs;
	wire alert_regwen_51_wd;
	wire alert_regwen_52_we;
	wire alert_regwen_52_qs;
	wire alert_regwen_52_wd;
	wire alert_regwen_53_we;
	wire alert_regwen_53_qs;
	wire alert_regwen_53_wd;
	wire alert_regwen_54_we;
	wire alert_regwen_54_qs;
	wire alert_regwen_54_wd;
	wire alert_regwen_55_we;
	wire alert_regwen_55_qs;
	wire alert_regwen_55_wd;
	wire alert_regwen_56_we;
	wire alert_regwen_56_qs;
	wire alert_regwen_56_wd;
	wire alert_regwen_57_we;
	wire alert_regwen_57_qs;
	wire alert_regwen_57_wd;
	wire alert_regwen_58_we;
	wire alert_regwen_58_qs;
	wire alert_regwen_58_wd;
	wire alert_regwen_59_we;
	wire alert_regwen_59_qs;
	wire alert_regwen_59_wd;
	wire alert_regwen_60_we;
	wire alert_regwen_60_qs;
	wire alert_regwen_60_wd;
	wire alert_regwen_61_we;
	wire alert_regwen_61_qs;
	wire alert_regwen_61_wd;
	wire alert_regwen_62_we;
	wire alert_regwen_62_qs;
	wire alert_regwen_62_wd;
	wire alert_regwen_63_we;
	wire alert_regwen_63_qs;
	wire alert_regwen_63_wd;
	wire alert_regwen_64_we;
	wire alert_regwen_64_qs;
	wire alert_regwen_64_wd;
	wire alert_en_shadowed_0_re;
	wire alert_en_shadowed_0_we;
	wire alert_en_shadowed_0_qs;
	wire alert_en_shadowed_0_wd;
	wire alert_en_shadowed_0_storage_err;
	wire alert_en_shadowed_0_update_err;
	wire alert_en_shadowed_1_re;
	wire alert_en_shadowed_1_we;
	wire alert_en_shadowed_1_qs;
	wire alert_en_shadowed_1_wd;
	wire alert_en_shadowed_1_storage_err;
	wire alert_en_shadowed_1_update_err;
	wire alert_en_shadowed_2_re;
	wire alert_en_shadowed_2_we;
	wire alert_en_shadowed_2_qs;
	wire alert_en_shadowed_2_wd;
	wire alert_en_shadowed_2_storage_err;
	wire alert_en_shadowed_2_update_err;
	wire alert_en_shadowed_3_re;
	wire alert_en_shadowed_3_we;
	wire alert_en_shadowed_3_qs;
	wire alert_en_shadowed_3_wd;
	wire alert_en_shadowed_3_storage_err;
	wire alert_en_shadowed_3_update_err;
	wire alert_en_shadowed_4_re;
	wire alert_en_shadowed_4_we;
	wire alert_en_shadowed_4_qs;
	wire alert_en_shadowed_4_wd;
	wire alert_en_shadowed_4_storage_err;
	wire alert_en_shadowed_4_update_err;
	wire alert_en_shadowed_5_re;
	wire alert_en_shadowed_5_we;
	wire alert_en_shadowed_5_qs;
	wire alert_en_shadowed_5_wd;
	wire alert_en_shadowed_5_storage_err;
	wire alert_en_shadowed_5_update_err;
	wire alert_en_shadowed_6_re;
	wire alert_en_shadowed_6_we;
	wire alert_en_shadowed_6_qs;
	wire alert_en_shadowed_6_wd;
	wire alert_en_shadowed_6_storage_err;
	wire alert_en_shadowed_6_update_err;
	wire alert_en_shadowed_7_re;
	wire alert_en_shadowed_7_we;
	wire alert_en_shadowed_7_qs;
	wire alert_en_shadowed_7_wd;
	wire alert_en_shadowed_7_storage_err;
	wire alert_en_shadowed_7_update_err;
	wire alert_en_shadowed_8_re;
	wire alert_en_shadowed_8_we;
	wire alert_en_shadowed_8_qs;
	wire alert_en_shadowed_8_wd;
	wire alert_en_shadowed_8_storage_err;
	wire alert_en_shadowed_8_update_err;
	wire alert_en_shadowed_9_re;
	wire alert_en_shadowed_9_we;
	wire alert_en_shadowed_9_qs;
	wire alert_en_shadowed_9_wd;
	wire alert_en_shadowed_9_storage_err;
	wire alert_en_shadowed_9_update_err;
	wire alert_en_shadowed_10_re;
	wire alert_en_shadowed_10_we;
	wire alert_en_shadowed_10_qs;
	wire alert_en_shadowed_10_wd;
	wire alert_en_shadowed_10_storage_err;
	wire alert_en_shadowed_10_update_err;
	wire alert_en_shadowed_11_re;
	wire alert_en_shadowed_11_we;
	wire alert_en_shadowed_11_qs;
	wire alert_en_shadowed_11_wd;
	wire alert_en_shadowed_11_storage_err;
	wire alert_en_shadowed_11_update_err;
	wire alert_en_shadowed_12_re;
	wire alert_en_shadowed_12_we;
	wire alert_en_shadowed_12_qs;
	wire alert_en_shadowed_12_wd;
	wire alert_en_shadowed_12_storage_err;
	wire alert_en_shadowed_12_update_err;
	wire alert_en_shadowed_13_re;
	wire alert_en_shadowed_13_we;
	wire alert_en_shadowed_13_qs;
	wire alert_en_shadowed_13_wd;
	wire alert_en_shadowed_13_storage_err;
	wire alert_en_shadowed_13_update_err;
	wire alert_en_shadowed_14_re;
	wire alert_en_shadowed_14_we;
	wire alert_en_shadowed_14_qs;
	wire alert_en_shadowed_14_wd;
	wire alert_en_shadowed_14_storage_err;
	wire alert_en_shadowed_14_update_err;
	wire alert_en_shadowed_15_re;
	wire alert_en_shadowed_15_we;
	wire alert_en_shadowed_15_qs;
	wire alert_en_shadowed_15_wd;
	wire alert_en_shadowed_15_storage_err;
	wire alert_en_shadowed_15_update_err;
	wire alert_en_shadowed_16_re;
	wire alert_en_shadowed_16_we;
	wire alert_en_shadowed_16_qs;
	wire alert_en_shadowed_16_wd;
	wire alert_en_shadowed_16_storage_err;
	wire alert_en_shadowed_16_update_err;
	wire alert_en_shadowed_17_re;
	wire alert_en_shadowed_17_we;
	wire alert_en_shadowed_17_qs;
	wire alert_en_shadowed_17_wd;
	wire alert_en_shadowed_17_storage_err;
	wire alert_en_shadowed_17_update_err;
	wire alert_en_shadowed_18_re;
	wire alert_en_shadowed_18_we;
	wire alert_en_shadowed_18_qs;
	wire alert_en_shadowed_18_wd;
	wire alert_en_shadowed_18_storage_err;
	wire alert_en_shadowed_18_update_err;
	wire alert_en_shadowed_19_re;
	wire alert_en_shadowed_19_we;
	wire alert_en_shadowed_19_qs;
	wire alert_en_shadowed_19_wd;
	wire alert_en_shadowed_19_storage_err;
	wire alert_en_shadowed_19_update_err;
	wire alert_en_shadowed_20_re;
	wire alert_en_shadowed_20_we;
	wire alert_en_shadowed_20_qs;
	wire alert_en_shadowed_20_wd;
	wire alert_en_shadowed_20_storage_err;
	wire alert_en_shadowed_20_update_err;
	wire alert_en_shadowed_21_re;
	wire alert_en_shadowed_21_we;
	wire alert_en_shadowed_21_qs;
	wire alert_en_shadowed_21_wd;
	wire alert_en_shadowed_21_storage_err;
	wire alert_en_shadowed_21_update_err;
	wire alert_en_shadowed_22_re;
	wire alert_en_shadowed_22_we;
	wire alert_en_shadowed_22_qs;
	wire alert_en_shadowed_22_wd;
	wire alert_en_shadowed_22_storage_err;
	wire alert_en_shadowed_22_update_err;
	wire alert_en_shadowed_23_re;
	wire alert_en_shadowed_23_we;
	wire alert_en_shadowed_23_qs;
	wire alert_en_shadowed_23_wd;
	wire alert_en_shadowed_23_storage_err;
	wire alert_en_shadowed_23_update_err;
	wire alert_en_shadowed_24_re;
	wire alert_en_shadowed_24_we;
	wire alert_en_shadowed_24_qs;
	wire alert_en_shadowed_24_wd;
	wire alert_en_shadowed_24_storage_err;
	wire alert_en_shadowed_24_update_err;
	wire alert_en_shadowed_25_re;
	wire alert_en_shadowed_25_we;
	wire alert_en_shadowed_25_qs;
	wire alert_en_shadowed_25_wd;
	wire alert_en_shadowed_25_storage_err;
	wire alert_en_shadowed_25_update_err;
	wire alert_en_shadowed_26_re;
	wire alert_en_shadowed_26_we;
	wire alert_en_shadowed_26_qs;
	wire alert_en_shadowed_26_wd;
	wire alert_en_shadowed_26_storage_err;
	wire alert_en_shadowed_26_update_err;
	wire alert_en_shadowed_27_re;
	wire alert_en_shadowed_27_we;
	wire alert_en_shadowed_27_qs;
	wire alert_en_shadowed_27_wd;
	wire alert_en_shadowed_27_storage_err;
	wire alert_en_shadowed_27_update_err;
	wire alert_en_shadowed_28_re;
	wire alert_en_shadowed_28_we;
	wire alert_en_shadowed_28_qs;
	wire alert_en_shadowed_28_wd;
	wire alert_en_shadowed_28_storage_err;
	wire alert_en_shadowed_28_update_err;
	wire alert_en_shadowed_29_re;
	wire alert_en_shadowed_29_we;
	wire alert_en_shadowed_29_qs;
	wire alert_en_shadowed_29_wd;
	wire alert_en_shadowed_29_storage_err;
	wire alert_en_shadowed_29_update_err;
	wire alert_en_shadowed_30_re;
	wire alert_en_shadowed_30_we;
	wire alert_en_shadowed_30_qs;
	wire alert_en_shadowed_30_wd;
	wire alert_en_shadowed_30_storage_err;
	wire alert_en_shadowed_30_update_err;
	wire alert_en_shadowed_31_re;
	wire alert_en_shadowed_31_we;
	wire alert_en_shadowed_31_qs;
	wire alert_en_shadowed_31_wd;
	wire alert_en_shadowed_31_storage_err;
	wire alert_en_shadowed_31_update_err;
	wire alert_en_shadowed_32_re;
	wire alert_en_shadowed_32_we;
	wire alert_en_shadowed_32_qs;
	wire alert_en_shadowed_32_wd;
	wire alert_en_shadowed_32_storage_err;
	wire alert_en_shadowed_32_update_err;
	wire alert_en_shadowed_33_re;
	wire alert_en_shadowed_33_we;
	wire alert_en_shadowed_33_qs;
	wire alert_en_shadowed_33_wd;
	wire alert_en_shadowed_33_storage_err;
	wire alert_en_shadowed_33_update_err;
	wire alert_en_shadowed_34_re;
	wire alert_en_shadowed_34_we;
	wire alert_en_shadowed_34_qs;
	wire alert_en_shadowed_34_wd;
	wire alert_en_shadowed_34_storage_err;
	wire alert_en_shadowed_34_update_err;
	wire alert_en_shadowed_35_re;
	wire alert_en_shadowed_35_we;
	wire alert_en_shadowed_35_qs;
	wire alert_en_shadowed_35_wd;
	wire alert_en_shadowed_35_storage_err;
	wire alert_en_shadowed_35_update_err;
	wire alert_en_shadowed_36_re;
	wire alert_en_shadowed_36_we;
	wire alert_en_shadowed_36_qs;
	wire alert_en_shadowed_36_wd;
	wire alert_en_shadowed_36_storage_err;
	wire alert_en_shadowed_36_update_err;
	wire alert_en_shadowed_37_re;
	wire alert_en_shadowed_37_we;
	wire alert_en_shadowed_37_qs;
	wire alert_en_shadowed_37_wd;
	wire alert_en_shadowed_37_storage_err;
	wire alert_en_shadowed_37_update_err;
	wire alert_en_shadowed_38_re;
	wire alert_en_shadowed_38_we;
	wire alert_en_shadowed_38_qs;
	wire alert_en_shadowed_38_wd;
	wire alert_en_shadowed_38_storage_err;
	wire alert_en_shadowed_38_update_err;
	wire alert_en_shadowed_39_re;
	wire alert_en_shadowed_39_we;
	wire alert_en_shadowed_39_qs;
	wire alert_en_shadowed_39_wd;
	wire alert_en_shadowed_39_storage_err;
	wire alert_en_shadowed_39_update_err;
	wire alert_en_shadowed_40_re;
	wire alert_en_shadowed_40_we;
	wire alert_en_shadowed_40_qs;
	wire alert_en_shadowed_40_wd;
	wire alert_en_shadowed_40_storage_err;
	wire alert_en_shadowed_40_update_err;
	wire alert_en_shadowed_41_re;
	wire alert_en_shadowed_41_we;
	wire alert_en_shadowed_41_qs;
	wire alert_en_shadowed_41_wd;
	wire alert_en_shadowed_41_storage_err;
	wire alert_en_shadowed_41_update_err;
	wire alert_en_shadowed_42_re;
	wire alert_en_shadowed_42_we;
	wire alert_en_shadowed_42_qs;
	wire alert_en_shadowed_42_wd;
	wire alert_en_shadowed_42_storage_err;
	wire alert_en_shadowed_42_update_err;
	wire alert_en_shadowed_43_re;
	wire alert_en_shadowed_43_we;
	wire alert_en_shadowed_43_qs;
	wire alert_en_shadowed_43_wd;
	wire alert_en_shadowed_43_storage_err;
	wire alert_en_shadowed_43_update_err;
	wire alert_en_shadowed_44_re;
	wire alert_en_shadowed_44_we;
	wire alert_en_shadowed_44_qs;
	wire alert_en_shadowed_44_wd;
	wire alert_en_shadowed_44_storage_err;
	wire alert_en_shadowed_44_update_err;
	wire alert_en_shadowed_45_re;
	wire alert_en_shadowed_45_we;
	wire alert_en_shadowed_45_qs;
	wire alert_en_shadowed_45_wd;
	wire alert_en_shadowed_45_storage_err;
	wire alert_en_shadowed_45_update_err;
	wire alert_en_shadowed_46_re;
	wire alert_en_shadowed_46_we;
	wire alert_en_shadowed_46_qs;
	wire alert_en_shadowed_46_wd;
	wire alert_en_shadowed_46_storage_err;
	wire alert_en_shadowed_46_update_err;
	wire alert_en_shadowed_47_re;
	wire alert_en_shadowed_47_we;
	wire alert_en_shadowed_47_qs;
	wire alert_en_shadowed_47_wd;
	wire alert_en_shadowed_47_storage_err;
	wire alert_en_shadowed_47_update_err;
	wire alert_en_shadowed_48_re;
	wire alert_en_shadowed_48_we;
	wire alert_en_shadowed_48_qs;
	wire alert_en_shadowed_48_wd;
	wire alert_en_shadowed_48_storage_err;
	wire alert_en_shadowed_48_update_err;
	wire alert_en_shadowed_49_re;
	wire alert_en_shadowed_49_we;
	wire alert_en_shadowed_49_qs;
	wire alert_en_shadowed_49_wd;
	wire alert_en_shadowed_49_storage_err;
	wire alert_en_shadowed_49_update_err;
	wire alert_en_shadowed_50_re;
	wire alert_en_shadowed_50_we;
	wire alert_en_shadowed_50_qs;
	wire alert_en_shadowed_50_wd;
	wire alert_en_shadowed_50_storage_err;
	wire alert_en_shadowed_50_update_err;
	wire alert_en_shadowed_51_re;
	wire alert_en_shadowed_51_we;
	wire alert_en_shadowed_51_qs;
	wire alert_en_shadowed_51_wd;
	wire alert_en_shadowed_51_storage_err;
	wire alert_en_shadowed_51_update_err;
	wire alert_en_shadowed_52_re;
	wire alert_en_shadowed_52_we;
	wire alert_en_shadowed_52_qs;
	wire alert_en_shadowed_52_wd;
	wire alert_en_shadowed_52_storage_err;
	wire alert_en_shadowed_52_update_err;
	wire alert_en_shadowed_53_re;
	wire alert_en_shadowed_53_we;
	wire alert_en_shadowed_53_qs;
	wire alert_en_shadowed_53_wd;
	wire alert_en_shadowed_53_storage_err;
	wire alert_en_shadowed_53_update_err;
	wire alert_en_shadowed_54_re;
	wire alert_en_shadowed_54_we;
	wire alert_en_shadowed_54_qs;
	wire alert_en_shadowed_54_wd;
	wire alert_en_shadowed_54_storage_err;
	wire alert_en_shadowed_54_update_err;
	wire alert_en_shadowed_55_re;
	wire alert_en_shadowed_55_we;
	wire alert_en_shadowed_55_qs;
	wire alert_en_shadowed_55_wd;
	wire alert_en_shadowed_55_storage_err;
	wire alert_en_shadowed_55_update_err;
	wire alert_en_shadowed_56_re;
	wire alert_en_shadowed_56_we;
	wire alert_en_shadowed_56_qs;
	wire alert_en_shadowed_56_wd;
	wire alert_en_shadowed_56_storage_err;
	wire alert_en_shadowed_56_update_err;
	wire alert_en_shadowed_57_re;
	wire alert_en_shadowed_57_we;
	wire alert_en_shadowed_57_qs;
	wire alert_en_shadowed_57_wd;
	wire alert_en_shadowed_57_storage_err;
	wire alert_en_shadowed_57_update_err;
	wire alert_en_shadowed_58_re;
	wire alert_en_shadowed_58_we;
	wire alert_en_shadowed_58_qs;
	wire alert_en_shadowed_58_wd;
	wire alert_en_shadowed_58_storage_err;
	wire alert_en_shadowed_58_update_err;
	wire alert_en_shadowed_59_re;
	wire alert_en_shadowed_59_we;
	wire alert_en_shadowed_59_qs;
	wire alert_en_shadowed_59_wd;
	wire alert_en_shadowed_59_storage_err;
	wire alert_en_shadowed_59_update_err;
	wire alert_en_shadowed_60_re;
	wire alert_en_shadowed_60_we;
	wire alert_en_shadowed_60_qs;
	wire alert_en_shadowed_60_wd;
	wire alert_en_shadowed_60_storage_err;
	wire alert_en_shadowed_60_update_err;
	wire alert_en_shadowed_61_re;
	wire alert_en_shadowed_61_we;
	wire alert_en_shadowed_61_qs;
	wire alert_en_shadowed_61_wd;
	wire alert_en_shadowed_61_storage_err;
	wire alert_en_shadowed_61_update_err;
	wire alert_en_shadowed_62_re;
	wire alert_en_shadowed_62_we;
	wire alert_en_shadowed_62_qs;
	wire alert_en_shadowed_62_wd;
	wire alert_en_shadowed_62_storage_err;
	wire alert_en_shadowed_62_update_err;
	wire alert_en_shadowed_63_re;
	wire alert_en_shadowed_63_we;
	wire alert_en_shadowed_63_qs;
	wire alert_en_shadowed_63_wd;
	wire alert_en_shadowed_63_storage_err;
	wire alert_en_shadowed_63_update_err;
	wire alert_en_shadowed_64_re;
	wire alert_en_shadowed_64_we;
	wire alert_en_shadowed_64_qs;
	wire alert_en_shadowed_64_wd;
	wire alert_en_shadowed_64_storage_err;
	wire alert_en_shadowed_64_update_err;
	wire alert_class_shadowed_0_re;
	wire alert_class_shadowed_0_we;
	wire [1:0] alert_class_shadowed_0_qs;
	wire [1:0] alert_class_shadowed_0_wd;
	wire alert_class_shadowed_0_storage_err;
	wire alert_class_shadowed_0_update_err;
	wire alert_class_shadowed_1_re;
	wire alert_class_shadowed_1_we;
	wire [1:0] alert_class_shadowed_1_qs;
	wire [1:0] alert_class_shadowed_1_wd;
	wire alert_class_shadowed_1_storage_err;
	wire alert_class_shadowed_1_update_err;
	wire alert_class_shadowed_2_re;
	wire alert_class_shadowed_2_we;
	wire [1:0] alert_class_shadowed_2_qs;
	wire [1:0] alert_class_shadowed_2_wd;
	wire alert_class_shadowed_2_storage_err;
	wire alert_class_shadowed_2_update_err;
	wire alert_class_shadowed_3_re;
	wire alert_class_shadowed_3_we;
	wire [1:0] alert_class_shadowed_3_qs;
	wire [1:0] alert_class_shadowed_3_wd;
	wire alert_class_shadowed_3_storage_err;
	wire alert_class_shadowed_3_update_err;
	wire alert_class_shadowed_4_re;
	wire alert_class_shadowed_4_we;
	wire [1:0] alert_class_shadowed_4_qs;
	wire [1:0] alert_class_shadowed_4_wd;
	wire alert_class_shadowed_4_storage_err;
	wire alert_class_shadowed_4_update_err;
	wire alert_class_shadowed_5_re;
	wire alert_class_shadowed_5_we;
	wire [1:0] alert_class_shadowed_5_qs;
	wire [1:0] alert_class_shadowed_5_wd;
	wire alert_class_shadowed_5_storage_err;
	wire alert_class_shadowed_5_update_err;
	wire alert_class_shadowed_6_re;
	wire alert_class_shadowed_6_we;
	wire [1:0] alert_class_shadowed_6_qs;
	wire [1:0] alert_class_shadowed_6_wd;
	wire alert_class_shadowed_6_storage_err;
	wire alert_class_shadowed_6_update_err;
	wire alert_class_shadowed_7_re;
	wire alert_class_shadowed_7_we;
	wire [1:0] alert_class_shadowed_7_qs;
	wire [1:0] alert_class_shadowed_7_wd;
	wire alert_class_shadowed_7_storage_err;
	wire alert_class_shadowed_7_update_err;
	wire alert_class_shadowed_8_re;
	wire alert_class_shadowed_8_we;
	wire [1:0] alert_class_shadowed_8_qs;
	wire [1:0] alert_class_shadowed_8_wd;
	wire alert_class_shadowed_8_storage_err;
	wire alert_class_shadowed_8_update_err;
	wire alert_class_shadowed_9_re;
	wire alert_class_shadowed_9_we;
	wire [1:0] alert_class_shadowed_9_qs;
	wire [1:0] alert_class_shadowed_9_wd;
	wire alert_class_shadowed_9_storage_err;
	wire alert_class_shadowed_9_update_err;
	wire alert_class_shadowed_10_re;
	wire alert_class_shadowed_10_we;
	wire [1:0] alert_class_shadowed_10_qs;
	wire [1:0] alert_class_shadowed_10_wd;
	wire alert_class_shadowed_10_storage_err;
	wire alert_class_shadowed_10_update_err;
	wire alert_class_shadowed_11_re;
	wire alert_class_shadowed_11_we;
	wire [1:0] alert_class_shadowed_11_qs;
	wire [1:0] alert_class_shadowed_11_wd;
	wire alert_class_shadowed_11_storage_err;
	wire alert_class_shadowed_11_update_err;
	wire alert_class_shadowed_12_re;
	wire alert_class_shadowed_12_we;
	wire [1:0] alert_class_shadowed_12_qs;
	wire [1:0] alert_class_shadowed_12_wd;
	wire alert_class_shadowed_12_storage_err;
	wire alert_class_shadowed_12_update_err;
	wire alert_class_shadowed_13_re;
	wire alert_class_shadowed_13_we;
	wire [1:0] alert_class_shadowed_13_qs;
	wire [1:0] alert_class_shadowed_13_wd;
	wire alert_class_shadowed_13_storage_err;
	wire alert_class_shadowed_13_update_err;
	wire alert_class_shadowed_14_re;
	wire alert_class_shadowed_14_we;
	wire [1:0] alert_class_shadowed_14_qs;
	wire [1:0] alert_class_shadowed_14_wd;
	wire alert_class_shadowed_14_storage_err;
	wire alert_class_shadowed_14_update_err;
	wire alert_class_shadowed_15_re;
	wire alert_class_shadowed_15_we;
	wire [1:0] alert_class_shadowed_15_qs;
	wire [1:0] alert_class_shadowed_15_wd;
	wire alert_class_shadowed_15_storage_err;
	wire alert_class_shadowed_15_update_err;
	wire alert_class_shadowed_16_re;
	wire alert_class_shadowed_16_we;
	wire [1:0] alert_class_shadowed_16_qs;
	wire [1:0] alert_class_shadowed_16_wd;
	wire alert_class_shadowed_16_storage_err;
	wire alert_class_shadowed_16_update_err;
	wire alert_class_shadowed_17_re;
	wire alert_class_shadowed_17_we;
	wire [1:0] alert_class_shadowed_17_qs;
	wire [1:0] alert_class_shadowed_17_wd;
	wire alert_class_shadowed_17_storage_err;
	wire alert_class_shadowed_17_update_err;
	wire alert_class_shadowed_18_re;
	wire alert_class_shadowed_18_we;
	wire [1:0] alert_class_shadowed_18_qs;
	wire [1:0] alert_class_shadowed_18_wd;
	wire alert_class_shadowed_18_storage_err;
	wire alert_class_shadowed_18_update_err;
	wire alert_class_shadowed_19_re;
	wire alert_class_shadowed_19_we;
	wire [1:0] alert_class_shadowed_19_qs;
	wire [1:0] alert_class_shadowed_19_wd;
	wire alert_class_shadowed_19_storage_err;
	wire alert_class_shadowed_19_update_err;
	wire alert_class_shadowed_20_re;
	wire alert_class_shadowed_20_we;
	wire [1:0] alert_class_shadowed_20_qs;
	wire [1:0] alert_class_shadowed_20_wd;
	wire alert_class_shadowed_20_storage_err;
	wire alert_class_shadowed_20_update_err;
	wire alert_class_shadowed_21_re;
	wire alert_class_shadowed_21_we;
	wire [1:0] alert_class_shadowed_21_qs;
	wire [1:0] alert_class_shadowed_21_wd;
	wire alert_class_shadowed_21_storage_err;
	wire alert_class_shadowed_21_update_err;
	wire alert_class_shadowed_22_re;
	wire alert_class_shadowed_22_we;
	wire [1:0] alert_class_shadowed_22_qs;
	wire [1:0] alert_class_shadowed_22_wd;
	wire alert_class_shadowed_22_storage_err;
	wire alert_class_shadowed_22_update_err;
	wire alert_class_shadowed_23_re;
	wire alert_class_shadowed_23_we;
	wire [1:0] alert_class_shadowed_23_qs;
	wire [1:0] alert_class_shadowed_23_wd;
	wire alert_class_shadowed_23_storage_err;
	wire alert_class_shadowed_23_update_err;
	wire alert_class_shadowed_24_re;
	wire alert_class_shadowed_24_we;
	wire [1:0] alert_class_shadowed_24_qs;
	wire [1:0] alert_class_shadowed_24_wd;
	wire alert_class_shadowed_24_storage_err;
	wire alert_class_shadowed_24_update_err;
	wire alert_class_shadowed_25_re;
	wire alert_class_shadowed_25_we;
	wire [1:0] alert_class_shadowed_25_qs;
	wire [1:0] alert_class_shadowed_25_wd;
	wire alert_class_shadowed_25_storage_err;
	wire alert_class_shadowed_25_update_err;
	wire alert_class_shadowed_26_re;
	wire alert_class_shadowed_26_we;
	wire [1:0] alert_class_shadowed_26_qs;
	wire [1:0] alert_class_shadowed_26_wd;
	wire alert_class_shadowed_26_storage_err;
	wire alert_class_shadowed_26_update_err;
	wire alert_class_shadowed_27_re;
	wire alert_class_shadowed_27_we;
	wire [1:0] alert_class_shadowed_27_qs;
	wire [1:0] alert_class_shadowed_27_wd;
	wire alert_class_shadowed_27_storage_err;
	wire alert_class_shadowed_27_update_err;
	wire alert_class_shadowed_28_re;
	wire alert_class_shadowed_28_we;
	wire [1:0] alert_class_shadowed_28_qs;
	wire [1:0] alert_class_shadowed_28_wd;
	wire alert_class_shadowed_28_storage_err;
	wire alert_class_shadowed_28_update_err;
	wire alert_class_shadowed_29_re;
	wire alert_class_shadowed_29_we;
	wire [1:0] alert_class_shadowed_29_qs;
	wire [1:0] alert_class_shadowed_29_wd;
	wire alert_class_shadowed_29_storage_err;
	wire alert_class_shadowed_29_update_err;
	wire alert_class_shadowed_30_re;
	wire alert_class_shadowed_30_we;
	wire [1:0] alert_class_shadowed_30_qs;
	wire [1:0] alert_class_shadowed_30_wd;
	wire alert_class_shadowed_30_storage_err;
	wire alert_class_shadowed_30_update_err;
	wire alert_class_shadowed_31_re;
	wire alert_class_shadowed_31_we;
	wire [1:0] alert_class_shadowed_31_qs;
	wire [1:0] alert_class_shadowed_31_wd;
	wire alert_class_shadowed_31_storage_err;
	wire alert_class_shadowed_31_update_err;
	wire alert_class_shadowed_32_re;
	wire alert_class_shadowed_32_we;
	wire [1:0] alert_class_shadowed_32_qs;
	wire [1:0] alert_class_shadowed_32_wd;
	wire alert_class_shadowed_32_storage_err;
	wire alert_class_shadowed_32_update_err;
	wire alert_class_shadowed_33_re;
	wire alert_class_shadowed_33_we;
	wire [1:0] alert_class_shadowed_33_qs;
	wire [1:0] alert_class_shadowed_33_wd;
	wire alert_class_shadowed_33_storage_err;
	wire alert_class_shadowed_33_update_err;
	wire alert_class_shadowed_34_re;
	wire alert_class_shadowed_34_we;
	wire [1:0] alert_class_shadowed_34_qs;
	wire [1:0] alert_class_shadowed_34_wd;
	wire alert_class_shadowed_34_storage_err;
	wire alert_class_shadowed_34_update_err;
	wire alert_class_shadowed_35_re;
	wire alert_class_shadowed_35_we;
	wire [1:0] alert_class_shadowed_35_qs;
	wire [1:0] alert_class_shadowed_35_wd;
	wire alert_class_shadowed_35_storage_err;
	wire alert_class_shadowed_35_update_err;
	wire alert_class_shadowed_36_re;
	wire alert_class_shadowed_36_we;
	wire [1:0] alert_class_shadowed_36_qs;
	wire [1:0] alert_class_shadowed_36_wd;
	wire alert_class_shadowed_36_storage_err;
	wire alert_class_shadowed_36_update_err;
	wire alert_class_shadowed_37_re;
	wire alert_class_shadowed_37_we;
	wire [1:0] alert_class_shadowed_37_qs;
	wire [1:0] alert_class_shadowed_37_wd;
	wire alert_class_shadowed_37_storage_err;
	wire alert_class_shadowed_37_update_err;
	wire alert_class_shadowed_38_re;
	wire alert_class_shadowed_38_we;
	wire [1:0] alert_class_shadowed_38_qs;
	wire [1:0] alert_class_shadowed_38_wd;
	wire alert_class_shadowed_38_storage_err;
	wire alert_class_shadowed_38_update_err;
	wire alert_class_shadowed_39_re;
	wire alert_class_shadowed_39_we;
	wire [1:0] alert_class_shadowed_39_qs;
	wire [1:0] alert_class_shadowed_39_wd;
	wire alert_class_shadowed_39_storage_err;
	wire alert_class_shadowed_39_update_err;
	wire alert_class_shadowed_40_re;
	wire alert_class_shadowed_40_we;
	wire [1:0] alert_class_shadowed_40_qs;
	wire [1:0] alert_class_shadowed_40_wd;
	wire alert_class_shadowed_40_storage_err;
	wire alert_class_shadowed_40_update_err;
	wire alert_class_shadowed_41_re;
	wire alert_class_shadowed_41_we;
	wire [1:0] alert_class_shadowed_41_qs;
	wire [1:0] alert_class_shadowed_41_wd;
	wire alert_class_shadowed_41_storage_err;
	wire alert_class_shadowed_41_update_err;
	wire alert_class_shadowed_42_re;
	wire alert_class_shadowed_42_we;
	wire [1:0] alert_class_shadowed_42_qs;
	wire [1:0] alert_class_shadowed_42_wd;
	wire alert_class_shadowed_42_storage_err;
	wire alert_class_shadowed_42_update_err;
	wire alert_class_shadowed_43_re;
	wire alert_class_shadowed_43_we;
	wire [1:0] alert_class_shadowed_43_qs;
	wire [1:0] alert_class_shadowed_43_wd;
	wire alert_class_shadowed_43_storage_err;
	wire alert_class_shadowed_43_update_err;
	wire alert_class_shadowed_44_re;
	wire alert_class_shadowed_44_we;
	wire [1:0] alert_class_shadowed_44_qs;
	wire [1:0] alert_class_shadowed_44_wd;
	wire alert_class_shadowed_44_storage_err;
	wire alert_class_shadowed_44_update_err;
	wire alert_class_shadowed_45_re;
	wire alert_class_shadowed_45_we;
	wire [1:0] alert_class_shadowed_45_qs;
	wire [1:0] alert_class_shadowed_45_wd;
	wire alert_class_shadowed_45_storage_err;
	wire alert_class_shadowed_45_update_err;
	wire alert_class_shadowed_46_re;
	wire alert_class_shadowed_46_we;
	wire [1:0] alert_class_shadowed_46_qs;
	wire [1:0] alert_class_shadowed_46_wd;
	wire alert_class_shadowed_46_storage_err;
	wire alert_class_shadowed_46_update_err;
	wire alert_class_shadowed_47_re;
	wire alert_class_shadowed_47_we;
	wire [1:0] alert_class_shadowed_47_qs;
	wire [1:0] alert_class_shadowed_47_wd;
	wire alert_class_shadowed_47_storage_err;
	wire alert_class_shadowed_47_update_err;
	wire alert_class_shadowed_48_re;
	wire alert_class_shadowed_48_we;
	wire [1:0] alert_class_shadowed_48_qs;
	wire [1:0] alert_class_shadowed_48_wd;
	wire alert_class_shadowed_48_storage_err;
	wire alert_class_shadowed_48_update_err;
	wire alert_class_shadowed_49_re;
	wire alert_class_shadowed_49_we;
	wire [1:0] alert_class_shadowed_49_qs;
	wire [1:0] alert_class_shadowed_49_wd;
	wire alert_class_shadowed_49_storage_err;
	wire alert_class_shadowed_49_update_err;
	wire alert_class_shadowed_50_re;
	wire alert_class_shadowed_50_we;
	wire [1:0] alert_class_shadowed_50_qs;
	wire [1:0] alert_class_shadowed_50_wd;
	wire alert_class_shadowed_50_storage_err;
	wire alert_class_shadowed_50_update_err;
	wire alert_class_shadowed_51_re;
	wire alert_class_shadowed_51_we;
	wire [1:0] alert_class_shadowed_51_qs;
	wire [1:0] alert_class_shadowed_51_wd;
	wire alert_class_shadowed_51_storage_err;
	wire alert_class_shadowed_51_update_err;
	wire alert_class_shadowed_52_re;
	wire alert_class_shadowed_52_we;
	wire [1:0] alert_class_shadowed_52_qs;
	wire [1:0] alert_class_shadowed_52_wd;
	wire alert_class_shadowed_52_storage_err;
	wire alert_class_shadowed_52_update_err;
	wire alert_class_shadowed_53_re;
	wire alert_class_shadowed_53_we;
	wire [1:0] alert_class_shadowed_53_qs;
	wire [1:0] alert_class_shadowed_53_wd;
	wire alert_class_shadowed_53_storage_err;
	wire alert_class_shadowed_53_update_err;
	wire alert_class_shadowed_54_re;
	wire alert_class_shadowed_54_we;
	wire [1:0] alert_class_shadowed_54_qs;
	wire [1:0] alert_class_shadowed_54_wd;
	wire alert_class_shadowed_54_storage_err;
	wire alert_class_shadowed_54_update_err;
	wire alert_class_shadowed_55_re;
	wire alert_class_shadowed_55_we;
	wire [1:0] alert_class_shadowed_55_qs;
	wire [1:0] alert_class_shadowed_55_wd;
	wire alert_class_shadowed_55_storage_err;
	wire alert_class_shadowed_55_update_err;
	wire alert_class_shadowed_56_re;
	wire alert_class_shadowed_56_we;
	wire [1:0] alert_class_shadowed_56_qs;
	wire [1:0] alert_class_shadowed_56_wd;
	wire alert_class_shadowed_56_storage_err;
	wire alert_class_shadowed_56_update_err;
	wire alert_class_shadowed_57_re;
	wire alert_class_shadowed_57_we;
	wire [1:0] alert_class_shadowed_57_qs;
	wire [1:0] alert_class_shadowed_57_wd;
	wire alert_class_shadowed_57_storage_err;
	wire alert_class_shadowed_57_update_err;
	wire alert_class_shadowed_58_re;
	wire alert_class_shadowed_58_we;
	wire [1:0] alert_class_shadowed_58_qs;
	wire [1:0] alert_class_shadowed_58_wd;
	wire alert_class_shadowed_58_storage_err;
	wire alert_class_shadowed_58_update_err;
	wire alert_class_shadowed_59_re;
	wire alert_class_shadowed_59_we;
	wire [1:0] alert_class_shadowed_59_qs;
	wire [1:0] alert_class_shadowed_59_wd;
	wire alert_class_shadowed_59_storage_err;
	wire alert_class_shadowed_59_update_err;
	wire alert_class_shadowed_60_re;
	wire alert_class_shadowed_60_we;
	wire [1:0] alert_class_shadowed_60_qs;
	wire [1:0] alert_class_shadowed_60_wd;
	wire alert_class_shadowed_60_storage_err;
	wire alert_class_shadowed_60_update_err;
	wire alert_class_shadowed_61_re;
	wire alert_class_shadowed_61_we;
	wire [1:0] alert_class_shadowed_61_qs;
	wire [1:0] alert_class_shadowed_61_wd;
	wire alert_class_shadowed_61_storage_err;
	wire alert_class_shadowed_61_update_err;
	wire alert_class_shadowed_62_re;
	wire alert_class_shadowed_62_we;
	wire [1:0] alert_class_shadowed_62_qs;
	wire [1:0] alert_class_shadowed_62_wd;
	wire alert_class_shadowed_62_storage_err;
	wire alert_class_shadowed_62_update_err;
	wire alert_class_shadowed_63_re;
	wire alert_class_shadowed_63_we;
	wire [1:0] alert_class_shadowed_63_qs;
	wire [1:0] alert_class_shadowed_63_wd;
	wire alert_class_shadowed_63_storage_err;
	wire alert_class_shadowed_63_update_err;
	wire alert_class_shadowed_64_re;
	wire alert_class_shadowed_64_we;
	wire [1:0] alert_class_shadowed_64_qs;
	wire [1:0] alert_class_shadowed_64_wd;
	wire alert_class_shadowed_64_storage_err;
	wire alert_class_shadowed_64_update_err;
	wire alert_cause_0_we;
	wire alert_cause_0_qs;
	wire alert_cause_0_wd;
	wire alert_cause_1_we;
	wire alert_cause_1_qs;
	wire alert_cause_1_wd;
	wire alert_cause_2_we;
	wire alert_cause_2_qs;
	wire alert_cause_2_wd;
	wire alert_cause_3_we;
	wire alert_cause_3_qs;
	wire alert_cause_3_wd;
	wire alert_cause_4_we;
	wire alert_cause_4_qs;
	wire alert_cause_4_wd;
	wire alert_cause_5_we;
	wire alert_cause_5_qs;
	wire alert_cause_5_wd;
	wire alert_cause_6_we;
	wire alert_cause_6_qs;
	wire alert_cause_6_wd;
	wire alert_cause_7_we;
	wire alert_cause_7_qs;
	wire alert_cause_7_wd;
	wire alert_cause_8_we;
	wire alert_cause_8_qs;
	wire alert_cause_8_wd;
	wire alert_cause_9_we;
	wire alert_cause_9_qs;
	wire alert_cause_9_wd;
	wire alert_cause_10_we;
	wire alert_cause_10_qs;
	wire alert_cause_10_wd;
	wire alert_cause_11_we;
	wire alert_cause_11_qs;
	wire alert_cause_11_wd;
	wire alert_cause_12_we;
	wire alert_cause_12_qs;
	wire alert_cause_12_wd;
	wire alert_cause_13_we;
	wire alert_cause_13_qs;
	wire alert_cause_13_wd;
	wire alert_cause_14_we;
	wire alert_cause_14_qs;
	wire alert_cause_14_wd;
	wire alert_cause_15_we;
	wire alert_cause_15_qs;
	wire alert_cause_15_wd;
	wire alert_cause_16_we;
	wire alert_cause_16_qs;
	wire alert_cause_16_wd;
	wire alert_cause_17_we;
	wire alert_cause_17_qs;
	wire alert_cause_17_wd;
	wire alert_cause_18_we;
	wire alert_cause_18_qs;
	wire alert_cause_18_wd;
	wire alert_cause_19_we;
	wire alert_cause_19_qs;
	wire alert_cause_19_wd;
	wire alert_cause_20_we;
	wire alert_cause_20_qs;
	wire alert_cause_20_wd;
	wire alert_cause_21_we;
	wire alert_cause_21_qs;
	wire alert_cause_21_wd;
	wire alert_cause_22_we;
	wire alert_cause_22_qs;
	wire alert_cause_22_wd;
	wire alert_cause_23_we;
	wire alert_cause_23_qs;
	wire alert_cause_23_wd;
	wire alert_cause_24_we;
	wire alert_cause_24_qs;
	wire alert_cause_24_wd;
	wire alert_cause_25_we;
	wire alert_cause_25_qs;
	wire alert_cause_25_wd;
	wire alert_cause_26_we;
	wire alert_cause_26_qs;
	wire alert_cause_26_wd;
	wire alert_cause_27_we;
	wire alert_cause_27_qs;
	wire alert_cause_27_wd;
	wire alert_cause_28_we;
	wire alert_cause_28_qs;
	wire alert_cause_28_wd;
	wire alert_cause_29_we;
	wire alert_cause_29_qs;
	wire alert_cause_29_wd;
	wire alert_cause_30_we;
	wire alert_cause_30_qs;
	wire alert_cause_30_wd;
	wire alert_cause_31_we;
	wire alert_cause_31_qs;
	wire alert_cause_31_wd;
	wire alert_cause_32_we;
	wire alert_cause_32_qs;
	wire alert_cause_32_wd;
	wire alert_cause_33_we;
	wire alert_cause_33_qs;
	wire alert_cause_33_wd;
	wire alert_cause_34_we;
	wire alert_cause_34_qs;
	wire alert_cause_34_wd;
	wire alert_cause_35_we;
	wire alert_cause_35_qs;
	wire alert_cause_35_wd;
	wire alert_cause_36_we;
	wire alert_cause_36_qs;
	wire alert_cause_36_wd;
	wire alert_cause_37_we;
	wire alert_cause_37_qs;
	wire alert_cause_37_wd;
	wire alert_cause_38_we;
	wire alert_cause_38_qs;
	wire alert_cause_38_wd;
	wire alert_cause_39_we;
	wire alert_cause_39_qs;
	wire alert_cause_39_wd;
	wire alert_cause_40_we;
	wire alert_cause_40_qs;
	wire alert_cause_40_wd;
	wire alert_cause_41_we;
	wire alert_cause_41_qs;
	wire alert_cause_41_wd;
	wire alert_cause_42_we;
	wire alert_cause_42_qs;
	wire alert_cause_42_wd;
	wire alert_cause_43_we;
	wire alert_cause_43_qs;
	wire alert_cause_43_wd;
	wire alert_cause_44_we;
	wire alert_cause_44_qs;
	wire alert_cause_44_wd;
	wire alert_cause_45_we;
	wire alert_cause_45_qs;
	wire alert_cause_45_wd;
	wire alert_cause_46_we;
	wire alert_cause_46_qs;
	wire alert_cause_46_wd;
	wire alert_cause_47_we;
	wire alert_cause_47_qs;
	wire alert_cause_47_wd;
	wire alert_cause_48_we;
	wire alert_cause_48_qs;
	wire alert_cause_48_wd;
	wire alert_cause_49_we;
	wire alert_cause_49_qs;
	wire alert_cause_49_wd;
	wire alert_cause_50_we;
	wire alert_cause_50_qs;
	wire alert_cause_50_wd;
	wire alert_cause_51_we;
	wire alert_cause_51_qs;
	wire alert_cause_51_wd;
	wire alert_cause_52_we;
	wire alert_cause_52_qs;
	wire alert_cause_52_wd;
	wire alert_cause_53_we;
	wire alert_cause_53_qs;
	wire alert_cause_53_wd;
	wire alert_cause_54_we;
	wire alert_cause_54_qs;
	wire alert_cause_54_wd;
	wire alert_cause_55_we;
	wire alert_cause_55_qs;
	wire alert_cause_55_wd;
	wire alert_cause_56_we;
	wire alert_cause_56_qs;
	wire alert_cause_56_wd;
	wire alert_cause_57_we;
	wire alert_cause_57_qs;
	wire alert_cause_57_wd;
	wire alert_cause_58_we;
	wire alert_cause_58_qs;
	wire alert_cause_58_wd;
	wire alert_cause_59_we;
	wire alert_cause_59_qs;
	wire alert_cause_59_wd;
	wire alert_cause_60_we;
	wire alert_cause_60_qs;
	wire alert_cause_60_wd;
	wire alert_cause_61_we;
	wire alert_cause_61_qs;
	wire alert_cause_61_wd;
	wire alert_cause_62_we;
	wire alert_cause_62_qs;
	wire alert_cause_62_wd;
	wire alert_cause_63_we;
	wire alert_cause_63_qs;
	wire alert_cause_63_wd;
	wire alert_cause_64_we;
	wire alert_cause_64_qs;
	wire alert_cause_64_wd;
	wire loc_alert_regwen_0_we;
	wire loc_alert_regwen_0_qs;
	wire loc_alert_regwen_0_wd;
	wire loc_alert_regwen_1_we;
	wire loc_alert_regwen_1_qs;
	wire loc_alert_regwen_1_wd;
	wire loc_alert_regwen_2_we;
	wire loc_alert_regwen_2_qs;
	wire loc_alert_regwen_2_wd;
	wire loc_alert_regwen_3_we;
	wire loc_alert_regwen_3_qs;
	wire loc_alert_regwen_3_wd;
	wire loc_alert_regwen_4_we;
	wire loc_alert_regwen_4_qs;
	wire loc_alert_regwen_4_wd;
	wire loc_alert_regwen_5_we;
	wire loc_alert_regwen_5_qs;
	wire loc_alert_regwen_5_wd;
	wire loc_alert_regwen_6_we;
	wire loc_alert_regwen_6_qs;
	wire loc_alert_regwen_6_wd;
	wire loc_alert_en_shadowed_0_re;
	wire loc_alert_en_shadowed_0_we;
	wire loc_alert_en_shadowed_0_qs;
	wire loc_alert_en_shadowed_0_wd;
	wire loc_alert_en_shadowed_0_storage_err;
	wire loc_alert_en_shadowed_0_update_err;
	wire loc_alert_en_shadowed_1_re;
	wire loc_alert_en_shadowed_1_we;
	wire loc_alert_en_shadowed_1_qs;
	wire loc_alert_en_shadowed_1_wd;
	wire loc_alert_en_shadowed_1_storage_err;
	wire loc_alert_en_shadowed_1_update_err;
	wire loc_alert_en_shadowed_2_re;
	wire loc_alert_en_shadowed_2_we;
	wire loc_alert_en_shadowed_2_qs;
	wire loc_alert_en_shadowed_2_wd;
	wire loc_alert_en_shadowed_2_storage_err;
	wire loc_alert_en_shadowed_2_update_err;
	wire loc_alert_en_shadowed_3_re;
	wire loc_alert_en_shadowed_3_we;
	wire loc_alert_en_shadowed_3_qs;
	wire loc_alert_en_shadowed_3_wd;
	wire loc_alert_en_shadowed_3_storage_err;
	wire loc_alert_en_shadowed_3_update_err;
	wire loc_alert_en_shadowed_4_re;
	wire loc_alert_en_shadowed_4_we;
	wire loc_alert_en_shadowed_4_qs;
	wire loc_alert_en_shadowed_4_wd;
	wire loc_alert_en_shadowed_4_storage_err;
	wire loc_alert_en_shadowed_4_update_err;
	wire loc_alert_en_shadowed_5_re;
	wire loc_alert_en_shadowed_5_we;
	wire loc_alert_en_shadowed_5_qs;
	wire loc_alert_en_shadowed_5_wd;
	wire loc_alert_en_shadowed_5_storage_err;
	wire loc_alert_en_shadowed_5_update_err;
	wire loc_alert_en_shadowed_6_re;
	wire loc_alert_en_shadowed_6_we;
	wire loc_alert_en_shadowed_6_qs;
	wire loc_alert_en_shadowed_6_wd;
	wire loc_alert_en_shadowed_6_storage_err;
	wire loc_alert_en_shadowed_6_update_err;
	wire loc_alert_class_shadowed_0_re;
	wire loc_alert_class_shadowed_0_we;
	wire [1:0] loc_alert_class_shadowed_0_qs;
	wire [1:0] loc_alert_class_shadowed_0_wd;
	wire loc_alert_class_shadowed_0_storage_err;
	wire loc_alert_class_shadowed_0_update_err;
	wire loc_alert_class_shadowed_1_re;
	wire loc_alert_class_shadowed_1_we;
	wire [1:0] loc_alert_class_shadowed_1_qs;
	wire [1:0] loc_alert_class_shadowed_1_wd;
	wire loc_alert_class_shadowed_1_storage_err;
	wire loc_alert_class_shadowed_1_update_err;
	wire loc_alert_class_shadowed_2_re;
	wire loc_alert_class_shadowed_2_we;
	wire [1:0] loc_alert_class_shadowed_2_qs;
	wire [1:0] loc_alert_class_shadowed_2_wd;
	wire loc_alert_class_shadowed_2_storage_err;
	wire loc_alert_class_shadowed_2_update_err;
	wire loc_alert_class_shadowed_3_re;
	wire loc_alert_class_shadowed_3_we;
	wire [1:0] loc_alert_class_shadowed_3_qs;
	wire [1:0] loc_alert_class_shadowed_3_wd;
	wire loc_alert_class_shadowed_3_storage_err;
	wire loc_alert_class_shadowed_3_update_err;
	wire loc_alert_class_shadowed_4_re;
	wire loc_alert_class_shadowed_4_we;
	wire [1:0] loc_alert_class_shadowed_4_qs;
	wire [1:0] loc_alert_class_shadowed_4_wd;
	wire loc_alert_class_shadowed_4_storage_err;
	wire loc_alert_class_shadowed_4_update_err;
	wire loc_alert_class_shadowed_5_re;
	wire loc_alert_class_shadowed_5_we;
	wire [1:0] loc_alert_class_shadowed_5_qs;
	wire [1:0] loc_alert_class_shadowed_5_wd;
	wire loc_alert_class_shadowed_5_storage_err;
	wire loc_alert_class_shadowed_5_update_err;
	wire loc_alert_class_shadowed_6_re;
	wire loc_alert_class_shadowed_6_we;
	wire [1:0] loc_alert_class_shadowed_6_qs;
	wire [1:0] loc_alert_class_shadowed_6_wd;
	wire loc_alert_class_shadowed_6_storage_err;
	wire loc_alert_class_shadowed_6_update_err;
	wire loc_alert_cause_0_we;
	wire loc_alert_cause_0_qs;
	wire loc_alert_cause_0_wd;
	wire loc_alert_cause_1_we;
	wire loc_alert_cause_1_qs;
	wire loc_alert_cause_1_wd;
	wire loc_alert_cause_2_we;
	wire loc_alert_cause_2_qs;
	wire loc_alert_cause_2_wd;
	wire loc_alert_cause_3_we;
	wire loc_alert_cause_3_qs;
	wire loc_alert_cause_3_wd;
	wire loc_alert_cause_4_we;
	wire loc_alert_cause_4_qs;
	wire loc_alert_cause_4_wd;
	wire loc_alert_cause_5_we;
	wire loc_alert_cause_5_qs;
	wire loc_alert_cause_5_wd;
	wire loc_alert_cause_6_we;
	wire loc_alert_cause_6_qs;
	wire loc_alert_cause_6_wd;
	wire classa_regwen_we;
	wire classa_regwen_qs;
	wire classa_regwen_wd;
	wire classa_ctrl_shadowed_re;
	wire classa_ctrl_shadowed_we;
	wire classa_ctrl_shadowed_en_qs;
	wire classa_ctrl_shadowed_en_wd;
	wire classa_ctrl_shadowed_en_storage_err;
	wire classa_ctrl_shadowed_en_update_err;
	wire classa_ctrl_shadowed_lock_qs;
	wire classa_ctrl_shadowed_lock_wd;
	wire classa_ctrl_shadowed_lock_storage_err;
	wire classa_ctrl_shadowed_lock_update_err;
	wire classa_ctrl_shadowed_en_e0_qs;
	wire classa_ctrl_shadowed_en_e0_wd;
	wire classa_ctrl_shadowed_en_e0_storage_err;
	wire classa_ctrl_shadowed_en_e0_update_err;
	wire classa_ctrl_shadowed_en_e1_qs;
	wire classa_ctrl_shadowed_en_e1_wd;
	wire classa_ctrl_shadowed_en_e1_storage_err;
	wire classa_ctrl_shadowed_en_e1_update_err;
	wire classa_ctrl_shadowed_en_e2_qs;
	wire classa_ctrl_shadowed_en_e2_wd;
	wire classa_ctrl_shadowed_en_e2_storage_err;
	wire classa_ctrl_shadowed_en_e2_update_err;
	wire classa_ctrl_shadowed_en_e3_qs;
	wire classa_ctrl_shadowed_en_e3_wd;
	wire classa_ctrl_shadowed_en_e3_storage_err;
	wire classa_ctrl_shadowed_en_e3_update_err;
	wire [1:0] classa_ctrl_shadowed_map_e0_qs;
	wire [1:0] classa_ctrl_shadowed_map_e0_wd;
	wire classa_ctrl_shadowed_map_e0_storage_err;
	wire classa_ctrl_shadowed_map_e0_update_err;
	wire [1:0] classa_ctrl_shadowed_map_e1_qs;
	wire [1:0] classa_ctrl_shadowed_map_e1_wd;
	wire classa_ctrl_shadowed_map_e1_storage_err;
	wire classa_ctrl_shadowed_map_e1_update_err;
	wire [1:0] classa_ctrl_shadowed_map_e2_qs;
	wire [1:0] classa_ctrl_shadowed_map_e2_wd;
	wire classa_ctrl_shadowed_map_e2_storage_err;
	wire classa_ctrl_shadowed_map_e2_update_err;
	wire [1:0] classa_ctrl_shadowed_map_e3_qs;
	wire [1:0] classa_ctrl_shadowed_map_e3_wd;
	wire classa_ctrl_shadowed_map_e3_storage_err;
	wire classa_ctrl_shadowed_map_e3_update_err;
	wire classa_clr_regwen_we;
	wire classa_clr_regwen_qs;
	wire classa_clr_regwen_wd;
	wire classa_clr_shadowed_re;
	wire classa_clr_shadowed_we;
	wire classa_clr_shadowed_qs;
	wire classa_clr_shadowed_wd;
	wire classa_clr_shadowed_storage_err;
	wire classa_clr_shadowed_update_err;
	wire classa_accum_cnt_re;
	wire [15:0] classa_accum_cnt_qs;
	wire classa_accum_thresh_shadowed_re;
	wire classa_accum_thresh_shadowed_we;
	wire [15:0] classa_accum_thresh_shadowed_qs;
	wire [15:0] classa_accum_thresh_shadowed_wd;
	wire classa_accum_thresh_shadowed_storage_err;
	wire classa_accum_thresh_shadowed_update_err;
	wire classa_timeout_cyc_shadowed_re;
	wire classa_timeout_cyc_shadowed_we;
	wire [31:0] classa_timeout_cyc_shadowed_qs;
	wire [31:0] classa_timeout_cyc_shadowed_wd;
	wire classa_timeout_cyc_shadowed_storage_err;
	wire classa_timeout_cyc_shadowed_update_err;
	wire classa_crashdump_trigger_shadowed_re;
	wire classa_crashdump_trigger_shadowed_we;
	wire [1:0] classa_crashdump_trigger_shadowed_qs;
	wire [1:0] classa_crashdump_trigger_shadowed_wd;
	wire classa_crashdump_trigger_shadowed_storage_err;
	wire classa_crashdump_trigger_shadowed_update_err;
	wire classa_phase0_cyc_shadowed_re;
	wire classa_phase0_cyc_shadowed_we;
	wire [31:0] classa_phase0_cyc_shadowed_qs;
	wire [31:0] classa_phase0_cyc_shadowed_wd;
	wire classa_phase0_cyc_shadowed_storage_err;
	wire classa_phase0_cyc_shadowed_update_err;
	wire classa_phase1_cyc_shadowed_re;
	wire classa_phase1_cyc_shadowed_we;
	wire [31:0] classa_phase1_cyc_shadowed_qs;
	wire [31:0] classa_phase1_cyc_shadowed_wd;
	wire classa_phase1_cyc_shadowed_storage_err;
	wire classa_phase1_cyc_shadowed_update_err;
	wire classa_phase2_cyc_shadowed_re;
	wire classa_phase2_cyc_shadowed_we;
	wire [31:0] classa_phase2_cyc_shadowed_qs;
	wire [31:0] classa_phase2_cyc_shadowed_wd;
	wire classa_phase2_cyc_shadowed_storage_err;
	wire classa_phase2_cyc_shadowed_update_err;
	wire classa_phase3_cyc_shadowed_re;
	wire classa_phase3_cyc_shadowed_we;
	wire [31:0] classa_phase3_cyc_shadowed_qs;
	wire [31:0] classa_phase3_cyc_shadowed_wd;
	wire classa_phase3_cyc_shadowed_storage_err;
	wire classa_phase3_cyc_shadowed_update_err;
	wire classa_esc_cnt_re;
	wire [31:0] classa_esc_cnt_qs;
	wire classa_state_re;
	wire [2:0] classa_state_qs;
	wire classb_regwen_we;
	wire classb_regwen_qs;
	wire classb_regwen_wd;
	wire classb_ctrl_shadowed_re;
	wire classb_ctrl_shadowed_we;
	wire classb_ctrl_shadowed_en_qs;
	wire classb_ctrl_shadowed_en_wd;
	wire classb_ctrl_shadowed_en_storage_err;
	wire classb_ctrl_shadowed_en_update_err;
	wire classb_ctrl_shadowed_lock_qs;
	wire classb_ctrl_shadowed_lock_wd;
	wire classb_ctrl_shadowed_lock_storage_err;
	wire classb_ctrl_shadowed_lock_update_err;
	wire classb_ctrl_shadowed_en_e0_qs;
	wire classb_ctrl_shadowed_en_e0_wd;
	wire classb_ctrl_shadowed_en_e0_storage_err;
	wire classb_ctrl_shadowed_en_e0_update_err;
	wire classb_ctrl_shadowed_en_e1_qs;
	wire classb_ctrl_shadowed_en_e1_wd;
	wire classb_ctrl_shadowed_en_e1_storage_err;
	wire classb_ctrl_shadowed_en_e1_update_err;
	wire classb_ctrl_shadowed_en_e2_qs;
	wire classb_ctrl_shadowed_en_e2_wd;
	wire classb_ctrl_shadowed_en_e2_storage_err;
	wire classb_ctrl_shadowed_en_e2_update_err;
	wire classb_ctrl_shadowed_en_e3_qs;
	wire classb_ctrl_shadowed_en_e3_wd;
	wire classb_ctrl_shadowed_en_e3_storage_err;
	wire classb_ctrl_shadowed_en_e3_update_err;
	wire [1:0] classb_ctrl_shadowed_map_e0_qs;
	wire [1:0] classb_ctrl_shadowed_map_e0_wd;
	wire classb_ctrl_shadowed_map_e0_storage_err;
	wire classb_ctrl_shadowed_map_e0_update_err;
	wire [1:0] classb_ctrl_shadowed_map_e1_qs;
	wire [1:0] classb_ctrl_shadowed_map_e1_wd;
	wire classb_ctrl_shadowed_map_e1_storage_err;
	wire classb_ctrl_shadowed_map_e1_update_err;
	wire [1:0] classb_ctrl_shadowed_map_e2_qs;
	wire [1:0] classb_ctrl_shadowed_map_e2_wd;
	wire classb_ctrl_shadowed_map_e2_storage_err;
	wire classb_ctrl_shadowed_map_e2_update_err;
	wire [1:0] classb_ctrl_shadowed_map_e3_qs;
	wire [1:0] classb_ctrl_shadowed_map_e3_wd;
	wire classb_ctrl_shadowed_map_e3_storage_err;
	wire classb_ctrl_shadowed_map_e3_update_err;
	wire classb_clr_regwen_we;
	wire classb_clr_regwen_qs;
	wire classb_clr_regwen_wd;
	wire classb_clr_shadowed_re;
	wire classb_clr_shadowed_we;
	wire classb_clr_shadowed_qs;
	wire classb_clr_shadowed_wd;
	wire classb_clr_shadowed_storage_err;
	wire classb_clr_shadowed_update_err;
	wire classb_accum_cnt_re;
	wire [15:0] classb_accum_cnt_qs;
	wire classb_accum_thresh_shadowed_re;
	wire classb_accum_thresh_shadowed_we;
	wire [15:0] classb_accum_thresh_shadowed_qs;
	wire [15:0] classb_accum_thresh_shadowed_wd;
	wire classb_accum_thresh_shadowed_storage_err;
	wire classb_accum_thresh_shadowed_update_err;
	wire classb_timeout_cyc_shadowed_re;
	wire classb_timeout_cyc_shadowed_we;
	wire [31:0] classb_timeout_cyc_shadowed_qs;
	wire [31:0] classb_timeout_cyc_shadowed_wd;
	wire classb_timeout_cyc_shadowed_storage_err;
	wire classb_timeout_cyc_shadowed_update_err;
	wire classb_crashdump_trigger_shadowed_re;
	wire classb_crashdump_trigger_shadowed_we;
	wire [1:0] classb_crashdump_trigger_shadowed_qs;
	wire [1:0] classb_crashdump_trigger_shadowed_wd;
	wire classb_crashdump_trigger_shadowed_storage_err;
	wire classb_crashdump_trigger_shadowed_update_err;
	wire classb_phase0_cyc_shadowed_re;
	wire classb_phase0_cyc_shadowed_we;
	wire [31:0] classb_phase0_cyc_shadowed_qs;
	wire [31:0] classb_phase0_cyc_shadowed_wd;
	wire classb_phase0_cyc_shadowed_storage_err;
	wire classb_phase0_cyc_shadowed_update_err;
	wire classb_phase1_cyc_shadowed_re;
	wire classb_phase1_cyc_shadowed_we;
	wire [31:0] classb_phase1_cyc_shadowed_qs;
	wire [31:0] classb_phase1_cyc_shadowed_wd;
	wire classb_phase1_cyc_shadowed_storage_err;
	wire classb_phase1_cyc_shadowed_update_err;
	wire classb_phase2_cyc_shadowed_re;
	wire classb_phase2_cyc_shadowed_we;
	wire [31:0] classb_phase2_cyc_shadowed_qs;
	wire [31:0] classb_phase2_cyc_shadowed_wd;
	wire classb_phase2_cyc_shadowed_storage_err;
	wire classb_phase2_cyc_shadowed_update_err;
	wire classb_phase3_cyc_shadowed_re;
	wire classb_phase3_cyc_shadowed_we;
	wire [31:0] classb_phase3_cyc_shadowed_qs;
	wire [31:0] classb_phase3_cyc_shadowed_wd;
	wire classb_phase3_cyc_shadowed_storage_err;
	wire classb_phase3_cyc_shadowed_update_err;
	wire classb_esc_cnt_re;
	wire [31:0] classb_esc_cnt_qs;
	wire classb_state_re;
	wire [2:0] classb_state_qs;
	wire classc_regwen_we;
	wire classc_regwen_qs;
	wire classc_regwen_wd;
	wire classc_ctrl_shadowed_re;
	wire classc_ctrl_shadowed_we;
	wire classc_ctrl_shadowed_en_qs;
	wire classc_ctrl_shadowed_en_wd;
	wire classc_ctrl_shadowed_en_storage_err;
	wire classc_ctrl_shadowed_en_update_err;
	wire classc_ctrl_shadowed_lock_qs;
	wire classc_ctrl_shadowed_lock_wd;
	wire classc_ctrl_shadowed_lock_storage_err;
	wire classc_ctrl_shadowed_lock_update_err;
	wire classc_ctrl_shadowed_en_e0_qs;
	wire classc_ctrl_shadowed_en_e0_wd;
	wire classc_ctrl_shadowed_en_e0_storage_err;
	wire classc_ctrl_shadowed_en_e0_update_err;
	wire classc_ctrl_shadowed_en_e1_qs;
	wire classc_ctrl_shadowed_en_e1_wd;
	wire classc_ctrl_shadowed_en_e1_storage_err;
	wire classc_ctrl_shadowed_en_e1_update_err;
	wire classc_ctrl_shadowed_en_e2_qs;
	wire classc_ctrl_shadowed_en_e2_wd;
	wire classc_ctrl_shadowed_en_e2_storage_err;
	wire classc_ctrl_shadowed_en_e2_update_err;
	wire classc_ctrl_shadowed_en_e3_qs;
	wire classc_ctrl_shadowed_en_e3_wd;
	wire classc_ctrl_shadowed_en_e3_storage_err;
	wire classc_ctrl_shadowed_en_e3_update_err;
	wire [1:0] classc_ctrl_shadowed_map_e0_qs;
	wire [1:0] classc_ctrl_shadowed_map_e0_wd;
	wire classc_ctrl_shadowed_map_e0_storage_err;
	wire classc_ctrl_shadowed_map_e0_update_err;
	wire [1:0] classc_ctrl_shadowed_map_e1_qs;
	wire [1:0] classc_ctrl_shadowed_map_e1_wd;
	wire classc_ctrl_shadowed_map_e1_storage_err;
	wire classc_ctrl_shadowed_map_e1_update_err;
	wire [1:0] classc_ctrl_shadowed_map_e2_qs;
	wire [1:0] classc_ctrl_shadowed_map_e2_wd;
	wire classc_ctrl_shadowed_map_e2_storage_err;
	wire classc_ctrl_shadowed_map_e2_update_err;
	wire [1:0] classc_ctrl_shadowed_map_e3_qs;
	wire [1:0] classc_ctrl_shadowed_map_e3_wd;
	wire classc_ctrl_shadowed_map_e3_storage_err;
	wire classc_ctrl_shadowed_map_e3_update_err;
	wire classc_clr_regwen_we;
	wire classc_clr_regwen_qs;
	wire classc_clr_regwen_wd;
	wire classc_clr_shadowed_re;
	wire classc_clr_shadowed_we;
	wire classc_clr_shadowed_qs;
	wire classc_clr_shadowed_wd;
	wire classc_clr_shadowed_storage_err;
	wire classc_clr_shadowed_update_err;
	wire classc_accum_cnt_re;
	wire [15:0] classc_accum_cnt_qs;
	wire classc_accum_thresh_shadowed_re;
	wire classc_accum_thresh_shadowed_we;
	wire [15:0] classc_accum_thresh_shadowed_qs;
	wire [15:0] classc_accum_thresh_shadowed_wd;
	wire classc_accum_thresh_shadowed_storage_err;
	wire classc_accum_thresh_shadowed_update_err;
	wire classc_timeout_cyc_shadowed_re;
	wire classc_timeout_cyc_shadowed_we;
	wire [31:0] classc_timeout_cyc_shadowed_qs;
	wire [31:0] classc_timeout_cyc_shadowed_wd;
	wire classc_timeout_cyc_shadowed_storage_err;
	wire classc_timeout_cyc_shadowed_update_err;
	wire classc_crashdump_trigger_shadowed_re;
	wire classc_crashdump_trigger_shadowed_we;
	wire [1:0] classc_crashdump_trigger_shadowed_qs;
	wire [1:0] classc_crashdump_trigger_shadowed_wd;
	wire classc_crashdump_trigger_shadowed_storage_err;
	wire classc_crashdump_trigger_shadowed_update_err;
	wire classc_phase0_cyc_shadowed_re;
	wire classc_phase0_cyc_shadowed_we;
	wire [31:0] classc_phase0_cyc_shadowed_qs;
	wire [31:0] classc_phase0_cyc_shadowed_wd;
	wire classc_phase0_cyc_shadowed_storage_err;
	wire classc_phase0_cyc_shadowed_update_err;
	wire classc_phase1_cyc_shadowed_re;
	wire classc_phase1_cyc_shadowed_we;
	wire [31:0] classc_phase1_cyc_shadowed_qs;
	wire [31:0] classc_phase1_cyc_shadowed_wd;
	wire classc_phase1_cyc_shadowed_storage_err;
	wire classc_phase1_cyc_shadowed_update_err;
	wire classc_phase2_cyc_shadowed_re;
	wire classc_phase2_cyc_shadowed_we;
	wire [31:0] classc_phase2_cyc_shadowed_qs;
	wire [31:0] classc_phase2_cyc_shadowed_wd;
	wire classc_phase2_cyc_shadowed_storage_err;
	wire classc_phase2_cyc_shadowed_update_err;
	wire classc_phase3_cyc_shadowed_re;
	wire classc_phase3_cyc_shadowed_we;
	wire [31:0] classc_phase3_cyc_shadowed_qs;
	wire [31:0] classc_phase3_cyc_shadowed_wd;
	wire classc_phase3_cyc_shadowed_storage_err;
	wire classc_phase3_cyc_shadowed_update_err;
	wire classc_esc_cnt_re;
	wire [31:0] classc_esc_cnt_qs;
	wire classc_state_re;
	wire [2:0] classc_state_qs;
	wire classd_regwen_we;
	wire classd_regwen_qs;
	wire classd_regwen_wd;
	wire classd_ctrl_shadowed_re;
	wire classd_ctrl_shadowed_we;
	wire classd_ctrl_shadowed_en_qs;
	wire classd_ctrl_shadowed_en_wd;
	wire classd_ctrl_shadowed_en_storage_err;
	wire classd_ctrl_shadowed_en_update_err;
	wire classd_ctrl_shadowed_lock_qs;
	wire classd_ctrl_shadowed_lock_wd;
	wire classd_ctrl_shadowed_lock_storage_err;
	wire classd_ctrl_shadowed_lock_update_err;
	wire classd_ctrl_shadowed_en_e0_qs;
	wire classd_ctrl_shadowed_en_e0_wd;
	wire classd_ctrl_shadowed_en_e0_storage_err;
	wire classd_ctrl_shadowed_en_e0_update_err;
	wire classd_ctrl_shadowed_en_e1_qs;
	wire classd_ctrl_shadowed_en_e1_wd;
	wire classd_ctrl_shadowed_en_e1_storage_err;
	wire classd_ctrl_shadowed_en_e1_update_err;
	wire classd_ctrl_shadowed_en_e2_qs;
	wire classd_ctrl_shadowed_en_e2_wd;
	wire classd_ctrl_shadowed_en_e2_storage_err;
	wire classd_ctrl_shadowed_en_e2_update_err;
	wire classd_ctrl_shadowed_en_e3_qs;
	wire classd_ctrl_shadowed_en_e3_wd;
	wire classd_ctrl_shadowed_en_e3_storage_err;
	wire classd_ctrl_shadowed_en_e3_update_err;
	wire [1:0] classd_ctrl_shadowed_map_e0_qs;
	wire [1:0] classd_ctrl_shadowed_map_e0_wd;
	wire classd_ctrl_shadowed_map_e0_storage_err;
	wire classd_ctrl_shadowed_map_e0_update_err;
	wire [1:0] classd_ctrl_shadowed_map_e1_qs;
	wire [1:0] classd_ctrl_shadowed_map_e1_wd;
	wire classd_ctrl_shadowed_map_e1_storage_err;
	wire classd_ctrl_shadowed_map_e1_update_err;
	wire [1:0] classd_ctrl_shadowed_map_e2_qs;
	wire [1:0] classd_ctrl_shadowed_map_e2_wd;
	wire classd_ctrl_shadowed_map_e2_storage_err;
	wire classd_ctrl_shadowed_map_e2_update_err;
	wire [1:0] classd_ctrl_shadowed_map_e3_qs;
	wire [1:0] classd_ctrl_shadowed_map_e3_wd;
	wire classd_ctrl_shadowed_map_e3_storage_err;
	wire classd_ctrl_shadowed_map_e3_update_err;
	wire classd_clr_regwen_we;
	wire classd_clr_regwen_qs;
	wire classd_clr_regwen_wd;
	wire classd_clr_shadowed_re;
	wire classd_clr_shadowed_we;
	wire classd_clr_shadowed_qs;
	wire classd_clr_shadowed_wd;
	wire classd_clr_shadowed_storage_err;
	wire classd_clr_shadowed_update_err;
	wire classd_accum_cnt_re;
	wire [15:0] classd_accum_cnt_qs;
	wire classd_accum_thresh_shadowed_re;
	wire classd_accum_thresh_shadowed_we;
	wire [15:0] classd_accum_thresh_shadowed_qs;
	wire [15:0] classd_accum_thresh_shadowed_wd;
	wire classd_accum_thresh_shadowed_storage_err;
	wire classd_accum_thresh_shadowed_update_err;
	wire classd_timeout_cyc_shadowed_re;
	wire classd_timeout_cyc_shadowed_we;
	wire [31:0] classd_timeout_cyc_shadowed_qs;
	wire [31:0] classd_timeout_cyc_shadowed_wd;
	wire classd_timeout_cyc_shadowed_storage_err;
	wire classd_timeout_cyc_shadowed_update_err;
	wire classd_crashdump_trigger_shadowed_re;
	wire classd_crashdump_trigger_shadowed_we;
	wire [1:0] classd_crashdump_trigger_shadowed_qs;
	wire [1:0] classd_crashdump_trigger_shadowed_wd;
	wire classd_crashdump_trigger_shadowed_storage_err;
	wire classd_crashdump_trigger_shadowed_update_err;
	wire classd_phase0_cyc_shadowed_re;
	wire classd_phase0_cyc_shadowed_we;
	wire [31:0] classd_phase0_cyc_shadowed_qs;
	wire [31:0] classd_phase0_cyc_shadowed_wd;
	wire classd_phase0_cyc_shadowed_storage_err;
	wire classd_phase0_cyc_shadowed_update_err;
	wire classd_phase1_cyc_shadowed_re;
	wire classd_phase1_cyc_shadowed_we;
	wire [31:0] classd_phase1_cyc_shadowed_qs;
	wire [31:0] classd_phase1_cyc_shadowed_wd;
	wire classd_phase1_cyc_shadowed_storage_err;
	wire classd_phase1_cyc_shadowed_update_err;
	wire classd_phase2_cyc_shadowed_re;
	wire classd_phase2_cyc_shadowed_we;
	wire [31:0] classd_phase2_cyc_shadowed_qs;
	wire [31:0] classd_phase2_cyc_shadowed_wd;
	wire classd_phase2_cyc_shadowed_storage_err;
	wire classd_phase2_cyc_shadowed_update_err;
	wire classd_phase3_cyc_shadowed_re;
	wire classd_phase3_cyc_shadowed_we;
	wire [31:0] classd_phase3_cyc_shadowed_qs;
	wire [31:0] classd_phase3_cyc_shadowed_wd;
	wire classd_phase3_cyc_shadowed_storage_err;
	wire classd_phase3_cyc_shadowed_update_err;
	wire classd_esc_cnt_re;
	wire [31:0] classd_esc_cnt_qs;
	wire classd_state_re;
	wire [2:0] classd_state_qs;
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_intr_state_classa(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_we),
		.wd(intr_state_classa_wd),
		.de(hw2reg[362]),
		.d(hw2reg[363]),
		.q(reg2hw[1161]),
		.qs(intr_state_classa_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_intr_state_classb(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_we),
		.wd(intr_state_classb_wd),
		.de(hw2reg[360]),
		.d(hw2reg[361]),
		.q(reg2hw[1160]),
		.qs(intr_state_classb_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_intr_state_classc(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_we),
		.wd(intr_state_classc_wd),
		.de(hw2reg[358]),
		.d(hw2reg[359]),
		.q(reg2hw[1159]),
		.qs(intr_state_classc_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_intr_state_classd(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_we),
		.wd(intr_state_classd_wd),
		.de(hw2reg[356]),
		.d(hw2reg[357]),
		.q(reg2hw[1158]),
		.qs(intr_state_classd_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_intr_enable_classa(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_we),
		.wd(intr_enable_classa_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1157]),
		.qs(intr_enable_classa_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_intr_enable_classb(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_we),
		.wd(intr_enable_classb_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1156]),
		.qs(intr_enable_classb_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_intr_enable_classc(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_we),
		.wd(intr_enable_classc_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1155]),
		.qs(intr_enable_classc_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_intr_enable_classd(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_we),
		.wd(intr_enable_classd_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1154]),
		.qs(intr_enable_classd_qs)
	);
	wire intr_test_qe;
	wire [3:0] intr_test_flds_we;
	assign intr_test_qe = &intr_test_flds_we;
	prim_subreg_ext #(.DW(1)) u_intr_test_classa(
		.re(1'b0),
		.we(intr_test_we),
		.wd(intr_test_classa_wd),
		.d(1'sb0),
		.qe(intr_test_flds_we[0]),
		.q(reg2hw[1153])
	);
	assign reg2hw[1152] = intr_test_qe;
	prim_subreg_ext #(.DW(1)) u_intr_test_classb(
		.re(1'b0),
		.we(intr_test_we),
		.wd(intr_test_classb_wd),
		.d(1'sb0),
		.qe(intr_test_flds_we[1]),
		.q(reg2hw[1151])
	);
	assign reg2hw[1150] = intr_test_qe;
	prim_subreg_ext #(.DW(1)) u_intr_test_classc(
		.re(1'b0),
		.we(intr_test_we),
		.wd(intr_test_classc_wd),
		.d(1'sb0),
		.qe(intr_test_flds_we[2]),
		.q(reg2hw[1149])
	);
	assign reg2hw[1148] = intr_test_qe;
	prim_subreg_ext #(.DW(1)) u_intr_test_classd(
		.re(1'b0),
		.we(intr_test_we),
		.wd(intr_test_classd_wd),
		.d(1'sb0),
		.qe(intr_test_flds_we[3]),
		.q(reg2hw[1147])
	);
	assign reg2hw[1146] = intr_test_qe;
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_ping_timer_regwen(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ping_timer_regwen_we),
		.wd(ping_timer_regwen_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(ping_timer_regwen_qs)
	);
	wire ping_timeout_cyc_shadowed_gated_we;
	assign ping_timeout_cyc_shadowed_gated_we = ping_timeout_cyc_shadowed_we & ping_timer_regwen_qs;
	prim_subreg_shadow #(
		.DW(16),
		.SwAccess(3'd0),
		.RESVAL(16'h0100)
	) u_ping_timeout_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(ping_timeout_cyc_shadowed_re),
		.we(ping_timeout_cyc_shadowed_gated_we),
		.wd(ping_timeout_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1145-:16]),
		.qs(ping_timeout_cyc_shadowed_qs),
		.err_update(ping_timeout_cyc_shadowed_update_err),
		.err_storage(ping_timeout_cyc_shadowed_storage_err)
	);
	wire ping_timer_en_shadowed_gated_we;
	assign ping_timer_en_shadowed_gated_we = ping_timer_en_shadowed_we & ping_timer_regwen_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd4),
		.RESVAL(1'h0)
	) u_ping_timer_en_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(ping_timer_en_shadowed_re),
		.we(ping_timer_en_shadowed_gated_we),
		.wd(ping_timer_en_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1129]),
		.qs(ping_timer_en_shadowed_qs),
		.err_update(ping_timer_en_shadowed_update_err),
		.err_storage(ping_timer_en_shadowed_storage_err)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_0_we),
		.wd(alert_regwen_0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1064]),
		.qs(alert_regwen_0_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_1_we),
		.wd(alert_regwen_1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1065]),
		.qs(alert_regwen_1_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_2_we),
		.wd(alert_regwen_2_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1066]),
		.qs(alert_regwen_2_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_3_we),
		.wd(alert_regwen_3_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1067]),
		.qs(alert_regwen_3_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_4_we),
		.wd(alert_regwen_4_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1068]),
		.qs(alert_regwen_4_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_5_we),
		.wd(alert_regwen_5_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1069]),
		.qs(alert_regwen_5_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_6_we),
		.wd(alert_regwen_6_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1070]),
		.qs(alert_regwen_6_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_7_we),
		.wd(alert_regwen_7_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1071]),
		.qs(alert_regwen_7_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_8_we),
		.wd(alert_regwen_8_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1072]),
		.qs(alert_regwen_8_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_9_we),
		.wd(alert_regwen_9_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1073]),
		.qs(alert_regwen_9_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_10_we),
		.wd(alert_regwen_10_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1074]),
		.qs(alert_regwen_10_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_11_we),
		.wd(alert_regwen_11_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1075]),
		.qs(alert_regwen_11_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_12_we),
		.wd(alert_regwen_12_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1076]),
		.qs(alert_regwen_12_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_13_we),
		.wd(alert_regwen_13_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1077]),
		.qs(alert_regwen_13_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_14_we),
		.wd(alert_regwen_14_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1078]),
		.qs(alert_regwen_14_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_15_we),
		.wd(alert_regwen_15_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1079]),
		.qs(alert_regwen_15_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_16_we),
		.wd(alert_regwen_16_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1080]),
		.qs(alert_regwen_16_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_17_we),
		.wd(alert_regwen_17_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1081]),
		.qs(alert_regwen_17_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_18_we),
		.wd(alert_regwen_18_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1082]),
		.qs(alert_regwen_18_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_19_we),
		.wd(alert_regwen_19_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1083]),
		.qs(alert_regwen_19_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_20_we),
		.wd(alert_regwen_20_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1084]),
		.qs(alert_regwen_20_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_21_we),
		.wd(alert_regwen_21_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1085]),
		.qs(alert_regwen_21_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_22_we),
		.wd(alert_regwen_22_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1086]),
		.qs(alert_regwen_22_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_23_we),
		.wd(alert_regwen_23_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1087]),
		.qs(alert_regwen_23_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_24_we),
		.wd(alert_regwen_24_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1088]),
		.qs(alert_regwen_24_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_25_we),
		.wd(alert_regwen_25_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1089]),
		.qs(alert_regwen_25_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_26_we),
		.wd(alert_regwen_26_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1090]),
		.qs(alert_regwen_26_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_27_we),
		.wd(alert_regwen_27_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1091]),
		.qs(alert_regwen_27_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_28_we),
		.wd(alert_regwen_28_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1092]),
		.qs(alert_regwen_28_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_29_we),
		.wd(alert_regwen_29_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1093]),
		.qs(alert_regwen_29_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_30_we),
		.wd(alert_regwen_30_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1094]),
		.qs(alert_regwen_30_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_31_we),
		.wd(alert_regwen_31_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1095]),
		.qs(alert_regwen_31_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_32(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_32_we),
		.wd(alert_regwen_32_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1096]),
		.qs(alert_regwen_32_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_33(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_33_we),
		.wd(alert_regwen_33_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1097]),
		.qs(alert_regwen_33_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_34(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_34_we),
		.wd(alert_regwen_34_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1098]),
		.qs(alert_regwen_34_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_35(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_35_we),
		.wd(alert_regwen_35_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1099]),
		.qs(alert_regwen_35_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_36(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_36_we),
		.wd(alert_regwen_36_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1100]),
		.qs(alert_regwen_36_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_37(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_37_we),
		.wd(alert_regwen_37_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1101]),
		.qs(alert_regwen_37_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_38(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_38_we),
		.wd(alert_regwen_38_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1102]),
		.qs(alert_regwen_38_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_39(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_39_we),
		.wd(alert_regwen_39_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1103]),
		.qs(alert_regwen_39_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_40(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_40_we),
		.wd(alert_regwen_40_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1104]),
		.qs(alert_regwen_40_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_41(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_41_we),
		.wd(alert_regwen_41_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1105]),
		.qs(alert_regwen_41_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_42(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_42_we),
		.wd(alert_regwen_42_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1106]),
		.qs(alert_regwen_42_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_43(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_43_we),
		.wd(alert_regwen_43_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1107]),
		.qs(alert_regwen_43_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_44(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_44_we),
		.wd(alert_regwen_44_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1108]),
		.qs(alert_regwen_44_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_45(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_45_we),
		.wd(alert_regwen_45_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1109]),
		.qs(alert_regwen_45_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_46(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_46_we),
		.wd(alert_regwen_46_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1110]),
		.qs(alert_regwen_46_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_47(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_47_we),
		.wd(alert_regwen_47_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1111]),
		.qs(alert_regwen_47_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_48(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_48_we),
		.wd(alert_regwen_48_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1112]),
		.qs(alert_regwen_48_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_49(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_49_we),
		.wd(alert_regwen_49_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1113]),
		.qs(alert_regwen_49_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_50(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_50_we),
		.wd(alert_regwen_50_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1114]),
		.qs(alert_regwen_50_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_51(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_51_we),
		.wd(alert_regwen_51_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1115]),
		.qs(alert_regwen_51_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_52(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_52_we),
		.wd(alert_regwen_52_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1116]),
		.qs(alert_regwen_52_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_53(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_53_we),
		.wd(alert_regwen_53_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1117]),
		.qs(alert_regwen_53_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_54(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_54_we),
		.wd(alert_regwen_54_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1118]),
		.qs(alert_regwen_54_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_55(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_55_we),
		.wd(alert_regwen_55_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1119]),
		.qs(alert_regwen_55_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_56(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_56_we),
		.wd(alert_regwen_56_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1120]),
		.qs(alert_regwen_56_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_57(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_57_we),
		.wd(alert_regwen_57_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1121]),
		.qs(alert_regwen_57_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_58(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_58_we),
		.wd(alert_regwen_58_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1122]),
		.qs(alert_regwen_58_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_59(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_59_we),
		.wd(alert_regwen_59_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1123]),
		.qs(alert_regwen_59_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_60(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_60_we),
		.wd(alert_regwen_60_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1124]),
		.qs(alert_regwen_60_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_61(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_61_we),
		.wd(alert_regwen_61_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1125]),
		.qs(alert_regwen_61_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_62(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_62_we),
		.wd(alert_regwen_62_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1126]),
		.qs(alert_regwen_62_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_63(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_63_we),
		.wd(alert_regwen_63_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1127]),
		.qs(alert_regwen_63_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_alert_regwen_64(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_regwen_64_we),
		.wd(alert_regwen_64_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1128]),
		.qs(alert_regwen_64_qs)
	);
	wire alert_en_shadowed_0_gated_we;
	assign alert_en_shadowed_0_gated_we = alert_en_shadowed_0_we & alert_regwen_0_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_0_re),
		.we(alert_en_shadowed_0_gated_we),
		.wd(alert_en_shadowed_0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[999]),
		.qs(alert_en_shadowed_0_qs),
		.err_update(alert_en_shadowed_0_update_err),
		.err_storage(alert_en_shadowed_0_storage_err)
	);
	wire alert_en_shadowed_1_gated_we;
	assign alert_en_shadowed_1_gated_we = alert_en_shadowed_1_we & alert_regwen_1_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_1_re),
		.we(alert_en_shadowed_1_gated_we),
		.wd(alert_en_shadowed_1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1000]),
		.qs(alert_en_shadowed_1_qs),
		.err_update(alert_en_shadowed_1_update_err),
		.err_storage(alert_en_shadowed_1_storage_err)
	);
	wire alert_en_shadowed_2_gated_we;
	assign alert_en_shadowed_2_gated_we = alert_en_shadowed_2_we & alert_regwen_2_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_2_re),
		.we(alert_en_shadowed_2_gated_we),
		.wd(alert_en_shadowed_2_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1001]),
		.qs(alert_en_shadowed_2_qs),
		.err_update(alert_en_shadowed_2_update_err),
		.err_storage(alert_en_shadowed_2_storage_err)
	);
	wire alert_en_shadowed_3_gated_we;
	assign alert_en_shadowed_3_gated_we = alert_en_shadowed_3_we & alert_regwen_3_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_3_re),
		.we(alert_en_shadowed_3_gated_we),
		.wd(alert_en_shadowed_3_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1002]),
		.qs(alert_en_shadowed_3_qs),
		.err_update(alert_en_shadowed_3_update_err),
		.err_storage(alert_en_shadowed_3_storage_err)
	);
	wire alert_en_shadowed_4_gated_we;
	assign alert_en_shadowed_4_gated_we = alert_en_shadowed_4_we & alert_regwen_4_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_4_re),
		.we(alert_en_shadowed_4_gated_we),
		.wd(alert_en_shadowed_4_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1003]),
		.qs(alert_en_shadowed_4_qs),
		.err_update(alert_en_shadowed_4_update_err),
		.err_storage(alert_en_shadowed_4_storage_err)
	);
	wire alert_en_shadowed_5_gated_we;
	assign alert_en_shadowed_5_gated_we = alert_en_shadowed_5_we & alert_regwen_5_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_5_re),
		.we(alert_en_shadowed_5_gated_we),
		.wd(alert_en_shadowed_5_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1004]),
		.qs(alert_en_shadowed_5_qs),
		.err_update(alert_en_shadowed_5_update_err),
		.err_storage(alert_en_shadowed_5_storage_err)
	);
	wire alert_en_shadowed_6_gated_we;
	assign alert_en_shadowed_6_gated_we = alert_en_shadowed_6_we & alert_regwen_6_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_6_re),
		.we(alert_en_shadowed_6_gated_we),
		.wd(alert_en_shadowed_6_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1005]),
		.qs(alert_en_shadowed_6_qs),
		.err_update(alert_en_shadowed_6_update_err),
		.err_storage(alert_en_shadowed_6_storage_err)
	);
	wire alert_en_shadowed_7_gated_we;
	assign alert_en_shadowed_7_gated_we = alert_en_shadowed_7_we & alert_regwen_7_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_7_re),
		.we(alert_en_shadowed_7_gated_we),
		.wd(alert_en_shadowed_7_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1006]),
		.qs(alert_en_shadowed_7_qs),
		.err_update(alert_en_shadowed_7_update_err),
		.err_storage(alert_en_shadowed_7_storage_err)
	);
	wire alert_en_shadowed_8_gated_we;
	assign alert_en_shadowed_8_gated_we = alert_en_shadowed_8_we & alert_regwen_8_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_8_re),
		.we(alert_en_shadowed_8_gated_we),
		.wd(alert_en_shadowed_8_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1007]),
		.qs(alert_en_shadowed_8_qs),
		.err_update(alert_en_shadowed_8_update_err),
		.err_storage(alert_en_shadowed_8_storage_err)
	);
	wire alert_en_shadowed_9_gated_we;
	assign alert_en_shadowed_9_gated_we = alert_en_shadowed_9_we & alert_regwen_9_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_9_re),
		.we(alert_en_shadowed_9_gated_we),
		.wd(alert_en_shadowed_9_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1008]),
		.qs(alert_en_shadowed_9_qs),
		.err_update(alert_en_shadowed_9_update_err),
		.err_storage(alert_en_shadowed_9_storage_err)
	);
	wire alert_en_shadowed_10_gated_we;
	assign alert_en_shadowed_10_gated_we = alert_en_shadowed_10_we & alert_regwen_10_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_10_re),
		.we(alert_en_shadowed_10_gated_we),
		.wd(alert_en_shadowed_10_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1009]),
		.qs(alert_en_shadowed_10_qs),
		.err_update(alert_en_shadowed_10_update_err),
		.err_storage(alert_en_shadowed_10_storage_err)
	);
	wire alert_en_shadowed_11_gated_we;
	assign alert_en_shadowed_11_gated_we = alert_en_shadowed_11_we & alert_regwen_11_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_11_re),
		.we(alert_en_shadowed_11_gated_we),
		.wd(alert_en_shadowed_11_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1010]),
		.qs(alert_en_shadowed_11_qs),
		.err_update(alert_en_shadowed_11_update_err),
		.err_storage(alert_en_shadowed_11_storage_err)
	);
	wire alert_en_shadowed_12_gated_we;
	assign alert_en_shadowed_12_gated_we = alert_en_shadowed_12_we & alert_regwen_12_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_12_re),
		.we(alert_en_shadowed_12_gated_we),
		.wd(alert_en_shadowed_12_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1011]),
		.qs(alert_en_shadowed_12_qs),
		.err_update(alert_en_shadowed_12_update_err),
		.err_storage(alert_en_shadowed_12_storage_err)
	);
	wire alert_en_shadowed_13_gated_we;
	assign alert_en_shadowed_13_gated_we = alert_en_shadowed_13_we & alert_regwen_13_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_13_re),
		.we(alert_en_shadowed_13_gated_we),
		.wd(alert_en_shadowed_13_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1012]),
		.qs(alert_en_shadowed_13_qs),
		.err_update(alert_en_shadowed_13_update_err),
		.err_storage(alert_en_shadowed_13_storage_err)
	);
	wire alert_en_shadowed_14_gated_we;
	assign alert_en_shadowed_14_gated_we = alert_en_shadowed_14_we & alert_regwen_14_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_14_re),
		.we(alert_en_shadowed_14_gated_we),
		.wd(alert_en_shadowed_14_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1013]),
		.qs(alert_en_shadowed_14_qs),
		.err_update(alert_en_shadowed_14_update_err),
		.err_storage(alert_en_shadowed_14_storage_err)
	);
	wire alert_en_shadowed_15_gated_we;
	assign alert_en_shadowed_15_gated_we = alert_en_shadowed_15_we & alert_regwen_15_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_15_re),
		.we(alert_en_shadowed_15_gated_we),
		.wd(alert_en_shadowed_15_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1014]),
		.qs(alert_en_shadowed_15_qs),
		.err_update(alert_en_shadowed_15_update_err),
		.err_storage(alert_en_shadowed_15_storage_err)
	);
	wire alert_en_shadowed_16_gated_we;
	assign alert_en_shadowed_16_gated_we = alert_en_shadowed_16_we & alert_regwen_16_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_16_re),
		.we(alert_en_shadowed_16_gated_we),
		.wd(alert_en_shadowed_16_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1015]),
		.qs(alert_en_shadowed_16_qs),
		.err_update(alert_en_shadowed_16_update_err),
		.err_storage(alert_en_shadowed_16_storage_err)
	);
	wire alert_en_shadowed_17_gated_we;
	assign alert_en_shadowed_17_gated_we = alert_en_shadowed_17_we & alert_regwen_17_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_17_re),
		.we(alert_en_shadowed_17_gated_we),
		.wd(alert_en_shadowed_17_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1016]),
		.qs(alert_en_shadowed_17_qs),
		.err_update(alert_en_shadowed_17_update_err),
		.err_storage(alert_en_shadowed_17_storage_err)
	);
	wire alert_en_shadowed_18_gated_we;
	assign alert_en_shadowed_18_gated_we = alert_en_shadowed_18_we & alert_regwen_18_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_18_re),
		.we(alert_en_shadowed_18_gated_we),
		.wd(alert_en_shadowed_18_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1017]),
		.qs(alert_en_shadowed_18_qs),
		.err_update(alert_en_shadowed_18_update_err),
		.err_storage(alert_en_shadowed_18_storage_err)
	);
	wire alert_en_shadowed_19_gated_we;
	assign alert_en_shadowed_19_gated_we = alert_en_shadowed_19_we & alert_regwen_19_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_19_re),
		.we(alert_en_shadowed_19_gated_we),
		.wd(alert_en_shadowed_19_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1018]),
		.qs(alert_en_shadowed_19_qs),
		.err_update(alert_en_shadowed_19_update_err),
		.err_storage(alert_en_shadowed_19_storage_err)
	);
	wire alert_en_shadowed_20_gated_we;
	assign alert_en_shadowed_20_gated_we = alert_en_shadowed_20_we & alert_regwen_20_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_20_re),
		.we(alert_en_shadowed_20_gated_we),
		.wd(alert_en_shadowed_20_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1019]),
		.qs(alert_en_shadowed_20_qs),
		.err_update(alert_en_shadowed_20_update_err),
		.err_storage(alert_en_shadowed_20_storage_err)
	);
	wire alert_en_shadowed_21_gated_we;
	assign alert_en_shadowed_21_gated_we = alert_en_shadowed_21_we & alert_regwen_21_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_21_re),
		.we(alert_en_shadowed_21_gated_we),
		.wd(alert_en_shadowed_21_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1020]),
		.qs(alert_en_shadowed_21_qs),
		.err_update(alert_en_shadowed_21_update_err),
		.err_storage(alert_en_shadowed_21_storage_err)
	);
	wire alert_en_shadowed_22_gated_we;
	assign alert_en_shadowed_22_gated_we = alert_en_shadowed_22_we & alert_regwen_22_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_22_re),
		.we(alert_en_shadowed_22_gated_we),
		.wd(alert_en_shadowed_22_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1021]),
		.qs(alert_en_shadowed_22_qs),
		.err_update(alert_en_shadowed_22_update_err),
		.err_storage(alert_en_shadowed_22_storage_err)
	);
	wire alert_en_shadowed_23_gated_we;
	assign alert_en_shadowed_23_gated_we = alert_en_shadowed_23_we & alert_regwen_23_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_23_re),
		.we(alert_en_shadowed_23_gated_we),
		.wd(alert_en_shadowed_23_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1022]),
		.qs(alert_en_shadowed_23_qs),
		.err_update(alert_en_shadowed_23_update_err),
		.err_storage(alert_en_shadowed_23_storage_err)
	);
	wire alert_en_shadowed_24_gated_we;
	assign alert_en_shadowed_24_gated_we = alert_en_shadowed_24_we & alert_regwen_24_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_24_re),
		.we(alert_en_shadowed_24_gated_we),
		.wd(alert_en_shadowed_24_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1023]),
		.qs(alert_en_shadowed_24_qs),
		.err_update(alert_en_shadowed_24_update_err),
		.err_storage(alert_en_shadowed_24_storage_err)
	);
	wire alert_en_shadowed_25_gated_we;
	assign alert_en_shadowed_25_gated_we = alert_en_shadowed_25_we & alert_regwen_25_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_25_re),
		.we(alert_en_shadowed_25_gated_we),
		.wd(alert_en_shadowed_25_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1024]),
		.qs(alert_en_shadowed_25_qs),
		.err_update(alert_en_shadowed_25_update_err),
		.err_storage(alert_en_shadowed_25_storage_err)
	);
	wire alert_en_shadowed_26_gated_we;
	assign alert_en_shadowed_26_gated_we = alert_en_shadowed_26_we & alert_regwen_26_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_26_re),
		.we(alert_en_shadowed_26_gated_we),
		.wd(alert_en_shadowed_26_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1025]),
		.qs(alert_en_shadowed_26_qs),
		.err_update(alert_en_shadowed_26_update_err),
		.err_storage(alert_en_shadowed_26_storage_err)
	);
	wire alert_en_shadowed_27_gated_we;
	assign alert_en_shadowed_27_gated_we = alert_en_shadowed_27_we & alert_regwen_27_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_27_re),
		.we(alert_en_shadowed_27_gated_we),
		.wd(alert_en_shadowed_27_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1026]),
		.qs(alert_en_shadowed_27_qs),
		.err_update(alert_en_shadowed_27_update_err),
		.err_storage(alert_en_shadowed_27_storage_err)
	);
	wire alert_en_shadowed_28_gated_we;
	assign alert_en_shadowed_28_gated_we = alert_en_shadowed_28_we & alert_regwen_28_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_28_re),
		.we(alert_en_shadowed_28_gated_we),
		.wd(alert_en_shadowed_28_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1027]),
		.qs(alert_en_shadowed_28_qs),
		.err_update(alert_en_shadowed_28_update_err),
		.err_storage(alert_en_shadowed_28_storage_err)
	);
	wire alert_en_shadowed_29_gated_we;
	assign alert_en_shadowed_29_gated_we = alert_en_shadowed_29_we & alert_regwen_29_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_29_re),
		.we(alert_en_shadowed_29_gated_we),
		.wd(alert_en_shadowed_29_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1028]),
		.qs(alert_en_shadowed_29_qs),
		.err_update(alert_en_shadowed_29_update_err),
		.err_storage(alert_en_shadowed_29_storage_err)
	);
	wire alert_en_shadowed_30_gated_we;
	assign alert_en_shadowed_30_gated_we = alert_en_shadowed_30_we & alert_regwen_30_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_30_re),
		.we(alert_en_shadowed_30_gated_we),
		.wd(alert_en_shadowed_30_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1029]),
		.qs(alert_en_shadowed_30_qs),
		.err_update(alert_en_shadowed_30_update_err),
		.err_storage(alert_en_shadowed_30_storage_err)
	);
	wire alert_en_shadowed_31_gated_we;
	assign alert_en_shadowed_31_gated_we = alert_en_shadowed_31_we & alert_regwen_31_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_31_re),
		.we(alert_en_shadowed_31_gated_we),
		.wd(alert_en_shadowed_31_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1030]),
		.qs(alert_en_shadowed_31_qs),
		.err_update(alert_en_shadowed_31_update_err),
		.err_storage(alert_en_shadowed_31_storage_err)
	);
	wire alert_en_shadowed_32_gated_we;
	assign alert_en_shadowed_32_gated_we = alert_en_shadowed_32_we & alert_regwen_32_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_32(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_32_re),
		.we(alert_en_shadowed_32_gated_we),
		.wd(alert_en_shadowed_32_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1031]),
		.qs(alert_en_shadowed_32_qs),
		.err_update(alert_en_shadowed_32_update_err),
		.err_storage(alert_en_shadowed_32_storage_err)
	);
	wire alert_en_shadowed_33_gated_we;
	assign alert_en_shadowed_33_gated_we = alert_en_shadowed_33_we & alert_regwen_33_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_33(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_33_re),
		.we(alert_en_shadowed_33_gated_we),
		.wd(alert_en_shadowed_33_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1032]),
		.qs(alert_en_shadowed_33_qs),
		.err_update(alert_en_shadowed_33_update_err),
		.err_storage(alert_en_shadowed_33_storage_err)
	);
	wire alert_en_shadowed_34_gated_we;
	assign alert_en_shadowed_34_gated_we = alert_en_shadowed_34_we & alert_regwen_34_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_34(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_34_re),
		.we(alert_en_shadowed_34_gated_we),
		.wd(alert_en_shadowed_34_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1033]),
		.qs(alert_en_shadowed_34_qs),
		.err_update(alert_en_shadowed_34_update_err),
		.err_storage(alert_en_shadowed_34_storage_err)
	);
	wire alert_en_shadowed_35_gated_we;
	assign alert_en_shadowed_35_gated_we = alert_en_shadowed_35_we & alert_regwen_35_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_35(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_35_re),
		.we(alert_en_shadowed_35_gated_we),
		.wd(alert_en_shadowed_35_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1034]),
		.qs(alert_en_shadowed_35_qs),
		.err_update(alert_en_shadowed_35_update_err),
		.err_storage(alert_en_shadowed_35_storage_err)
	);
	wire alert_en_shadowed_36_gated_we;
	assign alert_en_shadowed_36_gated_we = alert_en_shadowed_36_we & alert_regwen_36_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_36(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_36_re),
		.we(alert_en_shadowed_36_gated_we),
		.wd(alert_en_shadowed_36_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1035]),
		.qs(alert_en_shadowed_36_qs),
		.err_update(alert_en_shadowed_36_update_err),
		.err_storage(alert_en_shadowed_36_storage_err)
	);
	wire alert_en_shadowed_37_gated_we;
	assign alert_en_shadowed_37_gated_we = alert_en_shadowed_37_we & alert_regwen_37_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_37(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_37_re),
		.we(alert_en_shadowed_37_gated_we),
		.wd(alert_en_shadowed_37_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1036]),
		.qs(alert_en_shadowed_37_qs),
		.err_update(alert_en_shadowed_37_update_err),
		.err_storage(alert_en_shadowed_37_storage_err)
	);
	wire alert_en_shadowed_38_gated_we;
	assign alert_en_shadowed_38_gated_we = alert_en_shadowed_38_we & alert_regwen_38_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_38(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_38_re),
		.we(alert_en_shadowed_38_gated_we),
		.wd(alert_en_shadowed_38_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1037]),
		.qs(alert_en_shadowed_38_qs),
		.err_update(alert_en_shadowed_38_update_err),
		.err_storage(alert_en_shadowed_38_storage_err)
	);
	wire alert_en_shadowed_39_gated_we;
	assign alert_en_shadowed_39_gated_we = alert_en_shadowed_39_we & alert_regwen_39_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_39(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_39_re),
		.we(alert_en_shadowed_39_gated_we),
		.wd(alert_en_shadowed_39_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1038]),
		.qs(alert_en_shadowed_39_qs),
		.err_update(alert_en_shadowed_39_update_err),
		.err_storage(alert_en_shadowed_39_storage_err)
	);
	wire alert_en_shadowed_40_gated_we;
	assign alert_en_shadowed_40_gated_we = alert_en_shadowed_40_we & alert_regwen_40_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_40(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_40_re),
		.we(alert_en_shadowed_40_gated_we),
		.wd(alert_en_shadowed_40_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1039]),
		.qs(alert_en_shadowed_40_qs),
		.err_update(alert_en_shadowed_40_update_err),
		.err_storage(alert_en_shadowed_40_storage_err)
	);
	wire alert_en_shadowed_41_gated_we;
	assign alert_en_shadowed_41_gated_we = alert_en_shadowed_41_we & alert_regwen_41_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_41(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_41_re),
		.we(alert_en_shadowed_41_gated_we),
		.wd(alert_en_shadowed_41_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1040]),
		.qs(alert_en_shadowed_41_qs),
		.err_update(alert_en_shadowed_41_update_err),
		.err_storage(alert_en_shadowed_41_storage_err)
	);
	wire alert_en_shadowed_42_gated_we;
	assign alert_en_shadowed_42_gated_we = alert_en_shadowed_42_we & alert_regwen_42_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_42(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_42_re),
		.we(alert_en_shadowed_42_gated_we),
		.wd(alert_en_shadowed_42_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1041]),
		.qs(alert_en_shadowed_42_qs),
		.err_update(alert_en_shadowed_42_update_err),
		.err_storage(alert_en_shadowed_42_storage_err)
	);
	wire alert_en_shadowed_43_gated_we;
	assign alert_en_shadowed_43_gated_we = alert_en_shadowed_43_we & alert_regwen_43_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_43(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_43_re),
		.we(alert_en_shadowed_43_gated_we),
		.wd(alert_en_shadowed_43_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1042]),
		.qs(alert_en_shadowed_43_qs),
		.err_update(alert_en_shadowed_43_update_err),
		.err_storage(alert_en_shadowed_43_storage_err)
	);
	wire alert_en_shadowed_44_gated_we;
	assign alert_en_shadowed_44_gated_we = alert_en_shadowed_44_we & alert_regwen_44_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_44(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_44_re),
		.we(alert_en_shadowed_44_gated_we),
		.wd(alert_en_shadowed_44_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1043]),
		.qs(alert_en_shadowed_44_qs),
		.err_update(alert_en_shadowed_44_update_err),
		.err_storage(alert_en_shadowed_44_storage_err)
	);
	wire alert_en_shadowed_45_gated_we;
	assign alert_en_shadowed_45_gated_we = alert_en_shadowed_45_we & alert_regwen_45_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_45(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_45_re),
		.we(alert_en_shadowed_45_gated_we),
		.wd(alert_en_shadowed_45_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1044]),
		.qs(alert_en_shadowed_45_qs),
		.err_update(alert_en_shadowed_45_update_err),
		.err_storage(alert_en_shadowed_45_storage_err)
	);
	wire alert_en_shadowed_46_gated_we;
	assign alert_en_shadowed_46_gated_we = alert_en_shadowed_46_we & alert_regwen_46_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_46(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_46_re),
		.we(alert_en_shadowed_46_gated_we),
		.wd(alert_en_shadowed_46_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1045]),
		.qs(alert_en_shadowed_46_qs),
		.err_update(alert_en_shadowed_46_update_err),
		.err_storage(alert_en_shadowed_46_storage_err)
	);
	wire alert_en_shadowed_47_gated_we;
	assign alert_en_shadowed_47_gated_we = alert_en_shadowed_47_we & alert_regwen_47_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_47(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_47_re),
		.we(alert_en_shadowed_47_gated_we),
		.wd(alert_en_shadowed_47_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1046]),
		.qs(alert_en_shadowed_47_qs),
		.err_update(alert_en_shadowed_47_update_err),
		.err_storage(alert_en_shadowed_47_storage_err)
	);
	wire alert_en_shadowed_48_gated_we;
	assign alert_en_shadowed_48_gated_we = alert_en_shadowed_48_we & alert_regwen_48_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_48(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_48_re),
		.we(alert_en_shadowed_48_gated_we),
		.wd(alert_en_shadowed_48_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1047]),
		.qs(alert_en_shadowed_48_qs),
		.err_update(alert_en_shadowed_48_update_err),
		.err_storage(alert_en_shadowed_48_storage_err)
	);
	wire alert_en_shadowed_49_gated_we;
	assign alert_en_shadowed_49_gated_we = alert_en_shadowed_49_we & alert_regwen_49_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_49(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_49_re),
		.we(alert_en_shadowed_49_gated_we),
		.wd(alert_en_shadowed_49_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1048]),
		.qs(alert_en_shadowed_49_qs),
		.err_update(alert_en_shadowed_49_update_err),
		.err_storage(alert_en_shadowed_49_storage_err)
	);
	wire alert_en_shadowed_50_gated_we;
	assign alert_en_shadowed_50_gated_we = alert_en_shadowed_50_we & alert_regwen_50_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_50(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_50_re),
		.we(alert_en_shadowed_50_gated_we),
		.wd(alert_en_shadowed_50_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1049]),
		.qs(alert_en_shadowed_50_qs),
		.err_update(alert_en_shadowed_50_update_err),
		.err_storage(alert_en_shadowed_50_storage_err)
	);
	wire alert_en_shadowed_51_gated_we;
	assign alert_en_shadowed_51_gated_we = alert_en_shadowed_51_we & alert_regwen_51_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_51(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_51_re),
		.we(alert_en_shadowed_51_gated_we),
		.wd(alert_en_shadowed_51_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1050]),
		.qs(alert_en_shadowed_51_qs),
		.err_update(alert_en_shadowed_51_update_err),
		.err_storage(alert_en_shadowed_51_storage_err)
	);
	wire alert_en_shadowed_52_gated_we;
	assign alert_en_shadowed_52_gated_we = alert_en_shadowed_52_we & alert_regwen_52_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_52(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_52_re),
		.we(alert_en_shadowed_52_gated_we),
		.wd(alert_en_shadowed_52_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1051]),
		.qs(alert_en_shadowed_52_qs),
		.err_update(alert_en_shadowed_52_update_err),
		.err_storage(alert_en_shadowed_52_storage_err)
	);
	wire alert_en_shadowed_53_gated_we;
	assign alert_en_shadowed_53_gated_we = alert_en_shadowed_53_we & alert_regwen_53_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_53(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_53_re),
		.we(alert_en_shadowed_53_gated_we),
		.wd(alert_en_shadowed_53_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1052]),
		.qs(alert_en_shadowed_53_qs),
		.err_update(alert_en_shadowed_53_update_err),
		.err_storage(alert_en_shadowed_53_storage_err)
	);
	wire alert_en_shadowed_54_gated_we;
	assign alert_en_shadowed_54_gated_we = alert_en_shadowed_54_we & alert_regwen_54_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_54(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_54_re),
		.we(alert_en_shadowed_54_gated_we),
		.wd(alert_en_shadowed_54_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1053]),
		.qs(alert_en_shadowed_54_qs),
		.err_update(alert_en_shadowed_54_update_err),
		.err_storage(alert_en_shadowed_54_storage_err)
	);
	wire alert_en_shadowed_55_gated_we;
	assign alert_en_shadowed_55_gated_we = alert_en_shadowed_55_we & alert_regwen_55_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_55(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_55_re),
		.we(alert_en_shadowed_55_gated_we),
		.wd(alert_en_shadowed_55_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1054]),
		.qs(alert_en_shadowed_55_qs),
		.err_update(alert_en_shadowed_55_update_err),
		.err_storage(alert_en_shadowed_55_storage_err)
	);
	wire alert_en_shadowed_56_gated_we;
	assign alert_en_shadowed_56_gated_we = alert_en_shadowed_56_we & alert_regwen_56_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_56(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_56_re),
		.we(alert_en_shadowed_56_gated_we),
		.wd(alert_en_shadowed_56_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1055]),
		.qs(alert_en_shadowed_56_qs),
		.err_update(alert_en_shadowed_56_update_err),
		.err_storage(alert_en_shadowed_56_storage_err)
	);
	wire alert_en_shadowed_57_gated_we;
	assign alert_en_shadowed_57_gated_we = alert_en_shadowed_57_we & alert_regwen_57_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_57(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_57_re),
		.we(alert_en_shadowed_57_gated_we),
		.wd(alert_en_shadowed_57_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1056]),
		.qs(alert_en_shadowed_57_qs),
		.err_update(alert_en_shadowed_57_update_err),
		.err_storage(alert_en_shadowed_57_storage_err)
	);
	wire alert_en_shadowed_58_gated_we;
	assign alert_en_shadowed_58_gated_we = alert_en_shadowed_58_we & alert_regwen_58_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_58(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_58_re),
		.we(alert_en_shadowed_58_gated_we),
		.wd(alert_en_shadowed_58_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1057]),
		.qs(alert_en_shadowed_58_qs),
		.err_update(alert_en_shadowed_58_update_err),
		.err_storage(alert_en_shadowed_58_storage_err)
	);
	wire alert_en_shadowed_59_gated_we;
	assign alert_en_shadowed_59_gated_we = alert_en_shadowed_59_we & alert_regwen_59_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_59(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_59_re),
		.we(alert_en_shadowed_59_gated_we),
		.wd(alert_en_shadowed_59_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1058]),
		.qs(alert_en_shadowed_59_qs),
		.err_update(alert_en_shadowed_59_update_err),
		.err_storage(alert_en_shadowed_59_storage_err)
	);
	wire alert_en_shadowed_60_gated_we;
	assign alert_en_shadowed_60_gated_we = alert_en_shadowed_60_we & alert_regwen_60_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_60(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_60_re),
		.we(alert_en_shadowed_60_gated_we),
		.wd(alert_en_shadowed_60_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1059]),
		.qs(alert_en_shadowed_60_qs),
		.err_update(alert_en_shadowed_60_update_err),
		.err_storage(alert_en_shadowed_60_storage_err)
	);
	wire alert_en_shadowed_61_gated_we;
	assign alert_en_shadowed_61_gated_we = alert_en_shadowed_61_we & alert_regwen_61_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_61(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_61_re),
		.we(alert_en_shadowed_61_gated_we),
		.wd(alert_en_shadowed_61_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1060]),
		.qs(alert_en_shadowed_61_qs),
		.err_update(alert_en_shadowed_61_update_err),
		.err_storage(alert_en_shadowed_61_storage_err)
	);
	wire alert_en_shadowed_62_gated_we;
	assign alert_en_shadowed_62_gated_we = alert_en_shadowed_62_we & alert_regwen_62_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_62(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_62_re),
		.we(alert_en_shadowed_62_gated_we),
		.wd(alert_en_shadowed_62_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1061]),
		.qs(alert_en_shadowed_62_qs),
		.err_update(alert_en_shadowed_62_update_err),
		.err_storage(alert_en_shadowed_62_storage_err)
	);
	wire alert_en_shadowed_63_gated_we;
	assign alert_en_shadowed_63_gated_we = alert_en_shadowed_63_we & alert_regwen_63_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_63(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_63_re),
		.we(alert_en_shadowed_63_gated_we),
		.wd(alert_en_shadowed_63_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1062]),
		.qs(alert_en_shadowed_63_qs),
		.err_update(alert_en_shadowed_63_update_err),
		.err_storage(alert_en_shadowed_63_storage_err)
	);
	wire alert_en_shadowed_64_gated_we;
	assign alert_en_shadowed_64_gated_we = alert_en_shadowed_64_we & alert_regwen_64_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_alert_en_shadowed_64(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_en_shadowed_64_re),
		.we(alert_en_shadowed_64_gated_we),
		.wd(alert_en_shadowed_64_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[1063]),
		.qs(alert_en_shadowed_64_qs),
		.err_update(alert_en_shadowed_64_update_err),
		.err_storage(alert_en_shadowed_64_storage_err)
	);
	wire alert_class_shadowed_0_gated_we;
	assign alert_class_shadowed_0_gated_we = alert_class_shadowed_0_we & alert_regwen_0_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_0_re),
		.we(alert_class_shadowed_0_gated_we),
		.wd(alert_class_shadowed_0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[870-:2]),
		.qs(alert_class_shadowed_0_qs),
		.err_update(alert_class_shadowed_0_update_err),
		.err_storage(alert_class_shadowed_0_storage_err)
	);
	wire alert_class_shadowed_1_gated_we;
	assign alert_class_shadowed_1_gated_we = alert_class_shadowed_1_we & alert_regwen_1_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_1_re),
		.we(alert_class_shadowed_1_gated_we),
		.wd(alert_class_shadowed_1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[872-:2]),
		.qs(alert_class_shadowed_1_qs),
		.err_update(alert_class_shadowed_1_update_err),
		.err_storage(alert_class_shadowed_1_storage_err)
	);
	wire alert_class_shadowed_2_gated_we;
	assign alert_class_shadowed_2_gated_we = alert_class_shadowed_2_we & alert_regwen_2_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_2_re),
		.we(alert_class_shadowed_2_gated_we),
		.wd(alert_class_shadowed_2_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[874-:2]),
		.qs(alert_class_shadowed_2_qs),
		.err_update(alert_class_shadowed_2_update_err),
		.err_storage(alert_class_shadowed_2_storage_err)
	);
	wire alert_class_shadowed_3_gated_we;
	assign alert_class_shadowed_3_gated_we = alert_class_shadowed_3_we & alert_regwen_3_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_3_re),
		.we(alert_class_shadowed_3_gated_we),
		.wd(alert_class_shadowed_3_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[876-:2]),
		.qs(alert_class_shadowed_3_qs),
		.err_update(alert_class_shadowed_3_update_err),
		.err_storage(alert_class_shadowed_3_storage_err)
	);
	wire alert_class_shadowed_4_gated_we;
	assign alert_class_shadowed_4_gated_we = alert_class_shadowed_4_we & alert_regwen_4_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_4_re),
		.we(alert_class_shadowed_4_gated_we),
		.wd(alert_class_shadowed_4_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[878-:2]),
		.qs(alert_class_shadowed_4_qs),
		.err_update(alert_class_shadowed_4_update_err),
		.err_storage(alert_class_shadowed_4_storage_err)
	);
	wire alert_class_shadowed_5_gated_we;
	assign alert_class_shadowed_5_gated_we = alert_class_shadowed_5_we & alert_regwen_5_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_5_re),
		.we(alert_class_shadowed_5_gated_we),
		.wd(alert_class_shadowed_5_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[880-:2]),
		.qs(alert_class_shadowed_5_qs),
		.err_update(alert_class_shadowed_5_update_err),
		.err_storage(alert_class_shadowed_5_storage_err)
	);
	wire alert_class_shadowed_6_gated_we;
	assign alert_class_shadowed_6_gated_we = alert_class_shadowed_6_we & alert_regwen_6_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_6_re),
		.we(alert_class_shadowed_6_gated_we),
		.wd(alert_class_shadowed_6_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[882-:2]),
		.qs(alert_class_shadowed_6_qs),
		.err_update(alert_class_shadowed_6_update_err),
		.err_storage(alert_class_shadowed_6_storage_err)
	);
	wire alert_class_shadowed_7_gated_we;
	assign alert_class_shadowed_7_gated_we = alert_class_shadowed_7_we & alert_regwen_7_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_7_re),
		.we(alert_class_shadowed_7_gated_we),
		.wd(alert_class_shadowed_7_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[884-:2]),
		.qs(alert_class_shadowed_7_qs),
		.err_update(alert_class_shadowed_7_update_err),
		.err_storage(alert_class_shadowed_7_storage_err)
	);
	wire alert_class_shadowed_8_gated_we;
	assign alert_class_shadowed_8_gated_we = alert_class_shadowed_8_we & alert_regwen_8_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_8_re),
		.we(alert_class_shadowed_8_gated_we),
		.wd(alert_class_shadowed_8_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[886-:2]),
		.qs(alert_class_shadowed_8_qs),
		.err_update(alert_class_shadowed_8_update_err),
		.err_storage(alert_class_shadowed_8_storage_err)
	);
	wire alert_class_shadowed_9_gated_we;
	assign alert_class_shadowed_9_gated_we = alert_class_shadowed_9_we & alert_regwen_9_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_9_re),
		.we(alert_class_shadowed_9_gated_we),
		.wd(alert_class_shadowed_9_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[888-:2]),
		.qs(alert_class_shadowed_9_qs),
		.err_update(alert_class_shadowed_9_update_err),
		.err_storage(alert_class_shadowed_9_storage_err)
	);
	wire alert_class_shadowed_10_gated_we;
	assign alert_class_shadowed_10_gated_we = alert_class_shadowed_10_we & alert_regwen_10_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_10_re),
		.we(alert_class_shadowed_10_gated_we),
		.wd(alert_class_shadowed_10_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[890-:2]),
		.qs(alert_class_shadowed_10_qs),
		.err_update(alert_class_shadowed_10_update_err),
		.err_storage(alert_class_shadowed_10_storage_err)
	);
	wire alert_class_shadowed_11_gated_we;
	assign alert_class_shadowed_11_gated_we = alert_class_shadowed_11_we & alert_regwen_11_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_11_re),
		.we(alert_class_shadowed_11_gated_we),
		.wd(alert_class_shadowed_11_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[892-:2]),
		.qs(alert_class_shadowed_11_qs),
		.err_update(alert_class_shadowed_11_update_err),
		.err_storage(alert_class_shadowed_11_storage_err)
	);
	wire alert_class_shadowed_12_gated_we;
	assign alert_class_shadowed_12_gated_we = alert_class_shadowed_12_we & alert_regwen_12_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_12_re),
		.we(alert_class_shadowed_12_gated_we),
		.wd(alert_class_shadowed_12_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[894-:2]),
		.qs(alert_class_shadowed_12_qs),
		.err_update(alert_class_shadowed_12_update_err),
		.err_storage(alert_class_shadowed_12_storage_err)
	);
	wire alert_class_shadowed_13_gated_we;
	assign alert_class_shadowed_13_gated_we = alert_class_shadowed_13_we & alert_regwen_13_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_13_re),
		.we(alert_class_shadowed_13_gated_we),
		.wd(alert_class_shadowed_13_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[896-:2]),
		.qs(alert_class_shadowed_13_qs),
		.err_update(alert_class_shadowed_13_update_err),
		.err_storage(alert_class_shadowed_13_storage_err)
	);
	wire alert_class_shadowed_14_gated_we;
	assign alert_class_shadowed_14_gated_we = alert_class_shadowed_14_we & alert_regwen_14_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_14_re),
		.we(alert_class_shadowed_14_gated_we),
		.wd(alert_class_shadowed_14_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[898-:2]),
		.qs(alert_class_shadowed_14_qs),
		.err_update(alert_class_shadowed_14_update_err),
		.err_storage(alert_class_shadowed_14_storage_err)
	);
	wire alert_class_shadowed_15_gated_we;
	assign alert_class_shadowed_15_gated_we = alert_class_shadowed_15_we & alert_regwen_15_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_15_re),
		.we(alert_class_shadowed_15_gated_we),
		.wd(alert_class_shadowed_15_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[900-:2]),
		.qs(alert_class_shadowed_15_qs),
		.err_update(alert_class_shadowed_15_update_err),
		.err_storage(alert_class_shadowed_15_storage_err)
	);
	wire alert_class_shadowed_16_gated_we;
	assign alert_class_shadowed_16_gated_we = alert_class_shadowed_16_we & alert_regwen_16_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_16_re),
		.we(alert_class_shadowed_16_gated_we),
		.wd(alert_class_shadowed_16_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[902-:2]),
		.qs(alert_class_shadowed_16_qs),
		.err_update(alert_class_shadowed_16_update_err),
		.err_storage(alert_class_shadowed_16_storage_err)
	);
	wire alert_class_shadowed_17_gated_we;
	assign alert_class_shadowed_17_gated_we = alert_class_shadowed_17_we & alert_regwen_17_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_17_re),
		.we(alert_class_shadowed_17_gated_we),
		.wd(alert_class_shadowed_17_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[904-:2]),
		.qs(alert_class_shadowed_17_qs),
		.err_update(alert_class_shadowed_17_update_err),
		.err_storage(alert_class_shadowed_17_storage_err)
	);
	wire alert_class_shadowed_18_gated_we;
	assign alert_class_shadowed_18_gated_we = alert_class_shadowed_18_we & alert_regwen_18_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_18_re),
		.we(alert_class_shadowed_18_gated_we),
		.wd(alert_class_shadowed_18_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[906-:2]),
		.qs(alert_class_shadowed_18_qs),
		.err_update(alert_class_shadowed_18_update_err),
		.err_storage(alert_class_shadowed_18_storage_err)
	);
	wire alert_class_shadowed_19_gated_we;
	assign alert_class_shadowed_19_gated_we = alert_class_shadowed_19_we & alert_regwen_19_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_19_re),
		.we(alert_class_shadowed_19_gated_we),
		.wd(alert_class_shadowed_19_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[908-:2]),
		.qs(alert_class_shadowed_19_qs),
		.err_update(alert_class_shadowed_19_update_err),
		.err_storage(alert_class_shadowed_19_storage_err)
	);
	wire alert_class_shadowed_20_gated_we;
	assign alert_class_shadowed_20_gated_we = alert_class_shadowed_20_we & alert_regwen_20_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_20_re),
		.we(alert_class_shadowed_20_gated_we),
		.wd(alert_class_shadowed_20_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[910-:2]),
		.qs(alert_class_shadowed_20_qs),
		.err_update(alert_class_shadowed_20_update_err),
		.err_storage(alert_class_shadowed_20_storage_err)
	);
	wire alert_class_shadowed_21_gated_we;
	assign alert_class_shadowed_21_gated_we = alert_class_shadowed_21_we & alert_regwen_21_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_21_re),
		.we(alert_class_shadowed_21_gated_we),
		.wd(alert_class_shadowed_21_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[912-:2]),
		.qs(alert_class_shadowed_21_qs),
		.err_update(alert_class_shadowed_21_update_err),
		.err_storage(alert_class_shadowed_21_storage_err)
	);
	wire alert_class_shadowed_22_gated_we;
	assign alert_class_shadowed_22_gated_we = alert_class_shadowed_22_we & alert_regwen_22_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_22_re),
		.we(alert_class_shadowed_22_gated_we),
		.wd(alert_class_shadowed_22_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[914-:2]),
		.qs(alert_class_shadowed_22_qs),
		.err_update(alert_class_shadowed_22_update_err),
		.err_storage(alert_class_shadowed_22_storage_err)
	);
	wire alert_class_shadowed_23_gated_we;
	assign alert_class_shadowed_23_gated_we = alert_class_shadowed_23_we & alert_regwen_23_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_23_re),
		.we(alert_class_shadowed_23_gated_we),
		.wd(alert_class_shadowed_23_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[916-:2]),
		.qs(alert_class_shadowed_23_qs),
		.err_update(alert_class_shadowed_23_update_err),
		.err_storage(alert_class_shadowed_23_storage_err)
	);
	wire alert_class_shadowed_24_gated_we;
	assign alert_class_shadowed_24_gated_we = alert_class_shadowed_24_we & alert_regwen_24_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_24_re),
		.we(alert_class_shadowed_24_gated_we),
		.wd(alert_class_shadowed_24_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[918-:2]),
		.qs(alert_class_shadowed_24_qs),
		.err_update(alert_class_shadowed_24_update_err),
		.err_storage(alert_class_shadowed_24_storage_err)
	);
	wire alert_class_shadowed_25_gated_we;
	assign alert_class_shadowed_25_gated_we = alert_class_shadowed_25_we & alert_regwen_25_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_25_re),
		.we(alert_class_shadowed_25_gated_we),
		.wd(alert_class_shadowed_25_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[920-:2]),
		.qs(alert_class_shadowed_25_qs),
		.err_update(alert_class_shadowed_25_update_err),
		.err_storage(alert_class_shadowed_25_storage_err)
	);
	wire alert_class_shadowed_26_gated_we;
	assign alert_class_shadowed_26_gated_we = alert_class_shadowed_26_we & alert_regwen_26_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_26_re),
		.we(alert_class_shadowed_26_gated_we),
		.wd(alert_class_shadowed_26_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[922-:2]),
		.qs(alert_class_shadowed_26_qs),
		.err_update(alert_class_shadowed_26_update_err),
		.err_storage(alert_class_shadowed_26_storage_err)
	);
	wire alert_class_shadowed_27_gated_we;
	assign alert_class_shadowed_27_gated_we = alert_class_shadowed_27_we & alert_regwen_27_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_27_re),
		.we(alert_class_shadowed_27_gated_we),
		.wd(alert_class_shadowed_27_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[924-:2]),
		.qs(alert_class_shadowed_27_qs),
		.err_update(alert_class_shadowed_27_update_err),
		.err_storage(alert_class_shadowed_27_storage_err)
	);
	wire alert_class_shadowed_28_gated_we;
	assign alert_class_shadowed_28_gated_we = alert_class_shadowed_28_we & alert_regwen_28_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_28_re),
		.we(alert_class_shadowed_28_gated_we),
		.wd(alert_class_shadowed_28_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[926-:2]),
		.qs(alert_class_shadowed_28_qs),
		.err_update(alert_class_shadowed_28_update_err),
		.err_storage(alert_class_shadowed_28_storage_err)
	);
	wire alert_class_shadowed_29_gated_we;
	assign alert_class_shadowed_29_gated_we = alert_class_shadowed_29_we & alert_regwen_29_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_29_re),
		.we(alert_class_shadowed_29_gated_we),
		.wd(alert_class_shadowed_29_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[928-:2]),
		.qs(alert_class_shadowed_29_qs),
		.err_update(alert_class_shadowed_29_update_err),
		.err_storage(alert_class_shadowed_29_storage_err)
	);
	wire alert_class_shadowed_30_gated_we;
	assign alert_class_shadowed_30_gated_we = alert_class_shadowed_30_we & alert_regwen_30_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_30_re),
		.we(alert_class_shadowed_30_gated_we),
		.wd(alert_class_shadowed_30_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[930-:2]),
		.qs(alert_class_shadowed_30_qs),
		.err_update(alert_class_shadowed_30_update_err),
		.err_storage(alert_class_shadowed_30_storage_err)
	);
	wire alert_class_shadowed_31_gated_we;
	assign alert_class_shadowed_31_gated_we = alert_class_shadowed_31_we & alert_regwen_31_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_31_re),
		.we(alert_class_shadowed_31_gated_we),
		.wd(alert_class_shadowed_31_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[932-:2]),
		.qs(alert_class_shadowed_31_qs),
		.err_update(alert_class_shadowed_31_update_err),
		.err_storage(alert_class_shadowed_31_storage_err)
	);
	wire alert_class_shadowed_32_gated_we;
	assign alert_class_shadowed_32_gated_we = alert_class_shadowed_32_we & alert_regwen_32_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_32(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_32_re),
		.we(alert_class_shadowed_32_gated_we),
		.wd(alert_class_shadowed_32_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[934-:2]),
		.qs(alert_class_shadowed_32_qs),
		.err_update(alert_class_shadowed_32_update_err),
		.err_storage(alert_class_shadowed_32_storage_err)
	);
	wire alert_class_shadowed_33_gated_we;
	assign alert_class_shadowed_33_gated_we = alert_class_shadowed_33_we & alert_regwen_33_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_33(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_33_re),
		.we(alert_class_shadowed_33_gated_we),
		.wd(alert_class_shadowed_33_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[936-:2]),
		.qs(alert_class_shadowed_33_qs),
		.err_update(alert_class_shadowed_33_update_err),
		.err_storage(alert_class_shadowed_33_storage_err)
	);
	wire alert_class_shadowed_34_gated_we;
	assign alert_class_shadowed_34_gated_we = alert_class_shadowed_34_we & alert_regwen_34_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_34(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_34_re),
		.we(alert_class_shadowed_34_gated_we),
		.wd(alert_class_shadowed_34_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[938-:2]),
		.qs(alert_class_shadowed_34_qs),
		.err_update(alert_class_shadowed_34_update_err),
		.err_storage(alert_class_shadowed_34_storage_err)
	);
	wire alert_class_shadowed_35_gated_we;
	assign alert_class_shadowed_35_gated_we = alert_class_shadowed_35_we & alert_regwen_35_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_35(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_35_re),
		.we(alert_class_shadowed_35_gated_we),
		.wd(alert_class_shadowed_35_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[940-:2]),
		.qs(alert_class_shadowed_35_qs),
		.err_update(alert_class_shadowed_35_update_err),
		.err_storage(alert_class_shadowed_35_storage_err)
	);
	wire alert_class_shadowed_36_gated_we;
	assign alert_class_shadowed_36_gated_we = alert_class_shadowed_36_we & alert_regwen_36_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_36(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_36_re),
		.we(alert_class_shadowed_36_gated_we),
		.wd(alert_class_shadowed_36_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[942-:2]),
		.qs(alert_class_shadowed_36_qs),
		.err_update(alert_class_shadowed_36_update_err),
		.err_storage(alert_class_shadowed_36_storage_err)
	);
	wire alert_class_shadowed_37_gated_we;
	assign alert_class_shadowed_37_gated_we = alert_class_shadowed_37_we & alert_regwen_37_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_37(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_37_re),
		.we(alert_class_shadowed_37_gated_we),
		.wd(alert_class_shadowed_37_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[944-:2]),
		.qs(alert_class_shadowed_37_qs),
		.err_update(alert_class_shadowed_37_update_err),
		.err_storage(alert_class_shadowed_37_storage_err)
	);
	wire alert_class_shadowed_38_gated_we;
	assign alert_class_shadowed_38_gated_we = alert_class_shadowed_38_we & alert_regwen_38_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_38(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_38_re),
		.we(alert_class_shadowed_38_gated_we),
		.wd(alert_class_shadowed_38_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[946-:2]),
		.qs(alert_class_shadowed_38_qs),
		.err_update(alert_class_shadowed_38_update_err),
		.err_storage(alert_class_shadowed_38_storage_err)
	);
	wire alert_class_shadowed_39_gated_we;
	assign alert_class_shadowed_39_gated_we = alert_class_shadowed_39_we & alert_regwen_39_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_39(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_39_re),
		.we(alert_class_shadowed_39_gated_we),
		.wd(alert_class_shadowed_39_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[948-:2]),
		.qs(alert_class_shadowed_39_qs),
		.err_update(alert_class_shadowed_39_update_err),
		.err_storage(alert_class_shadowed_39_storage_err)
	);
	wire alert_class_shadowed_40_gated_we;
	assign alert_class_shadowed_40_gated_we = alert_class_shadowed_40_we & alert_regwen_40_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_40(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_40_re),
		.we(alert_class_shadowed_40_gated_we),
		.wd(alert_class_shadowed_40_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[950-:2]),
		.qs(alert_class_shadowed_40_qs),
		.err_update(alert_class_shadowed_40_update_err),
		.err_storage(alert_class_shadowed_40_storage_err)
	);
	wire alert_class_shadowed_41_gated_we;
	assign alert_class_shadowed_41_gated_we = alert_class_shadowed_41_we & alert_regwen_41_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_41(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_41_re),
		.we(alert_class_shadowed_41_gated_we),
		.wd(alert_class_shadowed_41_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[952-:2]),
		.qs(alert_class_shadowed_41_qs),
		.err_update(alert_class_shadowed_41_update_err),
		.err_storage(alert_class_shadowed_41_storage_err)
	);
	wire alert_class_shadowed_42_gated_we;
	assign alert_class_shadowed_42_gated_we = alert_class_shadowed_42_we & alert_regwen_42_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_42(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_42_re),
		.we(alert_class_shadowed_42_gated_we),
		.wd(alert_class_shadowed_42_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[954-:2]),
		.qs(alert_class_shadowed_42_qs),
		.err_update(alert_class_shadowed_42_update_err),
		.err_storage(alert_class_shadowed_42_storage_err)
	);
	wire alert_class_shadowed_43_gated_we;
	assign alert_class_shadowed_43_gated_we = alert_class_shadowed_43_we & alert_regwen_43_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_43(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_43_re),
		.we(alert_class_shadowed_43_gated_we),
		.wd(alert_class_shadowed_43_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[956-:2]),
		.qs(alert_class_shadowed_43_qs),
		.err_update(alert_class_shadowed_43_update_err),
		.err_storage(alert_class_shadowed_43_storage_err)
	);
	wire alert_class_shadowed_44_gated_we;
	assign alert_class_shadowed_44_gated_we = alert_class_shadowed_44_we & alert_regwen_44_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_44(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_44_re),
		.we(alert_class_shadowed_44_gated_we),
		.wd(alert_class_shadowed_44_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[958-:2]),
		.qs(alert_class_shadowed_44_qs),
		.err_update(alert_class_shadowed_44_update_err),
		.err_storage(alert_class_shadowed_44_storage_err)
	);
	wire alert_class_shadowed_45_gated_we;
	assign alert_class_shadowed_45_gated_we = alert_class_shadowed_45_we & alert_regwen_45_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_45(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_45_re),
		.we(alert_class_shadowed_45_gated_we),
		.wd(alert_class_shadowed_45_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[960-:2]),
		.qs(alert_class_shadowed_45_qs),
		.err_update(alert_class_shadowed_45_update_err),
		.err_storage(alert_class_shadowed_45_storage_err)
	);
	wire alert_class_shadowed_46_gated_we;
	assign alert_class_shadowed_46_gated_we = alert_class_shadowed_46_we & alert_regwen_46_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_46(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_46_re),
		.we(alert_class_shadowed_46_gated_we),
		.wd(alert_class_shadowed_46_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[962-:2]),
		.qs(alert_class_shadowed_46_qs),
		.err_update(alert_class_shadowed_46_update_err),
		.err_storage(alert_class_shadowed_46_storage_err)
	);
	wire alert_class_shadowed_47_gated_we;
	assign alert_class_shadowed_47_gated_we = alert_class_shadowed_47_we & alert_regwen_47_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_47(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_47_re),
		.we(alert_class_shadowed_47_gated_we),
		.wd(alert_class_shadowed_47_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[964-:2]),
		.qs(alert_class_shadowed_47_qs),
		.err_update(alert_class_shadowed_47_update_err),
		.err_storage(alert_class_shadowed_47_storage_err)
	);
	wire alert_class_shadowed_48_gated_we;
	assign alert_class_shadowed_48_gated_we = alert_class_shadowed_48_we & alert_regwen_48_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_48(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_48_re),
		.we(alert_class_shadowed_48_gated_we),
		.wd(alert_class_shadowed_48_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[966-:2]),
		.qs(alert_class_shadowed_48_qs),
		.err_update(alert_class_shadowed_48_update_err),
		.err_storage(alert_class_shadowed_48_storage_err)
	);
	wire alert_class_shadowed_49_gated_we;
	assign alert_class_shadowed_49_gated_we = alert_class_shadowed_49_we & alert_regwen_49_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_49(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_49_re),
		.we(alert_class_shadowed_49_gated_we),
		.wd(alert_class_shadowed_49_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[968-:2]),
		.qs(alert_class_shadowed_49_qs),
		.err_update(alert_class_shadowed_49_update_err),
		.err_storage(alert_class_shadowed_49_storage_err)
	);
	wire alert_class_shadowed_50_gated_we;
	assign alert_class_shadowed_50_gated_we = alert_class_shadowed_50_we & alert_regwen_50_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_50(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_50_re),
		.we(alert_class_shadowed_50_gated_we),
		.wd(alert_class_shadowed_50_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[970-:2]),
		.qs(alert_class_shadowed_50_qs),
		.err_update(alert_class_shadowed_50_update_err),
		.err_storage(alert_class_shadowed_50_storage_err)
	);
	wire alert_class_shadowed_51_gated_we;
	assign alert_class_shadowed_51_gated_we = alert_class_shadowed_51_we & alert_regwen_51_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_51(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_51_re),
		.we(alert_class_shadowed_51_gated_we),
		.wd(alert_class_shadowed_51_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[972-:2]),
		.qs(alert_class_shadowed_51_qs),
		.err_update(alert_class_shadowed_51_update_err),
		.err_storage(alert_class_shadowed_51_storage_err)
	);
	wire alert_class_shadowed_52_gated_we;
	assign alert_class_shadowed_52_gated_we = alert_class_shadowed_52_we & alert_regwen_52_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_52(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_52_re),
		.we(alert_class_shadowed_52_gated_we),
		.wd(alert_class_shadowed_52_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[974-:2]),
		.qs(alert_class_shadowed_52_qs),
		.err_update(alert_class_shadowed_52_update_err),
		.err_storage(alert_class_shadowed_52_storage_err)
	);
	wire alert_class_shadowed_53_gated_we;
	assign alert_class_shadowed_53_gated_we = alert_class_shadowed_53_we & alert_regwen_53_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_53(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_53_re),
		.we(alert_class_shadowed_53_gated_we),
		.wd(alert_class_shadowed_53_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[976-:2]),
		.qs(alert_class_shadowed_53_qs),
		.err_update(alert_class_shadowed_53_update_err),
		.err_storage(alert_class_shadowed_53_storage_err)
	);
	wire alert_class_shadowed_54_gated_we;
	assign alert_class_shadowed_54_gated_we = alert_class_shadowed_54_we & alert_regwen_54_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_54(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_54_re),
		.we(alert_class_shadowed_54_gated_we),
		.wd(alert_class_shadowed_54_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[978-:2]),
		.qs(alert_class_shadowed_54_qs),
		.err_update(alert_class_shadowed_54_update_err),
		.err_storage(alert_class_shadowed_54_storage_err)
	);
	wire alert_class_shadowed_55_gated_we;
	assign alert_class_shadowed_55_gated_we = alert_class_shadowed_55_we & alert_regwen_55_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_55(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_55_re),
		.we(alert_class_shadowed_55_gated_we),
		.wd(alert_class_shadowed_55_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[980-:2]),
		.qs(alert_class_shadowed_55_qs),
		.err_update(alert_class_shadowed_55_update_err),
		.err_storage(alert_class_shadowed_55_storage_err)
	);
	wire alert_class_shadowed_56_gated_we;
	assign alert_class_shadowed_56_gated_we = alert_class_shadowed_56_we & alert_regwen_56_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_56(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_56_re),
		.we(alert_class_shadowed_56_gated_we),
		.wd(alert_class_shadowed_56_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[982-:2]),
		.qs(alert_class_shadowed_56_qs),
		.err_update(alert_class_shadowed_56_update_err),
		.err_storage(alert_class_shadowed_56_storage_err)
	);
	wire alert_class_shadowed_57_gated_we;
	assign alert_class_shadowed_57_gated_we = alert_class_shadowed_57_we & alert_regwen_57_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_57(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_57_re),
		.we(alert_class_shadowed_57_gated_we),
		.wd(alert_class_shadowed_57_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[984-:2]),
		.qs(alert_class_shadowed_57_qs),
		.err_update(alert_class_shadowed_57_update_err),
		.err_storage(alert_class_shadowed_57_storage_err)
	);
	wire alert_class_shadowed_58_gated_we;
	assign alert_class_shadowed_58_gated_we = alert_class_shadowed_58_we & alert_regwen_58_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_58(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_58_re),
		.we(alert_class_shadowed_58_gated_we),
		.wd(alert_class_shadowed_58_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[986-:2]),
		.qs(alert_class_shadowed_58_qs),
		.err_update(alert_class_shadowed_58_update_err),
		.err_storage(alert_class_shadowed_58_storage_err)
	);
	wire alert_class_shadowed_59_gated_we;
	assign alert_class_shadowed_59_gated_we = alert_class_shadowed_59_we & alert_regwen_59_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_59(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_59_re),
		.we(alert_class_shadowed_59_gated_we),
		.wd(alert_class_shadowed_59_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[988-:2]),
		.qs(alert_class_shadowed_59_qs),
		.err_update(alert_class_shadowed_59_update_err),
		.err_storage(alert_class_shadowed_59_storage_err)
	);
	wire alert_class_shadowed_60_gated_we;
	assign alert_class_shadowed_60_gated_we = alert_class_shadowed_60_we & alert_regwen_60_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_60(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_60_re),
		.we(alert_class_shadowed_60_gated_we),
		.wd(alert_class_shadowed_60_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[990-:2]),
		.qs(alert_class_shadowed_60_qs),
		.err_update(alert_class_shadowed_60_update_err),
		.err_storage(alert_class_shadowed_60_storage_err)
	);
	wire alert_class_shadowed_61_gated_we;
	assign alert_class_shadowed_61_gated_we = alert_class_shadowed_61_we & alert_regwen_61_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_61(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_61_re),
		.we(alert_class_shadowed_61_gated_we),
		.wd(alert_class_shadowed_61_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[992-:2]),
		.qs(alert_class_shadowed_61_qs),
		.err_update(alert_class_shadowed_61_update_err),
		.err_storage(alert_class_shadowed_61_storage_err)
	);
	wire alert_class_shadowed_62_gated_we;
	assign alert_class_shadowed_62_gated_we = alert_class_shadowed_62_we & alert_regwen_62_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_62(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_62_re),
		.we(alert_class_shadowed_62_gated_we),
		.wd(alert_class_shadowed_62_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[994-:2]),
		.qs(alert_class_shadowed_62_qs),
		.err_update(alert_class_shadowed_62_update_err),
		.err_storage(alert_class_shadowed_62_storage_err)
	);
	wire alert_class_shadowed_63_gated_we;
	assign alert_class_shadowed_63_gated_we = alert_class_shadowed_63_we & alert_regwen_63_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_63(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_63_re),
		.we(alert_class_shadowed_63_gated_we),
		.wd(alert_class_shadowed_63_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[996-:2]),
		.qs(alert_class_shadowed_63_qs),
		.err_update(alert_class_shadowed_63_update_err),
		.err_storage(alert_class_shadowed_63_storage_err)
	);
	wire alert_class_shadowed_64_gated_we;
	assign alert_class_shadowed_64_gated_we = alert_class_shadowed_64_we & alert_regwen_64_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_alert_class_shadowed_64(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(alert_class_shadowed_64_re),
		.we(alert_class_shadowed_64_gated_we),
		.wd(alert_class_shadowed_64_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[998-:2]),
		.qs(alert_class_shadowed_64_qs),
		.err_update(alert_class_shadowed_64_update_err),
		.err_storage(alert_class_shadowed_64_storage_err)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_0_we),
		.wd(alert_cause_0_wd),
		.de(hw2reg[226]),
		.d(hw2reg[227]),
		.q(reg2hw[804]),
		.qs(alert_cause_0_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_1_we),
		.wd(alert_cause_1_wd),
		.de(hw2reg[228]),
		.d(hw2reg[229]),
		.q(reg2hw[805]),
		.qs(alert_cause_1_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_2_we),
		.wd(alert_cause_2_wd),
		.de(hw2reg[230]),
		.d(hw2reg[231]),
		.q(reg2hw[806]),
		.qs(alert_cause_2_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_3_we),
		.wd(alert_cause_3_wd),
		.de(hw2reg[232]),
		.d(hw2reg[233]),
		.q(reg2hw[807]),
		.qs(alert_cause_3_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_4_we),
		.wd(alert_cause_4_wd),
		.de(hw2reg[234]),
		.d(hw2reg[235]),
		.q(reg2hw[808]),
		.qs(alert_cause_4_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_5_we),
		.wd(alert_cause_5_wd),
		.de(hw2reg[236]),
		.d(hw2reg[237]),
		.q(reg2hw[809]),
		.qs(alert_cause_5_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_6_we),
		.wd(alert_cause_6_wd),
		.de(hw2reg[238]),
		.d(hw2reg[239]),
		.q(reg2hw[810]),
		.qs(alert_cause_6_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_7(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_7_we),
		.wd(alert_cause_7_wd),
		.de(hw2reg[240]),
		.d(hw2reg[241]),
		.q(reg2hw[811]),
		.qs(alert_cause_7_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_8(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_8_we),
		.wd(alert_cause_8_wd),
		.de(hw2reg[242]),
		.d(hw2reg[243]),
		.q(reg2hw[812]),
		.qs(alert_cause_8_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_9(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_9_we),
		.wd(alert_cause_9_wd),
		.de(hw2reg[244]),
		.d(hw2reg[245]),
		.q(reg2hw[813]),
		.qs(alert_cause_9_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_10(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_10_we),
		.wd(alert_cause_10_wd),
		.de(hw2reg[246]),
		.d(hw2reg[247]),
		.q(reg2hw[814]),
		.qs(alert_cause_10_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_11(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_11_we),
		.wd(alert_cause_11_wd),
		.de(hw2reg[248]),
		.d(hw2reg[249]),
		.q(reg2hw[815]),
		.qs(alert_cause_11_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_12(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_12_we),
		.wd(alert_cause_12_wd),
		.de(hw2reg[250]),
		.d(hw2reg[251]),
		.q(reg2hw[816]),
		.qs(alert_cause_12_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_13(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_13_we),
		.wd(alert_cause_13_wd),
		.de(hw2reg[252]),
		.d(hw2reg[253]),
		.q(reg2hw[817]),
		.qs(alert_cause_13_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_14(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_14_we),
		.wd(alert_cause_14_wd),
		.de(hw2reg[254]),
		.d(hw2reg[255]),
		.q(reg2hw[818]),
		.qs(alert_cause_14_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_15(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_15_we),
		.wd(alert_cause_15_wd),
		.de(hw2reg[256]),
		.d(hw2reg[257]),
		.q(reg2hw[819]),
		.qs(alert_cause_15_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_16(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_16_we),
		.wd(alert_cause_16_wd),
		.de(hw2reg[258]),
		.d(hw2reg[259]),
		.q(reg2hw[820]),
		.qs(alert_cause_16_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_17(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_17_we),
		.wd(alert_cause_17_wd),
		.de(hw2reg[260]),
		.d(hw2reg[261]),
		.q(reg2hw[821]),
		.qs(alert_cause_17_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_18(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_18_we),
		.wd(alert_cause_18_wd),
		.de(hw2reg[262]),
		.d(hw2reg[263]),
		.q(reg2hw[822]),
		.qs(alert_cause_18_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_19(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_19_we),
		.wd(alert_cause_19_wd),
		.de(hw2reg[264]),
		.d(hw2reg[265]),
		.q(reg2hw[823]),
		.qs(alert_cause_19_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_20(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_20_we),
		.wd(alert_cause_20_wd),
		.de(hw2reg[266]),
		.d(hw2reg[267]),
		.q(reg2hw[824]),
		.qs(alert_cause_20_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_21(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_21_we),
		.wd(alert_cause_21_wd),
		.de(hw2reg[268]),
		.d(hw2reg[269]),
		.q(reg2hw[825]),
		.qs(alert_cause_21_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_22(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_22_we),
		.wd(alert_cause_22_wd),
		.de(hw2reg[270]),
		.d(hw2reg[271]),
		.q(reg2hw[826]),
		.qs(alert_cause_22_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_23(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_23_we),
		.wd(alert_cause_23_wd),
		.de(hw2reg[272]),
		.d(hw2reg[273]),
		.q(reg2hw[827]),
		.qs(alert_cause_23_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_24(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_24_we),
		.wd(alert_cause_24_wd),
		.de(hw2reg[274]),
		.d(hw2reg[275]),
		.q(reg2hw[828]),
		.qs(alert_cause_24_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_25(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_25_we),
		.wd(alert_cause_25_wd),
		.de(hw2reg[276]),
		.d(hw2reg[277]),
		.q(reg2hw[829]),
		.qs(alert_cause_25_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_26(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_26_we),
		.wd(alert_cause_26_wd),
		.de(hw2reg[278]),
		.d(hw2reg[279]),
		.q(reg2hw[830]),
		.qs(alert_cause_26_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_27(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_27_we),
		.wd(alert_cause_27_wd),
		.de(hw2reg[280]),
		.d(hw2reg[281]),
		.q(reg2hw[831]),
		.qs(alert_cause_27_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_28(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_28_we),
		.wd(alert_cause_28_wd),
		.de(hw2reg[282]),
		.d(hw2reg[283]),
		.q(reg2hw[832]),
		.qs(alert_cause_28_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_29(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_29_we),
		.wd(alert_cause_29_wd),
		.de(hw2reg[284]),
		.d(hw2reg[285]),
		.q(reg2hw[833]),
		.qs(alert_cause_29_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_30(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_30_we),
		.wd(alert_cause_30_wd),
		.de(hw2reg[286]),
		.d(hw2reg[287]),
		.q(reg2hw[834]),
		.qs(alert_cause_30_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_31(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_31_we),
		.wd(alert_cause_31_wd),
		.de(hw2reg[288]),
		.d(hw2reg[289]),
		.q(reg2hw[835]),
		.qs(alert_cause_31_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_32(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_32_we),
		.wd(alert_cause_32_wd),
		.de(hw2reg[290]),
		.d(hw2reg[291]),
		.q(reg2hw[836]),
		.qs(alert_cause_32_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_33(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_33_we),
		.wd(alert_cause_33_wd),
		.de(hw2reg[292]),
		.d(hw2reg[293]),
		.q(reg2hw[837]),
		.qs(alert_cause_33_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_34(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_34_we),
		.wd(alert_cause_34_wd),
		.de(hw2reg[294]),
		.d(hw2reg[295]),
		.q(reg2hw[838]),
		.qs(alert_cause_34_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_35(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_35_we),
		.wd(alert_cause_35_wd),
		.de(hw2reg[296]),
		.d(hw2reg[297]),
		.q(reg2hw[839]),
		.qs(alert_cause_35_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_36(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_36_we),
		.wd(alert_cause_36_wd),
		.de(hw2reg[298]),
		.d(hw2reg[299]),
		.q(reg2hw[840]),
		.qs(alert_cause_36_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_37(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_37_we),
		.wd(alert_cause_37_wd),
		.de(hw2reg[300]),
		.d(hw2reg[301]),
		.q(reg2hw[841]),
		.qs(alert_cause_37_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_38(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_38_we),
		.wd(alert_cause_38_wd),
		.de(hw2reg[302]),
		.d(hw2reg[303]),
		.q(reg2hw[842]),
		.qs(alert_cause_38_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_39(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_39_we),
		.wd(alert_cause_39_wd),
		.de(hw2reg[304]),
		.d(hw2reg[305]),
		.q(reg2hw[843]),
		.qs(alert_cause_39_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_40(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_40_we),
		.wd(alert_cause_40_wd),
		.de(hw2reg[306]),
		.d(hw2reg[307]),
		.q(reg2hw[844]),
		.qs(alert_cause_40_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_41(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_41_we),
		.wd(alert_cause_41_wd),
		.de(hw2reg[308]),
		.d(hw2reg[309]),
		.q(reg2hw[845]),
		.qs(alert_cause_41_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_42(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_42_we),
		.wd(alert_cause_42_wd),
		.de(hw2reg[310]),
		.d(hw2reg[311]),
		.q(reg2hw[846]),
		.qs(alert_cause_42_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_43(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_43_we),
		.wd(alert_cause_43_wd),
		.de(hw2reg[312]),
		.d(hw2reg[313]),
		.q(reg2hw[847]),
		.qs(alert_cause_43_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_44(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_44_we),
		.wd(alert_cause_44_wd),
		.de(hw2reg[314]),
		.d(hw2reg[315]),
		.q(reg2hw[848]),
		.qs(alert_cause_44_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_45(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_45_we),
		.wd(alert_cause_45_wd),
		.de(hw2reg[316]),
		.d(hw2reg[317]),
		.q(reg2hw[849]),
		.qs(alert_cause_45_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_46(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_46_we),
		.wd(alert_cause_46_wd),
		.de(hw2reg[318]),
		.d(hw2reg[319]),
		.q(reg2hw[850]),
		.qs(alert_cause_46_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_47(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_47_we),
		.wd(alert_cause_47_wd),
		.de(hw2reg[320]),
		.d(hw2reg[321]),
		.q(reg2hw[851]),
		.qs(alert_cause_47_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_48(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_48_we),
		.wd(alert_cause_48_wd),
		.de(hw2reg[322]),
		.d(hw2reg[323]),
		.q(reg2hw[852]),
		.qs(alert_cause_48_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_49(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_49_we),
		.wd(alert_cause_49_wd),
		.de(hw2reg[324]),
		.d(hw2reg[325]),
		.q(reg2hw[853]),
		.qs(alert_cause_49_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_50(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_50_we),
		.wd(alert_cause_50_wd),
		.de(hw2reg[326]),
		.d(hw2reg[327]),
		.q(reg2hw[854]),
		.qs(alert_cause_50_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_51(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_51_we),
		.wd(alert_cause_51_wd),
		.de(hw2reg[328]),
		.d(hw2reg[329]),
		.q(reg2hw[855]),
		.qs(alert_cause_51_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_52(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_52_we),
		.wd(alert_cause_52_wd),
		.de(hw2reg[330]),
		.d(hw2reg[331]),
		.q(reg2hw[856]),
		.qs(alert_cause_52_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_53(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_53_we),
		.wd(alert_cause_53_wd),
		.de(hw2reg[332]),
		.d(hw2reg[333]),
		.q(reg2hw[857]),
		.qs(alert_cause_53_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_54(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_54_we),
		.wd(alert_cause_54_wd),
		.de(hw2reg[334]),
		.d(hw2reg[335]),
		.q(reg2hw[858]),
		.qs(alert_cause_54_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_55(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_55_we),
		.wd(alert_cause_55_wd),
		.de(hw2reg[336]),
		.d(hw2reg[337]),
		.q(reg2hw[859]),
		.qs(alert_cause_55_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_56(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_56_we),
		.wd(alert_cause_56_wd),
		.de(hw2reg[338]),
		.d(hw2reg[339]),
		.q(reg2hw[860]),
		.qs(alert_cause_56_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_57(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_57_we),
		.wd(alert_cause_57_wd),
		.de(hw2reg[340]),
		.d(hw2reg[341]),
		.q(reg2hw[861]),
		.qs(alert_cause_57_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_58(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_58_we),
		.wd(alert_cause_58_wd),
		.de(hw2reg[342]),
		.d(hw2reg[343]),
		.q(reg2hw[862]),
		.qs(alert_cause_58_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_59(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_59_we),
		.wd(alert_cause_59_wd),
		.de(hw2reg[344]),
		.d(hw2reg[345]),
		.q(reg2hw[863]),
		.qs(alert_cause_59_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_60(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_60_we),
		.wd(alert_cause_60_wd),
		.de(hw2reg[346]),
		.d(hw2reg[347]),
		.q(reg2hw[864]),
		.qs(alert_cause_60_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_61(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_61_we),
		.wd(alert_cause_61_wd),
		.de(hw2reg[348]),
		.d(hw2reg[349]),
		.q(reg2hw[865]),
		.qs(alert_cause_61_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_62(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_62_we),
		.wd(alert_cause_62_wd),
		.de(hw2reg[350]),
		.d(hw2reg[351]),
		.q(reg2hw[866]),
		.qs(alert_cause_62_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_63(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_63_we),
		.wd(alert_cause_63_wd),
		.de(hw2reg[352]),
		.d(hw2reg[353]),
		.q(reg2hw[867]),
		.qs(alert_cause_63_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_alert_cause_64(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(alert_cause_64_we),
		.wd(alert_cause_64_wd),
		.de(hw2reg[354]),
		.d(hw2reg[355]),
		.q(reg2hw[868]),
		.qs(alert_cause_64_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_loc_alert_regwen_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(loc_alert_regwen_0_we),
		.wd(loc_alert_regwen_0_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(loc_alert_regwen_0_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_loc_alert_regwen_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(loc_alert_regwen_1_we),
		.wd(loc_alert_regwen_1_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(loc_alert_regwen_1_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_loc_alert_regwen_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(loc_alert_regwen_2_we),
		.wd(loc_alert_regwen_2_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(loc_alert_regwen_2_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_loc_alert_regwen_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(loc_alert_regwen_3_we),
		.wd(loc_alert_regwen_3_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(loc_alert_regwen_3_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_loc_alert_regwen_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(loc_alert_regwen_4_we),
		.wd(loc_alert_regwen_4_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(loc_alert_regwen_4_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_loc_alert_regwen_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(loc_alert_regwen_5_we),
		.wd(loc_alert_regwen_5_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(loc_alert_regwen_5_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_loc_alert_regwen_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(loc_alert_regwen_6_we),
		.wd(loc_alert_regwen_6_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(loc_alert_regwen_6_qs)
	);
	wire loc_alert_en_shadowed_0_gated_we;
	assign loc_alert_en_shadowed_0_gated_we = loc_alert_en_shadowed_0_we & loc_alert_regwen_0_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_loc_alert_en_shadowed_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(loc_alert_en_shadowed_0_re),
		.we(loc_alert_en_shadowed_0_gated_we),
		.wd(loc_alert_en_shadowed_0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[797]),
		.qs(loc_alert_en_shadowed_0_qs),
		.err_update(loc_alert_en_shadowed_0_update_err),
		.err_storage(loc_alert_en_shadowed_0_storage_err)
	);
	wire loc_alert_en_shadowed_1_gated_we;
	assign loc_alert_en_shadowed_1_gated_we = loc_alert_en_shadowed_1_we & loc_alert_regwen_1_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_loc_alert_en_shadowed_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(loc_alert_en_shadowed_1_re),
		.we(loc_alert_en_shadowed_1_gated_we),
		.wd(loc_alert_en_shadowed_1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[798]),
		.qs(loc_alert_en_shadowed_1_qs),
		.err_update(loc_alert_en_shadowed_1_update_err),
		.err_storage(loc_alert_en_shadowed_1_storage_err)
	);
	wire loc_alert_en_shadowed_2_gated_we;
	assign loc_alert_en_shadowed_2_gated_we = loc_alert_en_shadowed_2_we & loc_alert_regwen_2_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_loc_alert_en_shadowed_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(loc_alert_en_shadowed_2_re),
		.we(loc_alert_en_shadowed_2_gated_we),
		.wd(loc_alert_en_shadowed_2_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[799]),
		.qs(loc_alert_en_shadowed_2_qs),
		.err_update(loc_alert_en_shadowed_2_update_err),
		.err_storage(loc_alert_en_shadowed_2_storage_err)
	);
	wire loc_alert_en_shadowed_3_gated_we;
	assign loc_alert_en_shadowed_3_gated_we = loc_alert_en_shadowed_3_we & loc_alert_regwen_3_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_loc_alert_en_shadowed_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(loc_alert_en_shadowed_3_re),
		.we(loc_alert_en_shadowed_3_gated_we),
		.wd(loc_alert_en_shadowed_3_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[800]),
		.qs(loc_alert_en_shadowed_3_qs),
		.err_update(loc_alert_en_shadowed_3_update_err),
		.err_storage(loc_alert_en_shadowed_3_storage_err)
	);
	wire loc_alert_en_shadowed_4_gated_we;
	assign loc_alert_en_shadowed_4_gated_we = loc_alert_en_shadowed_4_we & loc_alert_regwen_4_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_loc_alert_en_shadowed_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(loc_alert_en_shadowed_4_re),
		.we(loc_alert_en_shadowed_4_gated_we),
		.wd(loc_alert_en_shadowed_4_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[801]),
		.qs(loc_alert_en_shadowed_4_qs),
		.err_update(loc_alert_en_shadowed_4_update_err),
		.err_storage(loc_alert_en_shadowed_4_storage_err)
	);
	wire loc_alert_en_shadowed_5_gated_we;
	assign loc_alert_en_shadowed_5_gated_we = loc_alert_en_shadowed_5_we & loc_alert_regwen_5_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_loc_alert_en_shadowed_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(loc_alert_en_shadowed_5_re),
		.we(loc_alert_en_shadowed_5_gated_we),
		.wd(loc_alert_en_shadowed_5_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[802]),
		.qs(loc_alert_en_shadowed_5_qs),
		.err_update(loc_alert_en_shadowed_5_update_err),
		.err_storage(loc_alert_en_shadowed_5_storage_err)
	);
	wire loc_alert_en_shadowed_6_gated_we;
	assign loc_alert_en_shadowed_6_gated_we = loc_alert_en_shadowed_6_we & loc_alert_regwen_6_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_loc_alert_en_shadowed_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(loc_alert_en_shadowed_6_re),
		.we(loc_alert_en_shadowed_6_gated_we),
		.wd(loc_alert_en_shadowed_6_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[803]),
		.qs(loc_alert_en_shadowed_6_qs),
		.err_update(loc_alert_en_shadowed_6_update_err),
		.err_storage(loc_alert_en_shadowed_6_storage_err)
	);
	wire loc_alert_class_shadowed_0_gated_we;
	assign loc_alert_class_shadowed_0_gated_we = loc_alert_class_shadowed_0_we & loc_alert_regwen_0_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_loc_alert_class_shadowed_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(loc_alert_class_shadowed_0_re),
		.we(loc_alert_class_shadowed_0_gated_we),
		.wd(loc_alert_class_shadowed_0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[784-:2]),
		.qs(loc_alert_class_shadowed_0_qs),
		.err_update(loc_alert_class_shadowed_0_update_err),
		.err_storage(loc_alert_class_shadowed_0_storage_err)
	);
	wire loc_alert_class_shadowed_1_gated_we;
	assign loc_alert_class_shadowed_1_gated_we = loc_alert_class_shadowed_1_we & loc_alert_regwen_1_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_loc_alert_class_shadowed_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(loc_alert_class_shadowed_1_re),
		.we(loc_alert_class_shadowed_1_gated_we),
		.wd(loc_alert_class_shadowed_1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[786-:2]),
		.qs(loc_alert_class_shadowed_1_qs),
		.err_update(loc_alert_class_shadowed_1_update_err),
		.err_storage(loc_alert_class_shadowed_1_storage_err)
	);
	wire loc_alert_class_shadowed_2_gated_we;
	assign loc_alert_class_shadowed_2_gated_we = loc_alert_class_shadowed_2_we & loc_alert_regwen_2_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_loc_alert_class_shadowed_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(loc_alert_class_shadowed_2_re),
		.we(loc_alert_class_shadowed_2_gated_we),
		.wd(loc_alert_class_shadowed_2_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[788-:2]),
		.qs(loc_alert_class_shadowed_2_qs),
		.err_update(loc_alert_class_shadowed_2_update_err),
		.err_storage(loc_alert_class_shadowed_2_storage_err)
	);
	wire loc_alert_class_shadowed_3_gated_we;
	assign loc_alert_class_shadowed_3_gated_we = loc_alert_class_shadowed_3_we & loc_alert_regwen_3_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_loc_alert_class_shadowed_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(loc_alert_class_shadowed_3_re),
		.we(loc_alert_class_shadowed_3_gated_we),
		.wd(loc_alert_class_shadowed_3_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[790-:2]),
		.qs(loc_alert_class_shadowed_3_qs),
		.err_update(loc_alert_class_shadowed_3_update_err),
		.err_storage(loc_alert_class_shadowed_3_storage_err)
	);
	wire loc_alert_class_shadowed_4_gated_we;
	assign loc_alert_class_shadowed_4_gated_we = loc_alert_class_shadowed_4_we & loc_alert_regwen_4_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_loc_alert_class_shadowed_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(loc_alert_class_shadowed_4_re),
		.we(loc_alert_class_shadowed_4_gated_we),
		.wd(loc_alert_class_shadowed_4_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[792-:2]),
		.qs(loc_alert_class_shadowed_4_qs),
		.err_update(loc_alert_class_shadowed_4_update_err),
		.err_storage(loc_alert_class_shadowed_4_storage_err)
	);
	wire loc_alert_class_shadowed_5_gated_we;
	assign loc_alert_class_shadowed_5_gated_we = loc_alert_class_shadowed_5_we & loc_alert_regwen_5_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_loc_alert_class_shadowed_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(loc_alert_class_shadowed_5_re),
		.we(loc_alert_class_shadowed_5_gated_we),
		.wd(loc_alert_class_shadowed_5_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[794-:2]),
		.qs(loc_alert_class_shadowed_5_qs),
		.err_update(loc_alert_class_shadowed_5_update_err),
		.err_storage(loc_alert_class_shadowed_5_storage_err)
	);
	wire loc_alert_class_shadowed_6_gated_we;
	assign loc_alert_class_shadowed_6_gated_we = loc_alert_class_shadowed_6_we & loc_alert_regwen_6_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_loc_alert_class_shadowed_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(loc_alert_class_shadowed_6_re),
		.we(loc_alert_class_shadowed_6_gated_we),
		.wd(loc_alert_class_shadowed_6_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[796-:2]),
		.qs(loc_alert_class_shadowed_6_qs),
		.err_update(loc_alert_class_shadowed_6_update_err),
		.err_storage(loc_alert_class_shadowed_6_storage_err)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_loc_alert_cause_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(loc_alert_cause_0_we),
		.wd(loc_alert_cause_0_wd),
		.de(hw2reg[212]),
		.d(hw2reg[213]),
		.q(reg2hw[776]),
		.qs(loc_alert_cause_0_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_loc_alert_cause_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(loc_alert_cause_1_we),
		.wd(loc_alert_cause_1_wd),
		.de(hw2reg[214]),
		.d(hw2reg[215]),
		.q(reg2hw[777]),
		.qs(loc_alert_cause_1_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_loc_alert_cause_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(loc_alert_cause_2_we),
		.wd(loc_alert_cause_2_wd),
		.de(hw2reg[216]),
		.d(hw2reg[217]),
		.q(reg2hw[778]),
		.qs(loc_alert_cause_2_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_loc_alert_cause_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(loc_alert_cause_3_we),
		.wd(loc_alert_cause_3_wd),
		.de(hw2reg[218]),
		.d(hw2reg[219]),
		.q(reg2hw[779]),
		.qs(loc_alert_cause_3_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_loc_alert_cause_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(loc_alert_cause_4_we),
		.wd(loc_alert_cause_4_wd),
		.de(hw2reg[220]),
		.d(hw2reg[221]),
		.q(reg2hw[780]),
		.qs(loc_alert_cause_4_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_loc_alert_cause_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(loc_alert_cause_5_we),
		.wd(loc_alert_cause_5_wd),
		.de(hw2reg[222]),
		.d(hw2reg[223]),
		.q(reg2hw[781]),
		.qs(loc_alert_cause_5_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_loc_alert_cause_6(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(loc_alert_cause_6_we),
		.wd(loc_alert_cause_6_wd),
		.de(hw2reg[224]),
		.d(hw2reg[225]),
		.q(reg2hw[782]),
		.qs(loc_alert_cause_6_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_classa_regwen(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(classa_regwen_we),
		.wd(classa_regwen_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(classa_regwen_qs)
	);
	wire classa_ctrl_shadowed_gated_we;
	assign classa_ctrl_shadowed_gated_we = classa_ctrl_shadowed_we & classa_regwen_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_classa_ctrl_shadowed_en(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_ctrl_shadowed_re),
		.we(classa_ctrl_shadowed_gated_we),
		.wd(classa_ctrl_shadowed_en_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[775]),
		.qs(classa_ctrl_shadowed_en_qs),
		.err_update(classa_ctrl_shadowed_en_update_err),
		.err_storage(classa_ctrl_shadowed_en_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_classa_ctrl_shadowed_lock(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_ctrl_shadowed_re),
		.we(classa_ctrl_shadowed_gated_we),
		.wd(classa_ctrl_shadowed_lock_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[774]),
		.qs(classa_ctrl_shadowed_lock_qs),
		.err_update(classa_ctrl_shadowed_lock_update_err),
		.err_storage(classa_ctrl_shadowed_lock_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_classa_ctrl_shadowed_en_e0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_ctrl_shadowed_re),
		.we(classa_ctrl_shadowed_gated_we),
		.wd(classa_ctrl_shadowed_en_e0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[773]),
		.qs(classa_ctrl_shadowed_en_e0_qs),
		.err_update(classa_ctrl_shadowed_en_e0_update_err),
		.err_storage(classa_ctrl_shadowed_en_e0_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_classa_ctrl_shadowed_en_e1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_ctrl_shadowed_re),
		.we(classa_ctrl_shadowed_gated_we),
		.wd(classa_ctrl_shadowed_en_e1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[772]),
		.qs(classa_ctrl_shadowed_en_e1_qs),
		.err_update(classa_ctrl_shadowed_en_e1_update_err),
		.err_storage(classa_ctrl_shadowed_en_e1_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_classa_ctrl_shadowed_en_e2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_ctrl_shadowed_re),
		.we(classa_ctrl_shadowed_gated_we),
		.wd(classa_ctrl_shadowed_en_e2_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[771]),
		.qs(classa_ctrl_shadowed_en_e2_qs),
		.err_update(classa_ctrl_shadowed_en_e2_update_err),
		.err_storage(classa_ctrl_shadowed_en_e2_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_classa_ctrl_shadowed_en_e3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_ctrl_shadowed_re),
		.we(classa_ctrl_shadowed_gated_we),
		.wd(classa_ctrl_shadowed_en_e3_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[770]),
		.qs(classa_ctrl_shadowed_en_e3_qs),
		.err_update(classa_ctrl_shadowed_en_e3_update_err),
		.err_storage(classa_ctrl_shadowed_en_e3_storage_err)
	);
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_classa_ctrl_shadowed_map_e0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_ctrl_shadowed_re),
		.we(classa_ctrl_shadowed_gated_we),
		.wd(classa_ctrl_shadowed_map_e0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[769-:2]),
		.qs(classa_ctrl_shadowed_map_e0_qs),
		.err_update(classa_ctrl_shadowed_map_e0_update_err),
		.err_storage(classa_ctrl_shadowed_map_e0_storage_err)
	);
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h1)
	) u_classa_ctrl_shadowed_map_e1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_ctrl_shadowed_re),
		.we(classa_ctrl_shadowed_gated_we),
		.wd(classa_ctrl_shadowed_map_e1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[767-:2]),
		.qs(classa_ctrl_shadowed_map_e1_qs),
		.err_update(classa_ctrl_shadowed_map_e1_update_err),
		.err_storage(classa_ctrl_shadowed_map_e1_storage_err)
	);
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h2)
	) u_classa_ctrl_shadowed_map_e2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_ctrl_shadowed_re),
		.we(classa_ctrl_shadowed_gated_we),
		.wd(classa_ctrl_shadowed_map_e2_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[765-:2]),
		.qs(classa_ctrl_shadowed_map_e2_qs),
		.err_update(classa_ctrl_shadowed_map_e2_update_err),
		.err_storage(classa_ctrl_shadowed_map_e2_storage_err)
	);
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h3)
	) u_classa_ctrl_shadowed_map_e3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_ctrl_shadowed_re),
		.we(classa_ctrl_shadowed_gated_we),
		.wd(classa_ctrl_shadowed_map_e3_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[763-:2]),
		.qs(classa_ctrl_shadowed_map_e3_qs),
		.err_update(classa_ctrl_shadowed_map_e3_update_err),
		.err_storage(classa_ctrl_shadowed_map_e3_storage_err)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_classa_clr_regwen(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(classa_clr_regwen_we),
		.wd(classa_clr_regwen_wd),
		.de(hw2reg[210]),
		.d(hw2reg[211]),
		.qs(classa_clr_regwen_qs)
	);
	wire classa_clr_shadowed_qe;
	wire [0:0] classa_clr_shadowed_flds_we;
	prim_flop #(
		.Width(1),
		.ResetValue(0)
	) u_classa_clr_shadowed0_qe(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(&classa_clr_shadowed_flds_we),
		.q_o(classa_clr_shadowed_qe)
	);
	wire classa_clr_shadowed_gated_we;
	assign classa_clr_shadowed_gated_we = classa_clr_shadowed_we & classa_clr_regwen_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_classa_clr_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_clr_shadowed_re),
		.we(classa_clr_shadowed_gated_we),
		.wd(classa_clr_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.qe(classa_clr_shadowed_flds_we[0]),
		.q(reg2hw[761]),
		.qs(classa_clr_shadowed_qs),
		.err_update(classa_clr_shadowed_update_err),
		.err_storage(classa_clr_shadowed_storage_err)
	);
	assign reg2hw[760] = classa_clr_shadowed_qe;
	prim_subreg_ext #(.DW(16)) u_classa_accum_cnt(
		.re(classa_accum_cnt_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[209-:16]),
		.qs(classa_accum_cnt_qs)
	);
	wire classa_accum_thresh_shadowed_gated_we;
	assign classa_accum_thresh_shadowed_gated_we = classa_accum_thresh_shadowed_we & classa_regwen_qs;
	prim_subreg_shadow #(
		.DW(16),
		.SwAccess(3'd0),
		.RESVAL(16'h0000)
	) u_classa_accum_thresh_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_accum_thresh_shadowed_re),
		.we(classa_accum_thresh_shadowed_gated_we),
		.wd(classa_accum_thresh_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[759-:16]),
		.qs(classa_accum_thresh_shadowed_qs),
		.err_update(classa_accum_thresh_shadowed_update_err),
		.err_storage(classa_accum_thresh_shadowed_storage_err)
	);
	wire classa_timeout_cyc_shadowed_gated_we;
	assign classa_timeout_cyc_shadowed_gated_we = classa_timeout_cyc_shadowed_we & classa_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classa_timeout_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_timeout_cyc_shadowed_re),
		.we(classa_timeout_cyc_shadowed_gated_we),
		.wd(classa_timeout_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[743-:32]),
		.qs(classa_timeout_cyc_shadowed_qs),
		.err_update(classa_timeout_cyc_shadowed_update_err),
		.err_storage(classa_timeout_cyc_shadowed_storage_err)
	);
	wire classa_crashdump_trigger_shadowed_gated_we;
	assign classa_crashdump_trigger_shadowed_gated_we = classa_crashdump_trigger_shadowed_we & classa_regwen_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_classa_crashdump_trigger_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_crashdump_trigger_shadowed_re),
		.we(classa_crashdump_trigger_shadowed_gated_we),
		.wd(classa_crashdump_trigger_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[711-:2]),
		.qs(classa_crashdump_trigger_shadowed_qs),
		.err_update(classa_crashdump_trigger_shadowed_update_err),
		.err_storage(classa_crashdump_trigger_shadowed_storage_err)
	);
	wire classa_phase0_cyc_shadowed_gated_we;
	assign classa_phase0_cyc_shadowed_gated_we = classa_phase0_cyc_shadowed_we & classa_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classa_phase0_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_phase0_cyc_shadowed_re),
		.we(classa_phase0_cyc_shadowed_gated_we),
		.wd(classa_phase0_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[709-:32]),
		.qs(classa_phase0_cyc_shadowed_qs),
		.err_update(classa_phase0_cyc_shadowed_update_err),
		.err_storage(classa_phase0_cyc_shadowed_storage_err)
	);
	wire classa_phase1_cyc_shadowed_gated_we;
	assign classa_phase1_cyc_shadowed_gated_we = classa_phase1_cyc_shadowed_we & classa_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classa_phase1_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_phase1_cyc_shadowed_re),
		.we(classa_phase1_cyc_shadowed_gated_we),
		.wd(classa_phase1_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[677-:32]),
		.qs(classa_phase1_cyc_shadowed_qs),
		.err_update(classa_phase1_cyc_shadowed_update_err),
		.err_storage(classa_phase1_cyc_shadowed_storage_err)
	);
	wire classa_phase2_cyc_shadowed_gated_we;
	assign classa_phase2_cyc_shadowed_gated_we = classa_phase2_cyc_shadowed_we & classa_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classa_phase2_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_phase2_cyc_shadowed_re),
		.we(classa_phase2_cyc_shadowed_gated_we),
		.wd(classa_phase2_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[645-:32]),
		.qs(classa_phase2_cyc_shadowed_qs),
		.err_update(classa_phase2_cyc_shadowed_update_err),
		.err_storage(classa_phase2_cyc_shadowed_storage_err)
	);
	wire classa_phase3_cyc_shadowed_gated_we;
	assign classa_phase3_cyc_shadowed_gated_we = classa_phase3_cyc_shadowed_we & classa_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classa_phase3_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classa_phase3_cyc_shadowed_re),
		.we(classa_phase3_cyc_shadowed_gated_we),
		.wd(classa_phase3_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[613-:32]),
		.qs(classa_phase3_cyc_shadowed_qs),
		.err_update(classa_phase3_cyc_shadowed_update_err),
		.err_storage(classa_phase3_cyc_shadowed_storage_err)
	);
	prim_subreg_ext #(.DW(32)) u_classa_esc_cnt(
		.re(classa_esc_cnt_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[193-:32]),
		.qs(classa_esc_cnt_qs)
	);
	prim_subreg_ext #(.DW(3)) u_classa_state(
		.re(classa_state_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[161-:3]),
		.qs(classa_state_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_classb_regwen(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(classb_regwen_we),
		.wd(classb_regwen_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(classb_regwen_qs)
	);
	wire classb_ctrl_shadowed_gated_we;
	assign classb_ctrl_shadowed_gated_we = classb_ctrl_shadowed_we & classb_regwen_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_classb_ctrl_shadowed_en(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_ctrl_shadowed_re),
		.we(classb_ctrl_shadowed_gated_we),
		.wd(classb_ctrl_shadowed_en_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[581]),
		.qs(classb_ctrl_shadowed_en_qs),
		.err_update(classb_ctrl_shadowed_en_update_err),
		.err_storage(classb_ctrl_shadowed_en_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_classb_ctrl_shadowed_lock(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_ctrl_shadowed_re),
		.we(classb_ctrl_shadowed_gated_we),
		.wd(classb_ctrl_shadowed_lock_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[580]),
		.qs(classb_ctrl_shadowed_lock_qs),
		.err_update(classb_ctrl_shadowed_lock_update_err),
		.err_storage(classb_ctrl_shadowed_lock_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_classb_ctrl_shadowed_en_e0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_ctrl_shadowed_re),
		.we(classb_ctrl_shadowed_gated_we),
		.wd(classb_ctrl_shadowed_en_e0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[579]),
		.qs(classb_ctrl_shadowed_en_e0_qs),
		.err_update(classb_ctrl_shadowed_en_e0_update_err),
		.err_storage(classb_ctrl_shadowed_en_e0_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_classb_ctrl_shadowed_en_e1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_ctrl_shadowed_re),
		.we(classb_ctrl_shadowed_gated_we),
		.wd(classb_ctrl_shadowed_en_e1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[578]),
		.qs(classb_ctrl_shadowed_en_e1_qs),
		.err_update(classb_ctrl_shadowed_en_e1_update_err),
		.err_storage(classb_ctrl_shadowed_en_e1_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_classb_ctrl_shadowed_en_e2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_ctrl_shadowed_re),
		.we(classb_ctrl_shadowed_gated_we),
		.wd(classb_ctrl_shadowed_en_e2_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[577]),
		.qs(classb_ctrl_shadowed_en_e2_qs),
		.err_update(classb_ctrl_shadowed_en_e2_update_err),
		.err_storage(classb_ctrl_shadowed_en_e2_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_classb_ctrl_shadowed_en_e3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_ctrl_shadowed_re),
		.we(classb_ctrl_shadowed_gated_we),
		.wd(classb_ctrl_shadowed_en_e3_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[576]),
		.qs(classb_ctrl_shadowed_en_e3_qs),
		.err_update(classb_ctrl_shadowed_en_e3_update_err),
		.err_storage(classb_ctrl_shadowed_en_e3_storage_err)
	);
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_classb_ctrl_shadowed_map_e0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_ctrl_shadowed_re),
		.we(classb_ctrl_shadowed_gated_we),
		.wd(classb_ctrl_shadowed_map_e0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[575-:2]),
		.qs(classb_ctrl_shadowed_map_e0_qs),
		.err_update(classb_ctrl_shadowed_map_e0_update_err),
		.err_storage(classb_ctrl_shadowed_map_e0_storage_err)
	);
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h1)
	) u_classb_ctrl_shadowed_map_e1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_ctrl_shadowed_re),
		.we(classb_ctrl_shadowed_gated_we),
		.wd(classb_ctrl_shadowed_map_e1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[573-:2]),
		.qs(classb_ctrl_shadowed_map_e1_qs),
		.err_update(classb_ctrl_shadowed_map_e1_update_err),
		.err_storage(classb_ctrl_shadowed_map_e1_storage_err)
	);
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h2)
	) u_classb_ctrl_shadowed_map_e2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_ctrl_shadowed_re),
		.we(classb_ctrl_shadowed_gated_we),
		.wd(classb_ctrl_shadowed_map_e2_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[571-:2]),
		.qs(classb_ctrl_shadowed_map_e2_qs),
		.err_update(classb_ctrl_shadowed_map_e2_update_err),
		.err_storage(classb_ctrl_shadowed_map_e2_storage_err)
	);
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h3)
	) u_classb_ctrl_shadowed_map_e3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_ctrl_shadowed_re),
		.we(classb_ctrl_shadowed_gated_we),
		.wd(classb_ctrl_shadowed_map_e3_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[569-:2]),
		.qs(classb_ctrl_shadowed_map_e3_qs),
		.err_update(classb_ctrl_shadowed_map_e3_update_err),
		.err_storage(classb_ctrl_shadowed_map_e3_storage_err)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_classb_clr_regwen(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(classb_clr_regwen_we),
		.wd(classb_clr_regwen_wd),
		.de(hw2reg[157]),
		.d(hw2reg[158]),
		.qs(classb_clr_regwen_qs)
	);
	wire classb_clr_shadowed_qe;
	wire [0:0] classb_clr_shadowed_flds_we;
	prim_flop #(
		.Width(1),
		.ResetValue(0)
	) u_classb_clr_shadowed0_qe(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(&classb_clr_shadowed_flds_we),
		.q_o(classb_clr_shadowed_qe)
	);
	wire classb_clr_shadowed_gated_we;
	assign classb_clr_shadowed_gated_we = classb_clr_shadowed_we & classb_clr_regwen_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_classb_clr_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_clr_shadowed_re),
		.we(classb_clr_shadowed_gated_we),
		.wd(classb_clr_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.qe(classb_clr_shadowed_flds_we[0]),
		.q(reg2hw[567]),
		.qs(classb_clr_shadowed_qs),
		.err_update(classb_clr_shadowed_update_err),
		.err_storage(classb_clr_shadowed_storage_err)
	);
	assign reg2hw[566] = classb_clr_shadowed_qe;
	prim_subreg_ext #(.DW(16)) u_classb_accum_cnt(
		.re(classb_accum_cnt_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[156-:16]),
		.qs(classb_accum_cnt_qs)
	);
	wire classb_accum_thresh_shadowed_gated_we;
	assign classb_accum_thresh_shadowed_gated_we = classb_accum_thresh_shadowed_we & classb_regwen_qs;
	prim_subreg_shadow #(
		.DW(16),
		.SwAccess(3'd0),
		.RESVAL(16'h0000)
	) u_classb_accum_thresh_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_accum_thresh_shadowed_re),
		.we(classb_accum_thresh_shadowed_gated_we),
		.wd(classb_accum_thresh_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[565-:16]),
		.qs(classb_accum_thresh_shadowed_qs),
		.err_update(classb_accum_thresh_shadowed_update_err),
		.err_storage(classb_accum_thresh_shadowed_storage_err)
	);
	wire classb_timeout_cyc_shadowed_gated_we;
	assign classb_timeout_cyc_shadowed_gated_we = classb_timeout_cyc_shadowed_we & classb_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classb_timeout_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_timeout_cyc_shadowed_re),
		.we(classb_timeout_cyc_shadowed_gated_we),
		.wd(classb_timeout_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[549-:32]),
		.qs(classb_timeout_cyc_shadowed_qs),
		.err_update(classb_timeout_cyc_shadowed_update_err),
		.err_storage(classb_timeout_cyc_shadowed_storage_err)
	);
	wire classb_crashdump_trigger_shadowed_gated_we;
	assign classb_crashdump_trigger_shadowed_gated_we = classb_crashdump_trigger_shadowed_we & classb_regwen_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_classb_crashdump_trigger_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_crashdump_trigger_shadowed_re),
		.we(classb_crashdump_trigger_shadowed_gated_we),
		.wd(classb_crashdump_trigger_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[517-:2]),
		.qs(classb_crashdump_trigger_shadowed_qs),
		.err_update(classb_crashdump_trigger_shadowed_update_err),
		.err_storage(classb_crashdump_trigger_shadowed_storage_err)
	);
	wire classb_phase0_cyc_shadowed_gated_we;
	assign classb_phase0_cyc_shadowed_gated_we = classb_phase0_cyc_shadowed_we & classb_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classb_phase0_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_phase0_cyc_shadowed_re),
		.we(classb_phase0_cyc_shadowed_gated_we),
		.wd(classb_phase0_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[515-:32]),
		.qs(classb_phase0_cyc_shadowed_qs),
		.err_update(classb_phase0_cyc_shadowed_update_err),
		.err_storage(classb_phase0_cyc_shadowed_storage_err)
	);
	wire classb_phase1_cyc_shadowed_gated_we;
	assign classb_phase1_cyc_shadowed_gated_we = classb_phase1_cyc_shadowed_we & classb_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classb_phase1_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_phase1_cyc_shadowed_re),
		.we(classb_phase1_cyc_shadowed_gated_we),
		.wd(classb_phase1_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[483-:32]),
		.qs(classb_phase1_cyc_shadowed_qs),
		.err_update(classb_phase1_cyc_shadowed_update_err),
		.err_storage(classb_phase1_cyc_shadowed_storage_err)
	);
	wire classb_phase2_cyc_shadowed_gated_we;
	assign classb_phase2_cyc_shadowed_gated_we = classb_phase2_cyc_shadowed_we & classb_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classb_phase2_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_phase2_cyc_shadowed_re),
		.we(classb_phase2_cyc_shadowed_gated_we),
		.wd(classb_phase2_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[451-:32]),
		.qs(classb_phase2_cyc_shadowed_qs),
		.err_update(classb_phase2_cyc_shadowed_update_err),
		.err_storage(classb_phase2_cyc_shadowed_storage_err)
	);
	wire classb_phase3_cyc_shadowed_gated_we;
	assign classb_phase3_cyc_shadowed_gated_we = classb_phase3_cyc_shadowed_we & classb_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classb_phase3_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classb_phase3_cyc_shadowed_re),
		.we(classb_phase3_cyc_shadowed_gated_we),
		.wd(classb_phase3_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[419-:32]),
		.qs(classb_phase3_cyc_shadowed_qs),
		.err_update(classb_phase3_cyc_shadowed_update_err),
		.err_storage(classb_phase3_cyc_shadowed_storage_err)
	);
	prim_subreg_ext #(.DW(32)) u_classb_esc_cnt(
		.re(classb_esc_cnt_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[140-:32]),
		.qs(classb_esc_cnt_qs)
	);
	prim_subreg_ext #(.DW(3)) u_classb_state(
		.re(classb_state_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[108-:3]),
		.qs(classb_state_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_classc_regwen(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(classc_regwen_we),
		.wd(classc_regwen_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(classc_regwen_qs)
	);
	wire classc_ctrl_shadowed_gated_we;
	assign classc_ctrl_shadowed_gated_we = classc_ctrl_shadowed_we & classc_regwen_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_classc_ctrl_shadowed_en(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_ctrl_shadowed_re),
		.we(classc_ctrl_shadowed_gated_we),
		.wd(classc_ctrl_shadowed_en_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[387]),
		.qs(classc_ctrl_shadowed_en_qs),
		.err_update(classc_ctrl_shadowed_en_update_err),
		.err_storage(classc_ctrl_shadowed_en_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_classc_ctrl_shadowed_lock(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_ctrl_shadowed_re),
		.we(classc_ctrl_shadowed_gated_we),
		.wd(classc_ctrl_shadowed_lock_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[386]),
		.qs(classc_ctrl_shadowed_lock_qs),
		.err_update(classc_ctrl_shadowed_lock_update_err),
		.err_storage(classc_ctrl_shadowed_lock_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_classc_ctrl_shadowed_en_e0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_ctrl_shadowed_re),
		.we(classc_ctrl_shadowed_gated_we),
		.wd(classc_ctrl_shadowed_en_e0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[385]),
		.qs(classc_ctrl_shadowed_en_e0_qs),
		.err_update(classc_ctrl_shadowed_en_e0_update_err),
		.err_storage(classc_ctrl_shadowed_en_e0_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_classc_ctrl_shadowed_en_e1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_ctrl_shadowed_re),
		.we(classc_ctrl_shadowed_gated_we),
		.wd(classc_ctrl_shadowed_en_e1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[384]),
		.qs(classc_ctrl_shadowed_en_e1_qs),
		.err_update(classc_ctrl_shadowed_en_e1_update_err),
		.err_storage(classc_ctrl_shadowed_en_e1_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_classc_ctrl_shadowed_en_e2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_ctrl_shadowed_re),
		.we(classc_ctrl_shadowed_gated_we),
		.wd(classc_ctrl_shadowed_en_e2_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[383]),
		.qs(classc_ctrl_shadowed_en_e2_qs),
		.err_update(classc_ctrl_shadowed_en_e2_update_err),
		.err_storage(classc_ctrl_shadowed_en_e2_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_classc_ctrl_shadowed_en_e3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_ctrl_shadowed_re),
		.we(classc_ctrl_shadowed_gated_we),
		.wd(classc_ctrl_shadowed_en_e3_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[382]),
		.qs(classc_ctrl_shadowed_en_e3_qs),
		.err_update(classc_ctrl_shadowed_en_e3_update_err),
		.err_storage(classc_ctrl_shadowed_en_e3_storage_err)
	);
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_classc_ctrl_shadowed_map_e0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_ctrl_shadowed_re),
		.we(classc_ctrl_shadowed_gated_we),
		.wd(classc_ctrl_shadowed_map_e0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[381-:2]),
		.qs(classc_ctrl_shadowed_map_e0_qs),
		.err_update(classc_ctrl_shadowed_map_e0_update_err),
		.err_storage(classc_ctrl_shadowed_map_e0_storage_err)
	);
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h1)
	) u_classc_ctrl_shadowed_map_e1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_ctrl_shadowed_re),
		.we(classc_ctrl_shadowed_gated_we),
		.wd(classc_ctrl_shadowed_map_e1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[379-:2]),
		.qs(classc_ctrl_shadowed_map_e1_qs),
		.err_update(classc_ctrl_shadowed_map_e1_update_err),
		.err_storage(classc_ctrl_shadowed_map_e1_storage_err)
	);
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h2)
	) u_classc_ctrl_shadowed_map_e2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_ctrl_shadowed_re),
		.we(classc_ctrl_shadowed_gated_we),
		.wd(classc_ctrl_shadowed_map_e2_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[377-:2]),
		.qs(classc_ctrl_shadowed_map_e2_qs),
		.err_update(classc_ctrl_shadowed_map_e2_update_err),
		.err_storage(classc_ctrl_shadowed_map_e2_storage_err)
	);
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h3)
	) u_classc_ctrl_shadowed_map_e3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_ctrl_shadowed_re),
		.we(classc_ctrl_shadowed_gated_we),
		.wd(classc_ctrl_shadowed_map_e3_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[375-:2]),
		.qs(classc_ctrl_shadowed_map_e3_qs),
		.err_update(classc_ctrl_shadowed_map_e3_update_err),
		.err_storage(classc_ctrl_shadowed_map_e3_storage_err)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_classc_clr_regwen(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(classc_clr_regwen_we),
		.wd(classc_clr_regwen_wd),
		.de(hw2reg[104]),
		.d(hw2reg[105]),
		.qs(classc_clr_regwen_qs)
	);
	wire classc_clr_shadowed_qe;
	wire [0:0] classc_clr_shadowed_flds_we;
	prim_flop #(
		.Width(1),
		.ResetValue(0)
	) u_classc_clr_shadowed0_qe(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(&classc_clr_shadowed_flds_we),
		.q_o(classc_clr_shadowed_qe)
	);
	wire classc_clr_shadowed_gated_we;
	assign classc_clr_shadowed_gated_we = classc_clr_shadowed_we & classc_clr_regwen_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_classc_clr_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_clr_shadowed_re),
		.we(classc_clr_shadowed_gated_we),
		.wd(classc_clr_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.qe(classc_clr_shadowed_flds_we[0]),
		.q(reg2hw[373]),
		.qs(classc_clr_shadowed_qs),
		.err_update(classc_clr_shadowed_update_err),
		.err_storage(classc_clr_shadowed_storage_err)
	);
	assign reg2hw[372] = classc_clr_shadowed_qe;
	prim_subreg_ext #(.DW(16)) u_classc_accum_cnt(
		.re(classc_accum_cnt_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[103-:16]),
		.qs(classc_accum_cnt_qs)
	);
	wire classc_accum_thresh_shadowed_gated_we;
	assign classc_accum_thresh_shadowed_gated_we = classc_accum_thresh_shadowed_we & classc_regwen_qs;
	prim_subreg_shadow #(
		.DW(16),
		.SwAccess(3'd0),
		.RESVAL(16'h0000)
	) u_classc_accum_thresh_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_accum_thresh_shadowed_re),
		.we(classc_accum_thresh_shadowed_gated_we),
		.wd(classc_accum_thresh_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[371-:16]),
		.qs(classc_accum_thresh_shadowed_qs),
		.err_update(classc_accum_thresh_shadowed_update_err),
		.err_storage(classc_accum_thresh_shadowed_storage_err)
	);
	wire classc_timeout_cyc_shadowed_gated_we;
	assign classc_timeout_cyc_shadowed_gated_we = classc_timeout_cyc_shadowed_we & classc_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classc_timeout_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_timeout_cyc_shadowed_re),
		.we(classc_timeout_cyc_shadowed_gated_we),
		.wd(classc_timeout_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[355-:32]),
		.qs(classc_timeout_cyc_shadowed_qs),
		.err_update(classc_timeout_cyc_shadowed_update_err),
		.err_storage(classc_timeout_cyc_shadowed_storage_err)
	);
	wire classc_crashdump_trigger_shadowed_gated_we;
	assign classc_crashdump_trigger_shadowed_gated_we = classc_crashdump_trigger_shadowed_we & classc_regwen_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_classc_crashdump_trigger_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_crashdump_trigger_shadowed_re),
		.we(classc_crashdump_trigger_shadowed_gated_we),
		.wd(classc_crashdump_trigger_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[323-:2]),
		.qs(classc_crashdump_trigger_shadowed_qs),
		.err_update(classc_crashdump_trigger_shadowed_update_err),
		.err_storage(classc_crashdump_trigger_shadowed_storage_err)
	);
	wire classc_phase0_cyc_shadowed_gated_we;
	assign classc_phase0_cyc_shadowed_gated_we = classc_phase0_cyc_shadowed_we & classc_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classc_phase0_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_phase0_cyc_shadowed_re),
		.we(classc_phase0_cyc_shadowed_gated_we),
		.wd(classc_phase0_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[321-:32]),
		.qs(classc_phase0_cyc_shadowed_qs),
		.err_update(classc_phase0_cyc_shadowed_update_err),
		.err_storage(classc_phase0_cyc_shadowed_storage_err)
	);
	wire classc_phase1_cyc_shadowed_gated_we;
	assign classc_phase1_cyc_shadowed_gated_we = classc_phase1_cyc_shadowed_we & classc_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classc_phase1_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_phase1_cyc_shadowed_re),
		.we(classc_phase1_cyc_shadowed_gated_we),
		.wd(classc_phase1_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[289-:32]),
		.qs(classc_phase1_cyc_shadowed_qs),
		.err_update(classc_phase1_cyc_shadowed_update_err),
		.err_storage(classc_phase1_cyc_shadowed_storage_err)
	);
	wire classc_phase2_cyc_shadowed_gated_we;
	assign classc_phase2_cyc_shadowed_gated_we = classc_phase2_cyc_shadowed_we & classc_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classc_phase2_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_phase2_cyc_shadowed_re),
		.we(classc_phase2_cyc_shadowed_gated_we),
		.wd(classc_phase2_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[257-:32]),
		.qs(classc_phase2_cyc_shadowed_qs),
		.err_update(classc_phase2_cyc_shadowed_update_err),
		.err_storage(classc_phase2_cyc_shadowed_storage_err)
	);
	wire classc_phase3_cyc_shadowed_gated_we;
	assign classc_phase3_cyc_shadowed_gated_we = classc_phase3_cyc_shadowed_we & classc_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classc_phase3_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classc_phase3_cyc_shadowed_re),
		.we(classc_phase3_cyc_shadowed_gated_we),
		.wd(classc_phase3_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[225-:32]),
		.qs(classc_phase3_cyc_shadowed_qs),
		.err_update(classc_phase3_cyc_shadowed_update_err),
		.err_storage(classc_phase3_cyc_shadowed_storage_err)
	);
	prim_subreg_ext #(.DW(32)) u_classc_esc_cnt(
		.re(classc_esc_cnt_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[87-:32]),
		.qs(classc_esc_cnt_qs)
	);
	prim_subreg_ext #(.DW(3)) u_classc_state(
		.re(classc_state_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[55-:3]),
		.qs(classc_state_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_classd_regwen(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(classd_regwen_we),
		.wd(classd_regwen_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(classd_regwen_qs)
	);
	wire classd_ctrl_shadowed_gated_we;
	assign classd_ctrl_shadowed_gated_we = classd_ctrl_shadowed_we & classd_regwen_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_classd_ctrl_shadowed_en(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_ctrl_shadowed_re),
		.we(classd_ctrl_shadowed_gated_we),
		.wd(classd_ctrl_shadowed_en_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[193]),
		.qs(classd_ctrl_shadowed_en_qs),
		.err_update(classd_ctrl_shadowed_en_update_err),
		.err_storage(classd_ctrl_shadowed_en_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_classd_ctrl_shadowed_lock(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_ctrl_shadowed_re),
		.we(classd_ctrl_shadowed_gated_we),
		.wd(classd_ctrl_shadowed_lock_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[192]),
		.qs(classd_ctrl_shadowed_lock_qs),
		.err_update(classd_ctrl_shadowed_lock_update_err),
		.err_storage(classd_ctrl_shadowed_lock_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_classd_ctrl_shadowed_en_e0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_ctrl_shadowed_re),
		.we(classd_ctrl_shadowed_gated_we),
		.wd(classd_ctrl_shadowed_en_e0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[191]),
		.qs(classd_ctrl_shadowed_en_e0_qs),
		.err_update(classd_ctrl_shadowed_en_e0_update_err),
		.err_storage(classd_ctrl_shadowed_en_e0_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_classd_ctrl_shadowed_en_e1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_ctrl_shadowed_re),
		.we(classd_ctrl_shadowed_gated_we),
		.wd(classd_ctrl_shadowed_en_e1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[190]),
		.qs(classd_ctrl_shadowed_en_e1_qs),
		.err_update(classd_ctrl_shadowed_en_e1_update_err),
		.err_storage(classd_ctrl_shadowed_en_e1_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_classd_ctrl_shadowed_en_e2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_ctrl_shadowed_re),
		.we(classd_ctrl_shadowed_gated_we),
		.wd(classd_ctrl_shadowed_en_e2_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[189]),
		.qs(classd_ctrl_shadowed_en_e2_qs),
		.err_update(classd_ctrl_shadowed_en_e2_update_err),
		.err_storage(classd_ctrl_shadowed_en_e2_storage_err)
	);
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_classd_ctrl_shadowed_en_e3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_ctrl_shadowed_re),
		.we(classd_ctrl_shadowed_gated_we),
		.wd(classd_ctrl_shadowed_en_e3_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[188]),
		.qs(classd_ctrl_shadowed_en_e3_qs),
		.err_update(classd_ctrl_shadowed_en_e3_update_err),
		.err_storage(classd_ctrl_shadowed_en_e3_storage_err)
	);
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_classd_ctrl_shadowed_map_e0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_ctrl_shadowed_re),
		.we(classd_ctrl_shadowed_gated_we),
		.wd(classd_ctrl_shadowed_map_e0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[187-:2]),
		.qs(classd_ctrl_shadowed_map_e0_qs),
		.err_update(classd_ctrl_shadowed_map_e0_update_err),
		.err_storage(classd_ctrl_shadowed_map_e0_storage_err)
	);
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h1)
	) u_classd_ctrl_shadowed_map_e1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_ctrl_shadowed_re),
		.we(classd_ctrl_shadowed_gated_we),
		.wd(classd_ctrl_shadowed_map_e1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[185-:2]),
		.qs(classd_ctrl_shadowed_map_e1_qs),
		.err_update(classd_ctrl_shadowed_map_e1_update_err),
		.err_storage(classd_ctrl_shadowed_map_e1_storage_err)
	);
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h2)
	) u_classd_ctrl_shadowed_map_e2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_ctrl_shadowed_re),
		.we(classd_ctrl_shadowed_gated_we),
		.wd(classd_ctrl_shadowed_map_e2_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[183-:2]),
		.qs(classd_ctrl_shadowed_map_e2_qs),
		.err_update(classd_ctrl_shadowed_map_e2_update_err),
		.err_storage(classd_ctrl_shadowed_map_e2_storage_err)
	);
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h3)
	) u_classd_ctrl_shadowed_map_e3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_ctrl_shadowed_re),
		.we(classd_ctrl_shadowed_gated_we),
		.wd(classd_ctrl_shadowed_map_e3_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[181-:2]),
		.qs(classd_ctrl_shadowed_map_e3_qs),
		.err_update(classd_ctrl_shadowed_map_e3_update_err),
		.err_storage(classd_ctrl_shadowed_map_e3_storage_err)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_classd_clr_regwen(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(classd_clr_regwen_we),
		.wd(classd_clr_regwen_wd),
		.de(hw2reg[51]),
		.d(hw2reg[52]),
		.qs(classd_clr_regwen_qs)
	);
	wire classd_clr_shadowed_qe;
	wire [0:0] classd_clr_shadowed_flds_we;
	prim_flop #(
		.Width(1),
		.ResetValue(0)
	) u_classd_clr_shadowed0_qe(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(&classd_clr_shadowed_flds_we),
		.q_o(classd_clr_shadowed_qe)
	);
	wire classd_clr_shadowed_gated_we;
	assign classd_clr_shadowed_gated_we = classd_clr_shadowed_we & classd_clr_regwen_qs;
	prim_subreg_shadow #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_classd_clr_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_clr_shadowed_re),
		.we(classd_clr_shadowed_gated_we),
		.wd(classd_clr_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.qe(classd_clr_shadowed_flds_we[0]),
		.q(reg2hw[179]),
		.qs(classd_clr_shadowed_qs),
		.err_update(classd_clr_shadowed_update_err),
		.err_storage(classd_clr_shadowed_storage_err)
	);
	assign reg2hw[178] = classd_clr_shadowed_qe;
	prim_subreg_ext #(.DW(16)) u_classd_accum_cnt(
		.re(classd_accum_cnt_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[50-:16]),
		.qs(classd_accum_cnt_qs)
	);
	wire classd_accum_thresh_shadowed_gated_we;
	assign classd_accum_thresh_shadowed_gated_we = classd_accum_thresh_shadowed_we & classd_regwen_qs;
	prim_subreg_shadow #(
		.DW(16),
		.SwAccess(3'd0),
		.RESVAL(16'h0000)
	) u_classd_accum_thresh_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_accum_thresh_shadowed_re),
		.we(classd_accum_thresh_shadowed_gated_we),
		.wd(classd_accum_thresh_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[177-:16]),
		.qs(classd_accum_thresh_shadowed_qs),
		.err_update(classd_accum_thresh_shadowed_update_err),
		.err_storage(classd_accum_thresh_shadowed_storage_err)
	);
	wire classd_timeout_cyc_shadowed_gated_we;
	assign classd_timeout_cyc_shadowed_gated_we = classd_timeout_cyc_shadowed_we & classd_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classd_timeout_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_timeout_cyc_shadowed_re),
		.we(classd_timeout_cyc_shadowed_gated_we),
		.wd(classd_timeout_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[161-:32]),
		.qs(classd_timeout_cyc_shadowed_qs),
		.err_update(classd_timeout_cyc_shadowed_update_err),
		.err_storage(classd_timeout_cyc_shadowed_storage_err)
	);
	wire classd_crashdump_trigger_shadowed_gated_we;
	assign classd_crashdump_trigger_shadowed_gated_we = classd_crashdump_trigger_shadowed_we & classd_regwen_qs;
	prim_subreg_shadow #(
		.DW(2),
		.SwAccess(3'd0),
		.RESVAL(2'h0)
	) u_classd_crashdump_trigger_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_crashdump_trigger_shadowed_re),
		.we(classd_crashdump_trigger_shadowed_gated_we),
		.wd(classd_crashdump_trigger_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[129-:2]),
		.qs(classd_crashdump_trigger_shadowed_qs),
		.err_update(classd_crashdump_trigger_shadowed_update_err),
		.err_storage(classd_crashdump_trigger_shadowed_storage_err)
	);
	wire classd_phase0_cyc_shadowed_gated_we;
	assign classd_phase0_cyc_shadowed_gated_we = classd_phase0_cyc_shadowed_we & classd_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classd_phase0_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_phase0_cyc_shadowed_re),
		.we(classd_phase0_cyc_shadowed_gated_we),
		.wd(classd_phase0_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[127-:32]),
		.qs(classd_phase0_cyc_shadowed_qs),
		.err_update(classd_phase0_cyc_shadowed_update_err),
		.err_storage(classd_phase0_cyc_shadowed_storage_err)
	);
	wire classd_phase1_cyc_shadowed_gated_we;
	assign classd_phase1_cyc_shadowed_gated_we = classd_phase1_cyc_shadowed_we & classd_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classd_phase1_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_phase1_cyc_shadowed_re),
		.we(classd_phase1_cyc_shadowed_gated_we),
		.wd(classd_phase1_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[95-:32]),
		.qs(classd_phase1_cyc_shadowed_qs),
		.err_update(classd_phase1_cyc_shadowed_update_err),
		.err_storage(classd_phase1_cyc_shadowed_storage_err)
	);
	wire classd_phase2_cyc_shadowed_gated_we;
	assign classd_phase2_cyc_shadowed_gated_we = classd_phase2_cyc_shadowed_we & classd_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classd_phase2_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_phase2_cyc_shadowed_re),
		.we(classd_phase2_cyc_shadowed_gated_we),
		.wd(classd_phase2_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[63-:32]),
		.qs(classd_phase2_cyc_shadowed_qs),
		.err_update(classd_phase2_cyc_shadowed_update_err),
		.err_storage(classd_phase2_cyc_shadowed_storage_err)
	);
	wire classd_phase3_cyc_shadowed_gated_we;
	assign classd_phase3_cyc_shadowed_gated_we = classd_phase3_cyc_shadowed_we & classd_regwen_qs;
	prim_subreg_shadow #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_classd_phase3_cyc_shadowed(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rst_shadowed_ni(rst_shadowed_ni),
		.re(classd_phase3_cyc_shadowed_re),
		.we(classd_phase3_cyc_shadowed_gated_we),
		.wd(classd_phase3_cyc_shadowed_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[31-:32]),
		.qs(classd_phase3_cyc_shadowed_qs),
		.err_update(classd_phase3_cyc_shadowed_update_err),
		.err_storage(classd_phase3_cyc_shadowed_storage_err)
	);
	prim_subreg_ext #(.DW(32)) u_classd_esc_cnt(
		.re(classd_esc_cnt_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[34-:32]),
		.qs(classd_esc_cnt_qs)
	);
	prim_subreg_ext #(.DW(3)) u_classd_state(
		.re(classd_state_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[2-:3]),
		.qs(classd_state_qs)
	);
	reg [349:0] addr_hit;
	localparam signed [31:0] alert_handler_reg_pkg_BlockAw = 11;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_0_OFFSET = 11'h324;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_10_OFFSET = 11'h34c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_11_OFFSET = 11'h350;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_12_OFFSET = 11'h354;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_13_OFFSET = 11'h358;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_14_OFFSET = 11'h35c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_15_OFFSET = 11'h360;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_16_OFFSET = 11'h364;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_17_OFFSET = 11'h368;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_18_OFFSET = 11'h36c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_19_OFFSET = 11'h370;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_1_OFFSET = 11'h328;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_20_OFFSET = 11'h374;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_21_OFFSET = 11'h378;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_22_OFFSET = 11'h37c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_23_OFFSET = 11'h380;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_24_OFFSET = 11'h384;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_25_OFFSET = 11'h388;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_26_OFFSET = 11'h38c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_27_OFFSET = 11'h390;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_28_OFFSET = 11'h394;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_29_OFFSET = 11'h398;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_2_OFFSET = 11'h32c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_30_OFFSET = 11'h39c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_31_OFFSET = 11'h3a0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_32_OFFSET = 11'h3a4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_33_OFFSET = 11'h3a8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_34_OFFSET = 11'h3ac;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_35_OFFSET = 11'h3b0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_36_OFFSET = 11'h3b4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_37_OFFSET = 11'h3b8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_38_OFFSET = 11'h3bc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_39_OFFSET = 11'h3c0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_3_OFFSET = 11'h330;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_40_OFFSET = 11'h3c4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_41_OFFSET = 11'h3c8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_42_OFFSET = 11'h3cc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_43_OFFSET = 11'h3d0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_44_OFFSET = 11'h3d4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_45_OFFSET = 11'h3d8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_46_OFFSET = 11'h3dc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_47_OFFSET = 11'h3e0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_48_OFFSET = 11'h3e4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_49_OFFSET = 11'h3e8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_4_OFFSET = 11'h334;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_50_OFFSET = 11'h3ec;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_51_OFFSET = 11'h3f0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_52_OFFSET = 11'h3f4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_53_OFFSET = 11'h3f8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_54_OFFSET = 11'h3fc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_55_OFFSET = 11'h400;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_56_OFFSET = 11'h404;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_57_OFFSET = 11'h408;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_58_OFFSET = 11'h40c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_59_OFFSET = 11'h410;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_5_OFFSET = 11'h338;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_60_OFFSET = 11'h414;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_61_OFFSET = 11'h418;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_62_OFFSET = 11'h41c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_63_OFFSET = 11'h420;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_64_OFFSET = 11'h424;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_6_OFFSET = 11'h33c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_7_OFFSET = 11'h340;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_8_OFFSET = 11'h344;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_9_OFFSET = 11'h348;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_0_OFFSET = 11'h220;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_10_OFFSET = 11'h248;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_11_OFFSET = 11'h24c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_12_OFFSET = 11'h250;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_13_OFFSET = 11'h254;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_14_OFFSET = 11'h258;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_15_OFFSET = 11'h25c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_16_OFFSET = 11'h260;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_17_OFFSET = 11'h264;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_18_OFFSET = 11'h268;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_19_OFFSET = 11'h26c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_1_OFFSET = 11'h224;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_20_OFFSET = 11'h270;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_21_OFFSET = 11'h274;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_22_OFFSET = 11'h278;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_23_OFFSET = 11'h27c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_24_OFFSET = 11'h280;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_25_OFFSET = 11'h284;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_26_OFFSET = 11'h288;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_27_OFFSET = 11'h28c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_28_OFFSET = 11'h290;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_29_OFFSET = 11'h294;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_2_OFFSET = 11'h228;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_30_OFFSET = 11'h298;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_31_OFFSET = 11'h29c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_32_OFFSET = 11'h2a0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_33_OFFSET = 11'h2a4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_34_OFFSET = 11'h2a8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_35_OFFSET = 11'h2ac;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_36_OFFSET = 11'h2b0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_37_OFFSET = 11'h2b4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_38_OFFSET = 11'h2b8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_39_OFFSET = 11'h2bc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_3_OFFSET = 11'h22c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_40_OFFSET = 11'h2c0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_41_OFFSET = 11'h2c4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_42_OFFSET = 11'h2c8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_43_OFFSET = 11'h2cc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_44_OFFSET = 11'h2d0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_45_OFFSET = 11'h2d4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_46_OFFSET = 11'h2d8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_47_OFFSET = 11'h2dc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_48_OFFSET = 11'h2e0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_49_OFFSET = 11'h2e4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_4_OFFSET = 11'h230;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_50_OFFSET = 11'h2e8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_51_OFFSET = 11'h2ec;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_52_OFFSET = 11'h2f0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_53_OFFSET = 11'h2f4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_54_OFFSET = 11'h2f8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_55_OFFSET = 11'h2fc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_56_OFFSET = 11'h300;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_57_OFFSET = 11'h304;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_58_OFFSET = 11'h308;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_59_OFFSET = 11'h30c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_5_OFFSET = 11'h234;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_60_OFFSET = 11'h310;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_61_OFFSET = 11'h314;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_62_OFFSET = 11'h318;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_63_OFFSET = 11'h31c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_64_OFFSET = 11'h320;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_6_OFFSET = 11'h238;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_7_OFFSET = 11'h23c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_8_OFFSET = 11'h240;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_9_OFFSET = 11'h244;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_0_OFFSET = 11'h11c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_10_OFFSET = 11'h144;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_11_OFFSET = 11'h148;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_12_OFFSET = 11'h14c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_13_OFFSET = 11'h150;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_14_OFFSET = 11'h154;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_15_OFFSET = 11'h158;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_16_OFFSET = 11'h15c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_17_OFFSET = 11'h160;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_18_OFFSET = 11'h164;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_19_OFFSET = 11'h168;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_1_OFFSET = 11'h120;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_20_OFFSET = 11'h16c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_21_OFFSET = 11'h170;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_22_OFFSET = 11'h174;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_23_OFFSET = 11'h178;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_24_OFFSET = 11'h17c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_25_OFFSET = 11'h180;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_26_OFFSET = 11'h184;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_27_OFFSET = 11'h188;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_28_OFFSET = 11'h18c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_29_OFFSET = 11'h190;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_2_OFFSET = 11'h124;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_30_OFFSET = 11'h194;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_31_OFFSET = 11'h198;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_32_OFFSET = 11'h19c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_33_OFFSET = 11'h1a0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_34_OFFSET = 11'h1a4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_35_OFFSET = 11'h1a8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_36_OFFSET = 11'h1ac;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_37_OFFSET = 11'h1b0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_38_OFFSET = 11'h1b4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_39_OFFSET = 11'h1b8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_3_OFFSET = 11'h128;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_40_OFFSET = 11'h1bc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_41_OFFSET = 11'h1c0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_42_OFFSET = 11'h1c4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_43_OFFSET = 11'h1c8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_44_OFFSET = 11'h1cc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_45_OFFSET = 11'h1d0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_46_OFFSET = 11'h1d4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_47_OFFSET = 11'h1d8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_48_OFFSET = 11'h1dc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_49_OFFSET = 11'h1e0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_4_OFFSET = 11'h12c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_50_OFFSET = 11'h1e4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_51_OFFSET = 11'h1e8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_52_OFFSET = 11'h1ec;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_53_OFFSET = 11'h1f0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_54_OFFSET = 11'h1f4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_55_OFFSET = 11'h1f8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_56_OFFSET = 11'h1fc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_57_OFFSET = 11'h200;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_58_OFFSET = 11'h204;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_59_OFFSET = 11'h208;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_5_OFFSET = 11'h130;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_60_OFFSET = 11'h20c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_61_OFFSET = 11'h210;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_62_OFFSET = 11'h214;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_63_OFFSET = 11'h218;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_64_OFFSET = 11'h21c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_6_OFFSET = 11'h134;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_7_OFFSET = 11'h138;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_8_OFFSET = 11'h13c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_9_OFFSET = 11'h140;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_0_OFFSET = 11'h018;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_10_OFFSET = 11'h040;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_11_OFFSET = 11'h044;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_12_OFFSET = 11'h048;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_13_OFFSET = 11'h04c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_14_OFFSET = 11'h050;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_15_OFFSET = 11'h054;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_16_OFFSET = 11'h058;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_17_OFFSET = 11'h05c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_18_OFFSET = 11'h060;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_19_OFFSET = 11'h064;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_1_OFFSET = 11'h01c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_20_OFFSET = 11'h068;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_21_OFFSET = 11'h06c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_22_OFFSET = 11'h070;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_23_OFFSET = 11'h074;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_24_OFFSET = 11'h078;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_25_OFFSET = 11'h07c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_26_OFFSET = 11'h080;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_27_OFFSET = 11'h084;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_28_OFFSET = 11'h088;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_29_OFFSET = 11'h08c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_2_OFFSET = 11'h020;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_30_OFFSET = 11'h090;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_31_OFFSET = 11'h094;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_32_OFFSET = 11'h098;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_33_OFFSET = 11'h09c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_34_OFFSET = 11'h0a0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_35_OFFSET = 11'h0a4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_36_OFFSET = 11'h0a8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_37_OFFSET = 11'h0ac;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_38_OFFSET = 11'h0b0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_39_OFFSET = 11'h0b4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_3_OFFSET = 11'h024;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_40_OFFSET = 11'h0b8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_41_OFFSET = 11'h0bc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_42_OFFSET = 11'h0c0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_43_OFFSET = 11'h0c4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_44_OFFSET = 11'h0c8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_45_OFFSET = 11'h0cc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_46_OFFSET = 11'h0d0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_47_OFFSET = 11'h0d4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_48_OFFSET = 11'h0d8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_49_OFFSET = 11'h0dc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_4_OFFSET = 11'h028;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_50_OFFSET = 11'h0e0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_51_OFFSET = 11'h0e4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_52_OFFSET = 11'h0e8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_53_OFFSET = 11'h0ec;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_54_OFFSET = 11'h0f0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_55_OFFSET = 11'h0f4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_56_OFFSET = 11'h0f8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_57_OFFSET = 11'h0fc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_58_OFFSET = 11'h100;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_59_OFFSET = 11'h104;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_5_OFFSET = 11'h02c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_60_OFFSET = 11'h108;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_61_OFFSET = 11'h10c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_62_OFFSET = 11'h110;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_63_OFFSET = 11'h114;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_64_OFFSET = 11'h118;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_6_OFFSET = 11'h030;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_7_OFFSET = 11'h034;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_8_OFFSET = 11'h038;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_9_OFFSET = 11'h03c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_ACCUM_CNT_OFFSET = 11'h4a8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_ACCUM_THRESH_SHADOWED_OFFSET = 11'h4ac;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_CLR_REGWEN_OFFSET = 11'h4a0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_CLR_SHADOWED_OFFSET = 11'h4a4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_CRASHDUMP_TRIGGER_SHADOWED_OFFSET = 11'h4b4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_CTRL_SHADOWED_OFFSET = 11'h49c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_ESC_CNT_OFFSET = 11'h4c8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_PHASE0_CYC_SHADOWED_OFFSET = 11'h4b8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_PHASE1_CYC_SHADOWED_OFFSET = 11'h4bc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_PHASE2_CYC_SHADOWED_OFFSET = 11'h4c0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_PHASE3_CYC_SHADOWED_OFFSET = 11'h4c4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_REGWEN_OFFSET = 11'h498;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_STATE_OFFSET = 11'h4cc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_TIMEOUT_CYC_SHADOWED_OFFSET = 11'h4b0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_ACCUM_CNT_OFFSET = 11'h4e0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_ACCUM_THRESH_SHADOWED_OFFSET = 11'h4e4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_CLR_REGWEN_OFFSET = 11'h4d8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_CLR_SHADOWED_OFFSET = 11'h4dc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_CRASHDUMP_TRIGGER_SHADOWED_OFFSET = 11'h4ec;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_CTRL_SHADOWED_OFFSET = 11'h4d4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_ESC_CNT_OFFSET = 11'h500;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_PHASE0_CYC_SHADOWED_OFFSET = 11'h4f0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_PHASE1_CYC_SHADOWED_OFFSET = 11'h4f4;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_PHASE2_CYC_SHADOWED_OFFSET = 11'h4f8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_PHASE3_CYC_SHADOWED_OFFSET = 11'h4fc;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_REGWEN_OFFSET = 11'h4d0;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_STATE_OFFSET = 11'h504;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_TIMEOUT_CYC_SHADOWED_OFFSET = 11'h4e8;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_ACCUM_CNT_OFFSET = 11'h518;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_ACCUM_THRESH_SHADOWED_OFFSET = 11'h51c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_CLR_REGWEN_OFFSET = 11'h510;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_CLR_SHADOWED_OFFSET = 11'h514;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_CRASHDUMP_TRIGGER_SHADOWED_OFFSET = 11'h524;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_CTRL_SHADOWED_OFFSET = 11'h50c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_ESC_CNT_OFFSET = 11'h538;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_PHASE0_CYC_SHADOWED_OFFSET = 11'h528;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_PHASE1_CYC_SHADOWED_OFFSET = 11'h52c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_PHASE2_CYC_SHADOWED_OFFSET = 11'h530;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_PHASE3_CYC_SHADOWED_OFFSET = 11'h534;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_REGWEN_OFFSET = 11'h508;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_STATE_OFFSET = 11'h53c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_TIMEOUT_CYC_SHADOWED_OFFSET = 11'h520;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_ACCUM_CNT_OFFSET = 11'h550;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_ACCUM_THRESH_SHADOWED_OFFSET = 11'h554;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_CLR_REGWEN_OFFSET = 11'h548;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_CLR_SHADOWED_OFFSET = 11'h54c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_CRASHDUMP_TRIGGER_SHADOWED_OFFSET = 11'h55c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_CTRL_SHADOWED_OFFSET = 11'h544;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_ESC_CNT_OFFSET = 11'h570;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_PHASE0_CYC_SHADOWED_OFFSET = 11'h560;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_PHASE1_CYC_SHADOWED_OFFSET = 11'h564;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_PHASE2_CYC_SHADOWED_OFFSET = 11'h568;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_PHASE3_CYC_SHADOWED_OFFSET = 11'h56c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_REGWEN_OFFSET = 11'h540;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_STATE_OFFSET = 11'h574;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_TIMEOUT_CYC_SHADOWED_OFFSET = 11'h558;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_INTR_ENABLE_OFFSET = 11'h004;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_INTR_STATE_OFFSET = 11'h000;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_INTR_TEST_OFFSET = 11'h008;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CAUSE_0_OFFSET = 11'h47c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CAUSE_1_OFFSET = 11'h480;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CAUSE_2_OFFSET = 11'h484;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CAUSE_3_OFFSET = 11'h488;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CAUSE_4_OFFSET = 11'h48c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CAUSE_5_OFFSET = 11'h490;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CAUSE_6_OFFSET = 11'h494;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CLASS_SHADOWED_0_OFFSET = 11'h460;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CLASS_SHADOWED_1_OFFSET = 11'h464;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CLASS_SHADOWED_2_OFFSET = 11'h468;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CLASS_SHADOWED_3_OFFSET = 11'h46c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CLASS_SHADOWED_4_OFFSET = 11'h470;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CLASS_SHADOWED_5_OFFSET = 11'h474;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CLASS_SHADOWED_6_OFFSET = 11'h478;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_EN_SHADOWED_0_OFFSET = 11'h444;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_EN_SHADOWED_1_OFFSET = 11'h448;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_EN_SHADOWED_2_OFFSET = 11'h44c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_EN_SHADOWED_3_OFFSET = 11'h450;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_EN_SHADOWED_4_OFFSET = 11'h454;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_EN_SHADOWED_5_OFFSET = 11'h458;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_EN_SHADOWED_6_OFFSET = 11'h45c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_REGWEN_0_OFFSET = 11'h428;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_REGWEN_1_OFFSET = 11'h42c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_REGWEN_2_OFFSET = 11'h430;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_REGWEN_3_OFFSET = 11'h434;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_REGWEN_4_OFFSET = 11'h438;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_REGWEN_5_OFFSET = 11'h43c;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_REGWEN_6_OFFSET = 11'h440;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_PING_TIMEOUT_CYC_SHADOWED_OFFSET = 11'h010;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_PING_TIMER_EN_SHADOWED_OFFSET = 11'h014;
	localparam [10:0] alert_handler_reg_pkg_ALERT_HANDLER_PING_TIMER_REGWEN_OFFSET = 11'h00c;
	always @(*) begin
		addr_hit = 1'sb0;
		addr_hit[0] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_INTR_STATE_OFFSET;
		addr_hit[1] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_INTR_ENABLE_OFFSET;
		addr_hit[2] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_INTR_TEST_OFFSET;
		addr_hit[3] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_PING_TIMER_REGWEN_OFFSET;
		addr_hit[4] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_PING_TIMEOUT_CYC_SHADOWED_OFFSET;
		addr_hit[5] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_PING_TIMER_EN_SHADOWED_OFFSET;
		addr_hit[6] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_0_OFFSET;
		addr_hit[7] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_1_OFFSET;
		addr_hit[8] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_2_OFFSET;
		addr_hit[9] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_3_OFFSET;
		addr_hit[10] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_4_OFFSET;
		addr_hit[11] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_5_OFFSET;
		addr_hit[12] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_6_OFFSET;
		addr_hit[13] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_7_OFFSET;
		addr_hit[14] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_8_OFFSET;
		addr_hit[15] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_9_OFFSET;
		addr_hit[16] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_10_OFFSET;
		addr_hit[17] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_11_OFFSET;
		addr_hit[18] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_12_OFFSET;
		addr_hit[19] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_13_OFFSET;
		addr_hit[20] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_14_OFFSET;
		addr_hit[21] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_15_OFFSET;
		addr_hit[22] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_16_OFFSET;
		addr_hit[23] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_17_OFFSET;
		addr_hit[24] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_18_OFFSET;
		addr_hit[25] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_19_OFFSET;
		addr_hit[26] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_20_OFFSET;
		addr_hit[27] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_21_OFFSET;
		addr_hit[28] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_22_OFFSET;
		addr_hit[29] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_23_OFFSET;
		addr_hit[30] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_24_OFFSET;
		addr_hit[31] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_25_OFFSET;
		addr_hit[32] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_26_OFFSET;
		addr_hit[33] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_27_OFFSET;
		addr_hit[34] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_28_OFFSET;
		addr_hit[35] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_29_OFFSET;
		addr_hit[36] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_30_OFFSET;
		addr_hit[37] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_31_OFFSET;
		addr_hit[38] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_32_OFFSET;
		addr_hit[39] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_33_OFFSET;
		addr_hit[40] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_34_OFFSET;
		addr_hit[41] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_35_OFFSET;
		addr_hit[42] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_36_OFFSET;
		addr_hit[43] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_37_OFFSET;
		addr_hit[44] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_38_OFFSET;
		addr_hit[45] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_39_OFFSET;
		addr_hit[46] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_40_OFFSET;
		addr_hit[47] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_41_OFFSET;
		addr_hit[48] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_42_OFFSET;
		addr_hit[49] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_43_OFFSET;
		addr_hit[50] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_44_OFFSET;
		addr_hit[51] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_45_OFFSET;
		addr_hit[52] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_46_OFFSET;
		addr_hit[53] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_47_OFFSET;
		addr_hit[54] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_48_OFFSET;
		addr_hit[55] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_49_OFFSET;
		addr_hit[56] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_50_OFFSET;
		addr_hit[57] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_51_OFFSET;
		addr_hit[58] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_52_OFFSET;
		addr_hit[59] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_53_OFFSET;
		addr_hit[60] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_54_OFFSET;
		addr_hit[61] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_55_OFFSET;
		addr_hit[62] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_56_OFFSET;
		addr_hit[63] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_57_OFFSET;
		addr_hit[64] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_58_OFFSET;
		addr_hit[65] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_59_OFFSET;
		addr_hit[66] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_60_OFFSET;
		addr_hit[67] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_61_OFFSET;
		addr_hit[68] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_62_OFFSET;
		addr_hit[69] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_63_OFFSET;
		addr_hit[70] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_REGWEN_64_OFFSET;
		addr_hit[71] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_0_OFFSET;
		addr_hit[72] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_1_OFFSET;
		addr_hit[73] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_2_OFFSET;
		addr_hit[74] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_3_OFFSET;
		addr_hit[75] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_4_OFFSET;
		addr_hit[76] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_5_OFFSET;
		addr_hit[77] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_6_OFFSET;
		addr_hit[78] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_7_OFFSET;
		addr_hit[79] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_8_OFFSET;
		addr_hit[80] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_9_OFFSET;
		addr_hit[81] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_10_OFFSET;
		addr_hit[82] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_11_OFFSET;
		addr_hit[83] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_12_OFFSET;
		addr_hit[84] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_13_OFFSET;
		addr_hit[85] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_14_OFFSET;
		addr_hit[86] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_15_OFFSET;
		addr_hit[87] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_16_OFFSET;
		addr_hit[88] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_17_OFFSET;
		addr_hit[89] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_18_OFFSET;
		addr_hit[90] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_19_OFFSET;
		addr_hit[91] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_20_OFFSET;
		addr_hit[92] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_21_OFFSET;
		addr_hit[93] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_22_OFFSET;
		addr_hit[94] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_23_OFFSET;
		addr_hit[95] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_24_OFFSET;
		addr_hit[96] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_25_OFFSET;
		addr_hit[97] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_26_OFFSET;
		addr_hit[98] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_27_OFFSET;
		addr_hit[99] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_28_OFFSET;
		addr_hit[100] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_29_OFFSET;
		addr_hit[101] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_30_OFFSET;
		addr_hit[102] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_31_OFFSET;
		addr_hit[103] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_32_OFFSET;
		addr_hit[104] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_33_OFFSET;
		addr_hit[105] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_34_OFFSET;
		addr_hit[106] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_35_OFFSET;
		addr_hit[107] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_36_OFFSET;
		addr_hit[108] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_37_OFFSET;
		addr_hit[109] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_38_OFFSET;
		addr_hit[110] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_39_OFFSET;
		addr_hit[111] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_40_OFFSET;
		addr_hit[112] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_41_OFFSET;
		addr_hit[113] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_42_OFFSET;
		addr_hit[114] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_43_OFFSET;
		addr_hit[115] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_44_OFFSET;
		addr_hit[116] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_45_OFFSET;
		addr_hit[117] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_46_OFFSET;
		addr_hit[118] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_47_OFFSET;
		addr_hit[119] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_48_OFFSET;
		addr_hit[120] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_49_OFFSET;
		addr_hit[121] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_50_OFFSET;
		addr_hit[122] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_51_OFFSET;
		addr_hit[123] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_52_OFFSET;
		addr_hit[124] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_53_OFFSET;
		addr_hit[125] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_54_OFFSET;
		addr_hit[126] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_55_OFFSET;
		addr_hit[127] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_56_OFFSET;
		addr_hit[128] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_57_OFFSET;
		addr_hit[129] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_58_OFFSET;
		addr_hit[130] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_59_OFFSET;
		addr_hit[131] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_60_OFFSET;
		addr_hit[132] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_61_OFFSET;
		addr_hit[133] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_62_OFFSET;
		addr_hit[134] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_63_OFFSET;
		addr_hit[135] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_EN_SHADOWED_64_OFFSET;
		addr_hit[136] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_0_OFFSET;
		addr_hit[137] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_1_OFFSET;
		addr_hit[138] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_2_OFFSET;
		addr_hit[139] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_3_OFFSET;
		addr_hit[140] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_4_OFFSET;
		addr_hit[141] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_5_OFFSET;
		addr_hit[142] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_6_OFFSET;
		addr_hit[143] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_7_OFFSET;
		addr_hit[144] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_8_OFFSET;
		addr_hit[145] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_9_OFFSET;
		addr_hit[146] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_10_OFFSET;
		addr_hit[147] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_11_OFFSET;
		addr_hit[148] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_12_OFFSET;
		addr_hit[149] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_13_OFFSET;
		addr_hit[150] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_14_OFFSET;
		addr_hit[151] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_15_OFFSET;
		addr_hit[152] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_16_OFFSET;
		addr_hit[153] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_17_OFFSET;
		addr_hit[154] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_18_OFFSET;
		addr_hit[155] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_19_OFFSET;
		addr_hit[156] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_20_OFFSET;
		addr_hit[157] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_21_OFFSET;
		addr_hit[158] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_22_OFFSET;
		addr_hit[159] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_23_OFFSET;
		addr_hit[160] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_24_OFFSET;
		addr_hit[161] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_25_OFFSET;
		addr_hit[162] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_26_OFFSET;
		addr_hit[163] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_27_OFFSET;
		addr_hit[164] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_28_OFFSET;
		addr_hit[165] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_29_OFFSET;
		addr_hit[166] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_30_OFFSET;
		addr_hit[167] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_31_OFFSET;
		addr_hit[168] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_32_OFFSET;
		addr_hit[169] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_33_OFFSET;
		addr_hit[170] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_34_OFFSET;
		addr_hit[171] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_35_OFFSET;
		addr_hit[172] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_36_OFFSET;
		addr_hit[173] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_37_OFFSET;
		addr_hit[174] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_38_OFFSET;
		addr_hit[175] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_39_OFFSET;
		addr_hit[176] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_40_OFFSET;
		addr_hit[177] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_41_OFFSET;
		addr_hit[178] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_42_OFFSET;
		addr_hit[179] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_43_OFFSET;
		addr_hit[180] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_44_OFFSET;
		addr_hit[181] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_45_OFFSET;
		addr_hit[182] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_46_OFFSET;
		addr_hit[183] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_47_OFFSET;
		addr_hit[184] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_48_OFFSET;
		addr_hit[185] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_49_OFFSET;
		addr_hit[186] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_50_OFFSET;
		addr_hit[187] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_51_OFFSET;
		addr_hit[188] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_52_OFFSET;
		addr_hit[189] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_53_OFFSET;
		addr_hit[190] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_54_OFFSET;
		addr_hit[191] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_55_OFFSET;
		addr_hit[192] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_56_OFFSET;
		addr_hit[193] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_57_OFFSET;
		addr_hit[194] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_58_OFFSET;
		addr_hit[195] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_59_OFFSET;
		addr_hit[196] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_60_OFFSET;
		addr_hit[197] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_61_OFFSET;
		addr_hit[198] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_62_OFFSET;
		addr_hit[199] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_63_OFFSET;
		addr_hit[200] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CLASS_SHADOWED_64_OFFSET;
		addr_hit[201] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_0_OFFSET;
		addr_hit[202] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_1_OFFSET;
		addr_hit[203] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_2_OFFSET;
		addr_hit[204] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_3_OFFSET;
		addr_hit[205] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_4_OFFSET;
		addr_hit[206] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_5_OFFSET;
		addr_hit[207] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_6_OFFSET;
		addr_hit[208] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_7_OFFSET;
		addr_hit[209] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_8_OFFSET;
		addr_hit[210] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_9_OFFSET;
		addr_hit[211] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_10_OFFSET;
		addr_hit[212] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_11_OFFSET;
		addr_hit[213] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_12_OFFSET;
		addr_hit[214] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_13_OFFSET;
		addr_hit[215] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_14_OFFSET;
		addr_hit[216] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_15_OFFSET;
		addr_hit[217] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_16_OFFSET;
		addr_hit[218] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_17_OFFSET;
		addr_hit[219] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_18_OFFSET;
		addr_hit[220] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_19_OFFSET;
		addr_hit[221] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_20_OFFSET;
		addr_hit[222] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_21_OFFSET;
		addr_hit[223] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_22_OFFSET;
		addr_hit[224] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_23_OFFSET;
		addr_hit[225] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_24_OFFSET;
		addr_hit[226] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_25_OFFSET;
		addr_hit[227] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_26_OFFSET;
		addr_hit[228] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_27_OFFSET;
		addr_hit[229] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_28_OFFSET;
		addr_hit[230] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_29_OFFSET;
		addr_hit[231] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_30_OFFSET;
		addr_hit[232] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_31_OFFSET;
		addr_hit[233] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_32_OFFSET;
		addr_hit[234] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_33_OFFSET;
		addr_hit[235] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_34_OFFSET;
		addr_hit[236] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_35_OFFSET;
		addr_hit[237] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_36_OFFSET;
		addr_hit[238] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_37_OFFSET;
		addr_hit[239] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_38_OFFSET;
		addr_hit[240] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_39_OFFSET;
		addr_hit[241] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_40_OFFSET;
		addr_hit[242] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_41_OFFSET;
		addr_hit[243] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_42_OFFSET;
		addr_hit[244] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_43_OFFSET;
		addr_hit[245] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_44_OFFSET;
		addr_hit[246] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_45_OFFSET;
		addr_hit[247] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_46_OFFSET;
		addr_hit[248] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_47_OFFSET;
		addr_hit[249] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_48_OFFSET;
		addr_hit[250] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_49_OFFSET;
		addr_hit[251] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_50_OFFSET;
		addr_hit[252] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_51_OFFSET;
		addr_hit[253] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_52_OFFSET;
		addr_hit[254] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_53_OFFSET;
		addr_hit[255] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_54_OFFSET;
		addr_hit[256] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_55_OFFSET;
		addr_hit[257] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_56_OFFSET;
		addr_hit[258] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_57_OFFSET;
		addr_hit[259] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_58_OFFSET;
		addr_hit[260] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_59_OFFSET;
		addr_hit[261] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_60_OFFSET;
		addr_hit[262] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_61_OFFSET;
		addr_hit[263] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_62_OFFSET;
		addr_hit[264] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_63_OFFSET;
		addr_hit[265] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_ALERT_CAUSE_64_OFFSET;
		addr_hit[266] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_REGWEN_0_OFFSET;
		addr_hit[267] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_REGWEN_1_OFFSET;
		addr_hit[268] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_REGWEN_2_OFFSET;
		addr_hit[269] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_REGWEN_3_OFFSET;
		addr_hit[270] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_REGWEN_4_OFFSET;
		addr_hit[271] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_REGWEN_5_OFFSET;
		addr_hit[272] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_REGWEN_6_OFFSET;
		addr_hit[273] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_EN_SHADOWED_0_OFFSET;
		addr_hit[274] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_EN_SHADOWED_1_OFFSET;
		addr_hit[275] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_EN_SHADOWED_2_OFFSET;
		addr_hit[276] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_EN_SHADOWED_3_OFFSET;
		addr_hit[277] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_EN_SHADOWED_4_OFFSET;
		addr_hit[278] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_EN_SHADOWED_5_OFFSET;
		addr_hit[279] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_EN_SHADOWED_6_OFFSET;
		addr_hit[280] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CLASS_SHADOWED_0_OFFSET;
		addr_hit[281] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CLASS_SHADOWED_1_OFFSET;
		addr_hit[282] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CLASS_SHADOWED_2_OFFSET;
		addr_hit[283] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CLASS_SHADOWED_3_OFFSET;
		addr_hit[284] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CLASS_SHADOWED_4_OFFSET;
		addr_hit[285] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CLASS_SHADOWED_5_OFFSET;
		addr_hit[286] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CLASS_SHADOWED_6_OFFSET;
		addr_hit[287] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CAUSE_0_OFFSET;
		addr_hit[288] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CAUSE_1_OFFSET;
		addr_hit[289] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CAUSE_2_OFFSET;
		addr_hit[290] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CAUSE_3_OFFSET;
		addr_hit[291] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CAUSE_4_OFFSET;
		addr_hit[292] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CAUSE_5_OFFSET;
		addr_hit[293] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_LOC_ALERT_CAUSE_6_OFFSET;
		addr_hit[294] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_REGWEN_OFFSET;
		addr_hit[295] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_CTRL_SHADOWED_OFFSET;
		addr_hit[296] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_CLR_REGWEN_OFFSET;
		addr_hit[297] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_CLR_SHADOWED_OFFSET;
		addr_hit[298] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_ACCUM_CNT_OFFSET;
		addr_hit[299] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_ACCUM_THRESH_SHADOWED_OFFSET;
		addr_hit[300] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_TIMEOUT_CYC_SHADOWED_OFFSET;
		addr_hit[301] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_CRASHDUMP_TRIGGER_SHADOWED_OFFSET;
		addr_hit[302] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_PHASE0_CYC_SHADOWED_OFFSET;
		addr_hit[303] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_PHASE1_CYC_SHADOWED_OFFSET;
		addr_hit[304] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_PHASE2_CYC_SHADOWED_OFFSET;
		addr_hit[305] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_PHASE3_CYC_SHADOWED_OFFSET;
		addr_hit[306] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_ESC_CNT_OFFSET;
		addr_hit[307] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSA_STATE_OFFSET;
		addr_hit[308] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_REGWEN_OFFSET;
		addr_hit[309] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_CTRL_SHADOWED_OFFSET;
		addr_hit[310] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_CLR_REGWEN_OFFSET;
		addr_hit[311] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_CLR_SHADOWED_OFFSET;
		addr_hit[312] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_ACCUM_CNT_OFFSET;
		addr_hit[313] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_ACCUM_THRESH_SHADOWED_OFFSET;
		addr_hit[314] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_TIMEOUT_CYC_SHADOWED_OFFSET;
		addr_hit[315] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_CRASHDUMP_TRIGGER_SHADOWED_OFFSET;
		addr_hit[316] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_PHASE0_CYC_SHADOWED_OFFSET;
		addr_hit[317] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_PHASE1_CYC_SHADOWED_OFFSET;
		addr_hit[318] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_PHASE2_CYC_SHADOWED_OFFSET;
		addr_hit[319] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_PHASE3_CYC_SHADOWED_OFFSET;
		addr_hit[320] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_ESC_CNT_OFFSET;
		addr_hit[321] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSB_STATE_OFFSET;
		addr_hit[322] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_REGWEN_OFFSET;
		addr_hit[323] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_CTRL_SHADOWED_OFFSET;
		addr_hit[324] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_CLR_REGWEN_OFFSET;
		addr_hit[325] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_CLR_SHADOWED_OFFSET;
		addr_hit[326] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_ACCUM_CNT_OFFSET;
		addr_hit[327] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_ACCUM_THRESH_SHADOWED_OFFSET;
		addr_hit[328] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_TIMEOUT_CYC_SHADOWED_OFFSET;
		addr_hit[329] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_CRASHDUMP_TRIGGER_SHADOWED_OFFSET;
		addr_hit[330] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_PHASE0_CYC_SHADOWED_OFFSET;
		addr_hit[331] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_PHASE1_CYC_SHADOWED_OFFSET;
		addr_hit[332] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_PHASE2_CYC_SHADOWED_OFFSET;
		addr_hit[333] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_PHASE3_CYC_SHADOWED_OFFSET;
		addr_hit[334] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_ESC_CNT_OFFSET;
		addr_hit[335] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSC_STATE_OFFSET;
		addr_hit[336] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_REGWEN_OFFSET;
		addr_hit[337] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_CTRL_SHADOWED_OFFSET;
		addr_hit[338] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_CLR_REGWEN_OFFSET;
		addr_hit[339] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_CLR_SHADOWED_OFFSET;
		addr_hit[340] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_ACCUM_CNT_OFFSET;
		addr_hit[341] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_ACCUM_THRESH_SHADOWED_OFFSET;
		addr_hit[342] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_TIMEOUT_CYC_SHADOWED_OFFSET;
		addr_hit[343] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_CRASHDUMP_TRIGGER_SHADOWED_OFFSET;
		addr_hit[344] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_PHASE0_CYC_SHADOWED_OFFSET;
		addr_hit[345] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_PHASE1_CYC_SHADOWED_OFFSET;
		addr_hit[346] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_PHASE2_CYC_SHADOWED_OFFSET;
		addr_hit[347] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_PHASE3_CYC_SHADOWED_OFFSET;
		addr_hit[348] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_ESC_CNT_OFFSET;
		addr_hit[349] = reg_addr == alert_handler_reg_pkg_ALERT_HANDLER_CLASSD_STATE_OFFSET;
	end
	assign addrmiss = (reg_re || reg_we ? ~|addr_hit : 1'b0);
	localparam [1399:0] alert_handler_reg_pkg_ALERT_HANDLER_PERMIT = 1400'b10001000100010011000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010011000100010011001111110001111111111111111111110001000100110001000100110011111100011111111111111111111100010001001100010001001100111111000111111111111111111111000100010011000100010011001111110001111111111111111111110001;
	always @(*) wr_err = reg_we & ((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((addr_hit[0] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1396+:4] & ~reg_be)) | (addr_hit[1] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1392+:4] & ~reg_be))) | (addr_hit[2] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1388+:4] & ~reg_be))) | (addr_hit[3] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1384+:4] & ~reg_be))) | (addr_hit[4] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1380+:4] & ~reg_be))) | (addr_hit[5] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1376+:4] & ~reg_be))) | (addr_hit[6] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1372+:4] & ~reg_be))) | (addr_hit[7] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1368+:4] & ~reg_be))) | (addr_hit[8] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1364+:4] & ~reg_be))) | (addr_hit[9] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1360+:4] & ~reg_be))) | (addr_hit[10] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1356+:4] & ~reg_be))) | (addr_hit[11] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1352+:4] & ~reg_be))) | (addr_hit[12] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1348+:4] & ~reg_be))) | (addr_hit[13] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1344+:4] & ~reg_be))) | (addr_hit[14] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1340+:4] & ~reg_be))) | (addr_hit[15] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1336+:4] & ~reg_be))) | (addr_hit[16] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1332+:4] & ~reg_be))) | (addr_hit[17] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1328+:4] & ~reg_be))) | (addr_hit[18] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1324+:4] & ~reg_be))) | (addr_hit[19] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1320+:4] & ~reg_be))) | (addr_hit[20] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1316+:4] & ~reg_be))) | (addr_hit[21] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1312+:4] & ~reg_be))) | (addr_hit[22] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1308+:4] & ~reg_be))) | (addr_hit[23] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1304+:4] & ~reg_be))) | (addr_hit[24] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1300+:4] & ~reg_be))) | (addr_hit[25] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1296+:4] & ~reg_be))) | (addr_hit[26] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1292+:4] & ~reg_be))) | (addr_hit[27] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1288+:4] & ~reg_be))) | (addr_hit[28] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1284+:4] & ~reg_be))) | (addr_hit[29] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1280+:4] & ~reg_be))) | (addr_hit[30] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1276+:4] & ~reg_be))) | (addr_hit[31] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1272+:4] & ~reg_be))) | (addr_hit[32] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1268+:4] & ~reg_be))) | (addr_hit[33] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1264+:4] & ~reg_be))) | (addr_hit[34] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1260+:4] & ~reg_be))) | (addr_hit[35] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1256+:4] & ~reg_be))) | (addr_hit[36] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1252+:4] & ~reg_be))) | (addr_hit[37] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1248+:4] & ~reg_be))) | (addr_hit[38] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1244+:4] & ~reg_be))) | (addr_hit[39] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1240+:4] & ~reg_be))) | (addr_hit[40] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1236+:4] & ~reg_be))) | (addr_hit[41] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1232+:4] & ~reg_be))) | (addr_hit[42] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1228+:4] & ~reg_be))) | (addr_hit[43] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1224+:4] & ~reg_be))) | (addr_hit[44] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1220+:4] & ~reg_be))) | (addr_hit[45] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1216+:4] & ~reg_be))) | (addr_hit[46] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1212+:4] & ~reg_be))) | (addr_hit[47] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1208+:4] & ~reg_be))) | (addr_hit[48] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1204+:4] & ~reg_be))) | (addr_hit[49] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1200+:4] & ~reg_be))) | (addr_hit[50] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1196+:4] & ~reg_be))) | (addr_hit[51] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1192+:4] & ~reg_be))) | (addr_hit[52] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1188+:4] & ~reg_be))) | (addr_hit[53] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1184+:4] & ~reg_be))) | (addr_hit[54] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1180+:4] & ~reg_be))) | (addr_hit[55] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1176+:4] & ~reg_be))) | (addr_hit[56] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1172+:4] & ~reg_be))) | (addr_hit[57] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1168+:4] & ~reg_be))) | (addr_hit[58] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1164+:4] & ~reg_be))) | (addr_hit[59] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1160+:4] & ~reg_be))) | (addr_hit[60] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1156+:4] & ~reg_be))) | (addr_hit[61] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1152+:4] & ~reg_be))) | (addr_hit[62] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1148+:4] & ~reg_be))) | (addr_hit[63] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1144+:4] & ~reg_be))) | (addr_hit[64] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1140+:4] & ~reg_be))) | (addr_hit[65] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1136+:4] & ~reg_be))) | (addr_hit[66] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1132+:4] & ~reg_be))) | (addr_hit[67] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1128+:4] & ~reg_be))) | (addr_hit[68] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1124+:4] & ~reg_be))) | (addr_hit[69] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1120+:4] & ~reg_be))) | (addr_hit[70] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1116+:4] & ~reg_be))) | (addr_hit[71] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1112+:4] & ~reg_be))) | (addr_hit[72] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1108+:4] & ~reg_be))) | (addr_hit[73] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1104+:4] & ~reg_be))) | (addr_hit[74] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1100+:4] & ~reg_be))) | (addr_hit[75] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1096+:4] & ~reg_be))) | (addr_hit[76] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1092+:4] & ~reg_be))) | (addr_hit[77] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1088+:4] & ~reg_be))) | (addr_hit[78] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1084+:4] & ~reg_be))) | (addr_hit[79] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1080+:4] & ~reg_be))) | (addr_hit[80] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1076+:4] & ~reg_be))) | (addr_hit[81] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1072+:4] & ~reg_be))) | (addr_hit[82] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1068+:4] & ~reg_be))) | (addr_hit[83] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1064+:4] & ~reg_be))) | (addr_hit[84] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1060+:4] & ~reg_be))) | (addr_hit[85] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1056+:4] & ~reg_be))) | (addr_hit[86] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1052+:4] & ~reg_be))) | (addr_hit[87] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1048+:4] & ~reg_be))) | (addr_hit[88] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1044+:4] & ~reg_be))) | (addr_hit[89] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1040+:4] & ~reg_be))) | (addr_hit[90] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1036+:4] & ~reg_be))) | (addr_hit[91] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1032+:4] & ~reg_be))) | (addr_hit[92] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1028+:4] & ~reg_be))) | (addr_hit[93] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1024+:4] & ~reg_be))) | (addr_hit[94] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1020+:4] & ~reg_be))) | (addr_hit[95] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1016+:4] & ~reg_be))) | (addr_hit[96] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1012+:4] & ~reg_be))) | (addr_hit[97] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1008+:4] & ~reg_be))) | (addr_hit[98] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1004+:4] & ~reg_be))) | (addr_hit[99] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[1000+:4] & ~reg_be))) | (addr_hit[100] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[996+:4] & ~reg_be))) | (addr_hit[101] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[992+:4] & ~reg_be))) | (addr_hit[102] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[988+:4] & ~reg_be))) | (addr_hit[103] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[984+:4] & ~reg_be))) | (addr_hit[104] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[980+:4] & ~reg_be))) | (addr_hit[105] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[976+:4] & ~reg_be))) | (addr_hit[106] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[972+:4] & ~reg_be))) | (addr_hit[107] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[968+:4] & ~reg_be))) | (addr_hit[108] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[964+:4] & ~reg_be))) | (addr_hit[109] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[960+:4] & ~reg_be))) | (addr_hit[110] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[956+:4] & ~reg_be))) | (addr_hit[111] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[952+:4] & ~reg_be))) | (addr_hit[112] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[948+:4] & ~reg_be))) | (addr_hit[113] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[944+:4] & ~reg_be))) | (addr_hit[114] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[940+:4] & ~reg_be))) | (addr_hit[115] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[936+:4] & ~reg_be))) | (addr_hit[116] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[932+:4] & ~reg_be))) | (addr_hit[117] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[928+:4] & ~reg_be))) | (addr_hit[118] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[924+:4] & ~reg_be))) | (addr_hit[119] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[920+:4] & ~reg_be))) | (addr_hit[120] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[916+:4] & ~reg_be))) | (addr_hit[121] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[912+:4] & ~reg_be))) | (addr_hit[122] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[908+:4] & ~reg_be))) | (addr_hit[123] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[904+:4] & ~reg_be))) | (addr_hit[124] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[900+:4] & ~reg_be))) | (addr_hit[125] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[896+:4] & ~reg_be))) | (addr_hit[126] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[892+:4] & ~reg_be))) | (addr_hit[127] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[888+:4] & ~reg_be))) | (addr_hit[128] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[884+:4] & ~reg_be))) | (addr_hit[129] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[880+:4] & ~reg_be))) | (addr_hit[130] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[876+:4] & ~reg_be))) | (addr_hit[131] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[872+:4] & ~reg_be))) | (addr_hit[132] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[868+:4] & ~reg_be))) | (addr_hit[133] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[864+:4] & ~reg_be))) | (addr_hit[134] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[860+:4] & ~reg_be))) | (addr_hit[135] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[856+:4] & ~reg_be))) | (addr_hit[136] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[852+:4] & ~reg_be))) | (addr_hit[137] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[848+:4] & ~reg_be))) | (addr_hit[138] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[844+:4] & ~reg_be))) | (addr_hit[139] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[840+:4] & ~reg_be))) | (addr_hit[140] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[836+:4] & ~reg_be))) | (addr_hit[141] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[832+:4] & ~reg_be))) | (addr_hit[142] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[828+:4] & ~reg_be))) | (addr_hit[143] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[824+:4] & ~reg_be))) | (addr_hit[144] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[820+:4] & ~reg_be))) | (addr_hit[145] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[816+:4] & ~reg_be))) | (addr_hit[146] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[812+:4] & ~reg_be))) | (addr_hit[147] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[808+:4] & ~reg_be))) | (addr_hit[148] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[804+:4] & ~reg_be))) | (addr_hit[149] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[800+:4] & ~reg_be))) | (addr_hit[150] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[796+:4] & ~reg_be))) | (addr_hit[151] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[792+:4] & ~reg_be))) | (addr_hit[152] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[788+:4] & ~reg_be))) | (addr_hit[153] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[784+:4] & ~reg_be))) | (addr_hit[154] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[780+:4] & ~reg_be))) | (addr_hit[155] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[776+:4] & ~reg_be))) | (addr_hit[156] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[772+:4] & ~reg_be))) | (addr_hit[157] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[768+:4] & ~reg_be))) | (addr_hit[158] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[764+:4] & ~reg_be))) | (addr_hit[159] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[760+:4] & ~reg_be))) | (addr_hit[160] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[756+:4] & ~reg_be))) | (addr_hit[161] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[752+:4] & ~reg_be))) | (addr_hit[162] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[748+:4] & ~reg_be))) | (addr_hit[163] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[744+:4] & ~reg_be))) | (addr_hit[164] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[740+:4] & ~reg_be))) | (addr_hit[165] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[736+:4] & ~reg_be))) | (addr_hit[166] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[732+:4] & ~reg_be))) | (addr_hit[167] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[728+:4] & ~reg_be))) | (addr_hit[168] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[724+:4] & ~reg_be))) | (addr_hit[169] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[720+:4] & ~reg_be))) | (addr_hit[170] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[716+:4] & ~reg_be))) | (addr_hit[171] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[712+:4] & ~reg_be))) | (addr_hit[172] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[708+:4] & ~reg_be))) | (addr_hit[173] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[704+:4] & ~reg_be))) | (addr_hit[174] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[700+:4] & ~reg_be))) | (addr_hit[175] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[696+:4] & ~reg_be))) | (addr_hit[176] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[692+:4] & ~reg_be))) | (addr_hit[177] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[688+:4] & ~reg_be))) | (addr_hit[178] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[684+:4] & ~reg_be))) | (addr_hit[179] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[680+:4] & ~reg_be))) | (addr_hit[180] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[676+:4] & ~reg_be))) | (addr_hit[181] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[672+:4] & ~reg_be))) | (addr_hit[182] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[668+:4] & ~reg_be))) | (addr_hit[183] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[664+:4] & ~reg_be))) | (addr_hit[184] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[660+:4] & ~reg_be))) | (addr_hit[185] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[656+:4] & ~reg_be))) | (addr_hit[186] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[652+:4] & ~reg_be))) | (addr_hit[187] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[648+:4] & ~reg_be))) | (addr_hit[188] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[644+:4] & ~reg_be))) | (addr_hit[189] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[640+:4] & ~reg_be))) | (addr_hit[190] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[636+:4] & ~reg_be))) | (addr_hit[191] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[632+:4] & ~reg_be))) | (addr_hit[192] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[628+:4] & ~reg_be))) | (addr_hit[193] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[624+:4] & ~reg_be))) | (addr_hit[194] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[620+:4] & ~reg_be))) | (addr_hit[195] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[616+:4] & ~reg_be))) | (addr_hit[196] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[612+:4] & ~reg_be))) | (addr_hit[197] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[608+:4] & ~reg_be))) | (addr_hit[198] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[604+:4] & ~reg_be))) | (addr_hit[199] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[600+:4] & ~reg_be))) | (addr_hit[200] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[596+:4] & ~reg_be))) | (addr_hit[201] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[592+:4] & ~reg_be))) | (addr_hit[202] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[588+:4] & ~reg_be))) | (addr_hit[203] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[584+:4] & ~reg_be))) | (addr_hit[204] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[580+:4] & ~reg_be))) | (addr_hit[205] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[576+:4] & ~reg_be))) | (addr_hit[206] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[572+:4] & ~reg_be))) | (addr_hit[207] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[568+:4] & ~reg_be))) | (addr_hit[208] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[564+:4] & ~reg_be))) | (addr_hit[209] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[560+:4] & ~reg_be))) | (addr_hit[210] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[556+:4] & ~reg_be))) | (addr_hit[211] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[552+:4] & ~reg_be))) | (addr_hit[212] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[548+:4] & ~reg_be))) | (addr_hit[213] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[544+:4] & ~reg_be))) | (addr_hit[214] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[540+:4] & ~reg_be))) | (addr_hit[215] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[536+:4] & ~reg_be))) | (addr_hit[216] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[532+:4] & ~reg_be))) | (addr_hit[217] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[528+:4] & ~reg_be))) | (addr_hit[218] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[524+:4] & ~reg_be))) | (addr_hit[219] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[520+:4] & ~reg_be))) | (addr_hit[220] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[516+:4] & ~reg_be))) | (addr_hit[221] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[512+:4] & ~reg_be))) | (addr_hit[222] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[508+:4] & ~reg_be))) | (addr_hit[223] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[504+:4] & ~reg_be))) | (addr_hit[224] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[500+:4] & ~reg_be))) | (addr_hit[225] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[496+:4] & ~reg_be))) | (addr_hit[226] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[492+:4] & ~reg_be))) | (addr_hit[227] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[488+:4] & ~reg_be))) | (addr_hit[228] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[484+:4] & ~reg_be))) | (addr_hit[229] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[480+:4] & ~reg_be))) | (addr_hit[230] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[476+:4] & ~reg_be))) | (addr_hit[231] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[472+:4] & ~reg_be))) | (addr_hit[232] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[468+:4] & ~reg_be))) | (addr_hit[233] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[464+:4] & ~reg_be))) | (addr_hit[234] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[460+:4] & ~reg_be))) | (addr_hit[235] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[456+:4] & ~reg_be))) | (addr_hit[236] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[452+:4] & ~reg_be))) | (addr_hit[237] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[448+:4] & ~reg_be))) | (addr_hit[238] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[444+:4] & ~reg_be))) | (addr_hit[239] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[440+:4] & ~reg_be))) | (addr_hit[240] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[436+:4] & ~reg_be))) | (addr_hit[241] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[432+:4] & ~reg_be))) | (addr_hit[242] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[428+:4] & ~reg_be))) | (addr_hit[243] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[424+:4] & ~reg_be))) | (addr_hit[244] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[420+:4] & ~reg_be))) | (addr_hit[245] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[416+:4] & ~reg_be))) | (addr_hit[246] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[412+:4] & ~reg_be))) | (addr_hit[247] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[408+:4] & ~reg_be))) | (addr_hit[248] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[404+:4] & ~reg_be))) | (addr_hit[249] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[400+:4] & ~reg_be))) | (addr_hit[250] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[396+:4] & ~reg_be))) | (addr_hit[251] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[392+:4] & ~reg_be))) | (addr_hit[252] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[388+:4] & ~reg_be))) | (addr_hit[253] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[384+:4] & ~reg_be))) | (addr_hit[254] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[380+:4] & ~reg_be))) | (addr_hit[255] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[376+:4] & ~reg_be))) | (addr_hit[256] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[372+:4] & ~reg_be))) | (addr_hit[257] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[368+:4] & ~reg_be))) | (addr_hit[258] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[364+:4] & ~reg_be))) | (addr_hit[259] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[360+:4] & ~reg_be))) | (addr_hit[260] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[356+:4] & ~reg_be))) | (addr_hit[261] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[352+:4] & ~reg_be))) | (addr_hit[262] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[348+:4] & ~reg_be))) | (addr_hit[263] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[344+:4] & ~reg_be))) | (addr_hit[264] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[340+:4] & ~reg_be))) | (addr_hit[265] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[336+:4] & ~reg_be))) | (addr_hit[266] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[332+:4] & ~reg_be))) | (addr_hit[267] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[328+:4] & ~reg_be))) | (addr_hit[268] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[324+:4] & ~reg_be))) | (addr_hit[269] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[320+:4] & ~reg_be))) | (addr_hit[270] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[316+:4] & ~reg_be))) | (addr_hit[271] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[312+:4] & ~reg_be))) | (addr_hit[272] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[308+:4] & ~reg_be))) | (addr_hit[273] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[304+:4] & ~reg_be))) | (addr_hit[274] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[300+:4] & ~reg_be))) | (addr_hit[275] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[296+:4] & ~reg_be))) | (addr_hit[276] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[292+:4] & ~reg_be))) | (addr_hit[277] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[288+:4] & ~reg_be))) | (addr_hit[278] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[284+:4] & ~reg_be))) | (addr_hit[279] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[280+:4] & ~reg_be))) | (addr_hit[280] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[276+:4] & ~reg_be))) | (addr_hit[281] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[272+:4] & ~reg_be))) | (addr_hit[282] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[268+:4] & ~reg_be))) | (addr_hit[283] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[264+:4] & ~reg_be))) | (addr_hit[284] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[260+:4] & ~reg_be))) | (addr_hit[285] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[256+:4] & ~reg_be))) | (addr_hit[286] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[252+:4] & ~reg_be))) | (addr_hit[287] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[248+:4] & ~reg_be))) | (addr_hit[288] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[244+:4] & ~reg_be))) | (addr_hit[289] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[240+:4] & ~reg_be))) | (addr_hit[290] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[236+:4] & ~reg_be))) | (addr_hit[291] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[232+:4] & ~reg_be))) | (addr_hit[292] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[228+:4] & ~reg_be))) | (addr_hit[293] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[224+:4] & ~reg_be))) | (addr_hit[294] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[220+:4] & ~reg_be))) | (addr_hit[295] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[216+:4] & ~reg_be))) | (addr_hit[296] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[212+:4] & ~reg_be))) | (addr_hit[297] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[208+:4] & ~reg_be))) | (addr_hit[298] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[204+:4] & ~reg_be))) | (addr_hit[299] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[200+:4] & ~reg_be))) | (addr_hit[300] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[196+:4] & ~reg_be))) | (addr_hit[301] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[192+:4] & ~reg_be))) | (addr_hit[302] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[188+:4] & ~reg_be))) | (addr_hit[303] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[184+:4] & ~reg_be))) | (addr_hit[304] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[180+:4] & ~reg_be))) | (addr_hit[305] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[176+:4] & ~reg_be))) | (addr_hit[306] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[172+:4] & ~reg_be))) | (addr_hit[307] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[168+:4] & ~reg_be))) | (addr_hit[308] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[164+:4] & ~reg_be))) | (addr_hit[309] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[160+:4] & ~reg_be))) | (addr_hit[310] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[156+:4] & ~reg_be))) | (addr_hit[311] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[152+:4] & ~reg_be))) | (addr_hit[312] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[148+:4] & ~reg_be))) | (addr_hit[313] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[144+:4] & ~reg_be))) | (addr_hit[314] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[140+:4] & ~reg_be))) | (addr_hit[315] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[136+:4] & ~reg_be))) | (addr_hit[316] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[132+:4] & ~reg_be))) | (addr_hit[317] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[128+:4] & ~reg_be))) | (addr_hit[318] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[124+:4] & ~reg_be))) | (addr_hit[319] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[120+:4] & ~reg_be))) | (addr_hit[320] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[116+:4] & ~reg_be))) | (addr_hit[321] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[112+:4] & ~reg_be))) | (addr_hit[322] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[108+:4] & ~reg_be))) | (addr_hit[323] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[104+:4] & ~reg_be))) | (addr_hit[324] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[100+:4] & ~reg_be))) | (addr_hit[325] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[96+:4] & ~reg_be))) | (addr_hit[326] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[92+:4] & ~reg_be))) | (addr_hit[327] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[88+:4] & ~reg_be))) | (addr_hit[328] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[84+:4] & ~reg_be))) | (addr_hit[329] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[80+:4] & ~reg_be))) | (addr_hit[330] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[76+:4] & ~reg_be))) | (addr_hit[331] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[72+:4] & ~reg_be))) | (addr_hit[332] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[68+:4] & ~reg_be))) | (addr_hit[333] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[64+:4] & ~reg_be))) | (addr_hit[334] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[60+:4] & ~reg_be))) | (addr_hit[335] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[56+:4] & ~reg_be))) | (addr_hit[336] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[52+:4] & ~reg_be))) | (addr_hit[337] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[48+:4] & ~reg_be))) | (addr_hit[338] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[44+:4] & ~reg_be))) | (addr_hit[339] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[40+:4] & ~reg_be))) | (addr_hit[340] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[36+:4] & ~reg_be))) | (addr_hit[341] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[32+:4] & ~reg_be))) | (addr_hit[342] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[28+:4] & ~reg_be))) | (addr_hit[343] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[24+:4] & ~reg_be))) | (addr_hit[344] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[20+:4] & ~reg_be))) | (addr_hit[345] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[16+:4] & ~reg_be))) | (addr_hit[346] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[12+:4] & ~reg_be))) | (addr_hit[347] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[8+:4] & ~reg_be))) | (addr_hit[348] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[4+:4] & ~reg_be))) | (addr_hit[349] & |(alert_handler_reg_pkg_ALERT_HANDLER_PERMIT[0+:4] & ~reg_be)));
	assign intr_state_we = (addr_hit[0] & reg_we) & !reg_error;
	assign intr_state_classa_wd = reg_wdata[0];
	assign intr_state_classb_wd = reg_wdata[1];
	assign intr_state_classc_wd = reg_wdata[2];
	assign intr_state_classd_wd = reg_wdata[3];
	assign intr_enable_we = (addr_hit[1] & reg_we) & !reg_error;
	assign intr_enable_classa_wd = reg_wdata[0];
	assign intr_enable_classb_wd = reg_wdata[1];
	assign intr_enable_classc_wd = reg_wdata[2];
	assign intr_enable_classd_wd = reg_wdata[3];
	assign intr_test_we = (addr_hit[2] & reg_we) & !reg_error;
	assign intr_test_classa_wd = reg_wdata[0];
	assign intr_test_classb_wd = reg_wdata[1];
	assign intr_test_classc_wd = reg_wdata[2];
	assign intr_test_classd_wd = reg_wdata[3];
	assign ping_timer_regwen_we = (addr_hit[3] & reg_we) & !reg_error;
	assign ping_timer_regwen_wd = reg_wdata[0];
	assign ping_timeout_cyc_shadowed_re = (addr_hit[4] & reg_re) & !reg_error;
	assign ping_timeout_cyc_shadowed_we = (addr_hit[4] & reg_we) & !reg_error;
	assign ping_timeout_cyc_shadowed_wd = reg_wdata[15:0];
	assign ping_timer_en_shadowed_re = (addr_hit[5] & reg_re) & !reg_error;
	assign ping_timer_en_shadowed_we = (addr_hit[5] & reg_we) & !reg_error;
	assign ping_timer_en_shadowed_wd = reg_wdata[0];
	assign alert_regwen_0_we = (addr_hit[6] & reg_we) & !reg_error;
	assign alert_regwen_0_wd = reg_wdata[0];
	assign alert_regwen_1_we = (addr_hit[7] & reg_we) & !reg_error;
	assign alert_regwen_1_wd = reg_wdata[0];
	assign alert_regwen_2_we = (addr_hit[8] & reg_we) & !reg_error;
	assign alert_regwen_2_wd = reg_wdata[0];
	assign alert_regwen_3_we = (addr_hit[9] & reg_we) & !reg_error;
	assign alert_regwen_3_wd = reg_wdata[0];
	assign alert_regwen_4_we = (addr_hit[10] & reg_we) & !reg_error;
	assign alert_regwen_4_wd = reg_wdata[0];
	assign alert_regwen_5_we = (addr_hit[11] & reg_we) & !reg_error;
	assign alert_regwen_5_wd = reg_wdata[0];
	assign alert_regwen_6_we = (addr_hit[12] & reg_we) & !reg_error;
	assign alert_regwen_6_wd = reg_wdata[0];
	assign alert_regwen_7_we = (addr_hit[13] & reg_we) & !reg_error;
	assign alert_regwen_7_wd = reg_wdata[0];
	assign alert_regwen_8_we = (addr_hit[14] & reg_we) & !reg_error;
	assign alert_regwen_8_wd = reg_wdata[0];
	assign alert_regwen_9_we = (addr_hit[15] & reg_we) & !reg_error;
	assign alert_regwen_9_wd = reg_wdata[0];
	assign alert_regwen_10_we = (addr_hit[16] & reg_we) & !reg_error;
	assign alert_regwen_10_wd = reg_wdata[0];
	assign alert_regwen_11_we = (addr_hit[17] & reg_we) & !reg_error;
	assign alert_regwen_11_wd = reg_wdata[0];
	assign alert_regwen_12_we = (addr_hit[18] & reg_we) & !reg_error;
	assign alert_regwen_12_wd = reg_wdata[0];
	assign alert_regwen_13_we = (addr_hit[19] & reg_we) & !reg_error;
	assign alert_regwen_13_wd = reg_wdata[0];
	assign alert_regwen_14_we = (addr_hit[20] & reg_we) & !reg_error;
	assign alert_regwen_14_wd = reg_wdata[0];
	assign alert_regwen_15_we = (addr_hit[21] & reg_we) & !reg_error;
	assign alert_regwen_15_wd = reg_wdata[0];
	assign alert_regwen_16_we = (addr_hit[22] & reg_we) & !reg_error;
	assign alert_regwen_16_wd = reg_wdata[0];
	assign alert_regwen_17_we = (addr_hit[23] & reg_we) & !reg_error;
	assign alert_regwen_17_wd = reg_wdata[0];
	assign alert_regwen_18_we = (addr_hit[24] & reg_we) & !reg_error;
	assign alert_regwen_18_wd = reg_wdata[0];
	assign alert_regwen_19_we = (addr_hit[25] & reg_we) & !reg_error;
	assign alert_regwen_19_wd = reg_wdata[0];
	assign alert_regwen_20_we = (addr_hit[26] & reg_we) & !reg_error;
	assign alert_regwen_20_wd = reg_wdata[0];
	assign alert_regwen_21_we = (addr_hit[27] & reg_we) & !reg_error;
	assign alert_regwen_21_wd = reg_wdata[0];
	assign alert_regwen_22_we = (addr_hit[28] & reg_we) & !reg_error;
	assign alert_regwen_22_wd = reg_wdata[0];
	assign alert_regwen_23_we = (addr_hit[29] & reg_we) & !reg_error;
	assign alert_regwen_23_wd = reg_wdata[0];
	assign alert_regwen_24_we = (addr_hit[30] & reg_we) & !reg_error;
	assign alert_regwen_24_wd = reg_wdata[0];
	assign alert_regwen_25_we = (addr_hit[31] & reg_we) & !reg_error;
	assign alert_regwen_25_wd = reg_wdata[0];
	assign alert_regwen_26_we = (addr_hit[32] & reg_we) & !reg_error;
	assign alert_regwen_26_wd = reg_wdata[0];
	assign alert_regwen_27_we = (addr_hit[33] & reg_we) & !reg_error;
	assign alert_regwen_27_wd = reg_wdata[0];
	assign alert_regwen_28_we = (addr_hit[34] & reg_we) & !reg_error;
	assign alert_regwen_28_wd = reg_wdata[0];
	assign alert_regwen_29_we = (addr_hit[35] & reg_we) & !reg_error;
	assign alert_regwen_29_wd = reg_wdata[0];
	assign alert_regwen_30_we = (addr_hit[36] & reg_we) & !reg_error;
	assign alert_regwen_30_wd = reg_wdata[0];
	assign alert_regwen_31_we = (addr_hit[37] & reg_we) & !reg_error;
	assign alert_regwen_31_wd = reg_wdata[0];
	assign alert_regwen_32_we = (addr_hit[38] & reg_we) & !reg_error;
	assign alert_regwen_32_wd = reg_wdata[0];
	assign alert_regwen_33_we = (addr_hit[39] & reg_we) & !reg_error;
	assign alert_regwen_33_wd = reg_wdata[0];
	assign alert_regwen_34_we = (addr_hit[40] & reg_we) & !reg_error;
	assign alert_regwen_34_wd = reg_wdata[0];
	assign alert_regwen_35_we = (addr_hit[41] & reg_we) & !reg_error;
	assign alert_regwen_35_wd = reg_wdata[0];
	assign alert_regwen_36_we = (addr_hit[42] & reg_we) & !reg_error;
	assign alert_regwen_36_wd = reg_wdata[0];
	assign alert_regwen_37_we = (addr_hit[43] & reg_we) & !reg_error;
	assign alert_regwen_37_wd = reg_wdata[0];
	assign alert_regwen_38_we = (addr_hit[44] & reg_we) & !reg_error;
	assign alert_regwen_38_wd = reg_wdata[0];
	assign alert_regwen_39_we = (addr_hit[45] & reg_we) & !reg_error;
	assign alert_regwen_39_wd = reg_wdata[0];
	assign alert_regwen_40_we = (addr_hit[46] & reg_we) & !reg_error;
	assign alert_regwen_40_wd = reg_wdata[0];
	assign alert_regwen_41_we = (addr_hit[47] & reg_we) & !reg_error;
	assign alert_regwen_41_wd = reg_wdata[0];
	assign alert_regwen_42_we = (addr_hit[48] & reg_we) & !reg_error;
	assign alert_regwen_42_wd = reg_wdata[0];
	assign alert_regwen_43_we = (addr_hit[49] & reg_we) & !reg_error;
	assign alert_regwen_43_wd = reg_wdata[0];
	assign alert_regwen_44_we = (addr_hit[50] & reg_we) & !reg_error;
	assign alert_regwen_44_wd = reg_wdata[0];
	assign alert_regwen_45_we = (addr_hit[51] & reg_we) & !reg_error;
	assign alert_regwen_45_wd = reg_wdata[0];
	assign alert_regwen_46_we = (addr_hit[52] & reg_we) & !reg_error;
	assign alert_regwen_46_wd = reg_wdata[0];
	assign alert_regwen_47_we = (addr_hit[53] & reg_we) & !reg_error;
	assign alert_regwen_47_wd = reg_wdata[0];
	assign alert_regwen_48_we = (addr_hit[54] & reg_we) & !reg_error;
	assign alert_regwen_48_wd = reg_wdata[0];
	assign alert_regwen_49_we = (addr_hit[55] & reg_we) & !reg_error;
	assign alert_regwen_49_wd = reg_wdata[0];
	assign alert_regwen_50_we = (addr_hit[56] & reg_we) & !reg_error;
	assign alert_regwen_50_wd = reg_wdata[0];
	assign alert_regwen_51_we = (addr_hit[57] & reg_we) & !reg_error;
	assign alert_regwen_51_wd = reg_wdata[0];
	assign alert_regwen_52_we = (addr_hit[58] & reg_we) & !reg_error;
	assign alert_regwen_52_wd = reg_wdata[0];
	assign alert_regwen_53_we = (addr_hit[59] & reg_we) & !reg_error;
	assign alert_regwen_53_wd = reg_wdata[0];
	assign alert_regwen_54_we = (addr_hit[60] & reg_we) & !reg_error;
	assign alert_regwen_54_wd = reg_wdata[0];
	assign alert_regwen_55_we = (addr_hit[61] & reg_we) & !reg_error;
	assign alert_regwen_55_wd = reg_wdata[0];
	assign alert_regwen_56_we = (addr_hit[62] & reg_we) & !reg_error;
	assign alert_regwen_56_wd = reg_wdata[0];
	assign alert_regwen_57_we = (addr_hit[63] & reg_we) & !reg_error;
	assign alert_regwen_57_wd = reg_wdata[0];
	assign alert_regwen_58_we = (addr_hit[64] & reg_we) & !reg_error;
	assign alert_regwen_58_wd = reg_wdata[0];
	assign alert_regwen_59_we = (addr_hit[65] & reg_we) & !reg_error;
	assign alert_regwen_59_wd = reg_wdata[0];
	assign alert_regwen_60_we = (addr_hit[66] & reg_we) & !reg_error;
	assign alert_regwen_60_wd = reg_wdata[0];
	assign alert_regwen_61_we = (addr_hit[67] & reg_we) & !reg_error;
	assign alert_regwen_61_wd = reg_wdata[0];
	assign alert_regwen_62_we = (addr_hit[68] & reg_we) & !reg_error;
	assign alert_regwen_62_wd = reg_wdata[0];
	assign alert_regwen_63_we = (addr_hit[69] & reg_we) & !reg_error;
	assign alert_regwen_63_wd = reg_wdata[0];
	assign alert_regwen_64_we = (addr_hit[70] & reg_we) & !reg_error;
	assign alert_regwen_64_wd = reg_wdata[0];
	assign alert_en_shadowed_0_re = (addr_hit[71] & reg_re) & !reg_error;
	assign alert_en_shadowed_0_we = (addr_hit[71] & reg_we) & !reg_error;
	assign alert_en_shadowed_0_wd = reg_wdata[0];
	assign alert_en_shadowed_1_re = (addr_hit[72] & reg_re) & !reg_error;
	assign alert_en_shadowed_1_we = (addr_hit[72] & reg_we) & !reg_error;
	assign alert_en_shadowed_1_wd = reg_wdata[0];
	assign alert_en_shadowed_2_re = (addr_hit[73] & reg_re) & !reg_error;
	assign alert_en_shadowed_2_we = (addr_hit[73] & reg_we) & !reg_error;
	assign alert_en_shadowed_2_wd = reg_wdata[0];
	assign alert_en_shadowed_3_re = (addr_hit[74] & reg_re) & !reg_error;
	assign alert_en_shadowed_3_we = (addr_hit[74] & reg_we) & !reg_error;
	assign alert_en_shadowed_3_wd = reg_wdata[0];
	assign alert_en_shadowed_4_re = (addr_hit[75] & reg_re) & !reg_error;
	assign alert_en_shadowed_4_we = (addr_hit[75] & reg_we) & !reg_error;
	assign alert_en_shadowed_4_wd = reg_wdata[0];
	assign alert_en_shadowed_5_re = (addr_hit[76] & reg_re) & !reg_error;
	assign alert_en_shadowed_5_we = (addr_hit[76] & reg_we) & !reg_error;
	assign alert_en_shadowed_5_wd = reg_wdata[0];
	assign alert_en_shadowed_6_re = (addr_hit[77] & reg_re) & !reg_error;
	assign alert_en_shadowed_6_we = (addr_hit[77] & reg_we) & !reg_error;
	assign alert_en_shadowed_6_wd = reg_wdata[0];
	assign alert_en_shadowed_7_re = (addr_hit[78] & reg_re) & !reg_error;
	assign alert_en_shadowed_7_we = (addr_hit[78] & reg_we) & !reg_error;
	assign alert_en_shadowed_7_wd = reg_wdata[0];
	assign alert_en_shadowed_8_re = (addr_hit[79] & reg_re) & !reg_error;
	assign alert_en_shadowed_8_we = (addr_hit[79] & reg_we) & !reg_error;
	assign alert_en_shadowed_8_wd = reg_wdata[0];
	assign alert_en_shadowed_9_re = (addr_hit[80] & reg_re) & !reg_error;
	assign alert_en_shadowed_9_we = (addr_hit[80] & reg_we) & !reg_error;
	assign alert_en_shadowed_9_wd = reg_wdata[0];
	assign alert_en_shadowed_10_re = (addr_hit[81] & reg_re) & !reg_error;
	assign alert_en_shadowed_10_we = (addr_hit[81] & reg_we) & !reg_error;
	assign alert_en_shadowed_10_wd = reg_wdata[0];
	assign alert_en_shadowed_11_re = (addr_hit[82] & reg_re) & !reg_error;
	assign alert_en_shadowed_11_we = (addr_hit[82] & reg_we) & !reg_error;
	assign alert_en_shadowed_11_wd = reg_wdata[0];
	assign alert_en_shadowed_12_re = (addr_hit[83] & reg_re) & !reg_error;
	assign alert_en_shadowed_12_we = (addr_hit[83] & reg_we) & !reg_error;
	assign alert_en_shadowed_12_wd = reg_wdata[0];
	assign alert_en_shadowed_13_re = (addr_hit[84] & reg_re) & !reg_error;
	assign alert_en_shadowed_13_we = (addr_hit[84] & reg_we) & !reg_error;
	assign alert_en_shadowed_13_wd = reg_wdata[0];
	assign alert_en_shadowed_14_re = (addr_hit[85] & reg_re) & !reg_error;
	assign alert_en_shadowed_14_we = (addr_hit[85] & reg_we) & !reg_error;
	assign alert_en_shadowed_14_wd = reg_wdata[0];
	assign alert_en_shadowed_15_re = (addr_hit[86] & reg_re) & !reg_error;
	assign alert_en_shadowed_15_we = (addr_hit[86] & reg_we) & !reg_error;
	assign alert_en_shadowed_15_wd = reg_wdata[0];
	assign alert_en_shadowed_16_re = (addr_hit[87] & reg_re) & !reg_error;
	assign alert_en_shadowed_16_we = (addr_hit[87] & reg_we) & !reg_error;
	assign alert_en_shadowed_16_wd = reg_wdata[0];
	assign alert_en_shadowed_17_re = (addr_hit[88] & reg_re) & !reg_error;
	assign alert_en_shadowed_17_we = (addr_hit[88] & reg_we) & !reg_error;
	assign alert_en_shadowed_17_wd = reg_wdata[0];
	assign alert_en_shadowed_18_re = (addr_hit[89] & reg_re) & !reg_error;
	assign alert_en_shadowed_18_we = (addr_hit[89] & reg_we) & !reg_error;
	assign alert_en_shadowed_18_wd = reg_wdata[0];
	assign alert_en_shadowed_19_re = (addr_hit[90] & reg_re) & !reg_error;
	assign alert_en_shadowed_19_we = (addr_hit[90] & reg_we) & !reg_error;
	assign alert_en_shadowed_19_wd = reg_wdata[0];
	assign alert_en_shadowed_20_re = (addr_hit[91] & reg_re) & !reg_error;
	assign alert_en_shadowed_20_we = (addr_hit[91] & reg_we) & !reg_error;
	assign alert_en_shadowed_20_wd = reg_wdata[0];
	assign alert_en_shadowed_21_re = (addr_hit[92] & reg_re) & !reg_error;
	assign alert_en_shadowed_21_we = (addr_hit[92] & reg_we) & !reg_error;
	assign alert_en_shadowed_21_wd = reg_wdata[0];
	assign alert_en_shadowed_22_re = (addr_hit[93] & reg_re) & !reg_error;
	assign alert_en_shadowed_22_we = (addr_hit[93] & reg_we) & !reg_error;
	assign alert_en_shadowed_22_wd = reg_wdata[0];
	assign alert_en_shadowed_23_re = (addr_hit[94] & reg_re) & !reg_error;
	assign alert_en_shadowed_23_we = (addr_hit[94] & reg_we) & !reg_error;
	assign alert_en_shadowed_23_wd = reg_wdata[0];
	assign alert_en_shadowed_24_re = (addr_hit[95] & reg_re) & !reg_error;
	assign alert_en_shadowed_24_we = (addr_hit[95] & reg_we) & !reg_error;
	assign alert_en_shadowed_24_wd = reg_wdata[0];
	assign alert_en_shadowed_25_re = (addr_hit[96] & reg_re) & !reg_error;
	assign alert_en_shadowed_25_we = (addr_hit[96] & reg_we) & !reg_error;
	assign alert_en_shadowed_25_wd = reg_wdata[0];
	assign alert_en_shadowed_26_re = (addr_hit[97] & reg_re) & !reg_error;
	assign alert_en_shadowed_26_we = (addr_hit[97] & reg_we) & !reg_error;
	assign alert_en_shadowed_26_wd = reg_wdata[0];
	assign alert_en_shadowed_27_re = (addr_hit[98] & reg_re) & !reg_error;
	assign alert_en_shadowed_27_we = (addr_hit[98] & reg_we) & !reg_error;
	assign alert_en_shadowed_27_wd = reg_wdata[0];
	assign alert_en_shadowed_28_re = (addr_hit[99] & reg_re) & !reg_error;
	assign alert_en_shadowed_28_we = (addr_hit[99] & reg_we) & !reg_error;
	assign alert_en_shadowed_28_wd = reg_wdata[0];
	assign alert_en_shadowed_29_re = (addr_hit[100] & reg_re) & !reg_error;
	assign alert_en_shadowed_29_we = (addr_hit[100] & reg_we) & !reg_error;
	assign alert_en_shadowed_29_wd = reg_wdata[0];
	assign alert_en_shadowed_30_re = (addr_hit[101] & reg_re) & !reg_error;
	assign alert_en_shadowed_30_we = (addr_hit[101] & reg_we) & !reg_error;
	assign alert_en_shadowed_30_wd = reg_wdata[0];
	assign alert_en_shadowed_31_re = (addr_hit[102] & reg_re) & !reg_error;
	assign alert_en_shadowed_31_we = (addr_hit[102] & reg_we) & !reg_error;
	assign alert_en_shadowed_31_wd = reg_wdata[0];
	assign alert_en_shadowed_32_re = (addr_hit[103] & reg_re) & !reg_error;
	assign alert_en_shadowed_32_we = (addr_hit[103] & reg_we) & !reg_error;
	assign alert_en_shadowed_32_wd = reg_wdata[0];
	assign alert_en_shadowed_33_re = (addr_hit[104] & reg_re) & !reg_error;
	assign alert_en_shadowed_33_we = (addr_hit[104] & reg_we) & !reg_error;
	assign alert_en_shadowed_33_wd = reg_wdata[0];
	assign alert_en_shadowed_34_re = (addr_hit[105] & reg_re) & !reg_error;
	assign alert_en_shadowed_34_we = (addr_hit[105] & reg_we) & !reg_error;
	assign alert_en_shadowed_34_wd = reg_wdata[0];
	assign alert_en_shadowed_35_re = (addr_hit[106] & reg_re) & !reg_error;
	assign alert_en_shadowed_35_we = (addr_hit[106] & reg_we) & !reg_error;
	assign alert_en_shadowed_35_wd = reg_wdata[0];
	assign alert_en_shadowed_36_re = (addr_hit[107] & reg_re) & !reg_error;
	assign alert_en_shadowed_36_we = (addr_hit[107] & reg_we) & !reg_error;
	assign alert_en_shadowed_36_wd = reg_wdata[0];
	assign alert_en_shadowed_37_re = (addr_hit[108] & reg_re) & !reg_error;
	assign alert_en_shadowed_37_we = (addr_hit[108] & reg_we) & !reg_error;
	assign alert_en_shadowed_37_wd = reg_wdata[0];
	assign alert_en_shadowed_38_re = (addr_hit[109] & reg_re) & !reg_error;
	assign alert_en_shadowed_38_we = (addr_hit[109] & reg_we) & !reg_error;
	assign alert_en_shadowed_38_wd = reg_wdata[0];
	assign alert_en_shadowed_39_re = (addr_hit[110] & reg_re) & !reg_error;
	assign alert_en_shadowed_39_we = (addr_hit[110] & reg_we) & !reg_error;
	assign alert_en_shadowed_39_wd = reg_wdata[0];
	assign alert_en_shadowed_40_re = (addr_hit[111] & reg_re) & !reg_error;
	assign alert_en_shadowed_40_we = (addr_hit[111] & reg_we) & !reg_error;
	assign alert_en_shadowed_40_wd = reg_wdata[0];
	assign alert_en_shadowed_41_re = (addr_hit[112] & reg_re) & !reg_error;
	assign alert_en_shadowed_41_we = (addr_hit[112] & reg_we) & !reg_error;
	assign alert_en_shadowed_41_wd = reg_wdata[0];
	assign alert_en_shadowed_42_re = (addr_hit[113] & reg_re) & !reg_error;
	assign alert_en_shadowed_42_we = (addr_hit[113] & reg_we) & !reg_error;
	assign alert_en_shadowed_42_wd = reg_wdata[0];
	assign alert_en_shadowed_43_re = (addr_hit[114] & reg_re) & !reg_error;
	assign alert_en_shadowed_43_we = (addr_hit[114] & reg_we) & !reg_error;
	assign alert_en_shadowed_43_wd = reg_wdata[0];
	assign alert_en_shadowed_44_re = (addr_hit[115] & reg_re) & !reg_error;
	assign alert_en_shadowed_44_we = (addr_hit[115] & reg_we) & !reg_error;
	assign alert_en_shadowed_44_wd = reg_wdata[0];
	assign alert_en_shadowed_45_re = (addr_hit[116] & reg_re) & !reg_error;
	assign alert_en_shadowed_45_we = (addr_hit[116] & reg_we) & !reg_error;
	assign alert_en_shadowed_45_wd = reg_wdata[0];
	assign alert_en_shadowed_46_re = (addr_hit[117] & reg_re) & !reg_error;
	assign alert_en_shadowed_46_we = (addr_hit[117] & reg_we) & !reg_error;
	assign alert_en_shadowed_46_wd = reg_wdata[0];
	assign alert_en_shadowed_47_re = (addr_hit[118] & reg_re) & !reg_error;
	assign alert_en_shadowed_47_we = (addr_hit[118] & reg_we) & !reg_error;
	assign alert_en_shadowed_47_wd = reg_wdata[0];
	assign alert_en_shadowed_48_re = (addr_hit[119] & reg_re) & !reg_error;
	assign alert_en_shadowed_48_we = (addr_hit[119] & reg_we) & !reg_error;
	assign alert_en_shadowed_48_wd = reg_wdata[0];
	assign alert_en_shadowed_49_re = (addr_hit[120] & reg_re) & !reg_error;
	assign alert_en_shadowed_49_we = (addr_hit[120] & reg_we) & !reg_error;
	assign alert_en_shadowed_49_wd = reg_wdata[0];
	assign alert_en_shadowed_50_re = (addr_hit[121] & reg_re) & !reg_error;
	assign alert_en_shadowed_50_we = (addr_hit[121] & reg_we) & !reg_error;
	assign alert_en_shadowed_50_wd = reg_wdata[0];
	assign alert_en_shadowed_51_re = (addr_hit[122] & reg_re) & !reg_error;
	assign alert_en_shadowed_51_we = (addr_hit[122] & reg_we) & !reg_error;
	assign alert_en_shadowed_51_wd = reg_wdata[0];
	assign alert_en_shadowed_52_re = (addr_hit[123] & reg_re) & !reg_error;
	assign alert_en_shadowed_52_we = (addr_hit[123] & reg_we) & !reg_error;
	assign alert_en_shadowed_52_wd = reg_wdata[0];
	assign alert_en_shadowed_53_re = (addr_hit[124] & reg_re) & !reg_error;
	assign alert_en_shadowed_53_we = (addr_hit[124] & reg_we) & !reg_error;
	assign alert_en_shadowed_53_wd = reg_wdata[0];
	assign alert_en_shadowed_54_re = (addr_hit[125] & reg_re) & !reg_error;
	assign alert_en_shadowed_54_we = (addr_hit[125] & reg_we) & !reg_error;
	assign alert_en_shadowed_54_wd = reg_wdata[0];
	assign alert_en_shadowed_55_re = (addr_hit[126] & reg_re) & !reg_error;
	assign alert_en_shadowed_55_we = (addr_hit[126] & reg_we) & !reg_error;
	assign alert_en_shadowed_55_wd = reg_wdata[0];
	assign alert_en_shadowed_56_re = (addr_hit[127] & reg_re) & !reg_error;
	assign alert_en_shadowed_56_we = (addr_hit[127] & reg_we) & !reg_error;
	assign alert_en_shadowed_56_wd = reg_wdata[0];
	assign alert_en_shadowed_57_re = (addr_hit[128] & reg_re) & !reg_error;
	assign alert_en_shadowed_57_we = (addr_hit[128] & reg_we) & !reg_error;
	assign alert_en_shadowed_57_wd = reg_wdata[0];
	assign alert_en_shadowed_58_re = (addr_hit[129] & reg_re) & !reg_error;
	assign alert_en_shadowed_58_we = (addr_hit[129] & reg_we) & !reg_error;
	assign alert_en_shadowed_58_wd = reg_wdata[0];
	assign alert_en_shadowed_59_re = (addr_hit[130] & reg_re) & !reg_error;
	assign alert_en_shadowed_59_we = (addr_hit[130] & reg_we) & !reg_error;
	assign alert_en_shadowed_59_wd = reg_wdata[0];
	assign alert_en_shadowed_60_re = (addr_hit[131] & reg_re) & !reg_error;
	assign alert_en_shadowed_60_we = (addr_hit[131] & reg_we) & !reg_error;
	assign alert_en_shadowed_60_wd = reg_wdata[0];
	assign alert_en_shadowed_61_re = (addr_hit[132] & reg_re) & !reg_error;
	assign alert_en_shadowed_61_we = (addr_hit[132] & reg_we) & !reg_error;
	assign alert_en_shadowed_61_wd = reg_wdata[0];
	assign alert_en_shadowed_62_re = (addr_hit[133] & reg_re) & !reg_error;
	assign alert_en_shadowed_62_we = (addr_hit[133] & reg_we) & !reg_error;
	assign alert_en_shadowed_62_wd = reg_wdata[0];
	assign alert_en_shadowed_63_re = (addr_hit[134] & reg_re) & !reg_error;
	assign alert_en_shadowed_63_we = (addr_hit[134] & reg_we) & !reg_error;
	assign alert_en_shadowed_63_wd = reg_wdata[0];
	assign alert_en_shadowed_64_re = (addr_hit[135] & reg_re) & !reg_error;
	assign alert_en_shadowed_64_we = (addr_hit[135] & reg_we) & !reg_error;
	assign alert_en_shadowed_64_wd = reg_wdata[0];
	assign alert_class_shadowed_0_re = (addr_hit[136] & reg_re) & !reg_error;
	assign alert_class_shadowed_0_we = (addr_hit[136] & reg_we) & !reg_error;
	assign alert_class_shadowed_0_wd = reg_wdata[1:0];
	assign alert_class_shadowed_1_re = (addr_hit[137] & reg_re) & !reg_error;
	assign alert_class_shadowed_1_we = (addr_hit[137] & reg_we) & !reg_error;
	assign alert_class_shadowed_1_wd = reg_wdata[1:0];
	assign alert_class_shadowed_2_re = (addr_hit[138] & reg_re) & !reg_error;
	assign alert_class_shadowed_2_we = (addr_hit[138] & reg_we) & !reg_error;
	assign alert_class_shadowed_2_wd = reg_wdata[1:0];
	assign alert_class_shadowed_3_re = (addr_hit[139] & reg_re) & !reg_error;
	assign alert_class_shadowed_3_we = (addr_hit[139] & reg_we) & !reg_error;
	assign alert_class_shadowed_3_wd = reg_wdata[1:0];
	assign alert_class_shadowed_4_re = (addr_hit[140] & reg_re) & !reg_error;
	assign alert_class_shadowed_4_we = (addr_hit[140] & reg_we) & !reg_error;
	assign alert_class_shadowed_4_wd = reg_wdata[1:0];
	assign alert_class_shadowed_5_re = (addr_hit[141] & reg_re) & !reg_error;
	assign alert_class_shadowed_5_we = (addr_hit[141] & reg_we) & !reg_error;
	assign alert_class_shadowed_5_wd = reg_wdata[1:0];
	assign alert_class_shadowed_6_re = (addr_hit[142] & reg_re) & !reg_error;
	assign alert_class_shadowed_6_we = (addr_hit[142] & reg_we) & !reg_error;
	assign alert_class_shadowed_6_wd = reg_wdata[1:0];
	assign alert_class_shadowed_7_re = (addr_hit[143] & reg_re) & !reg_error;
	assign alert_class_shadowed_7_we = (addr_hit[143] & reg_we) & !reg_error;
	assign alert_class_shadowed_7_wd = reg_wdata[1:0];
	assign alert_class_shadowed_8_re = (addr_hit[144] & reg_re) & !reg_error;
	assign alert_class_shadowed_8_we = (addr_hit[144] & reg_we) & !reg_error;
	assign alert_class_shadowed_8_wd = reg_wdata[1:0];
	assign alert_class_shadowed_9_re = (addr_hit[145] & reg_re) & !reg_error;
	assign alert_class_shadowed_9_we = (addr_hit[145] & reg_we) & !reg_error;
	assign alert_class_shadowed_9_wd = reg_wdata[1:0];
	assign alert_class_shadowed_10_re = (addr_hit[146] & reg_re) & !reg_error;
	assign alert_class_shadowed_10_we = (addr_hit[146] & reg_we) & !reg_error;
	assign alert_class_shadowed_10_wd = reg_wdata[1:0];
	assign alert_class_shadowed_11_re = (addr_hit[147] & reg_re) & !reg_error;
	assign alert_class_shadowed_11_we = (addr_hit[147] & reg_we) & !reg_error;
	assign alert_class_shadowed_11_wd = reg_wdata[1:0];
	assign alert_class_shadowed_12_re = (addr_hit[148] & reg_re) & !reg_error;
	assign alert_class_shadowed_12_we = (addr_hit[148] & reg_we) & !reg_error;
	assign alert_class_shadowed_12_wd = reg_wdata[1:0];
	assign alert_class_shadowed_13_re = (addr_hit[149] & reg_re) & !reg_error;
	assign alert_class_shadowed_13_we = (addr_hit[149] & reg_we) & !reg_error;
	assign alert_class_shadowed_13_wd = reg_wdata[1:0];
	assign alert_class_shadowed_14_re = (addr_hit[150] & reg_re) & !reg_error;
	assign alert_class_shadowed_14_we = (addr_hit[150] & reg_we) & !reg_error;
	assign alert_class_shadowed_14_wd = reg_wdata[1:0];
	assign alert_class_shadowed_15_re = (addr_hit[151] & reg_re) & !reg_error;
	assign alert_class_shadowed_15_we = (addr_hit[151] & reg_we) & !reg_error;
	assign alert_class_shadowed_15_wd = reg_wdata[1:0];
	assign alert_class_shadowed_16_re = (addr_hit[152] & reg_re) & !reg_error;
	assign alert_class_shadowed_16_we = (addr_hit[152] & reg_we) & !reg_error;
	assign alert_class_shadowed_16_wd = reg_wdata[1:0];
	assign alert_class_shadowed_17_re = (addr_hit[153] & reg_re) & !reg_error;
	assign alert_class_shadowed_17_we = (addr_hit[153] & reg_we) & !reg_error;
	assign alert_class_shadowed_17_wd = reg_wdata[1:0];
	assign alert_class_shadowed_18_re = (addr_hit[154] & reg_re) & !reg_error;
	assign alert_class_shadowed_18_we = (addr_hit[154] & reg_we) & !reg_error;
	assign alert_class_shadowed_18_wd = reg_wdata[1:0];
	assign alert_class_shadowed_19_re = (addr_hit[155] & reg_re) & !reg_error;
	assign alert_class_shadowed_19_we = (addr_hit[155] & reg_we) & !reg_error;
	assign alert_class_shadowed_19_wd = reg_wdata[1:0];
	assign alert_class_shadowed_20_re = (addr_hit[156] & reg_re) & !reg_error;
	assign alert_class_shadowed_20_we = (addr_hit[156] & reg_we) & !reg_error;
	assign alert_class_shadowed_20_wd = reg_wdata[1:0];
	assign alert_class_shadowed_21_re = (addr_hit[157] & reg_re) & !reg_error;
	assign alert_class_shadowed_21_we = (addr_hit[157] & reg_we) & !reg_error;
	assign alert_class_shadowed_21_wd = reg_wdata[1:0];
	assign alert_class_shadowed_22_re = (addr_hit[158] & reg_re) & !reg_error;
	assign alert_class_shadowed_22_we = (addr_hit[158] & reg_we) & !reg_error;
	assign alert_class_shadowed_22_wd = reg_wdata[1:0];
	assign alert_class_shadowed_23_re = (addr_hit[159] & reg_re) & !reg_error;
	assign alert_class_shadowed_23_we = (addr_hit[159] & reg_we) & !reg_error;
	assign alert_class_shadowed_23_wd = reg_wdata[1:0];
	assign alert_class_shadowed_24_re = (addr_hit[160] & reg_re) & !reg_error;
	assign alert_class_shadowed_24_we = (addr_hit[160] & reg_we) & !reg_error;
	assign alert_class_shadowed_24_wd = reg_wdata[1:0];
	assign alert_class_shadowed_25_re = (addr_hit[161] & reg_re) & !reg_error;
	assign alert_class_shadowed_25_we = (addr_hit[161] & reg_we) & !reg_error;
	assign alert_class_shadowed_25_wd = reg_wdata[1:0];
	assign alert_class_shadowed_26_re = (addr_hit[162] & reg_re) & !reg_error;
	assign alert_class_shadowed_26_we = (addr_hit[162] & reg_we) & !reg_error;
	assign alert_class_shadowed_26_wd = reg_wdata[1:0];
	assign alert_class_shadowed_27_re = (addr_hit[163] & reg_re) & !reg_error;
	assign alert_class_shadowed_27_we = (addr_hit[163] & reg_we) & !reg_error;
	assign alert_class_shadowed_27_wd = reg_wdata[1:0];
	assign alert_class_shadowed_28_re = (addr_hit[164] & reg_re) & !reg_error;
	assign alert_class_shadowed_28_we = (addr_hit[164] & reg_we) & !reg_error;
	assign alert_class_shadowed_28_wd = reg_wdata[1:0];
	assign alert_class_shadowed_29_re = (addr_hit[165] & reg_re) & !reg_error;
	assign alert_class_shadowed_29_we = (addr_hit[165] & reg_we) & !reg_error;
	assign alert_class_shadowed_29_wd = reg_wdata[1:0];
	assign alert_class_shadowed_30_re = (addr_hit[166] & reg_re) & !reg_error;
	assign alert_class_shadowed_30_we = (addr_hit[166] & reg_we) & !reg_error;
	assign alert_class_shadowed_30_wd = reg_wdata[1:0];
	assign alert_class_shadowed_31_re = (addr_hit[167] & reg_re) & !reg_error;
	assign alert_class_shadowed_31_we = (addr_hit[167] & reg_we) & !reg_error;
	assign alert_class_shadowed_31_wd = reg_wdata[1:0];
	assign alert_class_shadowed_32_re = (addr_hit[168] & reg_re) & !reg_error;
	assign alert_class_shadowed_32_we = (addr_hit[168] & reg_we) & !reg_error;
	assign alert_class_shadowed_32_wd = reg_wdata[1:0];
	assign alert_class_shadowed_33_re = (addr_hit[169] & reg_re) & !reg_error;
	assign alert_class_shadowed_33_we = (addr_hit[169] & reg_we) & !reg_error;
	assign alert_class_shadowed_33_wd = reg_wdata[1:0];
	assign alert_class_shadowed_34_re = (addr_hit[170] & reg_re) & !reg_error;
	assign alert_class_shadowed_34_we = (addr_hit[170] & reg_we) & !reg_error;
	assign alert_class_shadowed_34_wd = reg_wdata[1:0];
	assign alert_class_shadowed_35_re = (addr_hit[171] & reg_re) & !reg_error;
	assign alert_class_shadowed_35_we = (addr_hit[171] & reg_we) & !reg_error;
	assign alert_class_shadowed_35_wd = reg_wdata[1:0];
	assign alert_class_shadowed_36_re = (addr_hit[172] & reg_re) & !reg_error;
	assign alert_class_shadowed_36_we = (addr_hit[172] & reg_we) & !reg_error;
	assign alert_class_shadowed_36_wd = reg_wdata[1:0];
	assign alert_class_shadowed_37_re = (addr_hit[173] & reg_re) & !reg_error;
	assign alert_class_shadowed_37_we = (addr_hit[173] & reg_we) & !reg_error;
	assign alert_class_shadowed_37_wd = reg_wdata[1:0];
	assign alert_class_shadowed_38_re = (addr_hit[174] & reg_re) & !reg_error;
	assign alert_class_shadowed_38_we = (addr_hit[174] & reg_we) & !reg_error;
	assign alert_class_shadowed_38_wd = reg_wdata[1:0];
	assign alert_class_shadowed_39_re = (addr_hit[175] & reg_re) & !reg_error;
	assign alert_class_shadowed_39_we = (addr_hit[175] & reg_we) & !reg_error;
	assign alert_class_shadowed_39_wd = reg_wdata[1:0];
	assign alert_class_shadowed_40_re = (addr_hit[176] & reg_re) & !reg_error;
	assign alert_class_shadowed_40_we = (addr_hit[176] & reg_we) & !reg_error;
	assign alert_class_shadowed_40_wd = reg_wdata[1:0];
	assign alert_class_shadowed_41_re = (addr_hit[177] & reg_re) & !reg_error;
	assign alert_class_shadowed_41_we = (addr_hit[177] & reg_we) & !reg_error;
	assign alert_class_shadowed_41_wd = reg_wdata[1:0];
	assign alert_class_shadowed_42_re = (addr_hit[178] & reg_re) & !reg_error;
	assign alert_class_shadowed_42_we = (addr_hit[178] & reg_we) & !reg_error;
	assign alert_class_shadowed_42_wd = reg_wdata[1:0];
	assign alert_class_shadowed_43_re = (addr_hit[179] & reg_re) & !reg_error;
	assign alert_class_shadowed_43_we = (addr_hit[179] & reg_we) & !reg_error;
	assign alert_class_shadowed_43_wd = reg_wdata[1:0];
	assign alert_class_shadowed_44_re = (addr_hit[180] & reg_re) & !reg_error;
	assign alert_class_shadowed_44_we = (addr_hit[180] & reg_we) & !reg_error;
	assign alert_class_shadowed_44_wd = reg_wdata[1:0];
	assign alert_class_shadowed_45_re = (addr_hit[181] & reg_re) & !reg_error;
	assign alert_class_shadowed_45_we = (addr_hit[181] & reg_we) & !reg_error;
	assign alert_class_shadowed_45_wd = reg_wdata[1:0];
	assign alert_class_shadowed_46_re = (addr_hit[182] & reg_re) & !reg_error;
	assign alert_class_shadowed_46_we = (addr_hit[182] & reg_we) & !reg_error;
	assign alert_class_shadowed_46_wd = reg_wdata[1:0];
	assign alert_class_shadowed_47_re = (addr_hit[183] & reg_re) & !reg_error;
	assign alert_class_shadowed_47_we = (addr_hit[183] & reg_we) & !reg_error;
	assign alert_class_shadowed_47_wd = reg_wdata[1:0];
	assign alert_class_shadowed_48_re = (addr_hit[184] & reg_re) & !reg_error;
	assign alert_class_shadowed_48_we = (addr_hit[184] & reg_we) & !reg_error;
	assign alert_class_shadowed_48_wd = reg_wdata[1:0];
	assign alert_class_shadowed_49_re = (addr_hit[185] & reg_re) & !reg_error;
	assign alert_class_shadowed_49_we = (addr_hit[185] & reg_we) & !reg_error;
	assign alert_class_shadowed_49_wd = reg_wdata[1:0];
	assign alert_class_shadowed_50_re = (addr_hit[186] & reg_re) & !reg_error;
	assign alert_class_shadowed_50_we = (addr_hit[186] & reg_we) & !reg_error;
	assign alert_class_shadowed_50_wd = reg_wdata[1:0];
	assign alert_class_shadowed_51_re = (addr_hit[187] & reg_re) & !reg_error;
	assign alert_class_shadowed_51_we = (addr_hit[187] & reg_we) & !reg_error;
	assign alert_class_shadowed_51_wd = reg_wdata[1:0];
	assign alert_class_shadowed_52_re = (addr_hit[188] & reg_re) & !reg_error;
	assign alert_class_shadowed_52_we = (addr_hit[188] & reg_we) & !reg_error;
	assign alert_class_shadowed_52_wd = reg_wdata[1:0];
	assign alert_class_shadowed_53_re = (addr_hit[189] & reg_re) & !reg_error;
	assign alert_class_shadowed_53_we = (addr_hit[189] & reg_we) & !reg_error;
	assign alert_class_shadowed_53_wd = reg_wdata[1:0];
	assign alert_class_shadowed_54_re = (addr_hit[190] & reg_re) & !reg_error;
	assign alert_class_shadowed_54_we = (addr_hit[190] & reg_we) & !reg_error;
	assign alert_class_shadowed_54_wd = reg_wdata[1:0];
	assign alert_class_shadowed_55_re = (addr_hit[191] & reg_re) & !reg_error;
	assign alert_class_shadowed_55_we = (addr_hit[191] & reg_we) & !reg_error;
	assign alert_class_shadowed_55_wd = reg_wdata[1:0];
	assign alert_class_shadowed_56_re = (addr_hit[192] & reg_re) & !reg_error;
	assign alert_class_shadowed_56_we = (addr_hit[192] & reg_we) & !reg_error;
	assign alert_class_shadowed_56_wd = reg_wdata[1:0];
	assign alert_class_shadowed_57_re = (addr_hit[193] & reg_re) & !reg_error;
	assign alert_class_shadowed_57_we = (addr_hit[193] & reg_we) & !reg_error;
	assign alert_class_shadowed_57_wd = reg_wdata[1:0];
	assign alert_class_shadowed_58_re = (addr_hit[194] & reg_re) & !reg_error;
	assign alert_class_shadowed_58_we = (addr_hit[194] & reg_we) & !reg_error;
	assign alert_class_shadowed_58_wd = reg_wdata[1:0];
	assign alert_class_shadowed_59_re = (addr_hit[195] & reg_re) & !reg_error;
	assign alert_class_shadowed_59_we = (addr_hit[195] & reg_we) & !reg_error;
	assign alert_class_shadowed_59_wd = reg_wdata[1:0];
	assign alert_class_shadowed_60_re = (addr_hit[196] & reg_re) & !reg_error;
	assign alert_class_shadowed_60_we = (addr_hit[196] & reg_we) & !reg_error;
	assign alert_class_shadowed_60_wd = reg_wdata[1:0];
	assign alert_class_shadowed_61_re = (addr_hit[197] & reg_re) & !reg_error;
	assign alert_class_shadowed_61_we = (addr_hit[197] & reg_we) & !reg_error;
	assign alert_class_shadowed_61_wd = reg_wdata[1:0];
	assign alert_class_shadowed_62_re = (addr_hit[198] & reg_re) & !reg_error;
	assign alert_class_shadowed_62_we = (addr_hit[198] & reg_we) & !reg_error;
	assign alert_class_shadowed_62_wd = reg_wdata[1:0];
	assign alert_class_shadowed_63_re = (addr_hit[199] & reg_re) & !reg_error;
	assign alert_class_shadowed_63_we = (addr_hit[199] & reg_we) & !reg_error;
	assign alert_class_shadowed_63_wd = reg_wdata[1:0];
	assign alert_class_shadowed_64_re = (addr_hit[200] & reg_re) & !reg_error;
	assign alert_class_shadowed_64_we = (addr_hit[200] & reg_we) & !reg_error;
	assign alert_class_shadowed_64_wd = reg_wdata[1:0];
	assign alert_cause_0_we = (addr_hit[201] & reg_we) & !reg_error;
	assign alert_cause_0_wd = reg_wdata[0];
	assign alert_cause_1_we = (addr_hit[202] & reg_we) & !reg_error;
	assign alert_cause_1_wd = reg_wdata[0];
	assign alert_cause_2_we = (addr_hit[203] & reg_we) & !reg_error;
	assign alert_cause_2_wd = reg_wdata[0];
	assign alert_cause_3_we = (addr_hit[204] & reg_we) & !reg_error;
	assign alert_cause_3_wd = reg_wdata[0];
	assign alert_cause_4_we = (addr_hit[205] & reg_we) & !reg_error;
	assign alert_cause_4_wd = reg_wdata[0];
	assign alert_cause_5_we = (addr_hit[206] & reg_we) & !reg_error;
	assign alert_cause_5_wd = reg_wdata[0];
	assign alert_cause_6_we = (addr_hit[207] & reg_we) & !reg_error;
	assign alert_cause_6_wd = reg_wdata[0];
	assign alert_cause_7_we = (addr_hit[208] & reg_we) & !reg_error;
	assign alert_cause_7_wd = reg_wdata[0];
	assign alert_cause_8_we = (addr_hit[209] & reg_we) & !reg_error;
	assign alert_cause_8_wd = reg_wdata[0];
	assign alert_cause_9_we = (addr_hit[210] & reg_we) & !reg_error;
	assign alert_cause_9_wd = reg_wdata[0];
	assign alert_cause_10_we = (addr_hit[211] & reg_we) & !reg_error;
	assign alert_cause_10_wd = reg_wdata[0];
	assign alert_cause_11_we = (addr_hit[212] & reg_we) & !reg_error;
	assign alert_cause_11_wd = reg_wdata[0];
	assign alert_cause_12_we = (addr_hit[213] & reg_we) & !reg_error;
	assign alert_cause_12_wd = reg_wdata[0];
	assign alert_cause_13_we = (addr_hit[214] & reg_we) & !reg_error;
	assign alert_cause_13_wd = reg_wdata[0];
	assign alert_cause_14_we = (addr_hit[215] & reg_we) & !reg_error;
	assign alert_cause_14_wd = reg_wdata[0];
	assign alert_cause_15_we = (addr_hit[216] & reg_we) & !reg_error;
	assign alert_cause_15_wd = reg_wdata[0];
	assign alert_cause_16_we = (addr_hit[217] & reg_we) & !reg_error;
	assign alert_cause_16_wd = reg_wdata[0];
	assign alert_cause_17_we = (addr_hit[218] & reg_we) & !reg_error;
	assign alert_cause_17_wd = reg_wdata[0];
	assign alert_cause_18_we = (addr_hit[219] & reg_we) & !reg_error;
	assign alert_cause_18_wd = reg_wdata[0];
	assign alert_cause_19_we = (addr_hit[220] & reg_we) & !reg_error;
	assign alert_cause_19_wd = reg_wdata[0];
	assign alert_cause_20_we = (addr_hit[221] & reg_we) & !reg_error;
	assign alert_cause_20_wd = reg_wdata[0];
	assign alert_cause_21_we = (addr_hit[222] & reg_we) & !reg_error;
	assign alert_cause_21_wd = reg_wdata[0];
	assign alert_cause_22_we = (addr_hit[223] & reg_we) & !reg_error;
	assign alert_cause_22_wd = reg_wdata[0];
	assign alert_cause_23_we = (addr_hit[224] & reg_we) & !reg_error;
	assign alert_cause_23_wd = reg_wdata[0];
	assign alert_cause_24_we = (addr_hit[225] & reg_we) & !reg_error;
	assign alert_cause_24_wd = reg_wdata[0];
	assign alert_cause_25_we = (addr_hit[226] & reg_we) & !reg_error;
	assign alert_cause_25_wd = reg_wdata[0];
	assign alert_cause_26_we = (addr_hit[227] & reg_we) & !reg_error;
	assign alert_cause_26_wd = reg_wdata[0];
	assign alert_cause_27_we = (addr_hit[228] & reg_we) & !reg_error;
	assign alert_cause_27_wd = reg_wdata[0];
	assign alert_cause_28_we = (addr_hit[229] & reg_we) & !reg_error;
	assign alert_cause_28_wd = reg_wdata[0];
	assign alert_cause_29_we = (addr_hit[230] & reg_we) & !reg_error;
	assign alert_cause_29_wd = reg_wdata[0];
	assign alert_cause_30_we = (addr_hit[231] & reg_we) & !reg_error;
	assign alert_cause_30_wd = reg_wdata[0];
	assign alert_cause_31_we = (addr_hit[232] & reg_we) & !reg_error;
	assign alert_cause_31_wd = reg_wdata[0];
	assign alert_cause_32_we = (addr_hit[233] & reg_we) & !reg_error;
	assign alert_cause_32_wd = reg_wdata[0];
	assign alert_cause_33_we = (addr_hit[234] & reg_we) & !reg_error;
	assign alert_cause_33_wd = reg_wdata[0];
	assign alert_cause_34_we = (addr_hit[235] & reg_we) & !reg_error;
	assign alert_cause_34_wd = reg_wdata[0];
	assign alert_cause_35_we = (addr_hit[236] & reg_we) & !reg_error;
	assign alert_cause_35_wd = reg_wdata[0];
	assign alert_cause_36_we = (addr_hit[237] & reg_we) & !reg_error;
	assign alert_cause_36_wd = reg_wdata[0];
	assign alert_cause_37_we = (addr_hit[238] & reg_we) & !reg_error;
	assign alert_cause_37_wd = reg_wdata[0];
	assign alert_cause_38_we = (addr_hit[239] & reg_we) & !reg_error;
	assign alert_cause_38_wd = reg_wdata[0];
	assign alert_cause_39_we = (addr_hit[240] & reg_we) & !reg_error;
	assign alert_cause_39_wd = reg_wdata[0];
	assign alert_cause_40_we = (addr_hit[241] & reg_we) & !reg_error;
	assign alert_cause_40_wd = reg_wdata[0];
	assign alert_cause_41_we = (addr_hit[242] & reg_we) & !reg_error;
	assign alert_cause_41_wd = reg_wdata[0];
	assign alert_cause_42_we = (addr_hit[243] & reg_we) & !reg_error;
	assign alert_cause_42_wd = reg_wdata[0];
	assign alert_cause_43_we = (addr_hit[244] & reg_we) & !reg_error;
	assign alert_cause_43_wd = reg_wdata[0];
	assign alert_cause_44_we = (addr_hit[245] & reg_we) & !reg_error;
	assign alert_cause_44_wd = reg_wdata[0];
	assign alert_cause_45_we = (addr_hit[246] & reg_we) & !reg_error;
	assign alert_cause_45_wd = reg_wdata[0];
	assign alert_cause_46_we = (addr_hit[247] & reg_we) & !reg_error;
	assign alert_cause_46_wd = reg_wdata[0];
	assign alert_cause_47_we = (addr_hit[248] & reg_we) & !reg_error;
	assign alert_cause_47_wd = reg_wdata[0];
	assign alert_cause_48_we = (addr_hit[249] & reg_we) & !reg_error;
	assign alert_cause_48_wd = reg_wdata[0];
	assign alert_cause_49_we = (addr_hit[250] & reg_we) & !reg_error;
	assign alert_cause_49_wd = reg_wdata[0];
	assign alert_cause_50_we = (addr_hit[251] & reg_we) & !reg_error;
	assign alert_cause_50_wd = reg_wdata[0];
	assign alert_cause_51_we = (addr_hit[252] & reg_we) & !reg_error;
	assign alert_cause_51_wd = reg_wdata[0];
	assign alert_cause_52_we = (addr_hit[253] & reg_we) & !reg_error;
	assign alert_cause_52_wd = reg_wdata[0];
	assign alert_cause_53_we = (addr_hit[254] & reg_we) & !reg_error;
	assign alert_cause_53_wd = reg_wdata[0];
	assign alert_cause_54_we = (addr_hit[255] & reg_we) & !reg_error;
	assign alert_cause_54_wd = reg_wdata[0];
	assign alert_cause_55_we = (addr_hit[256] & reg_we) & !reg_error;
	assign alert_cause_55_wd = reg_wdata[0];
	assign alert_cause_56_we = (addr_hit[257] & reg_we) & !reg_error;
	assign alert_cause_56_wd = reg_wdata[0];
	assign alert_cause_57_we = (addr_hit[258] & reg_we) & !reg_error;
	assign alert_cause_57_wd = reg_wdata[0];
	assign alert_cause_58_we = (addr_hit[259] & reg_we) & !reg_error;
	assign alert_cause_58_wd = reg_wdata[0];
	assign alert_cause_59_we = (addr_hit[260] & reg_we) & !reg_error;
	assign alert_cause_59_wd = reg_wdata[0];
	assign alert_cause_60_we = (addr_hit[261] & reg_we) & !reg_error;
	assign alert_cause_60_wd = reg_wdata[0];
	assign alert_cause_61_we = (addr_hit[262] & reg_we) & !reg_error;
	assign alert_cause_61_wd = reg_wdata[0];
	assign alert_cause_62_we = (addr_hit[263] & reg_we) & !reg_error;
	assign alert_cause_62_wd = reg_wdata[0];
	assign alert_cause_63_we = (addr_hit[264] & reg_we) & !reg_error;
	assign alert_cause_63_wd = reg_wdata[0];
	assign alert_cause_64_we = (addr_hit[265] & reg_we) & !reg_error;
	assign alert_cause_64_wd = reg_wdata[0];
	assign loc_alert_regwen_0_we = (addr_hit[266] & reg_we) & !reg_error;
	assign loc_alert_regwen_0_wd = reg_wdata[0];
	assign loc_alert_regwen_1_we = (addr_hit[267] & reg_we) & !reg_error;
	assign loc_alert_regwen_1_wd = reg_wdata[0];
	assign loc_alert_regwen_2_we = (addr_hit[268] & reg_we) & !reg_error;
	assign loc_alert_regwen_2_wd = reg_wdata[0];
	assign loc_alert_regwen_3_we = (addr_hit[269] & reg_we) & !reg_error;
	assign loc_alert_regwen_3_wd = reg_wdata[0];
	assign loc_alert_regwen_4_we = (addr_hit[270] & reg_we) & !reg_error;
	assign loc_alert_regwen_4_wd = reg_wdata[0];
	assign loc_alert_regwen_5_we = (addr_hit[271] & reg_we) & !reg_error;
	assign loc_alert_regwen_5_wd = reg_wdata[0];
	assign loc_alert_regwen_6_we = (addr_hit[272] & reg_we) & !reg_error;
	assign loc_alert_regwen_6_wd = reg_wdata[0];
	assign loc_alert_en_shadowed_0_re = (addr_hit[273] & reg_re) & !reg_error;
	assign loc_alert_en_shadowed_0_we = (addr_hit[273] & reg_we) & !reg_error;
	assign loc_alert_en_shadowed_0_wd = reg_wdata[0];
	assign loc_alert_en_shadowed_1_re = (addr_hit[274] & reg_re) & !reg_error;
	assign loc_alert_en_shadowed_1_we = (addr_hit[274] & reg_we) & !reg_error;
	assign loc_alert_en_shadowed_1_wd = reg_wdata[0];
	assign loc_alert_en_shadowed_2_re = (addr_hit[275] & reg_re) & !reg_error;
	assign loc_alert_en_shadowed_2_we = (addr_hit[275] & reg_we) & !reg_error;
	assign loc_alert_en_shadowed_2_wd = reg_wdata[0];
	assign loc_alert_en_shadowed_3_re = (addr_hit[276] & reg_re) & !reg_error;
	assign loc_alert_en_shadowed_3_we = (addr_hit[276] & reg_we) & !reg_error;
	assign loc_alert_en_shadowed_3_wd = reg_wdata[0];
	assign loc_alert_en_shadowed_4_re = (addr_hit[277] & reg_re) & !reg_error;
	assign loc_alert_en_shadowed_4_we = (addr_hit[277] & reg_we) & !reg_error;
	assign loc_alert_en_shadowed_4_wd = reg_wdata[0];
	assign loc_alert_en_shadowed_5_re = (addr_hit[278] & reg_re) & !reg_error;
	assign loc_alert_en_shadowed_5_we = (addr_hit[278] & reg_we) & !reg_error;
	assign loc_alert_en_shadowed_5_wd = reg_wdata[0];
	assign loc_alert_en_shadowed_6_re = (addr_hit[279] & reg_re) & !reg_error;
	assign loc_alert_en_shadowed_6_we = (addr_hit[279] & reg_we) & !reg_error;
	assign loc_alert_en_shadowed_6_wd = reg_wdata[0];
	assign loc_alert_class_shadowed_0_re = (addr_hit[280] & reg_re) & !reg_error;
	assign loc_alert_class_shadowed_0_we = (addr_hit[280] & reg_we) & !reg_error;
	assign loc_alert_class_shadowed_0_wd = reg_wdata[1:0];
	assign loc_alert_class_shadowed_1_re = (addr_hit[281] & reg_re) & !reg_error;
	assign loc_alert_class_shadowed_1_we = (addr_hit[281] & reg_we) & !reg_error;
	assign loc_alert_class_shadowed_1_wd = reg_wdata[1:0];
	assign loc_alert_class_shadowed_2_re = (addr_hit[282] & reg_re) & !reg_error;
	assign loc_alert_class_shadowed_2_we = (addr_hit[282] & reg_we) & !reg_error;
	assign loc_alert_class_shadowed_2_wd = reg_wdata[1:0];
	assign loc_alert_class_shadowed_3_re = (addr_hit[283] & reg_re) & !reg_error;
	assign loc_alert_class_shadowed_3_we = (addr_hit[283] & reg_we) & !reg_error;
	assign loc_alert_class_shadowed_3_wd = reg_wdata[1:0];
	assign loc_alert_class_shadowed_4_re = (addr_hit[284] & reg_re) & !reg_error;
	assign loc_alert_class_shadowed_4_we = (addr_hit[284] & reg_we) & !reg_error;
	assign loc_alert_class_shadowed_4_wd = reg_wdata[1:0];
	assign loc_alert_class_shadowed_5_re = (addr_hit[285] & reg_re) & !reg_error;
	assign loc_alert_class_shadowed_5_we = (addr_hit[285] & reg_we) & !reg_error;
	assign loc_alert_class_shadowed_5_wd = reg_wdata[1:0];
	assign loc_alert_class_shadowed_6_re = (addr_hit[286] & reg_re) & !reg_error;
	assign loc_alert_class_shadowed_6_we = (addr_hit[286] & reg_we) & !reg_error;
	assign loc_alert_class_shadowed_6_wd = reg_wdata[1:0];
	assign loc_alert_cause_0_we = (addr_hit[287] & reg_we) & !reg_error;
	assign loc_alert_cause_0_wd = reg_wdata[0];
	assign loc_alert_cause_1_we = (addr_hit[288] & reg_we) & !reg_error;
	assign loc_alert_cause_1_wd = reg_wdata[0];
	assign loc_alert_cause_2_we = (addr_hit[289] & reg_we) & !reg_error;
	assign loc_alert_cause_2_wd = reg_wdata[0];
	assign loc_alert_cause_3_we = (addr_hit[290] & reg_we) & !reg_error;
	assign loc_alert_cause_3_wd = reg_wdata[0];
	assign loc_alert_cause_4_we = (addr_hit[291] & reg_we) & !reg_error;
	assign loc_alert_cause_4_wd = reg_wdata[0];
	assign loc_alert_cause_5_we = (addr_hit[292] & reg_we) & !reg_error;
	assign loc_alert_cause_5_wd = reg_wdata[0];
	assign loc_alert_cause_6_we = (addr_hit[293] & reg_we) & !reg_error;
	assign loc_alert_cause_6_wd = reg_wdata[0];
	assign classa_regwen_we = (addr_hit[294] & reg_we) & !reg_error;
	assign classa_regwen_wd = reg_wdata[0];
	assign classa_ctrl_shadowed_re = (addr_hit[295] & reg_re) & !reg_error;
	assign classa_ctrl_shadowed_we = (addr_hit[295] & reg_we) & !reg_error;
	assign classa_ctrl_shadowed_en_wd = reg_wdata[0];
	assign classa_ctrl_shadowed_lock_wd = reg_wdata[1];
	assign classa_ctrl_shadowed_en_e0_wd = reg_wdata[2];
	assign classa_ctrl_shadowed_en_e1_wd = reg_wdata[3];
	assign classa_ctrl_shadowed_en_e2_wd = reg_wdata[4];
	assign classa_ctrl_shadowed_en_e3_wd = reg_wdata[5];
	assign classa_ctrl_shadowed_map_e0_wd = reg_wdata[7:6];
	assign classa_ctrl_shadowed_map_e1_wd = reg_wdata[9:8];
	assign classa_ctrl_shadowed_map_e2_wd = reg_wdata[11:10];
	assign classa_ctrl_shadowed_map_e3_wd = reg_wdata[13:12];
	assign classa_clr_regwen_we = (addr_hit[296] & reg_we) & !reg_error;
	assign classa_clr_regwen_wd = reg_wdata[0];
	assign classa_clr_shadowed_re = (addr_hit[297] & reg_re) & !reg_error;
	assign classa_clr_shadowed_we = (addr_hit[297] & reg_we) & !reg_error;
	assign classa_clr_shadowed_wd = reg_wdata[0];
	assign classa_accum_cnt_re = (addr_hit[298] & reg_re) & !reg_error;
	assign classa_accum_thresh_shadowed_re = (addr_hit[299] & reg_re) & !reg_error;
	assign classa_accum_thresh_shadowed_we = (addr_hit[299] & reg_we) & !reg_error;
	assign classa_accum_thresh_shadowed_wd = reg_wdata[15:0];
	assign classa_timeout_cyc_shadowed_re = (addr_hit[300] & reg_re) & !reg_error;
	assign classa_timeout_cyc_shadowed_we = (addr_hit[300] & reg_we) & !reg_error;
	assign classa_timeout_cyc_shadowed_wd = reg_wdata[31:0];
	assign classa_crashdump_trigger_shadowed_re = (addr_hit[301] & reg_re) & !reg_error;
	assign classa_crashdump_trigger_shadowed_we = (addr_hit[301] & reg_we) & !reg_error;
	assign classa_crashdump_trigger_shadowed_wd = reg_wdata[1:0];
	assign classa_phase0_cyc_shadowed_re = (addr_hit[302] & reg_re) & !reg_error;
	assign classa_phase0_cyc_shadowed_we = (addr_hit[302] & reg_we) & !reg_error;
	assign classa_phase0_cyc_shadowed_wd = reg_wdata[31:0];
	assign classa_phase1_cyc_shadowed_re = (addr_hit[303] & reg_re) & !reg_error;
	assign classa_phase1_cyc_shadowed_we = (addr_hit[303] & reg_we) & !reg_error;
	assign classa_phase1_cyc_shadowed_wd = reg_wdata[31:0];
	assign classa_phase2_cyc_shadowed_re = (addr_hit[304] & reg_re) & !reg_error;
	assign classa_phase2_cyc_shadowed_we = (addr_hit[304] & reg_we) & !reg_error;
	assign classa_phase2_cyc_shadowed_wd = reg_wdata[31:0];
	assign classa_phase3_cyc_shadowed_re = (addr_hit[305] & reg_re) & !reg_error;
	assign classa_phase3_cyc_shadowed_we = (addr_hit[305] & reg_we) & !reg_error;
	assign classa_phase3_cyc_shadowed_wd = reg_wdata[31:0];
	assign classa_esc_cnt_re = (addr_hit[306] & reg_re) & !reg_error;
	assign classa_state_re = (addr_hit[307] & reg_re) & !reg_error;
	assign classb_regwen_we = (addr_hit[308] & reg_we) & !reg_error;
	assign classb_regwen_wd = reg_wdata[0];
	assign classb_ctrl_shadowed_re = (addr_hit[309] & reg_re) & !reg_error;
	assign classb_ctrl_shadowed_we = (addr_hit[309] & reg_we) & !reg_error;
	assign classb_ctrl_shadowed_en_wd = reg_wdata[0];
	assign classb_ctrl_shadowed_lock_wd = reg_wdata[1];
	assign classb_ctrl_shadowed_en_e0_wd = reg_wdata[2];
	assign classb_ctrl_shadowed_en_e1_wd = reg_wdata[3];
	assign classb_ctrl_shadowed_en_e2_wd = reg_wdata[4];
	assign classb_ctrl_shadowed_en_e3_wd = reg_wdata[5];
	assign classb_ctrl_shadowed_map_e0_wd = reg_wdata[7:6];
	assign classb_ctrl_shadowed_map_e1_wd = reg_wdata[9:8];
	assign classb_ctrl_shadowed_map_e2_wd = reg_wdata[11:10];
	assign classb_ctrl_shadowed_map_e3_wd = reg_wdata[13:12];
	assign classb_clr_regwen_we = (addr_hit[310] & reg_we) & !reg_error;
	assign classb_clr_regwen_wd = reg_wdata[0];
	assign classb_clr_shadowed_re = (addr_hit[311] & reg_re) & !reg_error;
	assign classb_clr_shadowed_we = (addr_hit[311] & reg_we) & !reg_error;
	assign classb_clr_shadowed_wd = reg_wdata[0];
	assign classb_accum_cnt_re = (addr_hit[312] & reg_re) & !reg_error;
	assign classb_accum_thresh_shadowed_re = (addr_hit[313] & reg_re) & !reg_error;
	assign classb_accum_thresh_shadowed_we = (addr_hit[313] & reg_we) & !reg_error;
	assign classb_accum_thresh_shadowed_wd = reg_wdata[15:0];
	assign classb_timeout_cyc_shadowed_re = (addr_hit[314] & reg_re) & !reg_error;
	assign classb_timeout_cyc_shadowed_we = (addr_hit[314] & reg_we) & !reg_error;
	assign classb_timeout_cyc_shadowed_wd = reg_wdata[31:0];
	assign classb_crashdump_trigger_shadowed_re = (addr_hit[315] & reg_re) & !reg_error;
	assign classb_crashdump_trigger_shadowed_we = (addr_hit[315] & reg_we) & !reg_error;
	assign classb_crashdump_trigger_shadowed_wd = reg_wdata[1:0];
	assign classb_phase0_cyc_shadowed_re = (addr_hit[316] & reg_re) & !reg_error;
	assign classb_phase0_cyc_shadowed_we = (addr_hit[316] & reg_we) & !reg_error;
	assign classb_phase0_cyc_shadowed_wd = reg_wdata[31:0];
	assign classb_phase1_cyc_shadowed_re = (addr_hit[317] & reg_re) & !reg_error;
	assign classb_phase1_cyc_shadowed_we = (addr_hit[317] & reg_we) & !reg_error;
	assign classb_phase1_cyc_shadowed_wd = reg_wdata[31:0];
	assign classb_phase2_cyc_shadowed_re = (addr_hit[318] & reg_re) & !reg_error;
	assign classb_phase2_cyc_shadowed_we = (addr_hit[318] & reg_we) & !reg_error;
	assign classb_phase2_cyc_shadowed_wd = reg_wdata[31:0];
	assign classb_phase3_cyc_shadowed_re = (addr_hit[319] & reg_re) & !reg_error;
	assign classb_phase3_cyc_shadowed_we = (addr_hit[319] & reg_we) & !reg_error;
	assign classb_phase3_cyc_shadowed_wd = reg_wdata[31:0];
	assign classb_esc_cnt_re = (addr_hit[320] & reg_re) & !reg_error;
	assign classb_state_re = (addr_hit[321] & reg_re) & !reg_error;
	assign classc_regwen_we = (addr_hit[322] & reg_we) & !reg_error;
	assign classc_regwen_wd = reg_wdata[0];
	assign classc_ctrl_shadowed_re = (addr_hit[323] & reg_re) & !reg_error;
	assign classc_ctrl_shadowed_we = (addr_hit[323] & reg_we) & !reg_error;
	assign classc_ctrl_shadowed_en_wd = reg_wdata[0];
	assign classc_ctrl_shadowed_lock_wd = reg_wdata[1];
	assign classc_ctrl_shadowed_en_e0_wd = reg_wdata[2];
	assign classc_ctrl_shadowed_en_e1_wd = reg_wdata[3];
	assign classc_ctrl_shadowed_en_e2_wd = reg_wdata[4];
	assign classc_ctrl_shadowed_en_e3_wd = reg_wdata[5];
	assign classc_ctrl_shadowed_map_e0_wd = reg_wdata[7:6];
	assign classc_ctrl_shadowed_map_e1_wd = reg_wdata[9:8];
	assign classc_ctrl_shadowed_map_e2_wd = reg_wdata[11:10];
	assign classc_ctrl_shadowed_map_e3_wd = reg_wdata[13:12];
	assign classc_clr_regwen_we = (addr_hit[324] & reg_we) & !reg_error;
	assign classc_clr_regwen_wd = reg_wdata[0];
	assign classc_clr_shadowed_re = (addr_hit[325] & reg_re) & !reg_error;
	assign classc_clr_shadowed_we = (addr_hit[325] & reg_we) & !reg_error;
	assign classc_clr_shadowed_wd = reg_wdata[0];
	assign classc_accum_cnt_re = (addr_hit[326] & reg_re) & !reg_error;
	assign classc_accum_thresh_shadowed_re = (addr_hit[327] & reg_re) & !reg_error;
	assign classc_accum_thresh_shadowed_we = (addr_hit[327] & reg_we) & !reg_error;
	assign classc_accum_thresh_shadowed_wd = reg_wdata[15:0];
	assign classc_timeout_cyc_shadowed_re = (addr_hit[328] & reg_re) & !reg_error;
	assign classc_timeout_cyc_shadowed_we = (addr_hit[328] & reg_we) & !reg_error;
	assign classc_timeout_cyc_shadowed_wd = reg_wdata[31:0];
	assign classc_crashdump_trigger_shadowed_re = (addr_hit[329] & reg_re) & !reg_error;
	assign classc_crashdump_trigger_shadowed_we = (addr_hit[329] & reg_we) & !reg_error;
	assign classc_crashdump_trigger_shadowed_wd = reg_wdata[1:0];
	assign classc_phase0_cyc_shadowed_re = (addr_hit[330] & reg_re) & !reg_error;
	assign classc_phase0_cyc_shadowed_we = (addr_hit[330] & reg_we) & !reg_error;
	assign classc_phase0_cyc_shadowed_wd = reg_wdata[31:0];
	assign classc_phase1_cyc_shadowed_re = (addr_hit[331] & reg_re) & !reg_error;
	assign classc_phase1_cyc_shadowed_we = (addr_hit[331] & reg_we) & !reg_error;
	assign classc_phase1_cyc_shadowed_wd = reg_wdata[31:0];
	assign classc_phase2_cyc_shadowed_re = (addr_hit[332] & reg_re) & !reg_error;
	assign classc_phase2_cyc_shadowed_we = (addr_hit[332] & reg_we) & !reg_error;
	assign classc_phase2_cyc_shadowed_wd = reg_wdata[31:0];
	assign classc_phase3_cyc_shadowed_re = (addr_hit[333] & reg_re) & !reg_error;
	assign classc_phase3_cyc_shadowed_we = (addr_hit[333] & reg_we) & !reg_error;
	assign classc_phase3_cyc_shadowed_wd = reg_wdata[31:0];
	assign classc_esc_cnt_re = (addr_hit[334] & reg_re) & !reg_error;
	assign classc_state_re = (addr_hit[335] & reg_re) & !reg_error;
	assign classd_regwen_we = (addr_hit[336] & reg_we) & !reg_error;
	assign classd_regwen_wd = reg_wdata[0];
	assign classd_ctrl_shadowed_re = (addr_hit[337] & reg_re) & !reg_error;
	assign classd_ctrl_shadowed_we = (addr_hit[337] & reg_we) & !reg_error;
	assign classd_ctrl_shadowed_en_wd = reg_wdata[0];
	assign classd_ctrl_shadowed_lock_wd = reg_wdata[1];
	assign classd_ctrl_shadowed_en_e0_wd = reg_wdata[2];
	assign classd_ctrl_shadowed_en_e1_wd = reg_wdata[3];
	assign classd_ctrl_shadowed_en_e2_wd = reg_wdata[4];
	assign classd_ctrl_shadowed_en_e3_wd = reg_wdata[5];
	assign classd_ctrl_shadowed_map_e0_wd = reg_wdata[7:6];
	assign classd_ctrl_shadowed_map_e1_wd = reg_wdata[9:8];
	assign classd_ctrl_shadowed_map_e2_wd = reg_wdata[11:10];
	assign classd_ctrl_shadowed_map_e3_wd = reg_wdata[13:12];
	assign classd_clr_regwen_we = (addr_hit[338] & reg_we) & !reg_error;
	assign classd_clr_regwen_wd = reg_wdata[0];
	assign classd_clr_shadowed_re = (addr_hit[339] & reg_re) & !reg_error;
	assign classd_clr_shadowed_we = (addr_hit[339] & reg_we) & !reg_error;
	assign classd_clr_shadowed_wd = reg_wdata[0];
	assign classd_accum_cnt_re = (addr_hit[340] & reg_re) & !reg_error;
	assign classd_accum_thresh_shadowed_re = (addr_hit[341] & reg_re) & !reg_error;
	assign classd_accum_thresh_shadowed_we = (addr_hit[341] & reg_we) & !reg_error;
	assign classd_accum_thresh_shadowed_wd = reg_wdata[15:0];
	assign classd_timeout_cyc_shadowed_re = (addr_hit[342] & reg_re) & !reg_error;
	assign classd_timeout_cyc_shadowed_we = (addr_hit[342] & reg_we) & !reg_error;
	assign classd_timeout_cyc_shadowed_wd = reg_wdata[31:0];
	assign classd_crashdump_trigger_shadowed_re = (addr_hit[343] & reg_re) & !reg_error;
	assign classd_crashdump_trigger_shadowed_we = (addr_hit[343] & reg_we) & !reg_error;
	assign classd_crashdump_trigger_shadowed_wd = reg_wdata[1:0];
	assign classd_phase0_cyc_shadowed_re = (addr_hit[344] & reg_re) & !reg_error;
	assign classd_phase0_cyc_shadowed_we = (addr_hit[344] & reg_we) & !reg_error;
	assign classd_phase0_cyc_shadowed_wd = reg_wdata[31:0];
	assign classd_phase1_cyc_shadowed_re = (addr_hit[345] & reg_re) & !reg_error;
	assign classd_phase1_cyc_shadowed_we = (addr_hit[345] & reg_we) & !reg_error;
	assign classd_phase1_cyc_shadowed_wd = reg_wdata[31:0];
	assign classd_phase2_cyc_shadowed_re = (addr_hit[346] & reg_re) & !reg_error;
	assign classd_phase2_cyc_shadowed_we = (addr_hit[346] & reg_we) & !reg_error;
	assign classd_phase2_cyc_shadowed_wd = reg_wdata[31:0];
	assign classd_phase3_cyc_shadowed_re = (addr_hit[347] & reg_re) & !reg_error;
	assign classd_phase3_cyc_shadowed_we = (addr_hit[347] & reg_we) & !reg_error;
	assign classd_phase3_cyc_shadowed_wd = reg_wdata[31:0];
	assign classd_esc_cnt_re = (addr_hit[348] & reg_re) & !reg_error;
	assign classd_state_re = (addr_hit[349] & reg_re) & !reg_error;
	always @(*) begin
		reg_we_check = 1'sb0;
		reg_we_check[0] = intr_state_we;
		reg_we_check[1] = intr_enable_we;
		reg_we_check[2] = intr_test_we;
		reg_we_check[3] = ping_timer_regwen_we;
		reg_we_check[4] = ping_timeout_cyc_shadowed_gated_we;
		reg_we_check[5] = ping_timer_en_shadowed_gated_we;
		reg_we_check[6] = alert_regwen_0_we;
		reg_we_check[7] = alert_regwen_1_we;
		reg_we_check[8] = alert_regwen_2_we;
		reg_we_check[9] = alert_regwen_3_we;
		reg_we_check[10] = alert_regwen_4_we;
		reg_we_check[11] = alert_regwen_5_we;
		reg_we_check[12] = alert_regwen_6_we;
		reg_we_check[13] = alert_regwen_7_we;
		reg_we_check[14] = alert_regwen_8_we;
		reg_we_check[15] = alert_regwen_9_we;
		reg_we_check[16] = alert_regwen_10_we;
		reg_we_check[17] = alert_regwen_11_we;
		reg_we_check[18] = alert_regwen_12_we;
		reg_we_check[19] = alert_regwen_13_we;
		reg_we_check[20] = alert_regwen_14_we;
		reg_we_check[21] = alert_regwen_15_we;
		reg_we_check[22] = alert_regwen_16_we;
		reg_we_check[23] = alert_regwen_17_we;
		reg_we_check[24] = alert_regwen_18_we;
		reg_we_check[25] = alert_regwen_19_we;
		reg_we_check[26] = alert_regwen_20_we;
		reg_we_check[27] = alert_regwen_21_we;
		reg_we_check[28] = alert_regwen_22_we;
		reg_we_check[29] = alert_regwen_23_we;
		reg_we_check[30] = alert_regwen_24_we;
		reg_we_check[31] = alert_regwen_25_we;
		reg_we_check[32] = alert_regwen_26_we;
		reg_we_check[33] = alert_regwen_27_we;
		reg_we_check[34] = alert_regwen_28_we;
		reg_we_check[35] = alert_regwen_29_we;
		reg_we_check[36] = alert_regwen_30_we;
		reg_we_check[37] = alert_regwen_31_we;
		reg_we_check[38] = alert_regwen_32_we;
		reg_we_check[39] = alert_regwen_33_we;
		reg_we_check[40] = alert_regwen_34_we;
		reg_we_check[41] = alert_regwen_35_we;
		reg_we_check[42] = alert_regwen_36_we;
		reg_we_check[43] = alert_regwen_37_we;
		reg_we_check[44] = alert_regwen_38_we;
		reg_we_check[45] = alert_regwen_39_we;
		reg_we_check[46] = alert_regwen_40_we;
		reg_we_check[47] = alert_regwen_41_we;
		reg_we_check[48] = alert_regwen_42_we;
		reg_we_check[49] = alert_regwen_43_we;
		reg_we_check[50] = alert_regwen_44_we;
		reg_we_check[51] = alert_regwen_45_we;
		reg_we_check[52] = alert_regwen_46_we;
		reg_we_check[53] = alert_regwen_47_we;
		reg_we_check[54] = alert_regwen_48_we;
		reg_we_check[55] = alert_regwen_49_we;
		reg_we_check[56] = alert_regwen_50_we;
		reg_we_check[57] = alert_regwen_51_we;
		reg_we_check[58] = alert_regwen_52_we;
		reg_we_check[59] = alert_regwen_53_we;
		reg_we_check[60] = alert_regwen_54_we;
		reg_we_check[61] = alert_regwen_55_we;
		reg_we_check[62] = alert_regwen_56_we;
		reg_we_check[63] = alert_regwen_57_we;
		reg_we_check[64] = alert_regwen_58_we;
		reg_we_check[65] = alert_regwen_59_we;
		reg_we_check[66] = alert_regwen_60_we;
		reg_we_check[67] = alert_regwen_61_we;
		reg_we_check[68] = alert_regwen_62_we;
		reg_we_check[69] = alert_regwen_63_we;
		reg_we_check[70] = alert_regwen_64_we;
		reg_we_check[71] = alert_en_shadowed_0_gated_we;
		reg_we_check[72] = alert_en_shadowed_1_gated_we;
		reg_we_check[73] = alert_en_shadowed_2_gated_we;
		reg_we_check[74] = alert_en_shadowed_3_gated_we;
		reg_we_check[75] = alert_en_shadowed_4_gated_we;
		reg_we_check[76] = alert_en_shadowed_5_gated_we;
		reg_we_check[77] = alert_en_shadowed_6_gated_we;
		reg_we_check[78] = alert_en_shadowed_7_gated_we;
		reg_we_check[79] = alert_en_shadowed_8_gated_we;
		reg_we_check[80] = alert_en_shadowed_9_gated_we;
		reg_we_check[81] = alert_en_shadowed_10_gated_we;
		reg_we_check[82] = alert_en_shadowed_11_gated_we;
		reg_we_check[83] = alert_en_shadowed_12_gated_we;
		reg_we_check[84] = alert_en_shadowed_13_gated_we;
		reg_we_check[85] = alert_en_shadowed_14_gated_we;
		reg_we_check[86] = alert_en_shadowed_15_gated_we;
		reg_we_check[87] = alert_en_shadowed_16_gated_we;
		reg_we_check[88] = alert_en_shadowed_17_gated_we;
		reg_we_check[89] = alert_en_shadowed_18_gated_we;
		reg_we_check[90] = alert_en_shadowed_19_gated_we;
		reg_we_check[91] = alert_en_shadowed_20_gated_we;
		reg_we_check[92] = alert_en_shadowed_21_gated_we;
		reg_we_check[93] = alert_en_shadowed_22_gated_we;
		reg_we_check[94] = alert_en_shadowed_23_gated_we;
		reg_we_check[95] = alert_en_shadowed_24_gated_we;
		reg_we_check[96] = alert_en_shadowed_25_gated_we;
		reg_we_check[97] = alert_en_shadowed_26_gated_we;
		reg_we_check[98] = alert_en_shadowed_27_gated_we;
		reg_we_check[99] = alert_en_shadowed_28_gated_we;
		reg_we_check[100] = alert_en_shadowed_29_gated_we;
		reg_we_check[101] = alert_en_shadowed_30_gated_we;
		reg_we_check[102] = alert_en_shadowed_31_gated_we;
		reg_we_check[103] = alert_en_shadowed_32_gated_we;
		reg_we_check[104] = alert_en_shadowed_33_gated_we;
		reg_we_check[105] = alert_en_shadowed_34_gated_we;
		reg_we_check[106] = alert_en_shadowed_35_gated_we;
		reg_we_check[107] = alert_en_shadowed_36_gated_we;
		reg_we_check[108] = alert_en_shadowed_37_gated_we;
		reg_we_check[109] = alert_en_shadowed_38_gated_we;
		reg_we_check[110] = alert_en_shadowed_39_gated_we;
		reg_we_check[111] = alert_en_shadowed_40_gated_we;
		reg_we_check[112] = alert_en_shadowed_41_gated_we;
		reg_we_check[113] = alert_en_shadowed_42_gated_we;
		reg_we_check[114] = alert_en_shadowed_43_gated_we;
		reg_we_check[115] = alert_en_shadowed_44_gated_we;
		reg_we_check[116] = alert_en_shadowed_45_gated_we;
		reg_we_check[117] = alert_en_shadowed_46_gated_we;
		reg_we_check[118] = alert_en_shadowed_47_gated_we;
		reg_we_check[119] = alert_en_shadowed_48_gated_we;
		reg_we_check[120] = alert_en_shadowed_49_gated_we;
		reg_we_check[121] = alert_en_shadowed_50_gated_we;
		reg_we_check[122] = alert_en_shadowed_51_gated_we;
		reg_we_check[123] = alert_en_shadowed_52_gated_we;
		reg_we_check[124] = alert_en_shadowed_53_gated_we;
		reg_we_check[125] = alert_en_shadowed_54_gated_we;
		reg_we_check[126] = alert_en_shadowed_55_gated_we;
		reg_we_check[127] = alert_en_shadowed_56_gated_we;
		reg_we_check[128] = alert_en_shadowed_57_gated_we;
		reg_we_check[129] = alert_en_shadowed_58_gated_we;
		reg_we_check[130] = alert_en_shadowed_59_gated_we;
		reg_we_check[131] = alert_en_shadowed_60_gated_we;
		reg_we_check[132] = alert_en_shadowed_61_gated_we;
		reg_we_check[133] = alert_en_shadowed_62_gated_we;
		reg_we_check[134] = alert_en_shadowed_63_gated_we;
		reg_we_check[135] = alert_en_shadowed_64_gated_we;
		reg_we_check[136] = alert_class_shadowed_0_gated_we;
		reg_we_check[137] = alert_class_shadowed_1_gated_we;
		reg_we_check[138] = alert_class_shadowed_2_gated_we;
		reg_we_check[139] = alert_class_shadowed_3_gated_we;
		reg_we_check[140] = alert_class_shadowed_4_gated_we;
		reg_we_check[141] = alert_class_shadowed_5_gated_we;
		reg_we_check[142] = alert_class_shadowed_6_gated_we;
		reg_we_check[143] = alert_class_shadowed_7_gated_we;
		reg_we_check[144] = alert_class_shadowed_8_gated_we;
		reg_we_check[145] = alert_class_shadowed_9_gated_we;
		reg_we_check[146] = alert_class_shadowed_10_gated_we;
		reg_we_check[147] = alert_class_shadowed_11_gated_we;
		reg_we_check[148] = alert_class_shadowed_12_gated_we;
		reg_we_check[149] = alert_class_shadowed_13_gated_we;
		reg_we_check[150] = alert_class_shadowed_14_gated_we;
		reg_we_check[151] = alert_class_shadowed_15_gated_we;
		reg_we_check[152] = alert_class_shadowed_16_gated_we;
		reg_we_check[153] = alert_class_shadowed_17_gated_we;
		reg_we_check[154] = alert_class_shadowed_18_gated_we;
		reg_we_check[155] = alert_class_shadowed_19_gated_we;
		reg_we_check[156] = alert_class_shadowed_20_gated_we;
		reg_we_check[157] = alert_class_shadowed_21_gated_we;
		reg_we_check[158] = alert_class_shadowed_22_gated_we;
		reg_we_check[159] = alert_class_shadowed_23_gated_we;
		reg_we_check[160] = alert_class_shadowed_24_gated_we;
		reg_we_check[161] = alert_class_shadowed_25_gated_we;
		reg_we_check[162] = alert_class_shadowed_26_gated_we;
		reg_we_check[163] = alert_class_shadowed_27_gated_we;
		reg_we_check[164] = alert_class_shadowed_28_gated_we;
		reg_we_check[165] = alert_class_shadowed_29_gated_we;
		reg_we_check[166] = alert_class_shadowed_30_gated_we;
		reg_we_check[167] = alert_class_shadowed_31_gated_we;
		reg_we_check[168] = alert_class_shadowed_32_gated_we;
		reg_we_check[169] = alert_class_shadowed_33_gated_we;
		reg_we_check[170] = alert_class_shadowed_34_gated_we;
		reg_we_check[171] = alert_class_shadowed_35_gated_we;
		reg_we_check[172] = alert_class_shadowed_36_gated_we;
		reg_we_check[173] = alert_class_shadowed_37_gated_we;
		reg_we_check[174] = alert_class_shadowed_38_gated_we;
		reg_we_check[175] = alert_class_shadowed_39_gated_we;
		reg_we_check[176] = alert_class_shadowed_40_gated_we;
		reg_we_check[177] = alert_class_shadowed_41_gated_we;
		reg_we_check[178] = alert_class_shadowed_42_gated_we;
		reg_we_check[179] = alert_class_shadowed_43_gated_we;
		reg_we_check[180] = alert_class_shadowed_44_gated_we;
		reg_we_check[181] = alert_class_shadowed_45_gated_we;
		reg_we_check[182] = alert_class_shadowed_46_gated_we;
		reg_we_check[183] = alert_class_shadowed_47_gated_we;
		reg_we_check[184] = alert_class_shadowed_48_gated_we;
		reg_we_check[185] = alert_class_shadowed_49_gated_we;
		reg_we_check[186] = alert_class_shadowed_50_gated_we;
		reg_we_check[187] = alert_class_shadowed_51_gated_we;
		reg_we_check[188] = alert_class_shadowed_52_gated_we;
		reg_we_check[189] = alert_class_shadowed_53_gated_we;
		reg_we_check[190] = alert_class_shadowed_54_gated_we;
		reg_we_check[191] = alert_class_shadowed_55_gated_we;
		reg_we_check[192] = alert_class_shadowed_56_gated_we;
		reg_we_check[193] = alert_class_shadowed_57_gated_we;
		reg_we_check[194] = alert_class_shadowed_58_gated_we;
		reg_we_check[195] = alert_class_shadowed_59_gated_we;
		reg_we_check[196] = alert_class_shadowed_60_gated_we;
		reg_we_check[197] = alert_class_shadowed_61_gated_we;
		reg_we_check[198] = alert_class_shadowed_62_gated_we;
		reg_we_check[199] = alert_class_shadowed_63_gated_we;
		reg_we_check[200] = alert_class_shadowed_64_gated_we;
		reg_we_check[201] = alert_cause_0_we;
		reg_we_check[202] = alert_cause_1_we;
		reg_we_check[203] = alert_cause_2_we;
		reg_we_check[204] = alert_cause_3_we;
		reg_we_check[205] = alert_cause_4_we;
		reg_we_check[206] = alert_cause_5_we;
		reg_we_check[207] = alert_cause_6_we;
		reg_we_check[208] = alert_cause_7_we;
		reg_we_check[209] = alert_cause_8_we;
		reg_we_check[210] = alert_cause_9_we;
		reg_we_check[211] = alert_cause_10_we;
		reg_we_check[212] = alert_cause_11_we;
		reg_we_check[213] = alert_cause_12_we;
		reg_we_check[214] = alert_cause_13_we;
		reg_we_check[215] = alert_cause_14_we;
		reg_we_check[216] = alert_cause_15_we;
		reg_we_check[217] = alert_cause_16_we;
		reg_we_check[218] = alert_cause_17_we;
		reg_we_check[219] = alert_cause_18_we;
		reg_we_check[220] = alert_cause_19_we;
		reg_we_check[221] = alert_cause_20_we;
		reg_we_check[222] = alert_cause_21_we;
		reg_we_check[223] = alert_cause_22_we;
		reg_we_check[224] = alert_cause_23_we;
		reg_we_check[225] = alert_cause_24_we;
		reg_we_check[226] = alert_cause_25_we;
		reg_we_check[227] = alert_cause_26_we;
		reg_we_check[228] = alert_cause_27_we;
		reg_we_check[229] = alert_cause_28_we;
		reg_we_check[230] = alert_cause_29_we;
		reg_we_check[231] = alert_cause_30_we;
		reg_we_check[232] = alert_cause_31_we;
		reg_we_check[233] = alert_cause_32_we;
		reg_we_check[234] = alert_cause_33_we;
		reg_we_check[235] = alert_cause_34_we;
		reg_we_check[236] = alert_cause_35_we;
		reg_we_check[237] = alert_cause_36_we;
		reg_we_check[238] = alert_cause_37_we;
		reg_we_check[239] = alert_cause_38_we;
		reg_we_check[240] = alert_cause_39_we;
		reg_we_check[241] = alert_cause_40_we;
		reg_we_check[242] = alert_cause_41_we;
		reg_we_check[243] = alert_cause_42_we;
		reg_we_check[244] = alert_cause_43_we;
		reg_we_check[245] = alert_cause_44_we;
		reg_we_check[246] = alert_cause_45_we;
		reg_we_check[247] = alert_cause_46_we;
		reg_we_check[248] = alert_cause_47_we;
		reg_we_check[249] = alert_cause_48_we;
		reg_we_check[250] = alert_cause_49_we;
		reg_we_check[251] = alert_cause_50_we;
		reg_we_check[252] = alert_cause_51_we;
		reg_we_check[253] = alert_cause_52_we;
		reg_we_check[254] = alert_cause_53_we;
		reg_we_check[255] = alert_cause_54_we;
		reg_we_check[256] = alert_cause_55_we;
		reg_we_check[257] = alert_cause_56_we;
		reg_we_check[258] = alert_cause_57_we;
		reg_we_check[259] = alert_cause_58_we;
		reg_we_check[260] = alert_cause_59_we;
		reg_we_check[261] = alert_cause_60_we;
		reg_we_check[262] = alert_cause_61_we;
		reg_we_check[263] = alert_cause_62_we;
		reg_we_check[264] = alert_cause_63_we;
		reg_we_check[265] = alert_cause_64_we;
		reg_we_check[266] = loc_alert_regwen_0_we;
		reg_we_check[267] = loc_alert_regwen_1_we;
		reg_we_check[268] = loc_alert_regwen_2_we;
		reg_we_check[269] = loc_alert_regwen_3_we;
		reg_we_check[270] = loc_alert_regwen_4_we;
		reg_we_check[271] = loc_alert_regwen_5_we;
		reg_we_check[272] = loc_alert_regwen_6_we;
		reg_we_check[273] = loc_alert_en_shadowed_0_gated_we;
		reg_we_check[274] = loc_alert_en_shadowed_1_gated_we;
		reg_we_check[275] = loc_alert_en_shadowed_2_gated_we;
		reg_we_check[276] = loc_alert_en_shadowed_3_gated_we;
		reg_we_check[277] = loc_alert_en_shadowed_4_gated_we;
		reg_we_check[278] = loc_alert_en_shadowed_5_gated_we;
		reg_we_check[279] = loc_alert_en_shadowed_6_gated_we;
		reg_we_check[280] = loc_alert_class_shadowed_0_gated_we;
		reg_we_check[281] = loc_alert_class_shadowed_1_gated_we;
		reg_we_check[282] = loc_alert_class_shadowed_2_gated_we;
		reg_we_check[283] = loc_alert_class_shadowed_3_gated_we;
		reg_we_check[284] = loc_alert_class_shadowed_4_gated_we;
		reg_we_check[285] = loc_alert_class_shadowed_5_gated_we;
		reg_we_check[286] = loc_alert_class_shadowed_6_gated_we;
		reg_we_check[287] = loc_alert_cause_0_we;
		reg_we_check[288] = loc_alert_cause_1_we;
		reg_we_check[289] = loc_alert_cause_2_we;
		reg_we_check[290] = loc_alert_cause_3_we;
		reg_we_check[291] = loc_alert_cause_4_we;
		reg_we_check[292] = loc_alert_cause_5_we;
		reg_we_check[293] = loc_alert_cause_6_we;
		reg_we_check[294] = classa_regwen_we;
		reg_we_check[295] = classa_ctrl_shadowed_gated_we;
		reg_we_check[296] = classa_clr_regwen_we;
		reg_we_check[297] = classa_clr_shadowed_gated_we;
		reg_we_check[298] = 1'b0;
		reg_we_check[299] = classa_accum_thresh_shadowed_gated_we;
		reg_we_check[300] = classa_timeout_cyc_shadowed_gated_we;
		reg_we_check[301] = classa_crashdump_trigger_shadowed_gated_we;
		reg_we_check[302] = classa_phase0_cyc_shadowed_gated_we;
		reg_we_check[303] = classa_phase1_cyc_shadowed_gated_we;
		reg_we_check[304] = classa_phase2_cyc_shadowed_gated_we;
		reg_we_check[305] = classa_phase3_cyc_shadowed_gated_we;
		reg_we_check[306] = 1'b0;
		reg_we_check[307] = 1'b0;
		reg_we_check[308] = classb_regwen_we;
		reg_we_check[309] = classb_ctrl_shadowed_gated_we;
		reg_we_check[310] = classb_clr_regwen_we;
		reg_we_check[311] = classb_clr_shadowed_gated_we;
		reg_we_check[312] = 1'b0;
		reg_we_check[313] = classb_accum_thresh_shadowed_gated_we;
		reg_we_check[314] = classb_timeout_cyc_shadowed_gated_we;
		reg_we_check[315] = classb_crashdump_trigger_shadowed_gated_we;
		reg_we_check[316] = classb_phase0_cyc_shadowed_gated_we;
		reg_we_check[317] = classb_phase1_cyc_shadowed_gated_we;
		reg_we_check[318] = classb_phase2_cyc_shadowed_gated_we;
		reg_we_check[319] = classb_phase3_cyc_shadowed_gated_we;
		reg_we_check[320] = 1'b0;
		reg_we_check[321] = 1'b0;
		reg_we_check[322] = classc_regwen_we;
		reg_we_check[323] = classc_ctrl_shadowed_gated_we;
		reg_we_check[324] = classc_clr_regwen_we;
		reg_we_check[325] = classc_clr_shadowed_gated_we;
		reg_we_check[326] = 1'b0;
		reg_we_check[327] = classc_accum_thresh_shadowed_gated_we;
		reg_we_check[328] = classc_timeout_cyc_shadowed_gated_we;
		reg_we_check[329] = classc_crashdump_trigger_shadowed_gated_we;
		reg_we_check[330] = classc_phase0_cyc_shadowed_gated_we;
		reg_we_check[331] = classc_phase1_cyc_shadowed_gated_we;
		reg_we_check[332] = classc_phase2_cyc_shadowed_gated_we;
		reg_we_check[333] = classc_phase3_cyc_shadowed_gated_we;
		reg_we_check[334] = 1'b0;
		reg_we_check[335] = 1'b0;
		reg_we_check[336] = classd_regwen_we;
		reg_we_check[337] = classd_ctrl_shadowed_gated_we;
		reg_we_check[338] = classd_clr_regwen_we;
		reg_we_check[339] = classd_clr_shadowed_gated_we;
		reg_we_check[340] = 1'b0;
		reg_we_check[341] = classd_accum_thresh_shadowed_gated_we;
		reg_we_check[342] = classd_timeout_cyc_shadowed_gated_we;
		reg_we_check[343] = classd_crashdump_trigger_shadowed_gated_we;
		reg_we_check[344] = classd_phase0_cyc_shadowed_gated_we;
		reg_we_check[345] = classd_phase1_cyc_shadowed_gated_we;
		reg_we_check[346] = classd_phase2_cyc_shadowed_gated_we;
		reg_we_check[347] = classd_phase3_cyc_shadowed_gated_we;
		reg_we_check[348] = 1'b0;
		reg_we_check[349] = 1'b0;
	end
	always @(*) begin
		reg_rdata_next = 1'sb0;
		case (1'b1)
			addr_hit[0]: begin
				reg_rdata_next[0] = intr_state_classa_qs;
				reg_rdata_next[1] = intr_state_classb_qs;
				reg_rdata_next[2] = intr_state_classc_qs;
				reg_rdata_next[3] = intr_state_classd_qs;
			end
			addr_hit[1]: begin
				reg_rdata_next[0] = intr_enable_classa_qs;
				reg_rdata_next[1] = intr_enable_classb_qs;
				reg_rdata_next[2] = intr_enable_classc_qs;
				reg_rdata_next[3] = intr_enable_classd_qs;
			end
			addr_hit[2]: begin
				reg_rdata_next[0] = 1'sb0;
				reg_rdata_next[1] = 1'sb0;
				reg_rdata_next[2] = 1'sb0;
				reg_rdata_next[3] = 1'sb0;
			end
			addr_hit[3]: reg_rdata_next[0] = ping_timer_regwen_qs;
			addr_hit[4]: reg_rdata_next[15:0] = ping_timeout_cyc_shadowed_qs;
			addr_hit[5]: reg_rdata_next[0] = ping_timer_en_shadowed_qs;
			addr_hit[6]: reg_rdata_next[0] = alert_regwen_0_qs;
			addr_hit[7]: reg_rdata_next[0] = alert_regwen_1_qs;
			addr_hit[8]: reg_rdata_next[0] = alert_regwen_2_qs;
			addr_hit[9]: reg_rdata_next[0] = alert_regwen_3_qs;
			addr_hit[10]: reg_rdata_next[0] = alert_regwen_4_qs;
			addr_hit[11]: reg_rdata_next[0] = alert_regwen_5_qs;
			addr_hit[12]: reg_rdata_next[0] = alert_regwen_6_qs;
			addr_hit[13]: reg_rdata_next[0] = alert_regwen_7_qs;
			addr_hit[14]: reg_rdata_next[0] = alert_regwen_8_qs;
			addr_hit[15]: reg_rdata_next[0] = alert_regwen_9_qs;
			addr_hit[16]: reg_rdata_next[0] = alert_regwen_10_qs;
			addr_hit[17]: reg_rdata_next[0] = alert_regwen_11_qs;
			addr_hit[18]: reg_rdata_next[0] = alert_regwen_12_qs;
			addr_hit[19]: reg_rdata_next[0] = alert_regwen_13_qs;
			addr_hit[20]: reg_rdata_next[0] = alert_regwen_14_qs;
			addr_hit[21]: reg_rdata_next[0] = alert_regwen_15_qs;
			addr_hit[22]: reg_rdata_next[0] = alert_regwen_16_qs;
			addr_hit[23]: reg_rdata_next[0] = alert_regwen_17_qs;
			addr_hit[24]: reg_rdata_next[0] = alert_regwen_18_qs;
			addr_hit[25]: reg_rdata_next[0] = alert_regwen_19_qs;
			addr_hit[26]: reg_rdata_next[0] = alert_regwen_20_qs;
			addr_hit[27]: reg_rdata_next[0] = alert_regwen_21_qs;
			addr_hit[28]: reg_rdata_next[0] = alert_regwen_22_qs;
			addr_hit[29]: reg_rdata_next[0] = alert_regwen_23_qs;
			addr_hit[30]: reg_rdata_next[0] = alert_regwen_24_qs;
			addr_hit[31]: reg_rdata_next[0] = alert_regwen_25_qs;
			addr_hit[32]: reg_rdata_next[0] = alert_regwen_26_qs;
			addr_hit[33]: reg_rdata_next[0] = alert_regwen_27_qs;
			addr_hit[34]: reg_rdata_next[0] = alert_regwen_28_qs;
			addr_hit[35]: reg_rdata_next[0] = alert_regwen_29_qs;
			addr_hit[36]: reg_rdata_next[0] = alert_regwen_30_qs;
			addr_hit[37]: reg_rdata_next[0] = alert_regwen_31_qs;
			addr_hit[38]: reg_rdata_next[0] = alert_regwen_32_qs;
			addr_hit[39]: reg_rdata_next[0] = alert_regwen_33_qs;
			addr_hit[40]: reg_rdata_next[0] = alert_regwen_34_qs;
			addr_hit[41]: reg_rdata_next[0] = alert_regwen_35_qs;
			addr_hit[42]: reg_rdata_next[0] = alert_regwen_36_qs;
			addr_hit[43]: reg_rdata_next[0] = alert_regwen_37_qs;
			addr_hit[44]: reg_rdata_next[0] = alert_regwen_38_qs;
			addr_hit[45]: reg_rdata_next[0] = alert_regwen_39_qs;
			addr_hit[46]: reg_rdata_next[0] = alert_regwen_40_qs;
			addr_hit[47]: reg_rdata_next[0] = alert_regwen_41_qs;
			addr_hit[48]: reg_rdata_next[0] = alert_regwen_42_qs;
			addr_hit[49]: reg_rdata_next[0] = alert_regwen_43_qs;
			addr_hit[50]: reg_rdata_next[0] = alert_regwen_44_qs;
			addr_hit[51]: reg_rdata_next[0] = alert_regwen_45_qs;
			addr_hit[52]: reg_rdata_next[0] = alert_regwen_46_qs;
			addr_hit[53]: reg_rdata_next[0] = alert_regwen_47_qs;
			addr_hit[54]: reg_rdata_next[0] = alert_regwen_48_qs;
			addr_hit[55]: reg_rdata_next[0] = alert_regwen_49_qs;
			addr_hit[56]: reg_rdata_next[0] = alert_regwen_50_qs;
			addr_hit[57]: reg_rdata_next[0] = alert_regwen_51_qs;
			addr_hit[58]: reg_rdata_next[0] = alert_regwen_52_qs;
			addr_hit[59]: reg_rdata_next[0] = alert_regwen_53_qs;
			addr_hit[60]: reg_rdata_next[0] = alert_regwen_54_qs;
			addr_hit[61]: reg_rdata_next[0] = alert_regwen_55_qs;
			addr_hit[62]: reg_rdata_next[0] = alert_regwen_56_qs;
			addr_hit[63]: reg_rdata_next[0] = alert_regwen_57_qs;
			addr_hit[64]: reg_rdata_next[0] = alert_regwen_58_qs;
			addr_hit[65]: reg_rdata_next[0] = alert_regwen_59_qs;
			addr_hit[66]: reg_rdata_next[0] = alert_regwen_60_qs;
			addr_hit[67]: reg_rdata_next[0] = alert_regwen_61_qs;
			addr_hit[68]: reg_rdata_next[0] = alert_regwen_62_qs;
			addr_hit[69]: reg_rdata_next[0] = alert_regwen_63_qs;
			addr_hit[70]: reg_rdata_next[0] = alert_regwen_64_qs;
			addr_hit[71]: reg_rdata_next[0] = alert_en_shadowed_0_qs;
			addr_hit[72]: reg_rdata_next[0] = alert_en_shadowed_1_qs;
			addr_hit[73]: reg_rdata_next[0] = alert_en_shadowed_2_qs;
			addr_hit[74]: reg_rdata_next[0] = alert_en_shadowed_3_qs;
			addr_hit[75]: reg_rdata_next[0] = alert_en_shadowed_4_qs;
			addr_hit[76]: reg_rdata_next[0] = alert_en_shadowed_5_qs;
			addr_hit[77]: reg_rdata_next[0] = alert_en_shadowed_6_qs;
			addr_hit[78]: reg_rdata_next[0] = alert_en_shadowed_7_qs;
			addr_hit[79]: reg_rdata_next[0] = alert_en_shadowed_8_qs;
			addr_hit[80]: reg_rdata_next[0] = alert_en_shadowed_9_qs;
			addr_hit[81]: reg_rdata_next[0] = alert_en_shadowed_10_qs;
			addr_hit[82]: reg_rdata_next[0] = alert_en_shadowed_11_qs;
			addr_hit[83]: reg_rdata_next[0] = alert_en_shadowed_12_qs;
			addr_hit[84]: reg_rdata_next[0] = alert_en_shadowed_13_qs;
			addr_hit[85]: reg_rdata_next[0] = alert_en_shadowed_14_qs;
			addr_hit[86]: reg_rdata_next[0] = alert_en_shadowed_15_qs;
			addr_hit[87]: reg_rdata_next[0] = alert_en_shadowed_16_qs;
			addr_hit[88]: reg_rdata_next[0] = alert_en_shadowed_17_qs;
			addr_hit[89]: reg_rdata_next[0] = alert_en_shadowed_18_qs;
			addr_hit[90]: reg_rdata_next[0] = alert_en_shadowed_19_qs;
			addr_hit[91]: reg_rdata_next[0] = alert_en_shadowed_20_qs;
			addr_hit[92]: reg_rdata_next[0] = alert_en_shadowed_21_qs;
			addr_hit[93]: reg_rdata_next[0] = alert_en_shadowed_22_qs;
			addr_hit[94]: reg_rdata_next[0] = alert_en_shadowed_23_qs;
			addr_hit[95]: reg_rdata_next[0] = alert_en_shadowed_24_qs;
			addr_hit[96]: reg_rdata_next[0] = alert_en_shadowed_25_qs;
			addr_hit[97]: reg_rdata_next[0] = alert_en_shadowed_26_qs;
			addr_hit[98]: reg_rdata_next[0] = alert_en_shadowed_27_qs;
			addr_hit[99]: reg_rdata_next[0] = alert_en_shadowed_28_qs;
			addr_hit[100]: reg_rdata_next[0] = alert_en_shadowed_29_qs;
			addr_hit[101]: reg_rdata_next[0] = alert_en_shadowed_30_qs;
			addr_hit[102]: reg_rdata_next[0] = alert_en_shadowed_31_qs;
			addr_hit[103]: reg_rdata_next[0] = alert_en_shadowed_32_qs;
			addr_hit[104]: reg_rdata_next[0] = alert_en_shadowed_33_qs;
			addr_hit[105]: reg_rdata_next[0] = alert_en_shadowed_34_qs;
			addr_hit[106]: reg_rdata_next[0] = alert_en_shadowed_35_qs;
			addr_hit[107]: reg_rdata_next[0] = alert_en_shadowed_36_qs;
			addr_hit[108]: reg_rdata_next[0] = alert_en_shadowed_37_qs;
			addr_hit[109]: reg_rdata_next[0] = alert_en_shadowed_38_qs;
			addr_hit[110]: reg_rdata_next[0] = alert_en_shadowed_39_qs;
			addr_hit[111]: reg_rdata_next[0] = alert_en_shadowed_40_qs;
			addr_hit[112]: reg_rdata_next[0] = alert_en_shadowed_41_qs;
			addr_hit[113]: reg_rdata_next[0] = alert_en_shadowed_42_qs;
			addr_hit[114]: reg_rdata_next[0] = alert_en_shadowed_43_qs;
			addr_hit[115]: reg_rdata_next[0] = alert_en_shadowed_44_qs;
			addr_hit[116]: reg_rdata_next[0] = alert_en_shadowed_45_qs;
			addr_hit[117]: reg_rdata_next[0] = alert_en_shadowed_46_qs;
			addr_hit[118]: reg_rdata_next[0] = alert_en_shadowed_47_qs;
			addr_hit[119]: reg_rdata_next[0] = alert_en_shadowed_48_qs;
			addr_hit[120]: reg_rdata_next[0] = alert_en_shadowed_49_qs;
			addr_hit[121]: reg_rdata_next[0] = alert_en_shadowed_50_qs;
			addr_hit[122]: reg_rdata_next[0] = alert_en_shadowed_51_qs;
			addr_hit[123]: reg_rdata_next[0] = alert_en_shadowed_52_qs;
			addr_hit[124]: reg_rdata_next[0] = alert_en_shadowed_53_qs;
			addr_hit[125]: reg_rdata_next[0] = alert_en_shadowed_54_qs;
			addr_hit[126]: reg_rdata_next[0] = alert_en_shadowed_55_qs;
			addr_hit[127]: reg_rdata_next[0] = alert_en_shadowed_56_qs;
			addr_hit[128]: reg_rdata_next[0] = alert_en_shadowed_57_qs;
			addr_hit[129]: reg_rdata_next[0] = alert_en_shadowed_58_qs;
			addr_hit[130]: reg_rdata_next[0] = alert_en_shadowed_59_qs;
			addr_hit[131]: reg_rdata_next[0] = alert_en_shadowed_60_qs;
			addr_hit[132]: reg_rdata_next[0] = alert_en_shadowed_61_qs;
			addr_hit[133]: reg_rdata_next[0] = alert_en_shadowed_62_qs;
			addr_hit[134]: reg_rdata_next[0] = alert_en_shadowed_63_qs;
			addr_hit[135]: reg_rdata_next[0] = alert_en_shadowed_64_qs;
			addr_hit[136]: reg_rdata_next[1:0] = alert_class_shadowed_0_qs;
			addr_hit[137]: reg_rdata_next[1:0] = alert_class_shadowed_1_qs;
			addr_hit[138]: reg_rdata_next[1:0] = alert_class_shadowed_2_qs;
			addr_hit[139]: reg_rdata_next[1:0] = alert_class_shadowed_3_qs;
			addr_hit[140]: reg_rdata_next[1:0] = alert_class_shadowed_4_qs;
			addr_hit[141]: reg_rdata_next[1:0] = alert_class_shadowed_5_qs;
			addr_hit[142]: reg_rdata_next[1:0] = alert_class_shadowed_6_qs;
			addr_hit[143]: reg_rdata_next[1:0] = alert_class_shadowed_7_qs;
			addr_hit[144]: reg_rdata_next[1:0] = alert_class_shadowed_8_qs;
			addr_hit[145]: reg_rdata_next[1:0] = alert_class_shadowed_9_qs;
			addr_hit[146]: reg_rdata_next[1:0] = alert_class_shadowed_10_qs;
			addr_hit[147]: reg_rdata_next[1:0] = alert_class_shadowed_11_qs;
			addr_hit[148]: reg_rdata_next[1:0] = alert_class_shadowed_12_qs;
			addr_hit[149]: reg_rdata_next[1:0] = alert_class_shadowed_13_qs;
			addr_hit[150]: reg_rdata_next[1:0] = alert_class_shadowed_14_qs;
			addr_hit[151]: reg_rdata_next[1:0] = alert_class_shadowed_15_qs;
			addr_hit[152]: reg_rdata_next[1:0] = alert_class_shadowed_16_qs;
			addr_hit[153]: reg_rdata_next[1:0] = alert_class_shadowed_17_qs;
			addr_hit[154]: reg_rdata_next[1:0] = alert_class_shadowed_18_qs;
			addr_hit[155]: reg_rdata_next[1:0] = alert_class_shadowed_19_qs;
			addr_hit[156]: reg_rdata_next[1:0] = alert_class_shadowed_20_qs;
			addr_hit[157]: reg_rdata_next[1:0] = alert_class_shadowed_21_qs;
			addr_hit[158]: reg_rdata_next[1:0] = alert_class_shadowed_22_qs;
			addr_hit[159]: reg_rdata_next[1:0] = alert_class_shadowed_23_qs;
			addr_hit[160]: reg_rdata_next[1:0] = alert_class_shadowed_24_qs;
			addr_hit[161]: reg_rdata_next[1:0] = alert_class_shadowed_25_qs;
			addr_hit[162]: reg_rdata_next[1:0] = alert_class_shadowed_26_qs;
			addr_hit[163]: reg_rdata_next[1:0] = alert_class_shadowed_27_qs;
			addr_hit[164]: reg_rdata_next[1:0] = alert_class_shadowed_28_qs;
			addr_hit[165]: reg_rdata_next[1:0] = alert_class_shadowed_29_qs;
			addr_hit[166]: reg_rdata_next[1:0] = alert_class_shadowed_30_qs;
			addr_hit[167]: reg_rdata_next[1:0] = alert_class_shadowed_31_qs;
			addr_hit[168]: reg_rdata_next[1:0] = alert_class_shadowed_32_qs;
			addr_hit[169]: reg_rdata_next[1:0] = alert_class_shadowed_33_qs;
			addr_hit[170]: reg_rdata_next[1:0] = alert_class_shadowed_34_qs;
			addr_hit[171]: reg_rdata_next[1:0] = alert_class_shadowed_35_qs;
			addr_hit[172]: reg_rdata_next[1:0] = alert_class_shadowed_36_qs;
			addr_hit[173]: reg_rdata_next[1:0] = alert_class_shadowed_37_qs;
			addr_hit[174]: reg_rdata_next[1:0] = alert_class_shadowed_38_qs;
			addr_hit[175]: reg_rdata_next[1:0] = alert_class_shadowed_39_qs;
			addr_hit[176]: reg_rdata_next[1:0] = alert_class_shadowed_40_qs;
			addr_hit[177]: reg_rdata_next[1:0] = alert_class_shadowed_41_qs;
			addr_hit[178]: reg_rdata_next[1:0] = alert_class_shadowed_42_qs;
			addr_hit[179]: reg_rdata_next[1:0] = alert_class_shadowed_43_qs;
			addr_hit[180]: reg_rdata_next[1:0] = alert_class_shadowed_44_qs;
			addr_hit[181]: reg_rdata_next[1:0] = alert_class_shadowed_45_qs;
			addr_hit[182]: reg_rdata_next[1:0] = alert_class_shadowed_46_qs;
			addr_hit[183]: reg_rdata_next[1:0] = alert_class_shadowed_47_qs;
			addr_hit[184]: reg_rdata_next[1:0] = alert_class_shadowed_48_qs;
			addr_hit[185]: reg_rdata_next[1:0] = alert_class_shadowed_49_qs;
			addr_hit[186]: reg_rdata_next[1:0] = alert_class_shadowed_50_qs;
			addr_hit[187]: reg_rdata_next[1:0] = alert_class_shadowed_51_qs;
			addr_hit[188]: reg_rdata_next[1:0] = alert_class_shadowed_52_qs;
			addr_hit[189]: reg_rdata_next[1:0] = alert_class_shadowed_53_qs;
			addr_hit[190]: reg_rdata_next[1:0] = alert_class_shadowed_54_qs;
			addr_hit[191]: reg_rdata_next[1:0] = alert_class_shadowed_55_qs;
			addr_hit[192]: reg_rdata_next[1:0] = alert_class_shadowed_56_qs;
			addr_hit[193]: reg_rdata_next[1:0] = alert_class_shadowed_57_qs;
			addr_hit[194]: reg_rdata_next[1:0] = alert_class_shadowed_58_qs;
			addr_hit[195]: reg_rdata_next[1:0] = alert_class_shadowed_59_qs;
			addr_hit[196]: reg_rdata_next[1:0] = alert_class_shadowed_60_qs;
			addr_hit[197]: reg_rdata_next[1:0] = alert_class_shadowed_61_qs;
			addr_hit[198]: reg_rdata_next[1:0] = alert_class_shadowed_62_qs;
			addr_hit[199]: reg_rdata_next[1:0] = alert_class_shadowed_63_qs;
			addr_hit[200]: reg_rdata_next[1:0] = alert_class_shadowed_64_qs;
			addr_hit[201]: reg_rdata_next[0] = alert_cause_0_qs;
			addr_hit[202]: reg_rdata_next[0] = alert_cause_1_qs;
			addr_hit[203]: reg_rdata_next[0] = alert_cause_2_qs;
			addr_hit[204]: reg_rdata_next[0] = alert_cause_3_qs;
			addr_hit[205]: reg_rdata_next[0] = alert_cause_4_qs;
			addr_hit[206]: reg_rdata_next[0] = alert_cause_5_qs;
			addr_hit[207]: reg_rdata_next[0] = alert_cause_6_qs;
			addr_hit[208]: reg_rdata_next[0] = alert_cause_7_qs;
			addr_hit[209]: reg_rdata_next[0] = alert_cause_8_qs;
			addr_hit[210]: reg_rdata_next[0] = alert_cause_9_qs;
			addr_hit[211]: reg_rdata_next[0] = alert_cause_10_qs;
			addr_hit[212]: reg_rdata_next[0] = alert_cause_11_qs;
			addr_hit[213]: reg_rdata_next[0] = alert_cause_12_qs;
			addr_hit[214]: reg_rdata_next[0] = alert_cause_13_qs;
			addr_hit[215]: reg_rdata_next[0] = alert_cause_14_qs;
			addr_hit[216]: reg_rdata_next[0] = alert_cause_15_qs;
			addr_hit[217]: reg_rdata_next[0] = alert_cause_16_qs;
			addr_hit[218]: reg_rdata_next[0] = alert_cause_17_qs;
			addr_hit[219]: reg_rdata_next[0] = alert_cause_18_qs;
			addr_hit[220]: reg_rdata_next[0] = alert_cause_19_qs;
			addr_hit[221]: reg_rdata_next[0] = alert_cause_20_qs;
			addr_hit[222]: reg_rdata_next[0] = alert_cause_21_qs;
			addr_hit[223]: reg_rdata_next[0] = alert_cause_22_qs;
			addr_hit[224]: reg_rdata_next[0] = alert_cause_23_qs;
			addr_hit[225]: reg_rdata_next[0] = alert_cause_24_qs;
			addr_hit[226]: reg_rdata_next[0] = alert_cause_25_qs;
			addr_hit[227]: reg_rdata_next[0] = alert_cause_26_qs;
			addr_hit[228]: reg_rdata_next[0] = alert_cause_27_qs;
			addr_hit[229]: reg_rdata_next[0] = alert_cause_28_qs;
			addr_hit[230]: reg_rdata_next[0] = alert_cause_29_qs;
			addr_hit[231]: reg_rdata_next[0] = alert_cause_30_qs;
			addr_hit[232]: reg_rdata_next[0] = alert_cause_31_qs;
			addr_hit[233]: reg_rdata_next[0] = alert_cause_32_qs;
			addr_hit[234]: reg_rdata_next[0] = alert_cause_33_qs;
			addr_hit[235]: reg_rdata_next[0] = alert_cause_34_qs;
			addr_hit[236]: reg_rdata_next[0] = alert_cause_35_qs;
			addr_hit[237]: reg_rdata_next[0] = alert_cause_36_qs;
			addr_hit[238]: reg_rdata_next[0] = alert_cause_37_qs;
			addr_hit[239]: reg_rdata_next[0] = alert_cause_38_qs;
			addr_hit[240]: reg_rdata_next[0] = alert_cause_39_qs;
			addr_hit[241]: reg_rdata_next[0] = alert_cause_40_qs;
			addr_hit[242]: reg_rdata_next[0] = alert_cause_41_qs;
			addr_hit[243]: reg_rdata_next[0] = alert_cause_42_qs;
			addr_hit[244]: reg_rdata_next[0] = alert_cause_43_qs;
			addr_hit[245]: reg_rdata_next[0] = alert_cause_44_qs;
			addr_hit[246]: reg_rdata_next[0] = alert_cause_45_qs;
			addr_hit[247]: reg_rdata_next[0] = alert_cause_46_qs;
			addr_hit[248]: reg_rdata_next[0] = alert_cause_47_qs;
			addr_hit[249]: reg_rdata_next[0] = alert_cause_48_qs;
			addr_hit[250]: reg_rdata_next[0] = alert_cause_49_qs;
			addr_hit[251]: reg_rdata_next[0] = alert_cause_50_qs;
			addr_hit[252]: reg_rdata_next[0] = alert_cause_51_qs;
			addr_hit[253]: reg_rdata_next[0] = alert_cause_52_qs;
			addr_hit[254]: reg_rdata_next[0] = alert_cause_53_qs;
			addr_hit[255]: reg_rdata_next[0] = alert_cause_54_qs;
			addr_hit[256]: reg_rdata_next[0] = alert_cause_55_qs;
			addr_hit[257]: reg_rdata_next[0] = alert_cause_56_qs;
			addr_hit[258]: reg_rdata_next[0] = alert_cause_57_qs;
			addr_hit[259]: reg_rdata_next[0] = alert_cause_58_qs;
			addr_hit[260]: reg_rdata_next[0] = alert_cause_59_qs;
			addr_hit[261]: reg_rdata_next[0] = alert_cause_60_qs;
			addr_hit[262]: reg_rdata_next[0] = alert_cause_61_qs;
			addr_hit[263]: reg_rdata_next[0] = alert_cause_62_qs;
			addr_hit[264]: reg_rdata_next[0] = alert_cause_63_qs;
			addr_hit[265]: reg_rdata_next[0] = alert_cause_64_qs;
			addr_hit[266]: reg_rdata_next[0] = loc_alert_regwen_0_qs;
			addr_hit[267]: reg_rdata_next[0] = loc_alert_regwen_1_qs;
			addr_hit[268]: reg_rdata_next[0] = loc_alert_regwen_2_qs;
			addr_hit[269]: reg_rdata_next[0] = loc_alert_regwen_3_qs;
			addr_hit[270]: reg_rdata_next[0] = loc_alert_regwen_4_qs;
			addr_hit[271]: reg_rdata_next[0] = loc_alert_regwen_5_qs;
			addr_hit[272]: reg_rdata_next[0] = loc_alert_regwen_6_qs;
			addr_hit[273]: reg_rdata_next[0] = loc_alert_en_shadowed_0_qs;
			addr_hit[274]: reg_rdata_next[0] = loc_alert_en_shadowed_1_qs;
			addr_hit[275]: reg_rdata_next[0] = loc_alert_en_shadowed_2_qs;
			addr_hit[276]: reg_rdata_next[0] = loc_alert_en_shadowed_3_qs;
			addr_hit[277]: reg_rdata_next[0] = loc_alert_en_shadowed_4_qs;
			addr_hit[278]: reg_rdata_next[0] = loc_alert_en_shadowed_5_qs;
			addr_hit[279]: reg_rdata_next[0] = loc_alert_en_shadowed_6_qs;
			addr_hit[280]: reg_rdata_next[1:0] = loc_alert_class_shadowed_0_qs;
			addr_hit[281]: reg_rdata_next[1:0] = loc_alert_class_shadowed_1_qs;
			addr_hit[282]: reg_rdata_next[1:0] = loc_alert_class_shadowed_2_qs;
			addr_hit[283]: reg_rdata_next[1:0] = loc_alert_class_shadowed_3_qs;
			addr_hit[284]: reg_rdata_next[1:0] = loc_alert_class_shadowed_4_qs;
			addr_hit[285]: reg_rdata_next[1:0] = loc_alert_class_shadowed_5_qs;
			addr_hit[286]: reg_rdata_next[1:0] = loc_alert_class_shadowed_6_qs;
			addr_hit[287]: reg_rdata_next[0] = loc_alert_cause_0_qs;
			addr_hit[288]: reg_rdata_next[0] = loc_alert_cause_1_qs;
			addr_hit[289]: reg_rdata_next[0] = loc_alert_cause_2_qs;
			addr_hit[290]: reg_rdata_next[0] = loc_alert_cause_3_qs;
			addr_hit[291]: reg_rdata_next[0] = loc_alert_cause_4_qs;
			addr_hit[292]: reg_rdata_next[0] = loc_alert_cause_5_qs;
			addr_hit[293]: reg_rdata_next[0] = loc_alert_cause_6_qs;
			addr_hit[294]: reg_rdata_next[0] = classa_regwen_qs;
			addr_hit[295]: begin
				reg_rdata_next[0] = classa_ctrl_shadowed_en_qs;
				reg_rdata_next[1] = classa_ctrl_shadowed_lock_qs;
				reg_rdata_next[2] = classa_ctrl_shadowed_en_e0_qs;
				reg_rdata_next[3] = classa_ctrl_shadowed_en_e1_qs;
				reg_rdata_next[4] = classa_ctrl_shadowed_en_e2_qs;
				reg_rdata_next[5] = classa_ctrl_shadowed_en_e3_qs;
				reg_rdata_next[7:6] = classa_ctrl_shadowed_map_e0_qs;
				reg_rdata_next[9:8] = classa_ctrl_shadowed_map_e1_qs;
				reg_rdata_next[11:10] = classa_ctrl_shadowed_map_e2_qs;
				reg_rdata_next[13:12] = classa_ctrl_shadowed_map_e3_qs;
			end
			addr_hit[296]: reg_rdata_next[0] = classa_clr_regwen_qs;
			addr_hit[297]: reg_rdata_next[0] = classa_clr_shadowed_qs;
			addr_hit[298]: reg_rdata_next[15:0] = classa_accum_cnt_qs;
			addr_hit[299]: reg_rdata_next[15:0] = classa_accum_thresh_shadowed_qs;
			addr_hit[300]: reg_rdata_next[31:0] = classa_timeout_cyc_shadowed_qs;
			addr_hit[301]: reg_rdata_next[1:0] = classa_crashdump_trigger_shadowed_qs;
			addr_hit[302]: reg_rdata_next[31:0] = classa_phase0_cyc_shadowed_qs;
			addr_hit[303]: reg_rdata_next[31:0] = classa_phase1_cyc_shadowed_qs;
			addr_hit[304]: reg_rdata_next[31:0] = classa_phase2_cyc_shadowed_qs;
			addr_hit[305]: reg_rdata_next[31:0] = classa_phase3_cyc_shadowed_qs;
			addr_hit[306]: reg_rdata_next[31:0] = classa_esc_cnt_qs;
			addr_hit[307]: reg_rdata_next[2:0] = classa_state_qs;
			addr_hit[308]: reg_rdata_next[0] = classb_regwen_qs;
			addr_hit[309]: begin
				reg_rdata_next[0] = classb_ctrl_shadowed_en_qs;
				reg_rdata_next[1] = classb_ctrl_shadowed_lock_qs;
				reg_rdata_next[2] = classb_ctrl_shadowed_en_e0_qs;
				reg_rdata_next[3] = classb_ctrl_shadowed_en_e1_qs;
				reg_rdata_next[4] = classb_ctrl_shadowed_en_e2_qs;
				reg_rdata_next[5] = classb_ctrl_shadowed_en_e3_qs;
				reg_rdata_next[7:6] = classb_ctrl_shadowed_map_e0_qs;
				reg_rdata_next[9:8] = classb_ctrl_shadowed_map_e1_qs;
				reg_rdata_next[11:10] = classb_ctrl_shadowed_map_e2_qs;
				reg_rdata_next[13:12] = classb_ctrl_shadowed_map_e3_qs;
			end
			addr_hit[310]: reg_rdata_next[0] = classb_clr_regwen_qs;
			addr_hit[311]: reg_rdata_next[0] = classb_clr_shadowed_qs;
			addr_hit[312]: reg_rdata_next[15:0] = classb_accum_cnt_qs;
			addr_hit[313]: reg_rdata_next[15:0] = classb_accum_thresh_shadowed_qs;
			addr_hit[314]: reg_rdata_next[31:0] = classb_timeout_cyc_shadowed_qs;
			addr_hit[315]: reg_rdata_next[1:0] = classb_crashdump_trigger_shadowed_qs;
			addr_hit[316]: reg_rdata_next[31:0] = classb_phase0_cyc_shadowed_qs;
			addr_hit[317]: reg_rdata_next[31:0] = classb_phase1_cyc_shadowed_qs;
			addr_hit[318]: reg_rdata_next[31:0] = classb_phase2_cyc_shadowed_qs;
			addr_hit[319]: reg_rdata_next[31:0] = classb_phase3_cyc_shadowed_qs;
			addr_hit[320]: reg_rdata_next[31:0] = classb_esc_cnt_qs;
			addr_hit[321]: reg_rdata_next[2:0] = classb_state_qs;
			addr_hit[322]: reg_rdata_next[0] = classc_regwen_qs;
			addr_hit[323]: begin
				reg_rdata_next[0] = classc_ctrl_shadowed_en_qs;
				reg_rdata_next[1] = classc_ctrl_shadowed_lock_qs;
				reg_rdata_next[2] = classc_ctrl_shadowed_en_e0_qs;
				reg_rdata_next[3] = classc_ctrl_shadowed_en_e1_qs;
				reg_rdata_next[4] = classc_ctrl_shadowed_en_e2_qs;
				reg_rdata_next[5] = classc_ctrl_shadowed_en_e3_qs;
				reg_rdata_next[7:6] = classc_ctrl_shadowed_map_e0_qs;
				reg_rdata_next[9:8] = classc_ctrl_shadowed_map_e1_qs;
				reg_rdata_next[11:10] = classc_ctrl_shadowed_map_e2_qs;
				reg_rdata_next[13:12] = classc_ctrl_shadowed_map_e3_qs;
			end
			addr_hit[324]: reg_rdata_next[0] = classc_clr_regwen_qs;
			addr_hit[325]: reg_rdata_next[0] = classc_clr_shadowed_qs;
			addr_hit[326]: reg_rdata_next[15:0] = classc_accum_cnt_qs;
			addr_hit[327]: reg_rdata_next[15:0] = classc_accum_thresh_shadowed_qs;
			addr_hit[328]: reg_rdata_next[31:0] = classc_timeout_cyc_shadowed_qs;
			addr_hit[329]: reg_rdata_next[1:0] = classc_crashdump_trigger_shadowed_qs;
			addr_hit[330]: reg_rdata_next[31:0] = classc_phase0_cyc_shadowed_qs;
			addr_hit[331]: reg_rdata_next[31:0] = classc_phase1_cyc_shadowed_qs;
			addr_hit[332]: reg_rdata_next[31:0] = classc_phase2_cyc_shadowed_qs;
			addr_hit[333]: reg_rdata_next[31:0] = classc_phase3_cyc_shadowed_qs;
			addr_hit[334]: reg_rdata_next[31:0] = classc_esc_cnt_qs;
			addr_hit[335]: reg_rdata_next[2:0] = classc_state_qs;
			addr_hit[336]: reg_rdata_next[0] = classd_regwen_qs;
			addr_hit[337]: begin
				reg_rdata_next[0] = classd_ctrl_shadowed_en_qs;
				reg_rdata_next[1] = classd_ctrl_shadowed_lock_qs;
				reg_rdata_next[2] = classd_ctrl_shadowed_en_e0_qs;
				reg_rdata_next[3] = classd_ctrl_shadowed_en_e1_qs;
				reg_rdata_next[4] = classd_ctrl_shadowed_en_e2_qs;
				reg_rdata_next[5] = classd_ctrl_shadowed_en_e3_qs;
				reg_rdata_next[7:6] = classd_ctrl_shadowed_map_e0_qs;
				reg_rdata_next[9:8] = classd_ctrl_shadowed_map_e1_qs;
				reg_rdata_next[11:10] = classd_ctrl_shadowed_map_e2_qs;
				reg_rdata_next[13:12] = classd_ctrl_shadowed_map_e3_qs;
			end
			addr_hit[338]: reg_rdata_next[0] = classd_clr_regwen_qs;
			addr_hit[339]: reg_rdata_next[0] = classd_clr_shadowed_qs;
			addr_hit[340]: reg_rdata_next[15:0] = classd_accum_cnt_qs;
			addr_hit[341]: reg_rdata_next[15:0] = classd_accum_thresh_shadowed_qs;
			addr_hit[342]: reg_rdata_next[31:0] = classd_timeout_cyc_shadowed_qs;
			addr_hit[343]: reg_rdata_next[1:0] = classd_crashdump_trigger_shadowed_qs;
			addr_hit[344]: reg_rdata_next[31:0] = classd_phase0_cyc_shadowed_qs;
			addr_hit[345]: reg_rdata_next[31:0] = classd_phase1_cyc_shadowed_qs;
			addr_hit[346]: reg_rdata_next[31:0] = classd_phase2_cyc_shadowed_qs;
			addr_hit[347]: reg_rdata_next[31:0] = classd_phase3_cyc_shadowed_qs;
			addr_hit[348]: reg_rdata_next[31:0] = classd_esc_cnt_qs;
			addr_hit[349]: reg_rdata_next[2:0] = classd_state_qs;
			default: reg_rdata_next = 1'sb1;
		endcase
	end
	wire shadow_busy;
	reg rst_done;
	reg shadow_rst_done;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			rst_done <= 1'sb0;
		else
			rst_done <= 1'b1;
	always @(posedge clk_i or negedge rst_shadowed_ni)
		if (!rst_shadowed_ni)
			shadow_rst_done <= 1'sb0;
		else
			shadow_rst_done <= 1'b1;
	assign shadow_busy = ~(rst_done & shadow_rst_done);
	assign shadowed_storage_err_o = |{ping_timeout_cyc_shadowed_storage_err, ping_timer_en_shadowed_storage_err, alert_en_shadowed_0_storage_err, alert_en_shadowed_1_storage_err, alert_en_shadowed_2_storage_err, alert_en_shadowed_3_storage_err, alert_en_shadowed_4_storage_err, alert_en_shadowed_5_storage_err, alert_en_shadowed_6_storage_err, alert_en_shadowed_7_storage_err, alert_en_shadowed_8_storage_err, alert_en_shadowed_9_storage_err, alert_en_shadowed_10_storage_err, alert_en_shadowed_11_storage_err, alert_en_shadowed_12_storage_err, alert_en_shadowed_13_storage_err, alert_en_shadowed_14_storage_err, alert_en_shadowed_15_storage_err, alert_en_shadowed_16_storage_err, alert_en_shadowed_17_storage_err, alert_en_shadowed_18_storage_err, alert_en_shadowed_19_storage_err, alert_en_shadowed_20_storage_err, alert_en_shadowed_21_storage_err, alert_en_shadowed_22_storage_err, alert_en_shadowed_23_storage_err, alert_en_shadowed_24_storage_err, alert_en_shadowed_25_storage_err, alert_en_shadowed_26_storage_err, alert_en_shadowed_27_storage_err, alert_en_shadowed_28_storage_err, alert_en_shadowed_29_storage_err, alert_en_shadowed_30_storage_err, alert_en_shadowed_31_storage_err, alert_en_shadowed_32_storage_err, alert_en_shadowed_33_storage_err, alert_en_shadowed_34_storage_err, alert_en_shadowed_35_storage_err, alert_en_shadowed_36_storage_err, alert_en_shadowed_37_storage_err, alert_en_shadowed_38_storage_err, alert_en_shadowed_39_storage_err, alert_en_shadowed_40_storage_err, alert_en_shadowed_41_storage_err, alert_en_shadowed_42_storage_err, alert_en_shadowed_43_storage_err, alert_en_shadowed_44_storage_err, alert_en_shadowed_45_storage_err, alert_en_shadowed_46_storage_err, alert_en_shadowed_47_storage_err, alert_en_shadowed_48_storage_err, alert_en_shadowed_49_storage_err, alert_en_shadowed_50_storage_err, alert_en_shadowed_51_storage_err, alert_en_shadowed_52_storage_err, alert_en_shadowed_53_storage_err, alert_en_shadowed_54_storage_err, alert_en_shadowed_55_storage_err, alert_en_shadowed_56_storage_err, alert_en_shadowed_57_storage_err, alert_en_shadowed_58_storage_err, alert_en_shadowed_59_storage_err, alert_en_shadowed_60_storage_err, alert_en_shadowed_61_storage_err, alert_en_shadowed_62_storage_err, alert_en_shadowed_63_storage_err, alert_en_shadowed_64_storage_err, alert_class_shadowed_0_storage_err, alert_class_shadowed_1_storage_err, alert_class_shadowed_2_storage_err, alert_class_shadowed_3_storage_err, alert_class_shadowed_4_storage_err, alert_class_shadowed_5_storage_err, alert_class_shadowed_6_storage_err, alert_class_shadowed_7_storage_err, alert_class_shadowed_8_storage_err, alert_class_shadowed_9_storage_err, alert_class_shadowed_10_storage_err, alert_class_shadowed_11_storage_err, alert_class_shadowed_12_storage_err, alert_class_shadowed_13_storage_err, alert_class_shadowed_14_storage_err, alert_class_shadowed_15_storage_err, alert_class_shadowed_16_storage_err, alert_class_shadowed_17_storage_err, alert_class_shadowed_18_storage_err, alert_class_shadowed_19_storage_err, alert_class_shadowed_20_storage_err, alert_class_shadowed_21_storage_err, alert_class_shadowed_22_storage_err, alert_class_shadowed_23_storage_err, alert_class_shadowed_24_storage_err, alert_class_shadowed_25_storage_err, alert_class_shadowed_26_storage_err, alert_class_shadowed_27_storage_err, alert_class_shadowed_28_storage_err, alert_class_shadowed_29_storage_err, alert_class_shadowed_30_storage_err, alert_class_shadowed_31_storage_err, alert_class_shadowed_32_storage_err, alert_class_shadowed_33_storage_err, alert_class_shadowed_34_storage_err, alert_class_shadowed_35_storage_err, alert_class_shadowed_36_storage_err, alert_class_shadowed_37_storage_err, alert_class_shadowed_38_storage_err, alert_class_shadowed_39_storage_err, alert_class_shadowed_40_storage_err, alert_class_shadowed_41_storage_err, alert_class_shadowed_42_storage_err, alert_class_shadowed_43_storage_err, alert_class_shadowed_44_storage_err, alert_class_shadowed_45_storage_err, alert_class_shadowed_46_storage_err, alert_class_shadowed_47_storage_err, alert_class_shadowed_48_storage_err, alert_class_shadowed_49_storage_err, alert_class_shadowed_50_storage_err, alert_class_shadowed_51_storage_err, alert_class_shadowed_52_storage_err, alert_class_shadowed_53_storage_err, alert_class_shadowed_54_storage_err, alert_class_shadowed_55_storage_err, alert_class_shadowed_56_storage_err, alert_class_shadowed_57_storage_err, alert_class_shadowed_58_storage_err, alert_class_shadowed_59_storage_err, alert_class_shadowed_60_storage_err, alert_class_shadowed_61_storage_err, alert_class_shadowed_62_storage_err, alert_class_shadowed_63_storage_err, alert_class_shadowed_64_storage_err, loc_alert_en_shadowed_0_storage_err, loc_alert_en_shadowed_1_storage_err, loc_alert_en_shadowed_2_storage_err, loc_alert_en_shadowed_3_storage_err, loc_alert_en_shadowed_4_storage_err, loc_alert_en_shadowed_5_storage_err, loc_alert_en_shadowed_6_storage_err, loc_alert_class_shadowed_0_storage_err, loc_alert_class_shadowed_1_storage_err, loc_alert_class_shadowed_2_storage_err, loc_alert_class_shadowed_3_storage_err, loc_alert_class_shadowed_4_storage_err, loc_alert_class_shadowed_5_storage_err, loc_alert_class_shadowed_6_storage_err, classa_ctrl_shadowed_en_storage_err, classa_ctrl_shadowed_lock_storage_err, classa_ctrl_shadowed_en_e0_storage_err, classa_ctrl_shadowed_en_e1_storage_err, classa_ctrl_shadowed_en_e2_storage_err, classa_ctrl_shadowed_en_e3_storage_err, classa_ctrl_shadowed_map_e0_storage_err, classa_ctrl_shadowed_map_e1_storage_err, classa_ctrl_shadowed_map_e2_storage_err, classa_ctrl_shadowed_map_e3_storage_err, classa_clr_shadowed_storage_err, classa_accum_thresh_shadowed_storage_err, classa_timeout_cyc_shadowed_storage_err, classa_crashdump_trigger_shadowed_storage_err, classa_phase0_cyc_shadowed_storage_err, classa_phase1_cyc_shadowed_storage_err, classa_phase2_cyc_shadowed_storage_err, classa_phase3_cyc_shadowed_storage_err, classb_ctrl_shadowed_en_storage_err, classb_ctrl_shadowed_lock_storage_err, classb_ctrl_shadowed_en_e0_storage_err, classb_ctrl_shadowed_en_e1_storage_err, classb_ctrl_shadowed_en_e2_storage_err, classb_ctrl_shadowed_en_e3_storage_err, classb_ctrl_shadowed_map_e0_storage_err, classb_ctrl_shadowed_map_e1_storage_err, classb_ctrl_shadowed_map_e2_storage_err, classb_ctrl_shadowed_map_e3_storage_err, classb_clr_shadowed_storage_err, classb_accum_thresh_shadowed_storage_err, classb_timeout_cyc_shadowed_storage_err, classb_crashdump_trigger_shadowed_storage_err, classb_phase0_cyc_shadowed_storage_err, classb_phase1_cyc_shadowed_storage_err, classb_phase2_cyc_shadowed_storage_err, classb_phase3_cyc_shadowed_storage_err, classc_ctrl_shadowed_en_storage_err, classc_ctrl_shadowed_lock_storage_err, classc_ctrl_shadowed_en_e0_storage_err, classc_ctrl_shadowed_en_e1_storage_err, classc_ctrl_shadowed_en_e2_storage_err, classc_ctrl_shadowed_en_e3_storage_err, classc_ctrl_shadowed_map_e0_storage_err, classc_ctrl_shadowed_map_e1_storage_err, classc_ctrl_shadowed_map_e2_storage_err, classc_ctrl_shadowed_map_e3_storage_err, classc_clr_shadowed_storage_err, classc_accum_thresh_shadowed_storage_err, classc_timeout_cyc_shadowed_storage_err, classc_crashdump_trigger_shadowed_storage_err, classc_phase0_cyc_shadowed_storage_err, classc_phase1_cyc_shadowed_storage_err, classc_phase2_cyc_shadowed_storage_err, classc_phase3_cyc_shadowed_storage_err, classd_ctrl_shadowed_en_storage_err, classd_ctrl_shadowed_lock_storage_err, classd_ctrl_shadowed_en_e0_storage_err, classd_ctrl_shadowed_en_e1_storage_err, classd_ctrl_shadowed_en_e2_storage_err, classd_ctrl_shadowed_en_e3_storage_err, classd_ctrl_shadowed_map_e0_storage_err, classd_ctrl_shadowed_map_e1_storage_err, classd_ctrl_shadowed_map_e2_storage_err, classd_ctrl_shadowed_map_e3_storage_err, classd_clr_shadowed_storage_err, classd_accum_thresh_shadowed_storage_err, classd_timeout_cyc_shadowed_storage_err, classd_crashdump_trigger_shadowed_storage_err, classd_phase0_cyc_shadowed_storage_err, classd_phase1_cyc_shadowed_storage_err, classd_phase2_cyc_shadowed_storage_err, classd_phase3_cyc_shadowed_storage_err};
	assign shadowed_update_err_o = |{ping_timeout_cyc_shadowed_update_err, ping_timer_en_shadowed_update_err, alert_en_shadowed_0_update_err, alert_en_shadowed_1_update_err, alert_en_shadowed_2_update_err, alert_en_shadowed_3_update_err, alert_en_shadowed_4_update_err, alert_en_shadowed_5_update_err, alert_en_shadowed_6_update_err, alert_en_shadowed_7_update_err, alert_en_shadowed_8_update_err, alert_en_shadowed_9_update_err, alert_en_shadowed_10_update_err, alert_en_shadowed_11_update_err, alert_en_shadowed_12_update_err, alert_en_shadowed_13_update_err, alert_en_shadowed_14_update_err, alert_en_shadowed_15_update_err, alert_en_shadowed_16_update_err, alert_en_shadowed_17_update_err, alert_en_shadowed_18_update_err, alert_en_shadowed_19_update_err, alert_en_shadowed_20_update_err, alert_en_shadowed_21_update_err, alert_en_shadowed_22_update_err, alert_en_shadowed_23_update_err, alert_en_shadowed_24_update_err, alert_en_shadowed_25_update_err, alert_en_shadowed_26_update_err, alert_en_shadowed_27_update_err, alert_en_shadowed_28_update_err, alert_en_shadowed_29_update_err, alert_en_shadowed_30_update_err, alert_en_shadowed_31_update_err, alert_en_shadowed_32_update_err, alert_en_shadowed_33_update_err, alert_en_shadowed_34_update_err, alert_en_shadowed_35_update_err, alert_en_shadowed_36_update_err, alert_en_shadowed_37_update_err, alert_en_shadowed_38_update_err, alert_en_shadowed_39_update_err, alert_en_shadowed_40_update_err, alert_en_shadowed_41_update_err, alert_en_shadowed_42_update_err, alert_en_shadowed_43_update_err, alert_en_shadowed_44_update_err, alert_en_shadowed_45_update_err, alert_en_shadowed_46_update_err, alert_en_shadowed_47_update_err, alert_en_shadowed_48_update_err, alert_en_shadowed_49_update_err, alert_en_shadowed_50_update_err, alert_en_shadowed_51_update_err, alert_en_shadowed_52_update_err, alert_en_shadowed_53_update_err, alert_en_shadowed_54_update_err, alert_en_shadowed_55_update_err, alert_en_shadowed_56_update_err, alert_en_shadowed_57_update_err, alert_en_shadowed_58_update_err, alert_en_shadowed_59_update_err, alert_en_shadowed_60_update_err, alert_en_shadowed_61_update_err, alert_en_shadowed_62_update_err, alert_en_shadowed_63_update_err, alert_en_shadowed_64_update_err, alert_class_shadowed_0_update_err, alert_class_shadowed_1_update_err, alert_class_shadowed_2_update_err, alert_class_shadowed_3_update_err, alert_class_shadowed_4_update_err, alert_class_shadowed_5_update_err, alert_class_shadowed_6_update_err, alert_class_shadowed_7_update_err, alert_class_shadowed_8_update_err, alert_class_shadowed_9_update_err, alert_class_shadowed_10_update_err, alert_class_shadowed_11_update_err, alert_class_shadowed_12_update_err, alert_class_shadowed_13_update_err, alert_class_shadowed_14_update_err, alert_class_shadowed_15_update_err, alert_class_shadowed_16_update_err, alert_class_shadowed_17_update_err, alert_class_shadowed_18_update_err, alert_class_shadowed_19_update_err, alert_class_shadowed_20_update_err, alert_class_shadowed_21_update_err, alert_class_shadowed_22_update_err, alert_class_shadowed_23_update_err, alert_class_shadowed_24_update_err, alert_class_shadowed_25_update_err, alert_class_shadowed_26_update_err, alert_class_shadowed_27_update_err, alert_class_shadowed_28_update_err, alert_class_shadowed_29_update_err, alert_class_shadowed_30_update_err, alert_class_shadowed_31_update_err, alert_class_shadowed_32_update_err, alert_class_shadowed_33_update_err, alert_class_shadowed_34_update_err, alert_class_shadowed_35_update_err, alert_class_shadowed_36_update_err, alert_class_shadowed_37_update_err, alert_class_shadowed_38_update_err, alert_class_shadowed_39_update_err, alert_class_shadowed_40_update_err, alert_class_shadowed_41_update_err, alert_class_shadowed_42_update_err, alert_class_shadowed_43_update_err, alert_class_shadowed_44_update_err, alert_class_shadowed_45_update_err, alert_class_shadowed_46_update_err, alert_class_shadowed_47_update_err, alert_class_shadowed_48_update_err, alert_class_shadowed_49_update_err, alert_class_shadowed_50_update_err, alert_class_shadowed_51_update_err, alert_class_shadowed_52_update_err, alert_class_shadowed_53_update_err, alert_class_shadowed_54_update_err, alert_class_shadowed_55_update_err, alert_class_shadowed_56_update_err, alert_class_shadowed_57_update_err, alert_class_shadowed_58_update_err, alert_class_shadowed_59_update_err, alert_class_shadowed_60_update_err, alert_class_shadowed_61_update_err, alert_class_shadowed_62_update_err, alert_class_shadowed_63_update_err, alert_class_shadowed_64_update_err, loc_alert_en_shadowed_0_update_err, loc_alert_en_shadowed_1_update_err, loc_alert_en_shadowed_2_update_err, loc_alert_en_shadowed_3_update_err, loc_alert_en_shadowed_4_update_err, loc_alert_en_shadowed_5_update_err, loc_alert_en_shadowed_6_update_err, loc_alert_class_shadowed_0_update_err, loc_alert_class_shadowed_1_update_err, loc_alert_class_shadowed_2_update_err, loc_alert_class_shadowed_3_update_err, loc_alert_class_shadowed_4_update_err, loc_alert_class_shadowed_5_update_err, loc_alert_class_shadowed_6_update_err, classa_ctrl_shadowed_en_update_err, classa_ctrl_shadowed_lock_update_err, classa_ctrl_shadowed_en_e0_update_err, classa_ctrl_shadowed_en_e1_update_err, classa_ctrl_shadowed_en_e2_update_err, classa_ctrl_shadowed_en_e3_update_err, classa_ctrl_shadowed_map_e0_update_err, classa_ctrl_shadowed_map_e1_update_err, classa_ctrl_shadowed_map_e2_update_err, classa_ctrl_shadowed_map_e3_update_err, classa_clr_shadowed_update_err, classa_accum_thresh_shadowed_update_err, classa_timeout_cyc_shadowed_update_err, classa_crashdump_trigger_shadowed_update_err, classa_phase0_cyc_shadowed_update_err, classa_phase1_cyc_shadowed_update_err, classa_phase2_cyc_shadowed_update_err, classa_phase3_cyc_shadowed_update_err, classb_ctrl_shadowed_en_update_err, classb_ctrl_shadowed_lock_update_err, classb_ctrl_shadowed_en_e0_update_err, classb_ctrl_shadowed_en_e1_update_err, classb_ctrl_shadowed_en_e2_update_err, classb_ctrl_shadowed_en_e3_update_err, classb_ctrl_shadowed_map_e0_update_err, classb_ctrl_shadowed_map_e1_update_err, classb_ctrl_shadowed_map_e2_update_err, classb_ctrl_shadowed_map_e3_update_err, classb_clr_shadowed_update_err, classb_accum_thresh_shadowed_update_err, classb_timeout_cyc_shadowed_update_err, classb_crashdump_trigger_shadowed_update_err, classb_phase0_cyc_shadowed_update_err, classb_phase1_cyc_shadowed_update_err, classb_phase2_cyc_shadowed_update_err, classb_phase3_cyc_shadowed_update_err, classc_ctrl_shadowed_en_update_err, classc_ctrl_shadowed_lock_update_err, classc_ctrl_shadowed_en_e0_update_err, classc_ctrl_shadowed_en_e1_update_err, classc_ctrl_shadowed_en_e2_update_err, classc_ctrl_shadowed_en_e3_update_err, classc_ctrl_shadowed_map_e0_update_err, classc_ctrl_shadowed_map_e1_update_err, classc_ctrl_shadowed_map_e2_update_err, classc_ctrl_shadowed_map_e3_update_err, classc_clr_shadowed_update_err, classc_accum_thresh_shadowed_update_err, classc_timeout_cyc_shadowed_update_err, classc_crashdump_trigger_shadowed_update_err, classc_phase0_cyc_shadowed_update_err, classc_phase1_cyc_shadowed_update_err, classc_phase2_cyc_shadowed_update_err, classc_phase3_cyc_shadowed_update_err, classd_ctrl_shadowed_en_update_err, classd_ctrl_shadowed_lock_update_err, classd_ctrl_shadowed_en_e0_update_err, classd_ctrl_shadowed_en_e1_update_err, classd_ctrl_shadowed_en_e2_update_err, classd_ctrl_shadowed_en_e3_update_err, classd_ctrl_shadowed_map_e0_update_err, classd_ctrl_shadowed_map_e1_update_err, classd_ctrl_shadowed_map_e2_update_err, classd_ctrl_shadowed_map_e3_update_err, classd_clr_shadowed_update_err, classd_accum_thresh_shadowed_update_err, classd_timeout_cyc_shadowed_update_err, classd_crashdump_trigger_shadowed_update_err, classd_phase0_cyc_shadowed_update_err, classd_phase1_cyc_shadowed_update_err, classd_phase2_cyc_shadowed_update_err, classd_phase3_cyc_shadowed_update_err};
	assign reg_busy = shadow_busy;
	wire unused_wdata;
	wire unused_be;
	assign unused_wdata = ^reg_wdata;
	assign unused_be = ^reg_be;
endmodule
module cellift_rv_core_ibex_mem_top (
	clk_i,
	rst_ni,
	clk_edn_i,
	rst_edn_ni,
	clk_esc_i,
	rst_esc_ni,
	rst_cpu_n_o,
	ram_cfg_i,
	hart_id_i,
	boot_addr_i,
	instr_mem_req_o,
	instr_mem_gnt_i,
	instr_mem_addr_o,
	instr_mem_wdata_o,
	instr_mem_strb_o,
	instr_mem_we_o,
	instr_mem_rdata_i,
	data_mem_req_o,
	data_mem_gnt_i,
	data_mem_addr_o,
	data_mem_wdata_o,
	data_mem_strb_o,
	data_mem_we_o,
	data_mem_rdata_i,
	irq_software_i,
	irq_timer_i,
	irq_external_i,
	esc_tx_i,
	esc_rx_o,
	nmi_wdog_i,
	debug_req_i,
	crash_dump_o,
	pwrmgr_cpu_en_i,
	lc_cpu_en_i,
	pwrmgr_o,
	scan_rst_ni,
	scanmode_i,
	cfg_tl_d_i,
	cfg_tl_d_o,
	edn_o,
	edn_i,
	clk_otp_i,
	rst_otp_ni,
	icache_otp_key_o,
	icache_otp_key_i,
	fpga_info_i,
	alert_rx_i,
	alert_tx_o
);
	parameter [31:0] InstrMemAw = 20;
	parameter [31:0] DataMemAw = 20;
	input wire clk_i;
	input wire rst_ni;
	input wire clk_edn_i;
	input wire rst_edn_ni;
	input wire clk_esc_i;
	input wire rst_esc_ni;
	output wire rst_cpu_n_o;
	input wire [9:0] ram_cfg_i;
	input wire [31:0] hart_id_i;
	input wire [31:0] boot_addr_i;
	output wire instr_mem_req_o;
	input wire instr_mem_gnt_i;
	output wire [InstrMemAw:0] instr_mem_addr_o;
	output wire [31:0] instr_mem_wdata_o;
	output wire [31:0] instr_mem_strb_o;
	output wire instr_mem_we_o;
	input wire [31:0] instr_mem_rdata_i;
	output wire data_mem_req_o;
	input wire data_mem_gnt_i;
	output wire [InstrMemAw:0] data_mem_addr_o;
	output wire [31:0] data_mem_wdata_o;
	output wire [31:0] data_mem_strb_o;
	output wire data_mem_we_o;
	input wire [31:0] data_mem_rdata_i;
	input wire irq_software_i;
	input wire irq_timer_i;
	input wire irq_external_i;
	input wire [1:0] esc_tx_i;
	output wire [1:0] esc_rx_o;
	input wire nmi_wdog_i;
	input wire debug_req_i;
	output wire [159:0] crash_dump_o;
	localparam signed [31:0] lc_ctrl_pkg_TxWidth = 4;
	input wire [3:0] pwrmgr_cpu_en_i;
	input wire [3:0] lc_cpu_en_i;
	output wire [0:0] pwrmgr_o;
	input scan_rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	input wire [3:0] scanmode_i;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] cfg_tl_d_i;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] cfg_tl_d_o;
	output wire [0:0] edn_o;
	localparam [31:0] edn_pkg_ENDPOINT_BUS_WIDTH = 32;
	input wire [33:0] edn_i;
	input clk_otp_i;
	input rst_otp_ni;
	output wire [0:0] icache_otp_key_o;
	localparam signed [31:0] otp_ctrl_pkg_SramKeyWidth = 128;
	localparam signed [31:0] otp_ctrl_pkg_SramNonceWidth = 128;
	input wire [257:0] icache_otp_key_i;
	input [31:0] fpga_info_i;
	localparam signed [31:0] rv_core_ibex_reg_pkg_NumAlerts = 4;
	input wire [15:0] alert_rx_i;
	output wire [7:0] alert_tx_o;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_i_toibex;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_i_fromibex;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_d_toibex;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_d_fromibex;
	wire instr_rvalid_d;
	reg instr_rvalid_q;
	wire data_rvalid_d;
	reg data_rvalid_q;
	assign instr_rvalid_d = instr_mem_req_o & ~instr_mem_we_o;
	assign data_rvalid_d = data_mem_req_o & ~data_mem_we_o;
	always @(posedge clk_i)
		if (~rst_ni) begin
			instr_rvalid_q <= 1'sb0;
			data_rvalid_q <= 1'sb0;
		end
		else begin
			instr_rvalid_q <= instr_rvalid_d;
			data_rvalid_q <= data_rvalid_d;
		end
	function automatic [3:0] sv2v_cast_AC3DB;
		input reg [3:0] inp;
		sv2v_cast_AC3DB = inp;
	endfunction
	noerr_tlul_adapter_sram #(
		.SramAw(InstrMemAw),
		.SramDw(32),
		.Outstanding(1),
		.ByteAccess(1),
		.ErrOnWrite(0),
		.ErrOnRead(0),
		.CmdIntgCheck(0),
		.EnableRspIntgGen(0),
		.EnableDataIntgGen(0),
		.EnableDataIntgPt(0)
	) i_instr_tlul_adapter_sram(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_i_fromibex),
		.tl_o(tl_i_toibex),
		.en_ifetch_i(sv2v_cast_AC3DB(4'h6)),
		.req_o(instr_mem_req_o),
		.gnt_i(instr_mem_gnt_i),
		.we_o(instr_mem_we_o),
		.addr_o(instr_mem_addr_o),
		.wdata_o(instr_mem_wdata_o),
		.wmask_o(instr_mem_strb_o),
		.rdata_i(instr_mem_rdata_i),
		.rvalid_i(instr_rvalid_q),
		.rerror_i(2'b00)
	);
	noerr_tlul_adapter_sram #(
		.SramAw(DataMemAw),
		.SramDw(32),
		.Outstanding(1),
		.ByteAccess(1),
		.ErrOnWrite(0),
		.ErrOnRead(0),
		.CmdIntgCheck(0),
		.EnableRspIntgGen(0),
		.EnableDataIntgGen(0),
		.EnableDataIntgPt(0)
	) i_data_tlul_adapter_sram(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_d_fromibex),
		.tl_o(tl_d_toibex),
		.en_ifetch_i(sv2v_cast_AC3DB(4'h6)),
		.req_o(data_mem_req_o),
		.gnt_i(data_mem_gnt_i),
		.we_o(data_mem_we_o),
		.addr_o(data_mem_addr_o),
		.wdata_o(data_mem_wdata_o),
		.wmask_o(data_mem_strb_o),
		.rdata_i(data_mem_rdata_i),
		.rvalid_i(data_rvalid_q),
		.rerror_i(2'b00)
	);
	localparam signed [31:0] ibex_pkg_LfsrWidth = 32;
	localparam [159:0] ibex_pkg_RndCnstLfsrPermDefault = 160'h1e35ecba467fd1b12e958152c04fa43878a8daed;
	localparam [31:0] ibex_pkg_RndCnstLfsrSeedDefault = 32'hac533bf4;
	noerr_rv_core_ibex #(
		.PMPEnable(1'b0),
		.PMPGranularity(0),
		.PMPNumRegions(4),
		.MHPMCounterNum(0),
		.MHPMCounterWidth(40),
		.RV32E(1'b0),
		.RV32M(32'sd1),
		.RV32B(32'sd0),
		.BranchTargetALU(1'b0),
		.WritebackStage(1'b1),
		.ICache(1'b0),
		.ICacheECC(1'b0),
		.BranchPredictor(1'b0),
		.DbgTriggerEn(1'b0),
		.DbgHwBreakNum(1),
		.RndCnstLfsrSeed(ibex_pkg_RndCnstLfsrSeedDefault),
		.RndCnstLfsrPerm(ibex_pkg_RndCnstLfsrPermDefault),
		.SecureIbex(1'b0),
		.DmHaltAddr(32'h1a110800),
		.DmExceptionAddr(32'h01a11080)
	) i_rv_core_ibex(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clk_edn_i(clk_edn_i),
		.rst_edn_ni(rst_edn_ni),
		.clk_esc_i(clk_esc_i),
		.rst_esc_ni(rst_esc_ni),
		.rst_cpu_n_o(rst_cpu_n_o),
		.ram_cfg_i(ram_cfg_i),
		.hart_id_i(hart_id_i),
		.boot_addr_i(boot_addr_i),
		.corei_tl_h_o(tl_i_fromibex),
		.corei_tl_h_i(tl_i_toibex),
		.cored_tl_h_o(tl_d_fromibex),
		.cored_tl_h_i(tl_d_toibex),
		.irq_software_i(irq_software_i),
		.irq_timer_i(irq_timer_i),
		.irq_external_i(irq_external_i),
		.esc_tx_i(esc_tx_i),
		.esc_rx_o(esc_rx_o),
		.nmi_wdog_i(nmi_wdog_i),
		.debug_req_i(debug_req_i),
		.crash_dump_o(crash_dump_o),
		.lc_cpu_en_i(lc_cpu_en_i),
		.pwrmgr_cpu_en_i(pwrmgr_cpu_en_i),
		.pwrmgr_o(pwrmgr_o),
		.scan_rst_ni(scan_rst_ni),
		.scanmode_i(scanmode_i),
		.cfg_tl_d_i(cfg_tl_d_i),
		.cfg_tl_d_o(cfg_tl_d_o),
		.edn_o(edn_o),
		.edn_i(edn_i),
		.clk_otp_i(clk_otp_i),
		.rst_otp_ni(rst_otp_ni),
		.icache_otp_key_o(icache_otp_key_o),
		.icache_otp_key_i(icache_otp_key_i),
		.fpga_info_i(fpga_info_i),
		.alert_rx_i(alert_rx_i),
		.alert_tx_o(alert_tx_o)
	);
endmodule
module ibex_alu (
	operator_i,
	operand_a_i,
	operand_b_i,
	instr_first_cycle_i,
	multdiv_operand_a_i,
	multdiv_operand_b_i,
	multdiv_sel_i,
	imd_val_q_i,
	imd_val_d_o,
	imd_val_we_o,
	adder_result_o,
	adder_result_ext_o,
	result_o,
	comparison_result_o,
	is_equal_result_o
);
	parameter integer RV32B = 32'sd0;
	input wire [6:0] operator_i;
	input wire [31:0] operand_a_i;
	input wire [31:0] operand_b_i;
	input wire instr_first_cycle_i;
	input wire [32:0] multdiv_operand_a_i;
	input wire [32:0] multdiv_operand_b_i;
	input wire multdiv_sel_i;
	input wire [63:0] imd_val_q_i;
	output reg [63:0] imd_val_d_o;
	output reg [1:0] imd_val_we_o;
	output wire [31:0] adder_result_o;
	output wire [33:0] adder_result_ext_o;
	output reg [31:0] result_o;
	output wire comparison_result_o;
	output wire is_equal_result_o;
	wire [31:0] operand_a_rev;
	wire [32:0] operand_b_neg;
	genvar k;
	generate
		for (k = 0; k < 32; k = k + 1) begin : gen_rev_operand_a
			assign operand_a_rev[k] = operand_a_i[31 - k];
		end
	endgenerate
	reg adder_op_a_shift1;
	reg adder_op_a_shift2;
	reg adder_op_a_shift3;
	reg adder_op_b_negate;
	reg [32:0] adder_in_a;
	reg [32:0] adder_in_b;
	wire [31:0] adder_result;
	always @(*) begin
		adder_op_a_shift1 = 1'b0;
		adder_op_a_shift2 = 1'b0;
		adder_op_a_shift3 = 1'b0;
		adder_op_b_negate = 1'b0;
		case (operator_i)
			7'd1, 7'd29, 7'd30, 7'd27, 7'd28, 7'd25, 7'd26, 7'd43, 7'd44, 7'd31, 7'd32, 7'd33, 7'd34: adder_op_b_negate = 1'b1;
			7'd22:
				if (RV32B != 32'sd0)
					adder_op_a_shift1 = 1'b1;
			7'd23:
				if (RV32B != 32'sd0)
					adder_op_a_shift2 = 1'b1;
			7'd24:
				if (RV32B != 32'sd0)
					adder_op_a_shift3 = 1'b1;
			default:
				;
		endcase
	end
	always @(*)
		case (1'b1)
			multdiv_sel_i: adder_in_a = multdiv_operand_a_i;
			adder_op_a_shift1: adder_in_a = {operand_a_i[30:0], 2'b01};
			adder_op_a_shift2: adder_in_a = {operand_a_i[29:0], 3'b001};
			adder_op_a_shift3: adder_in_a = {operand_a_i[28:0], 4'b0001};
			default: adder_in_a = {operand_a_i, 1'b1};
		endcase
	assign operand_b_neg = {operand_b_i, 1'b0} ^ {33 {1'b1}};
	always @(*)
		case (1'b1)
			multdiv_sel_i: adder_in_b = multdiv_operand_b_i;
			adder_op_b_negate: adder_in_b = operand_b_neg;
			default: adder_in_b = {operand_b_i, 1'b0};
		endcase
	assign adder_result_ext_o = $unsigned(adder_in_a) + $unsigned(adder_in_b);
	assign adder_result = adder_result_ext_o[32:1];
	assign adder_result_o = adder_result;
	wire is_equal;
	reg is_greater_equal;
	reg cmp_signed;
	always @(*)
		case (operator_i)
			7'd27, 7'd25, 7'd43, 7'd31, 7'd33: cmp_signed = 1'b1;
			default: cmp_signed = 1'b0;
		endcase
	assign is_equal = adder_result == 32'b00000000000000000000000000000000;
	assign is_equal_result_o = is_equal;
	always @(*)
		if ((operand_a_i[31] ^ operand_b_i[31]) == 1'b0)
			is_greater_equal = adder_result[31] == 1'b0;
		else
			is_greater_equal = operand_a_i[31] ^ cmp_signed;
	reg cmp_result;
	always @(*)
		case (operator_i)
			7'd29: cmp_result = is_equal;
			7'd30: cmp_result = ~is_equal;
			7'd27, 7'd28, 7'd33, 7'd34: cmp_result = is_greater_equal;
			7'd25, 7'd26, 7'd31, 7'd32, 7'd43, 7'd44: cmp_result = ~is_greater_equal;
			default: cmp_result = is_equal;
		endcase
	assign comparison_result_o = cmp_result;
	reg shift_left;
	wire shift_ones;
	wire shift_arith;
	wire shift_funnel;
	wire shift_sbmode;
	reg [5:0] shift_amt;
	wire [5:0] shift_amt_compl;
	reg [31:0] shift_operand;
	reg signed [32:0] shift_result_ext_signed;
	reg [32:0] shift_result_ext;
	reg unused_shift_result_ext;
	reg [31:0] shift_result;
	reg [31:0] shift_result_rev;
	wire bfp_op;
	wire [4:0] bfp_len;
	wire [4:0] bfp_off;
	wire [31:0] bfp_mask;
	wire [31:0] bfp_mask_rev;
	wire [31:0] bfp_result;
	assign bfp_op = (RV32B != 32'sd0 ? operator_i == 7'd55 : 1'b0);
	assign bfp_len = {~(|operand_b_i[27:24]), operand_b_i[27:24]};
	assign bfp_off = operand_b_i[20:16];
	assign bfp_mask = (RV32B != 32'sd0 ? ~(32'hffffffff << bfp_len) : {32 {1'sb0}});
	genvar i;
	generate
		for (i = 0; i < 32; i = i + 1) begin : gen_rev_bfp_mask
			assign bfp_mask_rev[i] = bfp_mask[31 - i];
		end
	endgenerate
	assign bfp_result = (RV32B != 32'sd0 ? (~shift_result & operand_a_i) | ((operand_b_i & bfp_mask) << bfp_off) : {32 {1'sb0}});
	wire [1:1] sv2v_tmp_3EBA5;
	assign sv2v_tmp_3EBA5 = operand_b_i[5] & shift_funnel;
	always @(*) shift_amt[5] = sv2v_tmp_3EBA5;
	assign shift_amt_compl = 32 - operand_b_i[4:0];
	always @(*)
		if (bfp_op)
			shift_amt[4:0] = bfp_off;
		else
			shift_amt[4:0] = (instr_first_cycle_i ? (operand_b_i[5] && shift_funnel ? shift_amt_compl[4:0] : operand_b_i[4:0]) : (operand_b_i[5] && shift_funnel ? operand_b_i[4:0] : shift_amt_compl[4:0]));
	assign shift_sbmode = (RV32B != 32'sd0 ? ((operator_i == 7'd49) | (operator_i == 7'd50)) | (operator_i == 7'd51) : 1'b0);
	always @(*) begin
		case (operator_i)
			7'd10: shift_left = 1'b1;
			7'd12: shift_left = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? 1'b1 : 1'b0);
			7'd55: shift_left = (RV32B != 32'sd0 ? 1'b1 : 1'b0);
			7'd14: shift_left = (RV32B != 32'sd0 ? instr_first_cycle_i : 0);
			7'd13: shift_left = (RV32B != 32'sd0 ? ~instr_first_cycle_i : 0);
			7'd47: shift_left = (RV32B != 32'sd0 ? (shift_amt[5] ? ~instr_first_cycle_i : instr_first_cycle_i) : 1'b0);
			7'd48: shift_left = (RV32B != 32'sd0 ? (shift_amt[5] ? instr_first_cycle_i : ~instr_first_cycle_i) : 1'b0);
			default: shift_left = 1'b0;
		endcase
		if (shift_sbmode)
			shift_left = 1'b1;
	end
	assign shift_arith = operator_i == 7'd8;
	assign shift_ones = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? (operator_i == 7'd12) | (operator_i == 7'd11) : 1'b0);
	assign shift_funnel = (RV32B != 32'sd0 ? (operator_i == 7'd47) | (operator_i == 7'd48) : 1'b0);
	always @(*) begin
		if (RV32B == 32'sd0)
			shift_operand = (shift_left ? operand_a_rev : operand_a_i);
		else
			case (1'b1)
				bfp_op: shift_operand = bfp_mask_rev;
				shift_sbmode: shift_operand = 32'h80000000;
				default: shift_operand = (shift_left ? operand_a_rev : operand_a_i);
			endcase
		shift_result_ext_signed = $signed({shift_ones | (shift_arith & shift_operand[31]), shift_operand}) >>> shift_amt[4:0];
		shift_result_ext = $unsigned(shift_result_ext_signed);
		shift_result = shift_result_ext[31:0];
		unused_shift_result_ext = shift_result_ext[32];
		begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < 32; i = i + 1)
				shift_result_rev[i] = shift_result[31 - i];
		end
		shift_result = (shift_left ? shift_result_rev : shift_result);
	end
	wire bwlogic_or;
	wire bwlogic_and;
	wire [31:0] bwlogic_operand_b;
	wire [31:0] bwlogic_or_result;
	wire [31:0] bwlogic_and_result;
	wire [31:0] bwlogic_xor_result;
	reg [31:0] bwlogic_result;
	reg bwlogic_op_b_negate;
	always @(*)
		case (operator_i)
			7'd5, 7'd6, 7'd7: bwlogic_op_b_negate = (RV32B != 32'sd0 ? 1'b1 : 1'b0);
			7'd46: bwlogic_op_b_negate = (RV32B != 32'sd0 ? ~instr_first_cycle_i : 1'b0);
			default: bwlogic_op_b_negate = 1'b0;
		endcase
	assign bwlogic_operand_b = (bwlogic_op_b_negate ? operand_b_neg[32:1] : operand_b_i);
	assign bwlogic_or_result = operand_a_i | bwlogic_operand_b;
	assign bwlogic_and_result = operand_a_i & bwlogic_operand_b;
	assign bwlogic_xor_result = operand_a_i ^ bwlogic_operand_b;
	assign bwlogic_or = (operator_i == 7'd3) | (operator_i == 7'd6);
	assign bwlogic_and = (operator_i == 7'd4) | (operator_i == 7'd7);
	always @(*)
		case (1'b1)
			bwlogic_or: bwlogic_result = bwlogic_or_result;
			bwlogic_and: bwlogic_result = bwlogic_and_result;
			default: bwlogic_result = bwlogic_xor_result;
		endcase
	wire [5:0] bitcnt_result;
	wire [31:0] minmax_result;
	reg [31:0] pack_result;
	wire [31:0] sext_result;
	reg [31:0] singlebit_result;
	reg [31:0] rev_result;
	reg [31:0] shuffle_result;
	wire [31:0] xperm_result;
	reg [31:0] butterfly_result;
	reg [31:0] invbutterfly_result;
	reg [31:0] clmul_result;
	reg [31:0] multicycle_result;
	generate
		if (RV32B != 32'sd0) begin : g_alu_rvb
			wire zbe_op;
			wire bitcnt_ctz;
			wire bitcnt_clz;
			wire bitcnt_cz;
			reg [31:0] bitcnt_bits;
			wire [31:0] bitcnt_mask_op;
			reg [31:0] bitcnt_bit_mask;
			reg [191:0] bitcnt_partial;
			wire [31:0] bitcnt_partial_lsb_d;
			wire [31:0] bitcnt_partial_msb_d;
			assign bitcnt_ctz = operator_i == 7'd41;
			assign bitcnt_clz = operator_i == 7'd40;
			assign bitcnt_cz = bitcnt_ctz | bitcnt_clz;
			assign bitcnt_result = bitcnt_partial[0+:6];
			assign bitcnt_mask_op = (bitcnt_clz ? operand_a_rev : operand_a_i);
			always @(*) begin
				bitcnt_bit_mask = bitcnt_mask_op;
				bitcnt_bit_mask = bitcnt_bit_mask | (bitcnt_bit_mask << 1);
				bitcnt_bit_mask = bitcnt_bit_mask | (bitcnt_bit_mask << 2);
				bitcnt_bit_mask = bitcnt_bit_mask | (bitcnt_bit_mask << 4);
				bitcnt_bit_mask = bitcnt_bit_mask | (bitcnt_bit_mask << 8);
				bitcnt_bit_mask = bitcnt_bit_mask | (bitcnt_bit_mask << 16);
				bitcnt_bit_mask = ~bitcnt_bit_mask;
			end
			assign zbe_op = (operator_i == 7'd53) | (operator_i == 7'd54);
			always @(*)
				case (1'b1)
					zbe_op: bitcnt_bits = operand_b_i;
					bitcnt_cz: bitcnt_bits = bitcnt_bit_mask & ~bitcnt_mask_op;
					default: bitcnt_bits = operand_a_i;
				endcase
			always @(*) begin
				bitcnt_partial = {32 {6'b000000}};
				begin : sv2v_autoblock_2
					reg [31:0] i;
					for (i = 1; i < 32; i = i + 2)
						bitcnt_partial[(31 - i) * 6+:6] = {5'h00, bitcnt_bits[i]} + {5'h00, bitcnt_bits[i - 1]};
				end
				begin : sv2v_autoblock_3
					reg [31:0] i;
					for (i = 3; i < 32; i = i + 4)
						bitcnt_partial[(31 - i) * 6+:6] = bitcnt_partial[(33 - i) * 6+:6] + bitcnt_partial[(31 - i) * 6+:6];
				end
				begin : sv2v_autoblock_4
					reg [31:0] i;
					for (i = 7; i < 32; i = i + 8)
						bitcnt_partial[(31 - i) * 6+:6] = bitcnt_partial[(35 - i) * 6+:6] + bitcnt_partial[(31 - i) * 6+:6];
				end
				begin : sv2v_autoblock_5
					reg [31:0] i;
					for (i = 15; i < 32; i = i + 16)
						bitcnt_partial[(31 - i) * 6+:6] = bitcnt_partial[(39 - i) * 6+:6] + bitcnt_partial[(31 - i) * 6+:6];
				end
				bitcnt_partial[0+:6] = bitcnt_partial[96+:6] + bitcnt_partial[0+:6];
				bitcnt_partial[48+:6] = bitcnt_partial[96+:6] + bitcnt_partial[48+:6];
				begin : sv2v_autoblock_6
					reg [31:0] i;
					for (i = 11; i < 32; i = i + 8)
						bitcnt_partial[(31 - i) * 6+:6] = bitcnt_partial[(35 - i) * 6+:6] + bitcnt_partial[(31 - i) * 6+:6];
				end
				begin : sv2v_autoblock_7
					reg [31:0] i;
					for (i = 5; i < 32; i = i + 4)
						bitcnt_partial[(31 - i) * 6+:6] = bitcnt_partial[(33 - i) * 6+:6] + bitcnt_partial[(31 - i) * 6+:6];
				end
				bitcnt_partial[186+:6] = {5'h00, bitcnt_bits[0]};
				begin : sv2v_autoblock_8
					reg [31:0] i;
					for (i = 2; i < 32; i = i + 2)
						bitcnt_partial[(31 - i) * 6+:6] = bitcnt_partial[(32 - i) * 6+:6] + {5'h00, bitcnt_bits[i]};
				end
			end
			assign minmax_result = (cmp_result ? operand_a_i : operand_b_i);
			wire packu;
			wire packh;
			assign packu = operator_i == 7'd36;
			assign packh = operator_i == 7'd37;
			always @(*)
				case (1'b1)
					packu: pack_result = {operand_b_i[31:16], operand_a_i[31:16]};
					packh: pack_result = {16'h0000, operand_b_i[7:0], operand_a_i[7:0]};
					default: pack_result = {operand_b_i[15:0], operand_a_i[15:0]};
				endcase
			assign sext_result = (operator_i == 7'd38 ? {{24 {operand_a_i[7]}}, operand_a_i[7:0]} : {{16 {operand_a_i[15]}}, operand_a_i[15:0]});
			always @(*)
				case (operator_i)
					7'd49: singlebit_result = operand_a_i | shift_result;
					7'd50: singlebit_result = operand_a_i & ~shift_result;
					7'd51: singlebit_result = operand_a_i ^ shift_result;
					default: singlebit_result = {31'h00000000, shift_result[0]};
				endcase
			wire [4:0] zbp_shift_amt;
			wire gorc_op;
			assign gorc_op = operator_i == 7'd16;
			assign zbp_shift_amt[2:0] = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? shift_amt[2:0] : {3 {shift_amt[0]}});
			assign zbp_shift_amt[4:3] = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? shift_amt[4:3] : {2 {shift_amt[3]}});
			always @(*) begin
				rev_result = operand_a_i;
				if (zbp_shift_amt[0])
					rev_result = ((gorc_op ? rev_result : 32'h00000000) | ((rev_result & 32'h55555555) << 1)) | ((rev_result & 32'haaaaaaaa) >> 1);
				if (zbp_shift_amt[1])
					rev_result = ((gorc_op ? rev_result : 32'h00000000) | ((rev_result & 32'h33333333) << 2)) | ((rev_result & 32'hcccccccc) >> 2);
				if (zbp_shift_amt[2])
					rev_result = ((gorc_op ? rev_result : 32'h00000000) | ((rev_result & 32'h0f0f0f0f) << 4)) | ((rev_result & 32'hf0f0f0f0) >> 4);
				if (zbp_shift_amt[3])
					rev_result = ((((RV32B == 32'sd2) || (RV32B == 32'sd3)) && gorc_op ? rev_result : 32'h00000000) | ((rev_result & 32'h00ff00ff) << 8)) | ((rev_result & 32'hff00ff00) >> 8);
				if (zbp_shift_amt[4])
					rev_result = ((((RV32B == 32'sd2) || (RV32B == 32'sd3)) && gorc_op ? rev_result : 32'h00000000) | ((rev_result & 32'h0000ffff) << 16)) | ((rev_result & 32'hffff0000) >> 16);
			end
			wire crc_hmode;
			wire crc_bmode;
			wire [31:0] clmul_result_rev;
			if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin : gen_alu_rvb_otearlgrey_full
				localparam [127:0] SHUFFLE_MASK_L = 128'h00ff00000f000f003030303044444444;
				localparam [127:0] SHUFFLE_MASK_R = 128'h0000ff0000f000f00c0c0c0c22222222;
				localparam [127:0] FLIP_MASK_L = 128'h22001100004400004411000011000000;
				localparam [127:0] FLIP_MASK_R = 128'h00880044000022000000882200000088;
				wire [31:0] SHUFFLE_MASK_NOT [0:3];
				genvar i;
				for (i = 0; i < 4; i = i + 1) begin : gen_shuffle_mask_not
					assign SHUFFLE_MASK_NOT[i] = ~(SHUFFLE_MASK_L[(3 - i) * 32+:32] | SHUFFLE_MASK_R[(3 - i) * 32+:32]);
				end
				wire shuffle_flip;
				assign shuffle_flip = operator_i == 7'd18;
				reg [3:0] shuffle_mode;
				always @(*) begin
					shuffle_result = operand_a_i;
					if (shuffle_flip) begin
						shuffle_mode[3] = shift_amt[0];
						shuffle_mode[2] = shift_amt[1];
						shuffle_mode[1] = shift_amt[2];
						shuffle_mode[0] = shift_amt[3];
					end
					else
						shuffle_mode = shift_amt[3:0];
					if (shuffle_flip)
						shuffle_result = ((((((((shuffle_result & 32'h88224411) | ((shuffle_result << 6) & FLIP_MASK_L[96+:32])) | ((shuffle_result >> 6) & FLIP_MASK_R[96+:32])) | ((shuffle_result << 9) & FLIP_MASK_L[64+:32])) | ((shuffle_result >> 9) & FLIP_MASK_R[64+:32])) | ((shuffle_result << 15) & FLIP_MASK_L[32+:32])) | ((shuffle_result >> 15) & FLIP_MASK_R[32+:32])) | ((shuffle_result << 21) & FLIP_MASK_L[0+:32])) | ((shuffle_result >> 21) & FLIP_MASK_R[0+:32]);
					if (shuffle_mode[3])
						shuffle_result = (shuffle_result & SHUFFLE_MASK_NOT[0]) | (((shuffle_result << 8) & SHUFFLE_MASK_L[96+:32]) | ((shuffle_result >> 8) & SHUFFLE_MASK_R[96+:32]));
					if (shuffle_mode[2])
						shuffle_result = (shuffle_result & SHUFFLE_MASK_NOT[1]) | (((shuffle_result << 4) & SHUFFLE_MASK_L[64+:32]) | ((shuffle_result >> 4) & SHUFFLE_MASK_R[64+:32]));
					if (shuffle_mode[1])
						shuffle_result = (shuffle_result & SHUFFLE_MASK_NOT[2]) | (((shuffle_result << 2) & SHUFFLE_MASK_L[32+:32]) | ((shuffle_result >> 2) & SHUFFLE_MASK_R[32+:32]));
					if (shuffle_mode[0])
						shuffle_result = (shuffle_result & SHUFFLE_MASK_NOT[3]) | (((shuffle_result << 1) & SHUFFLE_MASK_L[0+:32]) | ((shuffle_result >> 1) & SHUFFLE_MASK_R[0+:32]));
					if (shuffle_flip)
						shuffle_result = ((((((((shuffle_result & 32'h88224411) | ((shuffle_result << 6) & FLIP_MASK_L[96+:32])) | ((shuffle_result >> 6) & FLIP_MASK_R[96+:32])) | ((shuffle_result << 9) & FLIP_MASK_L[64+:32])) | ((shuffle_result >> 9) & FLIP_MASK_R[64+:32])) | ((shuffle_result << 15) & FLIP_MASK_L[32+:32])) | ((shuffle_result >> 15) & FLIP_MASK_R[32+:32])) | ((shuffle_result << 21) & FLIP_MASK_L[0+:32])) | ((shuffle_result >> 21) & FLIP_MASK_R[0+:32]);
				end
				wire [23:0] sel_n;
				wire [7:0] vld_n;
				wire [7:0] sel_b;
				wire [3:0] vld_b;
				wire [1:0] sel_h;
				wire [1:0] vld_h;
				for (i = 0; i < 8; i = i + 1) begin : gen_sel_vld_n
					assign sel_n[i * 3+:3] = operand_b_i[i * 4+:3];
					assign vld_n[i] = ~|operand_b_i[(i * 4) + 3+:1];
				end
				for (i = 0; i < 4; i = i + 1) begin : gen_sel_vld_b
					assign sel_b[i * 2+:2] = operand_b_i[i * 8+:2];
					assign vld_b[i] = ~|operand_b_i[(i * 8) + 2+:6];
				end
				for (i = 0; i < 2; i = i + 1) begin : gen_sel_vld_h
					assign sel_h[i+:1] = operand_b_i[i * 16+:1];
					assign vld_h[i] = ~|operand_b_i[(i * 16) + 1+:15];
				end
				reg [23:0] sel;
				reg [7:0] vld;
				always @(*)
					case (operator_i)
						7'd19: begin
							sel = sel_n;
							vld = vld_n;
						end
						7'd20: begin : sv2v_autoblock_9
							reg signed [31:0] b;
							for (b = 0; b < 4; b = b + 1)
								begin
									sel[((b * 2) + 0) * 3+:3] = {sel_b[b * 2+:2], 1'b0};
									sel[((b * 2) + 1) * 3+:3] = {sel_b[b * 2+:2], 1'b1};
									vld[b * 2+:2] = {2 {vld_b[b]}};
								end
						end
						7'd21: begin : sv2v_autoblock_10
							reg signed [31:0] h;
							for (h = 0; h < 2; h = h + 1)
								begin
									sel[((h * 4) + 0) * 3+:3] = {sel_h[h+:1], 2'b00};
									sel[((h * 4) + 1) * 3+:3] = {sel_h[h+:1], 2'b01};
									sel[((h * 4) + 2) * 3+:3] = {sel_h[h+:1], 2'b10};
									sel[((h * 4) + 3) * 3+:3] = {sel_h[h+:1], 2'b11};
									vld[h * 4+:4] = {4 {vld_h[h]}};
								end
						end
						default: begin
							sel = sel_n;
							vld = 1'sb0;
						end
					endcase
				wire [31:0] val_n;
				wire [31:0] xperm_n;
				assign val_n = operand_a_i;
				for (i = 0; i < 8; i = i + 1) begin : gen_xperm_n
					assign xperm_n[i * 4+:4] = (vld[i] ? val_n[sel[i * 3+:3] * 4+:4] : {4 {1'sb0}});
				end
				assign xperm_result = xperm_n;
				wire clmul_rmode;
				wire clmul_hmode;
				reg [31:0] clmul_op_a;
				reg [31:0] clmul_op_b;
				wire [31:0] operand_b_rev;
				wire [31:0] clmul_and_stage [0:31];
				wire [31:0] clmul_xor_stage1 [0:15];
				wire [31:0] clmul_xor_stage2 [0:7];
				wire [31:0] clmul_xor_stage3 [0:3];
				wire [31:0] clmul_xor_stage4 [0:1];
				wire [31:0] clmul_result_raw;
				for (i = 0; i < 32; i = i + 1) begin : gen_rev_operand_b
					assign operand_b_rev[i] = operand_b_i[31 - i];
				end
				assign clmul_rmode = operator_i == 7'd57;
				assign clmul_hmode = operator_i == 7'd58;
				localparam [31:0] CRC32_POLYNOMIAL = 32'h04c11db7;
				localparam [31:0] CRC32_MU_REV = 32'hf7011641;
				localparam [31:0] CRC32C_POLYNOMIAL = 32'h1edc6f41;
				localparam [31:0] CRC32C_MU_REV = 32'hdea713f1;
				wire crc_op;
				wire crc_cpoly;
				reg [31:0] crc_operand;
				wire [31:0] crc_poly;
				wire [31:0] crc_mu_rev;
				assign crc_op = (((((operator_i == 7'd64) | (operator_i == 7'd63)) | (operator_i == 7'd62)) | (operator_i == 7'd61)) | (operator_i == 7'd60)) | (operator_i == 7'd59);
				assign crc_cpoly = ((operator_i == 7'd64) | (operator_i == 7'd62)) | (operator_i == 7'd60);
				assign crc_hmode = (operator_i == 7'd61) | (operator_i == 7'd62);
				assign crc_bmode = (operator_i == 7'd59) | (operator_i == 7'd60);
				assign crc_poly = (crc_cpoly ? CRC32C_POLYNOMIAL : CRC32_POLYNOMIAL);
				assign crc_mu_rev = (crc_cpoly ? CRC32C_MU_REV : CRC32_MU_REV);
				always @(*)
					case (1'b1)
						crc_bmode: crc_operand = {operand_a_i[7:0], 24'h000000};
						crc_hmode: crc_operand = {operand_a_i[15:0], 16'h0000};
						default: crc_operand = operand_a_i;
					endcase
				always @(*)
					if (crc_op) begin
						clmul_op_a = (instr_first_cycle_i ? crc_operand : imd_val_q_i[32+:32]);
						clmul_op_b = (instr_first_cycle_i ? crc_mu_rev : crc_poly);
					end
					else begin
						clmul_op_a = (clmul_rmode | clmul_hmode ? operand_a_rev : operand_a_i);
						clmul_op_b = (clmul_rmode | clmul_hmode ? operand_b_rev : operand_b_i);
					end
				for (i = 0; i < 32; i = i + 1) begin : gen_clmul_and_op
					assign clmul_and_stage[i] = (clmul_op_b[i] ? clmul_op_a << i : {32 {1'sb0}});
				end
				for (i = 0; i < 16; i = i + 1) begin : gen_clmul_xor_op_l1
					assign clmul_xor_stage1[i] = clmul_and_stage[2 * i] ^ clmul_and_stage[(2 * i) + 1];
				end
				for (i = 0; i < 8; i = i + 1) begin : gen_clmul_xor_op_l2
					assign clmul_xor_stage2[i] = clmul_xor_stage1[2 * i] ^ clmul_xor_stage1[(2 * i) + 1];
				end
				for (i = 0; i < 4; i = i + 1) begin : gen_clmul_xor_op_l3
					assign clmul_xor_stage3[i] = clmul_xor_stage2[2 * i] ^ clmul_xor_stage2[(2 * i) + 1];
				end
				for (i = 0; i < 2; i = i + 1) begin : gen_clmul_xor_op_l4
					assign clmul_xor_stage4[i] = clmul_xor_stage3[2 * i] ^ clmul_xor_stage3[(2 * i) + 1];
				end
				assign clmul_result_raw = clmul_xor_stage4[0] ^ clmul_xor_stage4[1];
				for (i = 0; i < 32; i = i + 1) begin : gen_rev_clmul_result
					assign clmul_result_rev[i] = clmul_result_raw[31 - i];
				end
				always @(*)
					case (1'b1)
						clmul_rmode: clmul_result = clmul_result_rev;
						clmul_hmode: clmul_result = {1'b0, clmul_result_rev[31:1]};
						default: clmul_result = clmul_result_raw;
					endcase
			end
			else begin : gen_alu_rvb_not_otearlgrey_full
				wire [32:1] sv2v_tmp_F189D;
				assign sv2v_tmp_F189D = 1'sb0;
				always @(*) shuffle_result = sv2v_tmp_F189D;
				assign xperm_result = 1'sb0;
				wire [32:1] sv2v_tmp_B9A55;
				assign sv2v_tmp_B9A55 = 1'sb0;
				always @(*) clmul_result = sv2v_tmp_B9A55;
				assign clmul_result_rev = 1'sb0;
				assign crc_bmode = 1'sb0;
				assign crc_hmode = 1'sb0;
			end
			if (RV32B == 32'sd3) begin : gen_alu_rvb_full
				reg [191:0] bitcnt_partial_q;
				genvar i;
				for (i = 0; i < 32; i = i + 1) begin : gen_bitcnt_reg_in_lsb
					assign bitcnt_partial_lsb_d[i] = bitcnt_partial[(31 - i) * 6];
				end
				for (i = 0; i < 16; i = i + 1) begin : gen_bitcnt_reg_in_b1
					assign bitcnt_partial_msb_d[i] = bitcnt_partial[((31 - ((2 * i) + 1)) * 6) + 1];
				end
				for (i = 0; i < 8; i = i + 1) begin : gen_bitcnt_reg_in_b2
					assign bitcnt_partial_msb_d[16 + i] = bitcnt_partial[((31 - ((4 * i) + 3)) * 6) + 2];
				end
				for (i = 0; i < 4; i = i + 1) begin : gen_bitcnt_reg_in_b3
					assign bitcnt_partial_msb_d[24 + i] = bitcnt_partial[((31 - ((8 * i) + 7)) * 6) + 3];
				end
				for (i = 0; i < 2; i = i + 1) begin : gen_bitcnt_reg_in_b4
					assign bitcnt_partial_msb_d[28 + i] = bitcnt_partial[((31 - ((16 * i) + 15)) * 6) + 4];
				end
				assign bitcnt_partial_msb_d[30] = bitcnt_partial[5];
				assign bitcnt_partial_msb_d[31] = 1'b0;
				always @(*) begin
					bitcnt_partial_q = {32 {6'b000000}};
					begin : sv2v_autoblock_11
						reg [31:0] i;
						for (i = 0; i < 32; i = i + 1)
							begin : gen_bitcnt_reg_out_lsb
								bitcnt_partial_q[(31 - i) * 6] = imd_val_q_i[32 + i];
							end
					end
					begin : sv2v_autoblock_12
						reg [31:0] i;
						for (i = 0; i < 16; i = i + 1)
							begin : gen_bitcnt_reg_out_b1
								bitcnt_partial_q[((31 - ((2 * i) + 1)) * 6) + 1] = imd_val_q_i[0 + i];
							end
					end
					begin : sv2v_autoblock_13
						reg [31:0] i;
						for (i = 0; i < 8; i = i + 1)
							begin : gen_bitcnt_reg_out_b2
								bitcnt_partial_q[((31 - ((4 * i) + 3)) * 6) + 2] = imd_val_q_i[16 + i];
							end
					end
					begin : sv2v_autoblock_14
						reg [31:0] i;
						for (i = 0; i < 4; i = i + 1)
							begin : gen_bitcnt_reg_out_b3
								bitcnt_partial_q[((31 - ((8 * i) + 7)) * 6) + 3] = imd_val_q_i[24 + i];
							end
					end
					begin : sv2v_autoblock_15
						reg [31:0] i;
						for (i = 0; i < 2; i = i + 1)
							begin : gen_bitcnt_reg_out_b4
								bitcnt_partial_q[((31 - ((16 * i) + 15)) * 6) + 4] = imd_val_q_i[28 + i];
							end
					end
					bitcnt_partial_q[5] = imd_val_q_i[30];
				end
				wire [31:0] butterfly_mask_l [0:4];
				wire [31:0] butterfly_mask_r [0:4];
				wire [31:0] butterfly_mask_not [0:4];
				wire [31:0] lrotc_stage [0:4];
				genvar stg;
				for (stg = 0; stg < 5; stg = stg + 1) begin : gen_butterfly_ctrl_stage
					genvar seg;
					for (seg = 0; seg < (2 ** stg); seg = seg + 1) begin : gen_butterfly_ctrl
						assign lrotc_stage[stg][((2 * (16 >> stg)) * (seg + 1)) - 1:(2 * (16 >> stg)) * seg] = {{16 >> stg {1'b0}}, {16 >> stg {1'b1}}} << bitcnt_partial_q[((32 - ((16 >> stg) * ((2 * seg) + 1))) * 6) + ($clog2(16 >> stg) >= 0 ? $clog2(16 >> stg) : ($clog2(16 >> stg) + ($clog2(16 >> stg) >= 0 ? $clog2(16 >> stg) + 1 : 1 - $clog2(16 >> stg))) - 1)-:($clog2(16 >> stg) >= 0 ? $clog2(16 >> stg) + 1 : 1 - $clog2(16 >> stg))];
						assign butterfly_mask_l[stg][((16 >> stg) * ((2 * seg) + 2)) - 1:(16 >> stg) * ((2 * seg) + 1)] = ~lrotc_stage[stg][((16 >> stg) * ((2 * seg) + 2)) - 1:(16 >> stg) * ((2 * seg) + 1)];
						assign butterfly_mask_r[stg][((16 >> stg) * ((2 * seg) + 1)) - 1:(16 >> stg) * (2 * seg)] = ~lrotc_stage[stg][((16 >> stg) * ((2 * seg) + 2)) - 1:(16 >> stg) * ((2 * seg) + 1)];
						assign butterfly_mask_l[stg][((16 >> stg) * ((2 * seg) + 1)) - 1:(16 >> stg) * (2 * seg)] = 1'sb0;
						assign butterfly_mask_r[stg][((16 >> stg) * ((2 * seg) + 2)) - 1:(16 >> stg) * ((2 * seg) + 1)] = 1'sb0;
					end
				end
				for (stg = 0; stg < 5; stg = stg + 1) begin : gen_butterfly_not
					assign butterfly_mask_not[stg] = ~(butterfly_mask_l[stg] | butterfly_mask_r[stg]);
				end
				always @(*) begin
					butterfly_result = operand_a_i;
					butterfly_result = ((butterfly_result & butterfly_mask_not[0]) | ((butterfly_result & butterfly_mask_l[0]) >> 16)) | ((butterfly_result & butterfly_mask_r[0]) << 16);
					butterfly_result = ((butterfly_result & butterfly_mask_not[1]) | ((butterfly_result & butterfly_mask_l[1]) >> 8)) | ((butterfly_result & butterfly_mask_r[1]) << 8);
					butterfly_result = ((butterfly_result & butterfly_mask_not[2]) | ((butterfly_result & butterfly_mask_l[2]) >> 4)) | ((butterfly_result & butterfly_mask_r[2]) << 4);
					butterfly_result = ((butterfly_result & butterfly_mask_not[3]) | ((butterfly_result & butterfly_mask_l[3]) >> 2)) | ((butterfly_result & butterfly_mask_r[3]) << 2);
					butterfly_result = ((butterfly_result & butterfly_mask_not[4]) | ((butterfly_result & butterfly_mask_l[4]) >> 1)) | ((butterfly_result & butterfly_mask_r[4]) << 1);
					butterfly_result = butterfly_result & operand_b_i;
				end
				always @(*) begin
					invbutterfly_result = operand_a_i & operand_b_i;
					invbutterfly_result = ((invbutterfly_result & butterfly_mask_not[4]) | ((invbutterfly_result & butterfly_mask_l[4]) >> 1)) | ((invbutterfly_result & butterfly_mask_r[4]) << 1);
					invbutterfly_result = ((invbutterfly_result & butterfly_mask_not[3]) | ((invbutterfly_result & butterfly_mask_l[3]) >> 2)) | ((invbutterfly_result & butterfly_mask_r[3]) << 2);
					invbutterfly_result = ((invbutterfly_result & butterfly_mask_not[2]) | ((invbutterfly_result & butterfly_mask_l[2]) >> 4)) | ((invbutterfly_result & butterfly_mask_r[2]) << 4);
					invbutterfly_result = ((invbutterfly_result & butterfly_mask_not[1]) | ((invbutterfly_result & butterfly_mask_l[1]) >> 8)) | ((invbutterfly_result & butterfly_mask_r[1]) << 8);
					invbutterfly_result = ((invbutterfly_result & butterfly_mask_not[0]) | ((invbutterfly_result & butterfly_mask_l[0]) >> 16)) | ((invbutterfly_result & butterfly_mask_r[0]) << 16);
				end
			end
			else begin : gen_alu_rvb_not_full
				wire [31:0] unused_imd_val_q_1;
				assign unused_imd_val_q_1 = imd_val_q_i[0+:32];
				wire [32:1] sv2v_tmp_F770D;
				assign sv2v_tmp_F770D = 1'sb0;
				always @(*) butterfly_result = sv2v_tmp_F770D;
				wire [32:1] sv2v_tmp_02B8B;
				assign sv2v_tmp_02B8B = 1'sb0;
				always @(*) invbutterfly_result = sv2v_tmp_02B8B;
				assign bitcnt_partial_lsb_d = 1'sb0;
				assign bitcnt_partial_msb_d = 1'sb0;
			end
			always @(*)
				case (operator_i)
					7'd45: begin
						multicycle_result = (operand_b_i == 32'h00000000 ? operand_a_i : imd_val_q_i[32+:32]);
						imd_val_d_o = {operand_a_i, 32'h00000000};
						if (instr_first_cycle_i)
							imd_val_we_o = 2'b01;
						else
							imd_val_we_o = 2'b00;
					end
					7'd46: begin
						multicycle_result = imd_val_q_i[32+:32] | bwlogic_and_result;
						imd_val_d_o = {bwlogic_and_result, 32'h00000000};
						if (instr_first_cycle_i)
							imd_val_we_o = 2'b01;
						else
							imd_val_we_o = 2'b00;
					end
					7'd48, 7'd47, 7'd14, 7'd13: begin
						if (shift_amt[4:0] == 5'h00)
							multicycle_result = (shift_amt[5] ? operand_a_i : imd_val_q_i[32+:32]);
						else
							multicycle_result = imd_val_q_i[32+:32] | shift_result;
						imd_val_d_o = {shift_result, 32'h00000000};
						if (instr_first_cycle_i)
							imd_val_we_o = 2'b01;
						else
							imd_val_we_o = 2'b00;
					end
					7'd63, 7'd64, 7'd61, 7'd62, 7'd59, 7'd60:
						if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin
							case (1'b1)
								crc_bmode: multicycle_result = clmul_result_rev ^ (operand_a_i >> 8);
								crc_hmode: multicycle_result = clmul_result_rev ^ (operand_a_i >> 16);
								default: multicycle_result = clmul_result_rev;
							endcase
							imd_val_d_o = {clmul_result_rev, 32'h00000000};
							if (instr_first_cycle_i)
								imd_val_we_o = 2'b01;
							else
								imd_val_we_o = 2'b00;
						end
						else begin
							imd_val_d_o = {operand_a_i, 32'h00000000};
							imd_val_we_o = 2'b00;
							multicycle_result = 1'sb0;
						end
					7'd53, 7'd54:
						if (RV32B == 32'sd3) begin
							multicycle_result = (operator_i == 7'd54 ? butterfly_result : invbutterfly_result);
							imd_val_d_o = {bitcnt_partial_lsb_d, bitcnt_partial_msb_d};
							if (instr_first_cycle_i)
								imd_val_we_o = 2'b11;
							else
								imd_val_we_o = 2'b00;
						end
						else begin
							imd_val_d_o = {operand_a_i, 32'h00000000};
							imd_val_we_o = 2'b00;
							multicycle_result = 1'sb0;
						end
					default: begin
						imd_val_d_o = {operand_a_i, 32'h00000000};
						imd_val_we_o = 2'b00;
						multicycle_result = 1'sb0;
					end
				endcase
		end
		else begin : g_no_alu_rvb
			wire [63:0] unused_imd_val_q;
			assign unused_imd_val_q = imd_val_q_i;
			wire [31:0] unused_butterfly_result;
			assign unused_butterfly_result = butterfly_result;
			wire [31:0] unused_invbutterfly_result;
			assign unused_invbutterfly_result = invbutterfly_result;
			assign bitcnt_result = 1'sb0;
			assign minmax_result = 1'sb0;
			wire [32:1] sv2v_tmp_B3EA0;
			assign sv2v_tmp_B3EA0 = 1'sb0;
			always @(*) pack_result = sv2v_tmp_B3EA0;
			assign sext_result = 1'sb0;
			wire [32:1] sv2v_tmp_C8829;
			assign sv2v_tmp_C8829 = 1'sb0;
			always @(*) singlebit_result = sv2v_tmp_C8829;
			wire [32:1] sv2v_tmp_F744D;
			assign sv2v_tmp_F744D = 1'sb0;
			always @(*) rev_result = sv2v_tmp_F744D;
			wire [32:1] sv2v_tmp_F189D;
			assign sv2v_tmp_F189D = 1'sb0;
			always @(*) shuffle_result = sv2v_tmp_F189D;
			assign xperm_result = 1'sb0;
			wire [32:1] sv2v_tmp_F770D;
			assign sv2v_tmp_F770D = 1'sb0;
			always @(*) butterfly_result = sv2v_tmp_F770D;
			wire [32:1] sv2v_tmp_02B8B;
			assign sv2v_tmp_02B8B = 1'sb0;
			always @(*) invbutterfly_result = sv2v_tmp_02B8B;
			wire [32:1] sv2v_tmp_B9A55;
			assign sv2v_tmp_B9A55 = 1'sb0;
			always @(*) clmul_result = sv2v_tmp_B9A55;
			wire [32:1] sv2v_tmp_8750A;
			assign sv2v_tmp_8750A = 1'sb0;
			always @(*) multicycle_result = sv2v_tmp_8750A;
			wire [64:1] sv2v_tmp_78BC2;
			assign sv2v_tmp_78BC2 = {2 {32'b00000000000000000000000000000000}};
			always @(*) imd_val_d_o = sv2v_tmp_78BC2;
			wire [2:1] sv2v_tmp_02FDF;
			assign sv2v_tmp_02FDF = {2 {1'b0}};
			always @(*) imd_val_we_o = sv2v_tmp_02FDF;
		end
	endgenerate
	always @(*) begin
		result_o = 1'sb0;
		case (operator_i)
			7'd2, 7'd5, 7'd3, 7'd6, 7'd4, 7'd7: result_o = bwlogic_result;
			7'd0, 7'd1, 7'd22, 7'd23, 7'd24: result_o = adder_result;
			7'd10, 7'd9, 7'd8, 7'd12, 7'd11: result_o = shift_result;
			7'd17, 7'd18: result_o = shuffle_result;
			7'd19, 7'd20, 7'd21: result_o = xperm_result;
			7'd29, 7'd30, 7'd27, 7'd28, 7'd25, 7'd26, 7'd43, 7'd44: result_o = {31'h00000000, cmp_result};
			7'd31, 7'd33, 7'd32, 7'd34: result_o = minmax_result;
			7'd40, 7'd41, 7'd42: result_o = {26'h0000000, bitcnt_result};
			7'd35, 7'd37, 7'd36: result_o = pack_result;
			7'd38, 7'd39: result_o = sext_result;
			7'd46, 7'd45, 7'd47, 7'd48, 7'd14, 7'd13, 7'd63, 7'd64, 7'd61, 7'd62, 7'd59, 7'd60, 7'd53, 7'd54: result_o = multicycle_result;
			7'd49, 7'd50, 7'd51, 7'd52: result_o = singlebit_result;
			7'd15, 7'd16: result_o = rev_result;
			7'd55: result_o = bfp_result;
			7'd56, 7'd57, 7'd58: result_o = clmul_result;
			default:
				;
		endcase
	end
	wire unused_shift_amt_compl;
	assign unused_shift_amt_compl = shift_amt_compl[5];
endmodule
module ibex_branch_predict (
	clk_i,
	rst_ni,
	fetch_rdata_i,
	fetch_pc_i,
	fetch_valid_i,
	predict_branch_taken_o,
	predict_branch_pc_o
);
	input wire clk_i;
	input wire rst_ni;
	input wire [31:0] fetch_rdata_i;
	input wire [31:0] fetch_pc_i;
	input wire fetch_valid_i;
	output wire predict_branch_taken_o;
	output wire [31:0] predict_branch_pc_o;
	wire [31:0] imm_j_type;
	wire [31:0] imm_b_type;
	wire [31:0] imm_cj_type;
	wire [31:0] imm_cb_type;
	reg [31:0] branch_imm;
	wire [31:0] instr;
	wire instr_j;
	wire instr_b;
	wire instr_cj;
	wire instr_cb;
	wire instr_b_taken;
	assign instr = fetch_rdata_i;
	assign imm_j_type = {{12 {instr[31]}}, instr[19:12], instr[20], instr[30:21], 1'b0};
	assign imm_b_type = {{19 {instr[31]}}, instr[31], instr[7], instr[30:25], instr[11:8], 1'b0};
	assign imm_cj_type = {{20 {instr[12]}}, instr[12], instr[8], instr[10:9], instr[6], instr[7], instr[2], instr[11], instr[5:3], 1'b0};
	assign imm_cb_type = {{23 {instr[12]}}, instr[12], instr[6:5], instr[2], instr[11:10], instr[4:3], 1'b0};
	assign instr_b = instr[6:0] == 7'h63;
	assign instr_j = instr[6:0] == 7'h6f;
	assign instr_cb = (instr[1:0] == 2'b01) & ((instr[15:13] == 3'b110) | (instr[15:13] == 3'b111));
	assign instr_cj = (instr[1:0] == 2'b01) & ((instr[15:13] == 3'b101) | (instr[15:13] == 3'b001));
	always @(*) begin
		branch_imm = imm_b_type;
		case (1'b1)
			instr_j: branch_imm = imm_j_type;
			instr_b: branch_imm = imm_b_type;
			instr_cj: branch_imm = imm_cj_type;
			instr_cb: branch_imm = imm_cb_type;
			default:
				;
		endcase
	end
	assign instr_b_taken = (instr_b & imm_b_type[31]) | (instr_cb & imm_cb_type[31]);
	assign predict_branch_taken_o = fetch_valid_i & ((instr_j | instr_cj) | instr_b_taken);
	assign predict_branch_pc_o = fetch_pc_i + branch_imm;
endmodule
module ibex_compressed_decoder (
	clk_i,
	rst_ni,
	valid_i,
	instr_i,
	instr_o,
	is_compressed_o,
	illegal_instr_o
);
	input wire clk_i;
	input wire rst_ni;
	input wire valid_i;
	input wire [31:0] instr_i;
	output reg [31:0] instr_o;
	output wire is_compressed_o;
	output reg illegal_instr_o;
	wire unused_valid;
	assign unused_valid = valid_i;
	always @(*) begin
		instr_o = instr_i;
		illegal_instr_o = 1'b0;
		case (instr_i[1:0])
			2'b00:
				case (instr_i[15:13])
					3'b000: begin
						instr_o = {2'b00, instr_i[10:7], instr_i[12:11], instr_i[5], instr_i[6], 2'b00, 5'h02, 3'b000, 2'b01, instr_i[4:2], 7'h13};
						if (instr_i[12:5] == 8'b00000000)
							illegal_instr_o = 1'b1;
					end
					3'b010: instr_o = {5'b00000, instr_i[5], instr_i[12:10], instr_i[6], 2'b00, 2'b01, instr_i[9:7], 3'b010, 2'b01, instr_i[4:2], 7'h03};
					3'b110: instr_o = {5'b00000, instr_i[5], instr_i[12], 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b010, instr_i[11:10], instr_i[6], 2'b00, 7'h23};
					3'b001, 3'b011, 3'b100, 3'b101, 3'b111: illegal_instr_o = 1'b1;
					default: illegal_instr_o = 1'b1;
				endcase
			2'b01:
				case (instr_i[15:13])
					3'b000: instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], instr_i[11:7], 3'b000, instr_i[11:7], 7'h13};
					3'b001, 3'b101: instr_o = {instr_i[12], instr_i[8], instr_i[10:9], instr_i[6], instr_i[7], instr_i[2], instr_i[11], instr_i[5:3], {9 {instr_i[12]}}, 4'b0000, ~instr_i[15], 7'h6f};
					3'b010: instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], 5'b00000, 3'b000, instr_i[11:7], 7'h13};
					3'b011: begin
						instr_o = {{15 {instr_i[12]}}, instr_i[6:2], instr_i[11:7], 7'h37};
						if (instr_i[11:7] == 5'h02)
							instr_o = {{3 {instr_i[12]}}, instr_i[4:3], instr_i[5], instr_i[2], instr_i[6], 4'b0000, 5'h02, 3'b000, 5'h02, 7'h13};
						if ({instr_i[12], instr_i[6:2]} == 6'b000000)
							illegal_instr_o = 1'b1;
					end
					3'b100:
						case (instr_i[11:10])
							2'b00, 2'b01: begin
								instr_o = {1'b0, instr_i[10], 5'b00000, instr_i[6:2], 2'b01, instr_i[9:7], 3'b101, 2'b01, instr_i[9:7], 7'h13};
								if (instr_i[12] == 1'b1)
									illegal_instr_o = 1'b1;
							end
							2'b10: instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], 2'b01, instr_i[9:7], 3'b111, 2'b01, instr_i[9:7], 7'h13};
							2'b11:
								case ({instr_i[12], instr_i[6:5]})
									3'b000: instr_o = {9'b010000001, instr_i[4:2], 2'b01, instr_i[9:7], 3'b000, 2'b01, instr_i[9:7], 7'h33};
									3'b001: instr_o = {9'b000000001, instr_i[4:2], 2'b01, instr_i[9:7], 3'b100, 2'b01, instr_i[9:7], 7'h33};
									3'b010: instr_o = {9'b000000001, instr_i[4:2], 2'b01, instr_i[9:7], 3'b110, 2'b01, instr_i[9:7], 7'h33};
									3'b011: instr_o = {9'b000000001, instr_i[4:2], 2'b01, instr_i[9:7], 3'b111, 2'b01, instr_i[9:7], 7'h33};
									3'b100, 3'b101, 3'b110, 3'b111: illegal_instr_o = 1'b1;
									default: illegal_instr_o = 1'b1;
								endcase
							default: illegal_instr_o = 1'b1;
						endcase
					3'b110, 3'b111: instr_o = {{4 {instr_i[12]}}, instr_i[6:5], instr_i[2], 5'b00000, 2'b01, instr_i[9:7], 2'b00, instr_i[13], instr_i[11:10], instr_i[4:3], instr_i[12], 7'h63};
					default: illegal_instr_o = 1'b1;
				endcase
			2'b10:
				case (instr_i[15:13])
					3'b000: begin
						instr_o = {7'b0000000, instr_i[6:2], instr_i[11:7], 3'b001, instr_i[11:7], 7'h13};
						if (instr_i[12] == 1'b1)
							illegal_instr_o = 1'b1;
					end
					3'b010: begin
						instr_o = {4'b0000, instr_i[3:2], instr_i[12], instr_i[6:4], 2'b00, 5'h02, 3'b010, instr_i[11:7], 7'h03};
						if (instr_i[11:7] == 5'b00000)
							illegal_instr_o = 1'b1;
					end
					3'b100:
						if (instr_i[12] == 1'b0) begin
							if (instr_i[6:2] != 5'b00000)
								instr_o = {7'b0000000, instr_i[6:2], 5'b00000, 3'b000, instr_i[11:7], 7'h33};
							else begin
								instr_o = {12'b000000000000, instr_i[11:7], 3'b000, 5'b00000, 7'h67};
								if (instr_i[11:7] == 5'b00000)
									illegal_instr_o = 1'b1;
							end
						end
						else if (instr_i[6:2] != 5'b00000)
							instr_o = {7'b0000000, instr_i[6:2], instr_i[11:7], 3'b000, instr_i[11:7], 7'h33};
						else if (instr_i[11:7] == 5'b00000)
							instr_o = 32'h00100073;
						else
							instr_o = {12'b000000000000, instr_i[11:7], 3'b000, 5'b00001, 7'h67};
					3'b110: instr_o = {4'b0000, instr_i[8:7], instr_i[12], instr_i[6:2], 5'h02, 3'b010, instr_i[11:9], 2'b00, 7'h23};
					3'b001, 3'b011, 3'b101, 3'b111: illegal_instr_o = 1'b1;
					default: illegal_instr_o = 1'b1;
				endcase
			2'b11:
				;
			default: illegal_instr_o = 1'b1;
		endcase
	end
	assign is_compressed_o = instr_i[1:0] != 2'b11;
endmodule
module ibex_controller (
	clk_i,
	rst_ni,
	ctrl_busy_o,
	illegal_insn_i,
	ecall_insn_i,
	mret_insn_i,
	dret_insn_i,
	wfi_insn_i,
	ebrk_insn_i,
	csr_pipe_flush_i,
	instr_valid_i,
	instr_i,
	instr_compressed_i,
	instr_is_compressed_i,
	instr_bp_taken_i,
	instr_fetch_err_i,
	instr_fetch_err_plus2_i,
	pc_id_i,
	instr_valid_clear_o,
	id_in_ready_o,
	controller_run_o,
	instr_exec_i,
	instr_req_o,
	pc_set_o,
	pc_mux_o,
	nt_branch_mispredict_o,
	exc_pc_mux_o,
	exc_cause_o,
	lsu_addr_last_i,
	load_err_i,
	store_err_i,
	mem_resp_intg_err_i,
	wb_exception_o,
	id_exception_o,
	branch_set_i,
	branch_not_set_i,
	jump_set_i,
	csr_mstatus_mie_i,
	irq_pending_i,
	irqs_i,
	irq_nm_ext_i,
	nmi_mode_o,
	debug_req_i,
	debug_cause_o,
	debug_csr_save_o,
	debug_mode_o,
	debug_mode_entering_o,
	debug_single_step_i,
	debug_ebreakm_i,
	debug_ebreaku_i,
	trigger_match_i,
	csr_save_if_o,
	csr_save_id_o,
	csr_save_wb_o,
	csr_restore_mret_id_o,
	csr_restore_dret_id_o,
	csr_save_cause_o,
	csr_mtval_o,
	priv_mode_i,
	stall_id_i,
	stall_wb_i,
	flush_id_o,
	ready_wb_i,
	perf_jump_o,
	perf_tbranch_o
);
	parameter [0:0] WritebackStage = 1'b0;
	parameter [0:0] BranchPredictor = 1'b0;
	parameter [0:0] MemECC = 1'b0;
	input wire clk_i;
	input wire rst_ni;
	output reg ctrl_busy_o;
	input wire illegal_insn_i;
	input wire ecall_insn_i;
	input wire mret_insn_i;
	input wire dret_insn_i;
	input wire wfi_insn_i;
	input wire ebrk_insn_i;
	input wire csr_pipe_flush_i;
	input wire instr_valid_i;
	input wire [31:0] instr_i;
	input wire [15:0] instr_compressed_i;
	input wire instr_is_compressed_i;
	input wire instr_bp_taken_i;
	input wire instr_fetch_err_i;
	input wire instr_fetch_err_plus2_i;
	input wire [31:0] pc_id_i;
	output wire instr_valid_clear_o;
	output wire id_in_ready_o;
	output reg controller_run_o;
	input wire instr_exec_i;
	output reg instr_req_o;
	output reg pc_set_o;
	output reg [2:0] pc_mux_o;
	output reg nt_branch_mispredict_o;
	output reg [1:0] exc_pc_mux_o;
	output reg [6:0] exc_cause_o;
	input wire [31:0] lsu_addr_last_i;
	input wire load_err_i;
	input wire store_err_i;
	input wire mem_resp_intg_err_i;
	output wire wb_exception_o;
	output wire id_exception_o;
	input wire branch_set_i;
	input wire branch_not_set_i;
	input wire jump_set_i;
	input wire csr_mstatus_mie_i;
	input wire irq_pending_i;
	input wire [17:0] irqs_i;
	input wire irq_nm_ext_i;
	output wire nmi_mode_o;
	input wire debug_req_i;
	output wire [2:0] debug_cause_o;
	output reg debug_csr_save_o;
	output wire debug_mode_o;
	output reg debug_mode_entering_o;
	input wire debug_single_step_i;
	input wire debug_ebreakm_i;
	input wire debug_ebreaku_i;
	input wire trigger_match_i;
	output reg csr_save_if_o;
	output reg csr_save_id_o;
	output reg csr_save_wb_o;
	output reg csr_restore_mret_id_o;
	output reg csr_restore_dret_id_o;
	output reg csr_save_cause_o;
	output reg [31:0] csr_mtval_o;
	input wire [1:0] priv_mode_i;
	input wire stall_id_i;
	input wire stall_wb_i;
	output wire flush_id_o;
	input wire ready_wb_i;
	output reg perf_jump_o;
	output reg perf_tbranch_o;
	reg [3:0] ctrl_fsm_cs;
	reg [3:0] ctrl_fsm_ns;
	reg nmi_mode_q;
	reg nmi_mode_d;
	reg debug_mode_q;
	reg debug_mode_d;
	wire [2:0] debug_cause_d;
	reg [2:0] debug_cause_q;
	reg load_err_q;
	wire load_err_d;
	reg store_err_q;
	wire store_err_d;
	reg exc_req_q;
	wire exc_req_d;
	reg illegal_insn_q;
	wire illegal_insn_d;
	reg instr_fetch_err_prio;
	reg illegal_insn_prio;
	reg ecall_insn_prio;
	reg ebrk_insn_prio;
	reg store_err_prio;
	reg load_err_prio;
	wire stall;
	reg halt_if;
	reg retain_id;
	reg flush_id;
	wire exc_req_lsu;
	wire special_req;
	wire special_req_pc_change;
	wire special_req_flush_only;
	wire do_single_step_d;
	reg do_single_step_q;
	wire enter_debug_mode_prio_d;
	reg enter_debug_mode_prio_q;
	wire enter_debug_mode;
	wire ebreak_into_debug;
	wire irq_enabled;
	wire handle_irq;
	wire id_wb_pending;
	wire irq_nm;
	wire irq_nm_int;
	wire [31:0] irq_nm_int_mtval;
	wire [4:0] irq_nm_int_cause;
	reg [3:0] mfip_id;
	wire unused_irq_timer;
	wire ecall_insn;
	wire mret_insn;
	wire dret_insn;
	wire wfi_insn;
	wire ebrk_insn;
	wire csr_pipe_flush;
	wire instr_fetch_err;
	assign load_err_d = load_err_i;
	assign store_err_d = store_err_i;
	assign ecall_insn = ecall_insn_i & instr_valid_i;
	assign mret_insn = mret_insn_i & instr_valid_i;
	assign dret_insn = dret_insn_i & instr_valid_i;
	assign wfi_insn = wfi_insn_i & instr_valid_i;
	assign ebrk_insn = ebrk_insn_i & instr_valid_i;
	assign csr_pipe_flush = csr_pipe_flush_i & instr_valid_i;
	assign instr_fetch_err = instr_fetch_err_i & instr_valid_i;
	assign illegal_insn_d = illegal_insn_i & (ctrl_fsm_cs != 4'd6);
	assign exc_req_d = (((ecall_insn | ebrk_insn) | illegal_insn_d) | instr_fetch_err) & (ctrl_fsm_cs != 4'd6);
	assign exc_req_lsu = store_err_i | load_err_i;
	assign id_exception_o = exc_req_d & ~wb_exception_o;
	assign special_req_flush_only = wfi_insn | csr_pipe_flush;
	assign special_req_pc_change = ((mret_insn | dret_insn) | exc_req_d) | exc_req_lsu;
	assign special_req = special_req_pc_change | special_req_flush_only;
	assign id_wb_pending = instr_valid_i | ~ready_wb_i;
	generate
		if (WritebackStage) begin : g_wb_exceptions
			always @(*) begin
				instr_fetch_err_prio = 0;
				illegal_insn_prio = 0;
				ecall_insn_prio = 0;
				ebrk_insn_prio = 0;
				store_err_prio = 0;
				load_err_prio = 0;
				if (store_err_q)
					store_err_prio = 1'b1;
				else if (load_err_q)
					load_err_prio = 1'b1;
				else if (instr_fetch_err)
					instr_fetch_err_prio = 1'b1;
				else if (illegal_insn_q)
					illegal_insn_prio = 1'b1;
				else if (ecall_insn)
					ecall_insn_prio = 1'b1;
				else if (ebrk_insn)
					ebrk_insn_prio = 1'b1;
			end
			assign wb_exception_o = ((load_err_q | store_err_q) | load_err_i) | store_err_i;
		end
		else begin : g_no_wb_exceptions
			always @(*) begin
				instr_fetch_err_prio = 0;
				illegal_insn_prio = 0;
				ecall_insn_prio = 0;
				ebrk_insn_prio = 0;
				store_err_prio = 0;
				load_err_prio = 0;
				if (instr_fetch_err)
					instr_fetch_err_prio = 1'b1;
				else if (illegal_insn_q)
					illegal_insn_prio = 1'b1;
				else if (ecall_insn)
					ecall_insn_prio = 1'b1;
				else if (ebrk_insn)
					ebrk_insn_prio = 1'b1;
				else if (store_err_q)
					store_err_prio = 1'b1;
				else if (load_err_q)
					load_err_prio = 1'b1;
			end
			assign wb_exception_o = 1'b0;
		end
		if (MemECC) begin : g_intg_irq_int
			reg mem_resp_intg_err_irq_pending_q;
			wire mem_resp_intg_err_irq_pending_d;
			reg [31:0] mem_resp_intg_err_addr_q;
			reg [31:0] mem_resp_intg_err_addr_d;
			reg mem_resp_intg_err_irq_set;
			reg mem_resp_intg_err_irq_clear;
			wire entering_nmi;
			assign entering_nmi = nmi_mode_d & ~nmi_mode_q;
			always @(*) begin
				mem_resp_intg_err_addr_d = mem_resp_intg_err_addr_q;
				mem_resp_intg_err_irq_set = 1'b0;
				mem_resp_intg_err_irq_clear = 1'b0;
				if (mem_resp_intg_err_irq_pending_q) begin
					if (entering_nmi & !irq_nm_ext_i)
						mem_resp_intg_err_irq_clear = 1'b1;
				end
				else if (mem_resp_intg_err_i) begin
					mem_resp_intg_err_addr_d = lsu_addr_last_i;
					mem_resp_intg_err_irq_set = 1'b1;
				end
			end
			assign mem_resp_intg_err_irq_pending_d = (mem_resp_intg_err_irq_pending_q & ~mem_resp_intg_err_irq_clear) | mem_resp_intg_err_irq_set;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni) begin
					mem_resp_intg_err_irq_pending_q <= 1'b0;
					mem_resp_intg_err_addr_q <= 1'sb0;
				end
				else begin
					mem_resp_intg_err_irq_pending_q <= mem_resp_intg_err_irq_pending_d;
					mem_resp_intg_err_addr_q <= mem_resp_intg_err_addr_d;
				end
			assign irq_nm_int = mem_resp_intg_err_irq_set | mem_resp_intg_err_irq_pending_q;
			assign irq_nm_int_cause = 5'b00000;
			assign irq_nm_int_mtval = mem_resp_intg_err_addr_q;
		end
		else begin : g_no_intg_irq_int
			wire unused_mem_resp_intg_err_i;
			assign unused_mem_resp_intg_err_i = mem_resp_intg_err_i;
			assign irq_nm_int = 1'b0;
			assign irq_nm_int_cause = 5'd0;
			assign irq_nm_int_mtval = 1'sb0;
		end
	endgenerate
	assign do_single_step_d = (instr_valid_i ? ~debug_mode_q & debug_single_step_i : do_single_step_q);
	assign enter_debug_mode_prio_d = (debug_req_i | do_single_step_d) & ~debug_mode_q;
	assign enter_debug_mode = enter_debug_mode_prio_d | (trigger_match_i & ~debug_mode_q);
	assign ebreak_into_debug = (priv_mode_i == 2'b11 ? debug_ebreakm_i : (priv_mode_i == 2'b00 ? debug_ebreaku_i : 1'b0));
	assign irq_nm = irq_nm_ext_i | irq_nm_int;
	assign irq_enabled = csr_mstatus_mie_i | (priv_mode_i == 2'b00);
	assign handle_irq = ((~debug_mode_q & ~debug_single_step_i) & ~nmi_mode_q) & (irq_nm | (irq_pending_i & irq_enabled));
	always @(*) begin : gen_mfip_id
		mfip_id = 4'd0;
		begin : sv2v_autoblock_1
			reg signed [31:0] i;
			for (i = 14; i >= 0; i = i - 1)
				if (irqs_i[0 + i])
					mfip_id = i[3:0];
		end
	end
	assign unused_irq_timer = irqs_i[16];
	assign debug_cause_d = (trigger_match_i ? 3'h2 : (ebrk_insn_prio & ebreak_into_debug ? 3'h1 : (debug_req_i ? 3'h3 : (do_single_step_d ? 3'h4 : 3'h0))));
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			debug_cause_q <= 3'h0;
		else
			debug_cause_q <= debug_cause_d;
	assign debug_cause_o = debug_cause_q;
	localparam [6:0] ibex_pkg_ExcCauseBreakpoint = 7'b0000011;
	localparam [6:0] ibex_pkg_ExcCauseEcallMMode = 7'b0001011;
	localparam [6:0] ibex_pkg_ExcCauseEcallUMode = 7'b0001000;
	localparam [6:0] ibex_pkg_ExcCauseIllegalInsn = 7'b0000010;
	localparam [6:0] ibex_pkg_ExcCauseInsnAddrMisa = 7'b0000000;
	localparam [6:0] ibex_pkg_ExcCauseInstrAccessFault = 7'b0000001;
	localparam [6:0] ibex_pkg_ExcCauseIrqExternalM = 7'b0101011;
	localparam [6:0] ibex_pkg_ExcCauseIrqNm = 7'b0111111;
	localparam [6:0] ibex_pkg_ExcCauseIrqSoftwareM = 7'b0100011;
	localparam [6:0] ibex_pkg_ExcCauseIrqTimerM = 7'b0100111;
	localparam [6:0] ibex_pkg_ExcCauseLoadAccessFault = 7'b0000101;
	localparam [6:0] ibex_pkg_ExcCauseStoreAccessFault = 7'b0000111;
	function automatic [4:0] sv2v_cast_5;
		input reg [4:0] inp;
		sv2v_cast_5 = inp;
	endfunction
	always @(*) begin
		instr_req_o = 1'b1;
		csr_save_if_o = 1'b0;
		csr_save_id_o = 1'b0;
		csr_save_wb_o = 1'b0;
		csr_restore_mret_id_o = 1'b0;
		csr_restore_dret_id_o = 1'b0;
		csr_save_cause_o = 1'b0;
		csr_mtval_o = 1'sb0;
		pc_mux_o = 3'd0;
		pc_set_o = 1'b0;
		nt_branch_mispredict_o = 1'b0;
		exc_pc_mux_o = 2'd1;
		exc_cause_o = ibex_pkg_ExcCauseInsnAddrMisa;
		ctrl_fsm_ns = ctrl_fsm_cs;
		ctrl_busy_o = 1'b1;
		halt_if = 1'b0;
		retain_id = 1'b0;
		flush_id = 1'b0;
		debug_csr_save_o = 1'b0;
		debug_mode_d = debug_mode_q;
		debug_mode_entering_o = 1'b0;
		nmi_mode_d = nmi_mode_q;
		perf_tbranch_o = 1'b0;
		perf_jump_o = 1'b0;
		controller_run_o = 1'b0;
		case (ctrl_fsm_cs)
			4'd0: begin
				instr_req_o = 1'b0;
				pc_mux_o = 3'd0;
				pc_set_o = 1'b1;
				ctrl_fsm_ns = 4'd1;
			end
			4'd1: begin
				instr_req_o = 1'b1;
				pc_mux_o = 3'd0;
				pc_set_o = 1'b1;
				ctrl_fsm_ns = 4'd4;
			end
			4'd2: begin
				ctrl_busy_o = 1'b0;
				instr_req_o = 1'b0;
				halt_if = 1'b1;
				flush_id = 1'b1;
				ctrl_fsm_ns = 4'd3;
			end
			4'd3: begin
				instr_req_o = 1'b0;
				halt_if = 1'b1;
				flush_id = 1'b1;
				if ((((irq_nm || irq_pending_i) || debug_req_i) || debug_mode_q) || debug_single_step_i)
					ctrl_fsm_ns = 4'd4;
				else
					ctrl_busy_o = 1'b0;
			end
			4'd4: begin
				if (id_in_ready_o)
					ctrl_fsm_ns = 4'd5;
				if (handle_irq) begin
					ctrl_fsm_ns = 4'd7;
					halt_if = 1'b1;
				end
				if (enter_debug_mode) begin
					ctrl_fsm_ns = 4'd8;
					halt_if = 1'b1;
				end
			end
			4'd5: begin
				controller_run_o = 1'b1;
				pc_mux_o = 3'd1;
				if (special_req) begin
					retain_id = 1'b1;
					if (ready_wb_i | wb_exception_o)
						ctrl_fsm_ns = 4'd6;
				end
				if (branch_set_i || jump_set_i) begin
					pc_set_o = (BranchPredictor ? ~instr_bp_taken_i : 1'b1);
					perf_tbranch_o = branch_set_i;
					perf_jump_o = jump_set_i;
				end
				if (BranchPredictor)
					if (instr_bp_taken_i & branch_not_set_i)
						nt_branch_mispredict_o = 1'b1;
				if ((enter_debug_mode || handle_irq) && (stall || id_wb_pending))
					halt_if = 1'b1;
				if ((!stall && !special_req) && !id_wb_pending)
					if (enter_debug_mode) begin
						ctrl_fsm_ns = 4'd8;
						halt_if = 1'b1;
					end
					else if (handle_irq) begin
						ctrl_fsm_ns = 4'd7;
						halt_if = 1'b1;
					end
			end
			4'd7: begin
				pc_mux_o = 3'd2;
				exc_pc_mux_o = 2'd1;
				if (handle_irq) begin
					pc_set_o = 1'b1;
					csr_save_if_o = 1'b1;
					csr_save_cause_o = 1'b1;
					if (irq_nm && !nmi_mode_q) begin
						exc_cause_o = (irq_nm_ext_i ? ibex_pkg_ExcCauseIrqNm : {2'b10, irq_nm_int_cause});
						if (irq_nm_int & !irq_nm_ext_i)
							csr_mtval_o = irq_nm_int_mtval;
						nmi_mode_d = 1'b1;
					end
					else if (irqs_i[14-:15] != 15'b000000000000000)
						exc_cause_o = {2'b01, sv2v_cast_5({1'b1, mfip_id})};
					else if (irqs_i[15])
						exc_cause_o = ibex_pkg_ExcCauseIrqExternalM;
					else if (irqs_i[17])
						exc_cause_o = ibex_pkg_ExcCauseIrqSoftwareM;
					else
						exc_cause_o = ibex_pkg_ExcCauseIrqTimerM;
				end
				ctrl_fsm_ns = 4'd5;
			end
			4'd8: begin
				pc_mux_o = 3'd2;
				exc_pc_mux_o = 2'd2;
				flush_id = 1'b1;
				pc_set_o = 1'b1;
				csr_save_if_o = 1'b1;
				debug_csr_save_o = 1'b1;
				csr_save_cause_o = 1'b1;
				debug_mode_d = 1'b1;
				debug_mode_entering_o = 1'b1;
				ctrl_fsm_ns = 4'd5;
			end
			4'd9: begin
				flush_id = 1'b1;
				pc_mux_o = 3'd2;
				pc_set_o = 1'b1;
				exc_pc_mux_o = 2'd2;
				if (ebreak_into_debug && !debug_mode_q) begin
					csr_save_cause_o = 1'b1;
					csr_save_id_o = 1'b1;
					debug_csr_save_o = 1'b1;
				end
				debug_mode_d = 1'b1;
				debug_mode_entering_o = 1'b1;
				ctrl_fsm_ns = 4'd5;
			end
			4'd6: begin
				halt_if = 1'b1;
				flush_id = 1'b1;
				ctrl_fsm_ns = 4'd5;
				if ((exc_req_q || store_err_q) || load_err_q) begin
					pc_set_o = 1'b1;
					pc_mux_o = 3'd2;
					exc_pc_mux_o = (debug_mode_q ? 2'd3 : 2'd0);
					if (WritebackStage) begin : g_writeback_mepc_save
						csr_save_id_o = ~(store_err_q | load_err_q);
						csr_save_wb_o = store_err_q | load_err_q;
					end
					else begin : g_no_writeback_mepc_save
						csr_save_id_o = 1'b0;
					end
					csr_save_cause_o = 1'b1;
					case (1'b1)
						instr_fetch_err_prio: begin
							exc_cause_o = ibex_pkg_ExcCauseInstrAccessFault;
							csr_mtval_o = (instr_fetch_err_plus2_i ? pc_id_i + 32'd2 : pc_id_i);
						end
						illegal_insn_prio: begin
							exc_cause_o = ibex_pkg_ExcCauseIllegalInsn;
							csr_mtval_o = (instr_is_compressed_i ? {16'b0000000000000000, instr_compressed_i} : instr_i);
						end
						ecall_insn_prio: exc_cause_o = (priv_mode_i == 2'b11 ? ibex_pkg_ExcCauseEcallMMode : ibex_pkg_ExcCauseEcallUMode);
						ebrk_insn_prio:
							if (debug_mode_q | ebreak_into_debug) begin
								pc_set_o = 1'b0;
								csr_save_id_o = 1'b0;
								csr_save_cause_o = 1'b0;
								ctrl_fsm_ns = 4'd9;
								flush_id = 1'b0;
							end
							else
								exc_cause_o = ibex_pkg_ExcCauseBreakpoint;
						store_err_prio: begin
							exc_cause_o = ibex_pkg_ExcCauseStoreAccessFault;
							csr_mtval_o = lsu_addr_last_i;
						end
						load_err_prio: begin
							exc_cause_o = ibex_pkg_ExcCauseLoadAccessFault;
							csr_mtval_o = lsu_addr_last_i;
						end
						default:
							;
					endcase
				end
				else if (mret_insn) begin
					pc_mux_o = 3'd3;
					pc_set_o = 1'b1;
					csr_restore_mret_id_o = 1'b1;
					if (nmi_mode_q)
						nmi_mode_d = 1'b0;
				end
				else if (dret_insn) begin
					pc_mux_o = 3'd4;
					pc_set_o = 1'b1;
					debug_mode_d = 1'b0;
					csr_restore_dret_id_o = 1'b1;
				end
				else if (wfi_insn)
					ctrl_fsm_ns = 4'd2;
				if (enter_debug_mode_prio_q && !(ebrk_insn_prio && ebreak_into_debug))
					ctrl_fsm_ns = 4'd8;
			end
			default: begin
				instr_req_o = 1'b0;
				ctrl_fsm_ns = 4'd0;
			end
		endcase
		if (~instr_exec_i)
			halt_if = 1'b1;
	end
	assign flush_id_o = flush_id;
	assign debug_mode_o = debug_mode_q;
	assign nmi_mode_o = nmi_mode_q;
	assign stall = stall_id_i | stall_wb_i;
	assign id_in_ready_o = (~stall & ~halt_if) & ~retain_id;
	assign instr_valid_clear_o = ~(stall | retain_id) | flush_id;
	always @(posedge clk_i or negedge rst_ni) begin : update_regs
		if (!rst_ni) begin
			ctrl_fsm_cs <= 4'd0;
			nmi_mode_q <= 1'b0;
			do_single_step_q <= 1'b0;
			debug_mode_q <= 1'b0;
			enter_debug_mode_prio_q <= 1'b0;
			load_err_q <= 1'b0;
			store_err_q <= 1'b0;
			exc_req_q <= 1'b0;
			illegal_insn_q <= 1'b0;
		end
		else begin
			ctrl_fsm_cs <= ctrl_fsm_ns;
			nmi_mode_q <= nmi_mode_d;
			do_single_step_q <= do_single_step_d;
			debug_mode_q <= debug_mode_d;
			enter_debug_mode_prio_q <= enter_debug_mode_prio_d;
			load_err_q <= load_err_d;
			store_err_q <= store_err_d;
			exc_req_q <= exc_req_d;
			illegal_insn_q <= illegal_insn_d;
		end
	end
endmodule
module ibex_core (
	clk_i,
	rst_ni,
	hart_id_i,
	boot_addr_i,
	instr_req_o,
	instr_gnt_i,
	instr_rvalid_i,
	instr_addr_o,
	instr_rdata_i,
	instr_err_i,
	data_req_o,
	data_gnt_i,
	data_rvalid_i,
	data_we_o,
	data_be_o,
	data_addr_o,
	data_wdata_o,
	data_rdata_i,
	data_err_i,
	dummy_instr_id_o,
	dummy_instr_wb_o,
	rf_raddr_a_o,
	rf_raddr_b_o,
	rf_waddr_wb_o,
	rf_we_wb_o,
	rf_wdata_wb_ecc_o,
	rf_rdata_a_ecc_i,
	rf_rdata_b_ecc_i,
	ic_tag_req_o,
	ic_tag_write_o,
	ic_tag_addr_o,
	ic_tag_wdata_o,
	ic_tag_rdata_i,
	ic_data_req_o,
	ic_data_write_o,
	ic_data_addr_o,
	ic_data_wdata_o,
	ic_data_rdata_i,
	ic_scr_key_valid_i,
	ic_scr_key_req_o,
	irq_software_i,
	irq_timer_i,
	irq_external_i,
	irq_fast_i,
	irq_nm_i,
	irq_pending_o,
	debug_req_i,
	crash_dump_o,
	double_fault_seen_o,
	fetch_enable_i,
	alert_minor_o,
	alert_major_internal_o,
	alert_major_bus_o,
	core_busy_o
);
	parameter [0:0] PMPEnable = 1'b0;
	parameter [31:0] PMPGranularity = 0;
	parameter [31:0] PMPNumRegions = 4;
	parameter [31:0] MHPMCounterNum = 0;
	parameter [31:0] MHPMCounterWidth = 40;
	parameter [0:0] RV32E = 1'b0;
	parameter integer RV32M = 32'sd1;
	parameter integer RV32B = 32'sd0;
	parameter [0:0] BranchTargetALU = 1'b0;
	parameter [0:0] WritebackStage = 1'b0;
	parameter [0:0] ICache = 1'b0;
	parameter [0:0] ICacheECC = 1'b0;
	localparam [31:0] ibex_pkg_BUS_SIZE = 32;
	parameter [31:0] BusSizeECC = ibex_pkg_BUS_SIZE;
	localparam [31:0] ibex_pkg_ADDR_W = 32;
	localparam [31:0] ibex_pkg_IC_LINE_SIZE = 64;
	localparam [31:0] ibex_pkg_IC_LINE_BYTES = 8;
	localparam [31:0] ibex_pkg_IC_NUM_WAYS = 2;
	localparam [31:0] ibex_pkg_IC_SIZE_BYTES = 4096;
	localparam [31:0] ibex_pkg_IC_NUM_LINES = (ibex_pkg_IC_SIZE_BYTES / ibex_pkg_IC_NUM_WAYS) / ibex_pkg_IC_LINE_BYTES;
	localparam [31:0] ibex_pkg_IC_INDEX_W = $clog2(ibex_pkg_IC_NUM_LINES);
	localparam [31:0] ibex_pkg_IC_LINE_W = 3;
	localparam [31:0] ibex_pkg_IC_TAG_SIZE = ((ibex_pkg_ADDR_W - ibex_pkg_IC_INDEX_W) - ibex_pkg_IC_LINE_W) + 1;
	parameter [31:0] TagSizeECC = ibex_pkg_IC_TAG_SIZE;
	parameter [31:0] LineSizeECC = ibex_pkg_IC_LINE_SIZE;
	parameter [0:0] BranchPredictor = 1'b0;
	parameter [0:0] DbgTriggerEn = 1'b0;
	parameter [31:0] DbgHwBreakNum = 1;
	parameter [0:0] ResetAll = 1'b0;
	localparam signed [31:0] ibex_pkg_LfsrWidth = 32;
	localparam [31:0] ibex_pkg_RndCnstLfsrSeedDefault = 32'hac533bf4;
	parameter [31:0] RndCnstLfsrSeed = ibex_pkg_RndCnstLfsrSeedDefault;
	localparam [159:0] ibex_pkg_RndCnstLfsrPermDefault = 160'h1e35ecba467fd1b12e958152c04fa43878a8daed;
	parameter [159:0] RndCnstLfsrPerm = ibex_pkg_RndCnstLfsrPermDefault;
	parameter [0:0] SecureIbex = 1'b0;
	parameter [0:0] DummyInstructions = 1'b0;
	parameter [0:0] RegFileECC = 1'b0;
	parameter [31:0] RegFileDataWidth = 32;
	parameter [0:0] MemECC = 1'b0;
	parameter [31:0] MemDataWidth = (MemECC ? 39 : 32);
	parameter [31:0] DmHaltAddr = 32'h1a110800;
	parameter [31:0] DmExceptionAddr = 32'h1a110808;
	input wire clk_i;
	input wire rst_ni;
	input wire [31:0] hart_id_i;
	input wire [31:0] boot_addr_i;
	output wire instr_req_o;
	input wire instr_gnt_i;
	input wire instr_rvalid_i;
	output wire [31:0] instr_addr_o;
	input wire [MemDataWidth - 1:0] instr_rdata_i;
	input wire instr_err_i;
	output wire data_req_o;
	input wire data_gnt_i;
	input wire data_rvalid_i;
	output wire data_we_o;
	output wire [3:0] data_be_o;
	output wire [31:0] data_addr_o;
	output wire [MemDataWidth - 1:0] data_wdata_o;
	input wire [MemDataWidth - 1:0] data_rdata_i;
	input wire data_err_i;
	output wire dummy_instr_id_o;
	output wire dummy_instr_wb_o;
	output wire [4:0] rf_raddr_a_o;
	output wire [4:0] rf_raddr_b_o;
	output wire [4:0] rf_waddr_wb_o;
	output wire rf_we_wb_o;
	output wire [RegFileDataWidth - 1:0] rf_wdata_wb_ecc_o;
	input wire [RegFileDataWidth - 1:0] rf_rdata_a_ecc_i;
	input wire [RegFileDataWidth - 1:0] rf_rdata_b_ecc_i;
	output wire [1:0] ic_tag_req_o;
	output wire ic_tag_write_o;
	output wire [ibex_pkg_IC_INDEX_W - 1:0] ic_tag_addr_o;
	output wire [TagSizeECC - 1:0] ic_tag_wdata_o;
	input wire [(ibex_pkg_IC_NUM_WAYS * TagSizeECC) - 1:0] ic_tag_rdata_i;
	output wire [1:0] ic_data_req_o;
	output wire ic_data_write_o;
	output wire [ibex_pkg_IC_INDEX_W - 1:0] ic_data_addr_o;
	output wire [LineSizeECC - 1:0] ic_data_wdata_o;
	input wire [(ibex_pkg_IC_NUM_WAYS * LineSizeECC) - 1:0] ic_data_rdata_i;
	input wire ic_scr_key_valid_i;
	output wire ic_scr_key_req_o;
	input wire irq_software_i;
	input wire irq_timer_i;
	input wire irq_external_i;
	input wire [14:0] irq_fast_i;
	input wire irq_nm_i;
	output wire irq_pending_o;
	input wire debug_req_i;
	output wire [159:0] crash_dump_o;
	output wire double_fault_seen_o;
	input wire [3:0] fetch_enable_i;
	output wire alert_minor_o;
	output wire alert_major_internal_o;
	output wire alert_major_bus_o;
	output wire [3:0] core_busy_o;
	localparam [31:0] PMPNumChan = 3;
	localparam [0:0] DataIndTiming = SecureIbex;
	localparam [0:0] PCIncrCheck = SecureIbex;
	localparam [0:0] ShadowCSR = 1'b0;
	wire dummy_instr_id;
	wire instr_valid_id;
	wire instr_new_id;
	wire [31:0] instr_rdata_id;
	wire [31:0] instr_rdata_alu_id;
	wire [15:0] instr_rdata_c_id;
	wire instr_is_compressed_id;
	wire instr_perf_count_id;
	wire instr_bp_taken_id;
	wire instr_fetch_err;
	wire instr_fetch_err_plus2;
	wire illegal_c_insn_id;
	wire [31:0] pc_if;
	wire [31:0] pc_id;
	wire [31:0] pc_wb;
	wire [67:0] imd_val_d_ex;
	wire [67:0] imd_val_q_ex;
	wire [1:0] imd_val_we_ex;
	wire data_ind_timing;
	wire dummy_instr_en;
	wire [2:0] dummy_instr_mask;
	wire dummy_instr_seed_en;
	wire [31:0] dummy_instr_seed;
	wire icache_enable;
	wire icache_inval;
	wire icache_ecc_error;
	wire pc_mismatch_alert;
	wire csr_shadow_err;
	wire instr_first_cycle_id;
	wire instr_valid_clear;
	wire pc_set;
	wire nt_branch_mispredict;
	wire [31:0] nt_branch_addr;
	wire [2:0] pc_mux_id;
	wire [1:0] exc_pc_mux_id;
	wire [6:0] exc_cause;
	wire instr_intg_err;
	wire lsu_load_err;
	wire lsu_store_err;
	wire lsu_load_resp_intg_err;
	wire lsu_store_resp_intg_err;
	wire lsu_addr_incr_req;
	wire [31:0] lsu_addr_last;
	wire [31:0] branch_target_ex;
	wire branch_decision;
	wire ctrl_busy;
	wire if_busy;
	wire lsu_busy;
	wire [4:0] rf_raddr_a;
	wire [31:0] rf_rdata_a;
	wire [4:0] rf_raddr_b;
	wire [31:0] rf_rdata_b;
	wire rf_ren_a;
	wire rf_ren_b;
	wire [4:0] rf_waddr_wb;
	wire [31:0] rf_wdata_wb;
	wire [31:0] rf_wdata_fwd_wb;
	wire [31:0] rf_wdata_lsu;
	wire rf_we_wb;
	wire rf_we_lsu;
	wire rf_ecc_err_comb;
	wire [4:0] rf_waddr_id;
	wire [31:0] rf_wdata_id;
	wire rf_we_id;
	wire rf_rd_a_wb_match;
	wire rf_rd_b_wb_match;
	wire [6:0] alu_operator_ex;
	wire [31:0] alu_operand_a_ex;
	wire [31:0] alu_operand_b_ex;
	wire [31:0] bt_a_operand;
	wire [31:0] bt_b_operand;
	wire [31:0] alu_adder_result_ex;
	wire [31:0] result_ex;
	wire mult_en_ex;
	wire div_en_ex;
	wire mult_sel_ex;
	wire div_sel_ex;
	wire [1:0] multdiv_operator_ex;
	wire [1:0] multdiv_signed_mode_ex;
	wire [31:0] multdiv_operand_a_ex;
	wire [31:0] multdiv_operand_b_ex;
	wire multdiv_ready_id;
	wire csr_access;
	wire [1:0] csr_op;
	wire csr_op_en;
	wire [11:0] csr_addr;
	wire [31:0] csr_rdata;
	wire [31:0] csr_wdata;
	wire illegal_csr_insn_id;
	wire lsu_we;
	wire [1:0] lsu_type;
	wire lsu_sign_ext;
	wire lsu_req;
	wire [31:0] lsu_wdata;
	wire lsu_req_done;
	wire id_in_ready;
	wire ex_valid;
	wire lsu_resp_valid;
	wire lsu_resp_err;
	wire instr_req_int;
	wire instr_req_gated;
	wire instr_exec;
	wire en_wb;
	wire [1:0] instr_type_wb;
	wire ready_wb;
	wire rf_write_wb;
	wire outstanding_load_wb;
	wire outstanding_store_wb;
	wire dummy_instr_wb;
	wire nmi_mode;
	wire [17:0] irqs;
	wire csr_mstatus_mie;
	wire [31:0] csr_mepc;
	wire [31:0] csr_depc;
	wire [(PMPNumRegions * 34) - 1:0] csr_pmp_addr;
	wire [(PMPNumRegions * 6) - 1:0] csr_pmp_cfg;
	wire [2:0] csr_pmp_mseccfg;
	wire [0:2] pmp_req_err;
	wire data_req_out;
	wire csr_save_if;
	wire csr_save_id;
	wire csr_save_wb;
	wire csr_restore_mret_id;
	wire csr_restore_dret_id;
	wire csr_save_cause;
	wire csr_mtvec_init;
	wire [31:0] csr_mtvec;
	wire [31:0] csr_mtval;
	wire csr_mstatus_tw;
	wire [1:0] priv_mode_id;
	wire [1:0] priv_mode_lsu;
	wire debug_mode;
	wire debug_mode_entering;
	wire [2:0] debug_cause;
	wire debug_csr_save;
	wire debug_single_step;
	wire debug_ebreakm;
	wire debug_ebreaku;
	wire trigger_match;
	wire instr_id_done;
	wire instr_done_wb;
	wire perf_instr_ret_wb;
	wire perf_instr_ret_compressed_wb;
	wire perf_instr_ret_wb_spec;
	wire perf_instr_ret_compressed_wb_spec;
	wire perf_iside_wait;
	wire perf_dside_wait;
	wire perf_mul_wait;
	wire perf_div_wait;
	wire perf_jump;
	wire perf_branch;
	wire perf_tbranch;
	wire perf_load;
	wire perf_store;
	wire illegal_insn_id;
	wire unused_illegal_insn_id;
	localparam [3:0] ibex_pkg_IbexMuBiOff = 4'b1010;
	localparam [3:0] ibex_pkg_IbexMuBiOn = 4'b0101;
	generate
		if (SecureIbex) begin : g_core_busy_secure
			localparam [31:0] NumBusySignals = 3;
			localparam [31:0] NumBusyBits = 12;
			wire [11:0] busy_bits_buf;
			prim_buf #(.Width(NumBusyBits)) u_fetch_enable_buf(
				.in_i({4 {ctrl_busy, if_busy, lsu_busy}}),
				.out_o(busy_bits_buf)
			);
			genvar i;
			for (i = 0; i < 4; i = i + 1) begin : g_core_busy_bits
				if (ibex_pkg_IbexMuBiOn[i] == 1'b1) begin : g_pos
					assign core_busy_o[i] = |busy_bits_buf[i * NumBusySignals+:NumBusySignals];
				end
				else begin : g_neg
					assign core_busy_o[i] = ~|busy_bits_buf[i * NumBusySignals+:NumBusySignals];
				end
			end
		end
		else begin : g_core_busy_non_secure
			assign core_busy_o = ((ctrl_busy || if_busy) || lsu_busy ? ibex_pkg_IbexMuBiOn : ibex_pkg_IbexMuBiOff);
		end
	endgenerate
	localparam [31:0] ibex_pkg_PMP_I = 0;
	localparam [31:0] ibex_pkg_PMP_I2 = 1;
	ibex_if_stage #(
		.DmHaltAddr(DmHaltAddr),
		.DmExceptionAddr(DmExceptionAddr),
		.DummyInstructions(DummyInstructions),
		.ICache(ICache),
		.ICacheECC(ICacheECC),
		.BusSizeECC(BusSizeECC),
		.TagSizeECC(TagSizeECC),
		.LineSizeECC(LineSizeECC),
		.PCIncrCheck(PCIncrCheck),
		.ResetAll(ResetAll),
		.RndCnstLfsrSeed(RndCnstLfsrSeed),
		.RndCnstLfsrPerm(RndCnstLfsrPerm),
		.BranchPredictor(BranchPredictor),
		.MemECC(MemECC),
		.MemDataWidth(MemDataWidth)
	) if_stage_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.boot_addr_i(boot_addr_i),
		.req_i(instr_req_gated),
		.instr_req_o(instr_req_o),
		.instr_addr_o(instr_addr_o),
		.instr_gnt_i(instr_gnt_i),
		.instr_rvalid_i(instr_rvalid_i),
		.instr_rdata_i(instr_rdata_i),
		.instr_bus_err_i(instr_err_i),
		.instr_intg_err_o(instr_intg_err),
		.ic_tag_req_o(ic_tag_req_o),
		.ic_tag_write_o(ic_tag_write_o),
		.ic_tag_addr_o(ic_tag_addr_o),
		.ic_tag_wdata_o(ic_tag_wdata_o),
		.ic_tag_rdata_i(ic_tag_rdata_i),
		.ic_data_req_o(ic_data_req_o),
		.ic_data_write_o(ic_data_write_o),
		.ic_data_addr_o(ic_data_addr_o),
		.ic_data_wdata_o(ic_data_wdata_o),
		.ic_data_rdata_i(ic_data_rdata_i),
		.ic_scr_key_valid_i(ic_scr_key_valid_i),
		.ic_scr_key_req_o(ic_scr_key_req_o),
		.instr_valid_id_o(instr_valid_id),
		.instr_new_id_o(instr_new_id),
		.instr_rdata_id_o(instr_rdata_id),
		.instr_rdata_alu_id_o(instr_rdata_alu_id),
		.instr_rdata_c_id_o(instr_rdata_c_id),
		.instr_is_compressed_id_o(instr_is_compressed_id),
		.instr_bp_taken_o(instr_bp_taken_id),
		.instr_fetch_err_o(instr_fetch_err),
		.instr_fetch_err_plus2_o(instr_fetch_err_plus2),
		.illegal_c_insn_id_o(illegal_c_insn_id),
		.dummy_instr_id_o(dummy_instr_id),
		.pc_if_o(pc_if),
		.pc_id_o(pc_id),
		.pmp_err_if_i(pmp_req_err[ibex_pkg_PMP_I]),
		.pmp_err_if_plus2_i(pmp_req_err[ibex_pkg_PMP_I2]),
		.instr_valid_clear_i(instr_valid_clear),
		.pc_set_i(pc_set),
		.pc_mux_i(pc_mux_id),
		.nt_branch_mispredict_i(nt_branch_mispredict),
		.exc_pc_mux_i(exc_pc_mux_id),
		.exc_cause(exc_cause),
		.dummy_instr_en_i(dummy_instr_en),
		.dummy_instr_mask_i(dummy_instr_mask),
		.dummy_instr_seed_en_i(dummy_instr_seed_en),
		.dummy_instr_seed_i(dummy_instr_seed),
		.icache_enable_i(icache_enable),
		.icache_inval_i(icache_inval),
		.icache_ecc_error_o(icache_ecc_error),
		.branch_target_ex_i(branch_target_ex),
		.nt_branch_addr_i(nt_branch_addr),
		.csr_mepc_i(csr_mepc),
		.csr_depc_i(csr_depc),
		.csr_mtvec_i(csr_mtvec),
		.csr_mtvec_init_o(csr_mtvec_init),
		.id_in_ready_i(id_in_ready),
		.pc_mismatch_alert_o(pc_mismatch_alert),
		.if_busy_o(if_busy)
	);
	assign perf_iside_wait = id_in_ready & ~instr_valid_id;
	generate
		if (SecureIbex) begin : g_instr_req_gated_secure
			assign instr_req_gated = instr_req_int & (fetch_enable_i == ibex_pkg_IbexMuBiOn);
			assign instr_exec = fetch_enable_i == ibex_pkg_IbexMuBiOn;
		end
		else begin : g_instr_req_gated_non_secure
			wire unused_fetch_enable;
			assign unused_fetch_enable = ^fetch_enable_i[3:1];
			assign instr_req_gated = instr_req_int & fetch_enable_i[0];
			assign instr_exec = fetch_enable_i[0];
		end
	endgenerate
	ibex_id_stage #(
		.RV32E(RV32E),
		.RV32M(RV32M),
		.RV32B(RV32B),
		.BranchTargetALU(BranchTargetALU),
		.DataIndTiming(DataIndTiming),
		.WritebackStage(WritebackStage),
		.BranchPredictor(BranchPredictor),
		.MemECC(MemECC)
	) id_stage_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.ctrl_busy_o(ctrl_busy),
		.illegal_insn_o(illegal_insn_id),
		.instr_valid_i(instr_valid_id),
		.instr_rdata_i(instr_rdata_id),
		.instr_rdata_alu_i(instr_rdata_alu_id),
		.instr_rdata_c_i(instr_rdata_c_id),
		.instr_is_compressed_i(instr_is_compressed_id),
		.instr_bp_taken_i(instr_bp_taken_id),
		.branch_decision_i(branch_decision),
		.instr_first_cycle_id_o(instr_first_cycle_id),
		.instr_valid_clear_o(instr_valid_clear),
		.id_in_ready_o(id_in_ready),
		.instr_exec_i(instr_exec),
		.instr_req_o(instr_req_int),
		.pc_set_o(pc_set),
		.pc_mux_o(pc_mux_id),
		.nt_branch_mispredict_o(nt_branch_mispredict),
		.nt_branch_addr_o(nt_branch_addr),
		.exc_pc_mux_o(exc_pc_mux_id),
		.exc_cause_o(exc_cause),
		.icache_inval_o(icache_inval),
		.instr_fetch_err_i(instr_fetch_err),
		.instr_fetch_err_plus2_i(instr_fetch_err_plus2),
		.illegal_c_insn_i(illegal_c_insn_id),
		.pc_id_i(pc_id),
		.ex_valid_i(ex_valid),
		.lsu_resp_valid_i(lsu_resp_valid),
		.alu_operator_ex_o(alu_operator_ex),
		.alu_operand_a_ex_o(alu_operand_a_ex),
		.alu_operand_b_ex_o(alu_operand_b_ex),
		.imd_val_q_ex_o(imd_val_q_ex),
		.imd_val_d_ex_i(imd_val_d_ex),
		.imd_val_we_ex_i(imd_val_we_ex),
		.bt_a_operand_o(bt_a_operand),
		.bt_b_operand_o(bt_b_operand),
		.mult_en_ex_o(mult_en_ex),
		.div_en_ex_o(div_en_ex),
		.mult_sel_ex_o(mult_sel_ex),
		.div_sel_ex_o(div_sel_ex),
		.multdiv_operator_ex_o(multdiv_operator_ex),
		.multdiv_signed_mode_ex_o(multdiv_signed_mode_ex),
		.multdiv_operand_a_ex_o(multdiv_operand_a_ex),
		.multdiv_operand_b_ex_o(multdiv_operand_b_ex),
		.multdiv_ready_id_o(multdiv_ready_id),
		.csr_access_o(csr_access),
		.csr_op_o(csr_op),
		.csr_op_en_o(csr_op_en),
		.csr_save_if_o(csr_save_if),
		.csr_save_id_o(csr_save_id),
		.csr_save_wb_o(csr_save_wb),
		.csr_restore_mret_id_o(csr_restore_mret_id),
		.csr_restore_dret_id_o(csr_restore_dret_id),
		.csr_save_cause_o(csr_save_cause),
		.csr_mtval_o(csr_mtval),
		.priv_mode_i(priv_mode_id),
		.csr_mstatus_tw_i(csr_mstatus_tw),
		.illegal_csr_insn_i(illegal_csr_insn_id),
		.data_ind_timing_i(data_ind_timing),
		.lsu_req_o(lsu_req),
		.lsu_we_o(lsu_we),
		.lsu_type_o(lsu_type),
		.lsu_sign_ext_o(lsu_sign_ext),
		.lsu_wdata_o(lsu_wdata),
		.lsu_req_done_i(lsu_req_done),
		.lsu_addr_incr_req_i(lsu_addr_incr_req),
		.lsu_addr_last_i(lsu_addr_last),
		.lsu_load_err_i(lsu_load_err),
		.lsu_load_resp_intg_err_i(lsu_load_resp_intg_err),
		.lsu_store_err_i(lsu_store_err),
		.lsu_store_resp_intg_err_i(lsu_store_resp_intg_err),
		.csr_mstatus_mie_i(csr_mstatus_mie),
		.irq_pending_i(irq_pending_o),
		.irqs_i(irqs),
		.irq_nm_i(irq_nm_i),
		.nmi_mode_o(nmi_mode),
		.debug_mode_o(debug_mode),
		.debug_mode_entering_o(debug_mode_entering),
		.debug_cause_o(debug_cause),
		.debug_csr_save_o(debug_csr_save),
		.debug_req_i(debug_req_i),
		.debug_single_step_i(debug_single_step),
		.debug_ebreakm_i(debug_ebreakm),
		.debug_ebreaku_i(debug_ebreaku),
		.trigger_match_i(trigger_match),
		.result_ex_i(result_ex),
		.csr_rdata_i(csr_rdata),
		.rf_raddr_a_o(rf_raddr_a),
		.rf_rdata_a_i(rf_rdata_a),
		.rf_raddr_b_o(rf_raddr_b),
		.rf_rdata_b_i(rf_rdata_b),
		.rf_ren_a_o(rf_ren_a),
		.rf_ren_b_o(rf_ren_b),
		.rf_waddr_id_o(rf_waddr_id),
		.rf_wdata_id_o(rf_wdata_id),
		.rf_we_id_o(rf_we_id),
		.rf_rd_a_wb_match_o(rf_rd_a_wb_match),
		.rf_rd_b_wb_match_o(rf_rd_b_wb_match),
		.rf_waddr_wb_i(rf_waddr_wb),
		.rf_wdata_fwd_wb_i(rf_wdata_fwd_wb),
		.rf_write_wb_i(rf_write_wb),
		.en_wb_o(en_wb),
		.instr_type_wb_o(instr_type_wb),
		.instr_perf_count_id_o(instr_perf_count_id),
		.ready_wb_i(ready_wb),
		.outstanding_load_wb_i(outstanding_load_wb),
		.outstanding_store_wb_i(outstanding_store_wb),
		.perf_jump_o(perf_jump),
		.perf_branch_o(perf_branch),
		.perf_tbranch_o(perf_tbranch),
		.perf_dside_wait_o(perf_dside_wait),
		.perf_mul_wait_o(perf_mul_wait),
		.perf_div_wait_o(perf_div_wait),
		.instr_id_done_o(instr_id_done)
	);
	assign unused_illegal_insn_id = illegal_insn_id;
	ibex_ex_block #(
		.RV32M(RV32M),
		.RV32B(RV32B),
		.BranchTargetALU(BranchTargetALU)
	) ex_block_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.alu_operator_i(alu_operator_ex),
		.alu_operand_a_i(alu_operand_a_ex),
		.alu_operand_b_i(alu_operand_b_ex),
		.alu_instr_first_cycle_i(instr_first_cycle_id),
		.bt_a_operand_i(bt_a_operand),
		.bt_b_operand_i(bt_b_operand),
		.multdiv_operator_i(multdiv_operator_ex),
		.mult_en_i(mult_en_ex),
		.div_en_i(div_en_ex),
		.mult_sel_i(mult_sel_ex),
		.div_sel_i(div_sel_ex),
		.multdiv_signed_mode_i(multdiv_signed_mode_ex),
		.multdiv_operand_a_i(multdiv_operand_a_ex),
		.multdiv_operand_b_i(multdiv_operand_b_ex),
		.multdiv_ready_id_i(multdiv_ready_id),
		.data_ind_timing_i(data_ind_timing),
		.imd_val_we_o(imd_val_we_ex),
		.imd_val_d_o(imd_val_d_ex),
		.imd_val_q_i(imd_val_q_ex),
		.alu_adder_result_ex_o(alu_adder_result_ex),
		.result_ex_o(result_ex),
		.branch_target_o(branch_target_ex),
		.branch_decision_o(branch_decision),
		.ex_valid_o(ex_valid)
	);
	localparam [31:0] ibex_pkg_PMP_D = 2;
	assign data_req_o = data_req_out & ~pmp_req_err[ibex_pkg_PMP_D];
	assign lsu_resp_err = lsu_load_err | lsu_store_err;
	ibex_load_store_unit #(
		.MemECC(MemECC),
		.MemDataWidth(MemDataWidth)
	) load_store_unit_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.data_req_o(data_req_out),
		.data_gnt_i(data_gnt_i),
		.data_rvalid_i(data_rvalid_i),
		.data_bus_err_i(data_err_i),
		.data_pmp_err_i(pmp_req_err[ibex_pkg_PMP_D]),
		.data_addr_o(data_addr_o),
		.data_we_o(data_we_o),
		.data_be_o(data_be_o),
		.data_wdata_o(data_wdata_o),
		.data_rdata_i(data_rdata_i),
		.lsu_we_i(lsu_we),
		.lsu_type_i(lsu_type),
		.lsu_wdata_i(lsu_wdata),
		.lsu_sign_ext_i(lsu_sign_ext),
		.lsu_rdata_o(rf_wdata_lsu),
		.lsu_rdata_valid_o(rf_we_lsu),
		.lsu_req_i(lsu_req),
		.lsu_req_done_o(lsu_req_done),
		.adder_result_ex_i(alu_adder_result_ex),
		.addr_incr_req_o(lsu_addr_incr_req),
		.addr_last_o(lsu_addr_last),
		.lsu_resp_valid_o(lsu_resp_valid),
		.load_err_o(lsu_load_err),
		.load_resp_intg_err_o(lsu_load_resp_intg_err),
		.store_err_o(lsu_store_err),
		.store_resp_intg_err_o(lsu_store_resp_intg_err),
		.busy_o(lsu_busy),
		.perf_load_o(perf_load),
		.perf_store_o(perf_store)
	);
	ibex_wb_stage #(
		.ResetAll(ResetAll),
		.WritebackStage(WritebackStage),
		.DummyInstructions(DummyInstructions)
	) wb_stage_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.en_wb_i(en_wb),
		.instr_type_wb_i(instr_type_wb),
		.pc_id_i(pc_id),
		.instr_is_compressed_id_i(instr_is_compressed_id),
		.instr_perf_count_id_i(instr_perf_count_id),
		.ready_wb_o(ready_wb),
		.rf_write_wb_o(rf_write_wb),
		.outstanding_load_wb_o(outstanding_load_wb),
		.outstanding_store_wb_o(outstanding_store_wb),
		.pc_wb_o(pc_wb),
		.perf_instr_ret_wb_o(perf_instr_ret_wb),
		.perf_instr_ret_compressed_wb_o(perf_instr_ret_compressed_wb),
		.perf_instr_ret_wb_spec_o(perf_instr_ret_wb_spec),
		.perf_instr_ret_compressed_wb_spec_o(perf_instr_ret_compressed_wb_spec),
		.rf_waddr_id_i(rf_waddr_id),
		.rf_wdata_id_i(rf_wdata_id),
		.rf_we_id_i(rf_we_id),
		.dummy_instr_id_i(dummy_instr_id),
		.rf_wdata_lsu_i(rf_wdata_lsu),
		.rf_we_lsu_i(rf_we_lsu),
		.rf_wdata_fwd_wb_o(rf_wdata_fwd_wb),
		.rf_waddr_wb_o(rf_waddr_wb),
		.rf_wdata_wb_o(rf_wdata_wb),
		.rf_we_wb_o(rf_we_wb),
		.dummy_instr_wb_o(dummy_instr_wb),
		.lsu_resp_valid_i(lsu_resp_valid),
		.lsu_resp_err_i(lsu_resp_err),
		.instr_done_wb_o(instr_done_wb)
	);
	assign dummy_instr_id_o = dummy_instr_id;
	assign dummy_instr_wb_o = dummy_instr_wb;
	assign rf_raddr_a_o = rf_raddr_a;
	assign rf_waddr_wb_o = rf_waddr_wb;
	assign rf_we_wb_o = rf_we_wb;
	assign rf_raddr_b_o = rf_raddr_b;
	generate
		if (RegFileECC) begin : gen_regfile_ecc
			wire [1:0] rf_ecc_err_a;
			wire [1:0] rf_ecc_err_b;
			wire rf_ecc_err_a_id;
			wire rf_ecc_err_b_id;
			prim_secded_inv_39_32_enc regfile_ecc_enc(
				.data_i(rf_wdata_wb),
				.data_o(rf_wdata_wb_ecc_o)
			);
			prim_secded_inv_39_32_dec regfile_ecc_dec_a(
				.data_i(rf_rdata_a_ecc_i),
				.err_o(rf_ecc_err_a)
			);
			prim_secded_inv_39_32_dec regfile_ecc_dec_b(
				.data_i(rf_rdata_b_ecc_i),
				.err_o(rf_ecc_err_b)
			);
			assign rf_rdata_a = rf_rdata_a_ecc_i[31:0];
			assign rf_rdata_b = rf_rdata_b_ecc_i[31:0];
			assign rf_ecc_err_a_id = (|rf_ecc_err_a & rf_ren_a) & ~rf_rd_a_wb_match;
			assign rf_ecc_err_b_id = (|rf_ecc_err_b & rf_ren_b) & ~rf_rd_b_wb_match;
			assign rf_ecc_err_comb = instr_valid_id & (rf_ecc_err_a_id | rf_ecc_err_b_id);
		end
		else begin : gen_no_regfile_ecc
			wire unused_rf_ren_a;
			wire unused_rf_ren_b;
			wire unused_rf_rd_a_wb_match;
			wire unused_rf_rd_b_wb_match;
			assign unused_rf_ren_a = rf_ren_a;
			assign unused_rf_ren_b = rf_ren_b;
			assign unused_rf_rd_a_wb_match = rf_rd_a_wb_match;
			assign unused_rf_rd_b_wb_match = rf_rd_b_wb_match;
			assign rf_wdata_wb_ecc_o = rf_wdata_wb;
			assign rf_rdata_a = rf_rdata_a_ecc_i;
			assign rf_rdata_b = rf_rdata_b_ecc_i;
			assign rf_ecc_err_comb = 1'b0;
		end
	endgenerate
	wire [31:0] crash_dump_mtval;
	assign crash_dump_o[159-:32] = pc_id;
	assign crash_dump_o[127-:32] = pc_if;
	assign crash_dump_o[95-:32] = lsu_addr_last;
	assign crash_dump_o[63-:32] = csr_mepc;
	assign crash_dump_o[31-:32] = crash_dump_mtval;
	assign alert_minor_o = icache_ecc_error;
	assign alert_major_internal_o = (rf_ecc_err_comb | pc_mismatch_alert) | csr_shadow_err;
	assign alert_major_bus_o = (lsu_load_resp_intg_err | lsu_store_resp_intg_err) | instr_intg_err;
	assign csr_wdata = alu_operand_a_ex;
	function automatic [11:0] sv2v_cast_12;
		input reg [11:0] inp;
		sv2v_cast_12 = inp;
	endfunction
	assign csr_addr = sv2v_cast_12((csr_access ? alu_operand_b_ex[11:0] : 12'b000000000000));
	ibex_cs_registers #(
		.DbgTriggerEn(DbgTriggerEn),
		.DbgHwBreakNum(DbgHwBreakNum),
		.DataIndTiming(DataIndTiming),
		.DummyInstructions(DummyInstructions),
		.ShadowCSR(ShadowCSR),
		.ICache(ICache),
		.MHPMCounterNum(MHPMCounterNum),
		.MHPMCounterWidth(MHPMCounterWidth),
		.PMPEnable(PMPEnable),
		.PMPGranularity(PMPGranularity),
		.PMPNumRegions(PMPNumRegions),
		.RV32E(RV32E),
		.RV32M(RV32M),
		.RV32B(RV32B)
	) cs_registers_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.hart_id_i(hart_id_i),
		.priv_mode_id_o(priv_mode_id),
		.priv_mode_lsu_o(priv_mode_lsu),
		.csr_mtvec_o(csr_mtvec),
		.csr_mtvec_init_i(csr_mtvec_init),
		.boot_addr_i(boot_addr_i),
		.csr_access_i(csr_access),
		.csr_addr_i(csr_addr),
		.csr_wdata_i(csr_wdata),
		.csr_op_i(csr_op),
		.csr_op_en_i(csr_op_en),
		.csr_rdata_o(csr_rdata),
		.irq_software_i(irq_software_i),
		.irq_timer_i(irq_timer_i),
		.irq_external_i(irq_external_i),
		.irq_fast_i(irq_fast_i),
		.nmi_mode_i(nmi_mode),
		.irq_pending_o(irq_pending_o),
		.irqs_o(irqs),
		.csr_mstatus_mie_o(csr_mstatus_mie),
		.csr_mstatus_tw_o(csr_mstatus_tw),
		.csr_mepc_o(csr_mepc),
		.csr_mtval_o(crash_dump_mtval),
		.csr_pmp_cfg_o(csr_pmp_cfg),
		.csr_pmp_addr_o(csr_pmp_addr),
		.csr_pmp_mseccfg_o(csr_pmp_mseccfg),
		.csr_depc_o(csr_depc),
		.debug_mode_i(debug_mode),
		.debug_mode_entering_i(debug_mode_entering),
		.debug_cause_i(debug_cause),
		.debug_csr_save_i(debug_csr_save),
		.debug_single_step_o(debug_single_step),
		.debug_ebreakm_o(debug_ebreakm),
		.debug_ebreaku_o(debug_ebreaku),
		.trigger_match_o(trigger_match),
		.pc_if_i(pc_if),
		.pc_id_i(pc_id),
		.pc_wb_i(pc_wb),
		.data_ind_timing_o(data_ind_timing),
		.dummy_instr_en_o(dummy_instr_en),
		.dummy_instr_mask_o(dummy_instr_mask),
		.dummy_instr_seed_en_o(dummy_instr_seed_en),
		.dummy_instr_seed_o(dummy_instr_seed),
		.icache_enable_o(icache_enable),
		.csr_shadow_err_o(csr_shadow_err),
		.ic_scr_key_valid_i(ic_scr_key_valid_i),
		.csr_save_if_i(csr_save_if),
		.csr_save_id_i(csr_save_id),
		.csr_save_wb_i(csr_save_wb),
		.csr_restore_mret_i(csr_restore_mret_id),
		.csr_restore_dret_i(csr_restore_dret_id),
		.csr_save_cause_i(csr_save_cause),
		.csr_mcause_i(exc_cause),
		.csr_mtval_i(csr_mtval),
		.illegal_csr_insn_o(illegal_csr_insn_id),
		.double_fault_seen_o(double_fault_seen_o),
		.instr_ret_i(perf_instr_ret_wb),
		.instr_ret_compressed_i(perf_instr_ret_compressed_wb),
		.instr_ret_spec_i(perf_instr_ret_wb_spec),
		.instr_ret_compressed_spec_i(perf_instr_ret_compressed_wb_spec),
		.iside_wait_i(perf_iside_wait),
		.jump_i(perf_jump),
		.branch_i(perf_branch),
		.branch_taken_i(perf_tbranch),
		.mem_load_i(perf_load),
		.mem_store_i(perf_store),
		.dside_wait_i(perf_dside_wait),
		.mul_wait_i(perf_mul_wait),
		.div_wait_i(perf_div_wait)
	);
	generate
		if (PMPEnable) begin : g_pmp
			wire [31:0] pc_if_inc;
			wire [101:0] pmp_req_addr;
			wire [5:0] pmp_req_type;
			wire [5:0] pmp_priv_lvl;
			assign pc_if_inc = pc_if + 32'd2;
			assign pmp_req_addr[68+:34] = {2'b00, pc_if};
			assign pmp_req_type[4+:2] = 2'b00;
			assign pmp_priv_lvl[4+:2] = priv_mode_id;
			assign pmp_req_addr[34+:34] = {2'b00, pc_if_inc};
			assign pmp_req_type[2+:2] = 2'b00;
			assign pmp_priv_lvl[2+:2] = priv_mode_id;
			assign pmp_req_addr[0+:34] = {2'b00, data_addr_o[31:0]};
			assign pmp_req_type[0+:2] = (data_we_o ? 2'b01 : 2'b10);
			assign pmp_priv_lvl[0+:2] = priv_mode_lsu;
			ibex_pmp #(
				.PMPGranularity(PMPGranularity),
				.PMPNumChan(PMPNumChan),
				.PMPNumRegions(PMPNumRegions)
			) pmp_i(
				.csr_pmp_cfg_i(csr_pmp_cfg),
				.csr_pmp_addr_i(csr_pmp_addr),
				.csr_pmp_mseccfg_i(csr_pmp_mseccfg),
				.priv_mode_i(pmp_priv_lvl),
				.pmp_req_addr_i(pmp_req_addr),
				.pmp_req_type_i(pmp_req_type),
				.pmp_req_err_o(pmp_req_err)
			);
		end
		else begin : g_no_pmp
			wire [1:0] unused_priv_lvl_ls;
			wire [(PMPNumRegions * 34) - 1:0] unused_csr_pmp_addr;
			wire [(PMPNumRegions * 6) - 1:0] unused_csr_pmp_cfg;
			wire [2:0] unused_csr_pmp_mseccfg;
			assign unused_priv_lvl_ls = priv_mode_lsu;
			assign unused_csr_pmp_addr = csr_pmp_addr;
			assign unused_csr_pmp_cfg = csr_pmp_cfg;
			assign unused_csr_pmp_mseccfg = csr_pmp_mseccfg;
			assign pmp_req_err[ibex_pkg_PMP_I] = 1'b0;
			assign pmp_req_err[ibex_pkg_PMP_I2] = 1'b0;
			assign pmp_req_err[ibex_pkg_PMP_D] = 1'b0;
		end
	endgenerate
	wire unused_instr_new_id;
	wire unused_instr_id_done;
	wire unused_instr_done_wb;
	assign unused_instr_id_done = instr_id_done;
	assign unused_instr_new_id = instr_new_id;
	assign unused_instr_done_wb = instr_done_wb;
endmodule
module ibex_counter (
	clk_i,
	rst_ni,
	counter_inc_i,
	counterh_we_i,
	counter_we_i,
	counter_val_i,
	counter_val_o,
	counter_val_upd_o
);
	parameter signed [31:0] CounterWidth = 32;
	parameter [0:0] ProvideValUpd = 0;
	input wire clk_i;
	input wire rst_ni;
	input wire counter_inc_i;
	input wire counterh_we_i;
	input wire counter_we_i;
	input wire [31:0] counter_val_i;
	output wire [63:0] counter_val_o;
	output wire [63:0] counter_val_upd_o;
	wire [63:0] counter;
	wire [CounterWidth - 1:0] counter_upd;
	reg [63:0] counter_load;
	reg we;
	reg [CounterWidth - 1:0] counter_d;
	assign counter_upd = counter[CounterWidth - 1:0] + {{CounterWidth - 1 {1'b0}}, 1'b1};
	always @(*) begin
		we = counter_we_i | counterh_we_i;
		counter_load[63:32] = counter[63:32];
		counter_load[31:0] = counter_val_i;
		if (counterh_we_i) begin
			counter_load[63:32] = counter_val_i;
			counter_load[31:0] = counter[31:0];
		end
		if (we)
			counter_d = counter_load[CounterWidth - 1:0];
		else if (counter_inc_i)
			counter_d = counter_upd[CounterWidth - 1:0];
		else
			counter_d = counter[CounterWidth - 1:0];
	end
	reg [CounterWidth - 1:0] counter_q;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			counter_q <= 1'sb0;
		else
			counter_q <= counter_d;
	generate
		if (CounterWidth < 64) begin : g_counter_narrow
			wire [63:CounterWidth] unused_counter_load;
			assign counter[CounterWidth - 1:0] = counter_q;
			assign counter[63:CounterWidth] = 1'sb0;
			if (ProvideValUpd) begin : g_counter_val_upd_o
				assign counter_val_upd_o[CounterWidth - 1:0] = counter_upd;
			end
			else begin : g_no_counter_val_upd_o
				assign counter_val_upd_o[CounterWidth - 1:0] = 1'sb0;
			end
			assign counter_val_upd_o[63:CounterWidth] = 1'sb0;
			assign unused_counter_load = counter_load[63:CounterWidth];
		end
		else begin : g_counter_full
			assign counter = counter_q;
			if (ProvideValUpd) begin : g_counter_val_upd_o
				assign counter_val_upd_o = counter_upd;
			end
			else begin : g_no_counter_val_upd_o
				assign counter_val_upd_o = 1'sb0;
			end
		end
	endgenerate
	assign counter_val_o = counter;
endmodule
module ibex_cs_registers (
	clk_i,
	rst_ni,
	hart_id_i,
	priv_mode_id_o,
	priv_mode_lsu_o,
	csr_mstatus_tw_o,
	csr_mtvec_o,
	csr_mtvec_init_i,
	boot_addr_i,
	csr_access_i,
	csr_addr_i,
	csr_wdata_i,
	csr_op_i,
	csr_op_en_i,
	csr_rdata_o,
	irq_software_i,
	irq_timer_i,
	irq_external_i,
	irq_fast_i,
	nmi_mode_i,
	irq_pending_o,
	irqs_o,
	csr_mstatus_mie_o,
	csr_mepc_o,
	csr_mtval_o,
	csr_pmp_cfg_o,
	csr_pmp_addr_o,
	csr_pmp_mseccfg_o,
	debug_mode_i,
	debug_mode_entering_i,
	debug_cause_i,
	debug_csr_save_i,
	csr_depc_o,
	debug_single_step_o,
	debug_ebreakm_o,
	debug_ebreaku_o,
	trigger_match_o,
	pc_if_i,
	pc_id_i,
	pc_wb_i,
	data_ind_timing_o,
	dummy_instr_en_o,
	dummy_instr_mask_o,
	dummy_instr_seed_en_o,
	dummy_instr_seed_o,
	icache_enable_o,
	csr_shadow_err_o,
	ic_scr_key_valid_i,
	csr_save_if_i,
	csr_save_id_i,
	csr_save_wb_i,
	csr_restore_mret_i,
	csr_restore_dret_i,
	csr_save_cause_i,
	csr_mcause_i,
	csr_mtval_i,
	illegal_csr_insn_o,
	double_fault_seen_o,
	instr_ret_i,
	instr_ret_compressed_i,
	instr_ret_spec_i,
	instr_ret_compressed_spec_i,
	iside_wait_i,
	jump_i,
	branch_i,
	branch_taken_i,
	mem_load_i,
	mem_store_i,
	dside_wait_i,
	mul_wait_i,
	div_wait_i
);
	parameter [0:0] DbgTriggerEn = 0;
	parameter [31:0] DbgHwBreakNum = 1;
	parameter [0:0] DataIndTiming = 1'b0;
	parameter [0:0] DummyInstructions = 1'b0;
	parameter [0:0] ShadowCSR = 1'b0;
	parameter [0:0] ICache = 1'b0;
	parameter [31:0] MHPMCounterNum = 10;
	parameter [31:0] MHPMCounterWidth = 40;
	parameter [0:0] PMPEnable = 0;
	parameter [31:0] PMPGranularity = 0;
	parameter [31:0] PMPNumRegions = 4;
	parameter [0:0] RV32E = 0;
	parameter integer RV32M = 32'sd2;
	parameter integer RV32B = 32'sd0;
	input wire clk_i;
	input wire rst_ni;
	input wire [31:0] hart_id_i;
	output wire [1:0] priv_mode_id_o;
	output wire [1:0] priv_mode_lsu_o;
	output wire csr_mstatus_tw_o;
	output wire [31:0] csr_mtvec_o;
	input wire csr_mtvec_init_i;
	input wire [31:0] boot_addr_i;
	input wire csr_access_i;
	input wire [11:0] csr_addr_i;
	input wire [31:0] csr_wdata_i;
	input wire [1:0] csr_op_i;
	input csr_op_en_i;
	output wire [31:0] csr_rdata_o;
	input wire irq_software_i;
	input wire irq_timer_i;
	input wire irq_external_i;
	input wire [14:0] irq_fast_i;
	input wire nmi_mode_i;
	output wire irq_pending_o;
	output wire [17:0] irqs_o;
	output wire csr_mstatus_mie_o;
	output wire [31:0] csr_mepc_o;
	output wire [31:0] csr_mtval_o;
	output wire [(PMPNumRegions * 6) - 1:0] csr_pmp_cfg_o;
	output wire [(PMPNumRegions * 34) - 1:0] csr_pmp_addr_o;
	output wire [2:0] csr_pmp_mseccfg_o;
	input wire debug_mode_i;
	input wire debug_mode_entering_i;
	input wire [2:0] debug_cause_i;
	input wire debug_csr_save_i;
	output wire [31:0] csr_depc_o;
	output wire debug_single_step_o;
	output wire debug_ebreakm_o;
	output wire debug_ebreaku_o;
	output wire trigger_match_o;
	input wire [31:0] pc_if_i;
	input wire [31:0] pc_id_i;
	input wire [31:0] pc_wb_i;
	output wire data_ind_timing_o;
	output wire dummy_instr_en_o;
	output wire [2:0] dummy_instr_mask_o;
	output wire dummy_instr_seed_en_o;
	output wire [31:0] dummy_instr_seed_o;
	output wire icache_enable_o;
	output wire csr_shadow_err_o;
	input wire ic_scr_key_valid_i;
	input wire csr_save_if_i;
	input wire csr_save_id_i;
	input wire csr_save_wb_i;
	input wire csr_restore_mret_i;
	input wire csr_restore_dret_i;
	input wire csr_save_cause_i;
	input wire [6:0] csr_mcause_i;
	input wire [31:0] csr_mtval_i;
	output wire illegal_csr_insn_o;
	output reg double_fault_seen_o;
	input wire instr_ret_i;
	input wire instr_ret_compressed_i;
	input wire instr_ret_spec_i;
	input wire instr_ret_compressed_spec_i;
	input wire iside_wait_i;
	input wire jump_i;
	input wire branch_i;
	input wire branch_taken_i;
	input wire mem_load_i;
	input wire mem_store_i;
	input wire dside_wait_i;
	input wire mul_wait_i;
	input wire div_wait_i;
	function automatic is_mml_m_exec_cfg;
		input reg [5:0] pmp_cfg;
		reg unused_cfg;
		reg value;
		begin
			unused_cfg = ^{pmp_cfg[4-:2]};
			value = 1'b0;
			if (pmp_cfg[5])
				case ({pmp_cfg[0], pmp_cfg[1], pmp_cfg[2]})
					3'b001, 3'b010, 3'b011, 3'b101: value = 1'b1;
					default: value = 1'b0;
				endcase
			is_mml_m_exec_cfg = value;
		end
	endfunction
	localparam [31:0] RV32BExtra = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? 1 : 0);
	localparam [31:0] RV32MEnabled = (RV32M == 32'sd0 ? 0 : 1);
	localparam [31:0] PMPAddrWidth = (PMPGranularity > 0 ? 33 - PMPGranularity : 32);
	localparam [1:0] ibex_pkg_CSR_MISA_MXL = 2'd1;
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	localparam [31:0] MISA_VALUE = (((((((((((0 | 0) | 4) | 0) | (sv2v_cast_32(RV32E) << 4)) | 0) | (sv2v_cast_32(!RV32E) << 8)) | (RV32MEnabled << 12)) | 0) | 0) | 1048576) | (RV32BExtra << 23)) | (sv2v_cast_32(ibex_pkg_CSR_MISA_MXL) << 30);
	reg [31:0] exception_pc;
	reg [1:0] priv_lvl_q;
	reg [1:0] priv_lvl_d;
	wire [5:0] mstatus_q;
	reg [5:0] mstatus_d;
	wire mstatus_err;
	reg mstatus_en;
	wire [17:0] mie_q;
	wire [17:0] mie_d;
	reg mie_en;
	wire [31:0] mscratch_q;
	reg mscratch_en;
	wire [31:0] mepc_q;
	reg [31:0] mepc_d;
	reg mepc_en;
	wire [6:0] mcause_q;
	reg [6:0] mcause_d;
	reg mcause_en;
	wire [31:0] mtval_q;
	reg [31:0] mtval_d;
	reg mtval_en;
	wire [31:0] mtvec_q;
	reg [31:0] mtvec_d;
	wire mtvec_err;
	reg mtvec_en;
	wire [17:0] mip;
	wire [31:0] dcsr_q;
	reg [31:0] dcsr_d;
	reg dcsr_en;
	wire [31:0] depc_q;
	reg [31:0] depc_d;
	reg depc_en;
	wire [31:0] dscratch0_q;
	wire [31:0] dscratch1_q;
	reg dscratch0_en;
	reg dscratch1_en;
	wire [2:0] mstack_q;
	reg [2:0] mstack_d;
	reg mstack_en;
	wire [31:0] mstack_epc_q;
	reg [31:0] mstack_epc_d;
	wire [6:0] mstack_cause_q;
	reg [6:0] mstack_cause_d;
	localparam [31:0] ibex_pkg_PMP_MAX_REGIONS = 16;
	reg [31:0] pmp_addr_rdata [0:15];
	localparam [31:0] ibex_pkg_PMP_CFG_W = 8;
	wire [7:0] pmp_cfg_rdata [0:15];
	wire pmp_csr_err;
	wire [2:0] pmp_mseccfg;
	wire [31:0] mcountinhibit;
	reg [MHPMCounterNum + 2:0] mcountinhibit_d;
	reg [MHPMCounterNum + 2:0] mcountinhibit_q;
	reg mcountinhibit_we;
	wire [63:0] mhpmcounter [0:31];
	reg [31:0] mhpmcounter_we;
	reg [31:0] mhpmcounterh_we;
	reg [31:0] mhpmcounter_incr;
	reg [31:0] mhpmevent [0:31];
	wire [4:0] mhpmcounter_idx;
	wire unused_mhpmcounter_we_1;
	wire unused_mhpmcounterh_we_1;
	wire unused_mhpmcounter_incr_1;
	wire [63:0] minstret_next;
	wire [63:0] minstret_raw;
	wire [31:0] tselect_rdata;
	wire [31:0] tmatch_control_rdata;
	wire [31:0] tmatch_value_rdata;
	wire [7:0] cpuctrlsts_part_q;
	reg [7:0] cpuctrlsts_part_d;
	wire [7:0] cpuctrlsts_part_wdata_raw;
	wire [7:0] cpuctrlsts_part_wdata;
	reg cpuctrlsts_part_we;
	wire cpuctrlsts_part_err;
	wire cpuctrlsts_ic_scr_key_valid_q;
	wire cpuctrlsts_ic_scr_key_err;
	reg [31:0] csr_wdata_int;
	reg [31:0] csr_rdata_int;
	wire csr_we_int;
	wire csr_wr;
	reg dbg_csr;
	reg illegal_csr;
	wire illegal_csr_priv;
	wire illegal_csr_dbg;
	wire illegal_csr_write;
	wire [7:0] unused_boot_addr;
	wire [2:0] unused_csr_addr;
	assign unused_boot_addr = boot_addr_i[7:0];
	wire [11:0] csr_addr;
	assign csr_addr = {csr_addr_i};
	assign unused_csr_addr = csr_addr[7:5];
	assign mhpmcounter_idx = csr_addr[4:0];
	assign illegal_csr_dbg = dbg_csr & ~debug_mode_i;
	assign illegal_csr_priv = csr_addr[9:8] > {priv_lvl_q};
	assign illegal_csr_write = (csr_addr[11:10] == 2'b11) && csr_wr;
	assign illegal_csr_insn_o = csr_access_i & (((illegal_csr | illegal_csr_write) | illegal_csr_priv) | illegal_csr_dbg);
	assign mip[17] = irq_software_i;
	assign mip[16] = irq_timer_i;
	assign mip[15] = irq_external_i;
	assign mip[14-:15] = irq_fast_i;
	localparam [31:0] ibex_pkg_CSR_MARCHID_VALUE = 32'b00000000000000000000000000010110;
	localparam [31:0] ibex_pkg_CSR_MCONFIGPTR_VALUE = 32'b00000000000000000000000000000000;
	localparam [31:0] ibex_pkg_CSR_MEIX_BIT = 11;
	localparam [31:0] ibex_pkg_CSR_MFIX_BIT_HIGH = 30;
	localparam [31:0] ibex_pkg_CSR_MFIX_BIT_LOW = 16;
	localparam [31:0] ibex_pkg_CSR_MIMPID_VALUE = 32'b00000000000000000000000000000000;
	localparam [31:0] ibex_pkg_CSR_MSECCFG_MML_BIT = 0;
	localparam [31:0] ibex_pkg_CSR_MSECCFG_MMWP_BIT = 1;
	localparam [31:0] ibex_pkg_CSR_MSECCFG_RLB_BIT = 2;
	localparam [31:0] ibex_pkg_CSR_MSIX_BIT = 3;
	localparam [31:0] ibex_pkg_CSR_MSTATUS_MIE_BIT = 3;
	localparam [31:0] ibex_pkg_CSR_MSTATUS_MPIE_BIT = 7;
	localparam [31:0] ibex_pkg_CSR_MSTATUS_MPP_BIT_HIGH = 12;
	localparam [31:0] ibex_pkg_CSR_MSTATUS_MPP_BIT_LOW = 11;
	localparam [31:0] ibex_pkg_CSR_MSTATUS_MPRV_BIT = 17;
	localparam [31:0] ibex_pkg_CSR_MSTATUS_TW_BIT = 21;
	localparam [31:0] ibex_pkg_CSR_MTIX_BIT = 7;
	localparam [31:0] ibex_pkg_CSR_MVENDORID_VALUE = 32'b00000000000000000000000000000000;
	always @(*) begin
		csr_rdata_int = 1'sb0;
		illegal_csr = 1'b0;
		dbg_csr = 1'b0;
		case (csr_addr_i)
			12'hf11: csr_rdata_int = ibex_pkg_CSR_MVENDORID_VALUE;
			12'hf12: csr_rdata_int = ibex_pkg_CSR_MARCHID_VALUE;
			12'hf13: csr_rdata_int = ibex_pkg_CSR_MIMPID_VALUE;
			12'hf14: csr_rdata_int = hart_id_i;
			12'hf15: csr_rdata_int = ibex_pkg_CSR_MCONFIGPTR_VALUE;
			12'h300: begin
				csr_rdata_int = 1'sb0;
				csr_rdata_int[ibex_pkg_CSR_MSTATUS_MIE_BIT] = mstatus_q[5];
				csr_rdata_int[ibex_pkg_CSR_MSTATUS_MPIE_BIT] = mstatus_q[4];
				csr_rdata_int[ibex_pkg_CSR_MSTATUS_MPP_BIT_HIGH:ibex_pkg_CSR_MSTATUS_MPP_BIT_LOW] = mstatus_q[3-:2];
				csr_rdata_int[ibex_pkg_CSR_MSTATUS_MPRV_BIT] = mstatus_q[1];
				csr_rdata_int[ibex_pkg_CSR_MSTATUS_TW_BIT] = mstatus_q[0];
			end
			12'h310: csr_rdata_int = 1'sb0;
			12'h30a, 12'h31a: csr_rdata_int = 1'sb0;
			12'h301: csr_rdata_int = MISA_VALUE;
			12'h304: begin
				csr_rdata_int = 1'sb0;
				csr_rdata_int[ibex_pkg_CSR_MSIX_BIT] = mie_q[17];
				csr_rdata_int[ibex_pkg_CSR_MTIX_BIT] = mie_q[16];
				csr_rdata_int[ibex_pkg_CSR_MEIX_BIT] = mie_q[15];
				csr_rdata_int[ibex_pkg_CSR_MFIX_BIT_HIGH:ibex_pkg_CSR_MFIX_BIT_LOW] = mie_q[14-:15];
			end
			12'h306: csr_rdata_int = 1'sb0;
			12'h340: csr_rdata_int = mscratch_q;
			12'h305: csr_rdata_int = mtvec_q;
			12'h341: csr_rdata_int = mepc_q;
			12'h342: csr_rdata_int = {mcause_q[5] | mcause_q[6], (mcause_q[6] ? {26 {1'b1}} : 26'b00000000000000000000000000), mcause_q[4:0]};
			12'h343: csr_rdata_int = mtval_q;
			12'h344: begin
				csr_rdata_int = 1'sb0;
				csr_rdata_int[ibex_pkg_CSR_MSIX_BIT] = mip[17];
				csr_rdata_int[ibex_pkg_CSR_MTIX_BIT] = mip[16];
				csr_rdata_int[ibex_pkg_CSR_MEIX_BIT] = mip[15];
				csr_rdata_int[ibex_pkg_CSR_MFIX_BIT_HIGH:ibex_pkg_CSR_MFIX_BIT_LOW] = mip[14-:15];
			end
			12'h747:
				if (PMPEnable) begin
					csr_rdata_int = 1'sb0;
					csr_rdata_int[ibex_pkg_CSR_MSECCFG_MML_BIT] = pmp_mseccfg[0];
					csr_rdata_int[ibex_pkg_CSR_MSECCFG_MMWP_BIT] = pmp_mseccfg[1];
					csr_rdata_int[ibex_pkg_CSR_MSECCFG_RLB_BIT] = pmp_mseccfg[2];
				end
				else
					illegal_csr = 1'b1;
			12'h757:
				if (PMPEnable)
					csr_rdata_int = 1'sb0;
				else
					illegal_csr = 1'b1;
			12'h3a0: csr_rdata_int = {pmp_cfg_rdata[3], pmp_cfg_rdata[2], pmp_cfg_rdata[1], pmp_cfg_rdata[0]};
			12'h3a1: csr_rdata_int = {pmp_cfg_rdata[7], pmp_cfg_rdata[6], pmp_cfg_rdata[5], pmp_cfg_rdata[4]};
			12'h3a2: csr_rdata_int = {pmp_cfg_rdata[11], pmp_cfg_rdata[10], pmp_cfg_rdata[9], pmp_cfg_rdata[8]};
			12'h3a3: csr_rdata_int = {pmp_cfg_rdata[15], pmp_cfg_rdata[14], pmp_cfg_rdata[13], pmp_cfg_rdata[12]};
			12'h3b0: csr_rdata_int = pmp_addr_rdata[0];
			12'h3b1: csr_rdata_int = pmp_addr_rdata[1];
			12'h3b2: csr_rdata_int = pmp_addr_rdata[2];
			12'h3b3: csr_rdata_int = pmp_addr_rdata[3];
			12'h3b4: csr_rdata_int = pmp_addr_rdata[4];
			12'h3b5: csr_rdata_int = pmp_addr_rdata[5];
			12'h3b6: csr_rdata_int = pmp_addr_rdata[6];
			12'h3b7: csr_rdata_int = pmp_addr_rdata[7];
			12'h3b8: csr_rdata_int = pmp_addr_rdata[8];
			12'h3b9: csr_rdata_int = pmp_addr_rdata[9];
			12'h3ba: csr_rdata_int = pmp_addr_rdata[10];
			12'h3bb: csr_rdata_int = pmp_addr_rdata[11];
			12'h3bc: csr_rdata_int = pmp_addr_rdata[12];
			12'h3bd: csr_rdata_int = pmp_addr_rdata[13];
			12'h3be: csr_rdata_int = pmp_addr_rdata[14];
			12'h3bf: csr_rdata_int = pmp_addr_rdata[15];
			12'h7b0: begin
				csr_rdata_int = dcsr_q;
				dbg_csr = 1'b1;
			end
			12'h7b1: begin
				csr_rdata_int = depc_q;
				dbg_csr = 1'b1;
			end
			12'h7b2: begin
				csr_rdata_int = dscratch0_q;
				dbg_csr = 1'b1;
			end
			12'h7b3: begin
				csr_rdata_int = dscratch1_q;
				dbg_csr = 1'b1;
			end
			12'h320: csr_rdata_int = mcountinhibit;
			12'h323, 12'h324, 12'h325, 12'h326, 12'h327, 12'h328, 12'h329, 12'h32a, 12'h32b, 12'h32c, 12'h32d, 12'h32e, 12'h32f, 12'h330, 12'h331, 12'h332, 12'h333, 12'h334, 12'h335, 12'h336, 12'h337, 12'h338, 12'h339, 12'h33a, 12'h33b, 12'h33c, 12'h33d, 12'h33e, 12'h33f: csr_rdata_int = mhpmevent[mhpmcounter_idx];
			12'hb00, 12'hb02, 12'hb03, 12'hb04, 12'hb05, 12'hb06, 12'hb07, 12'hb08, 12'hb09, 12'hb0a, 12'hb0b, 12'hb0c, 12'hb0d, 12'hb0e, 12'hb0f, 12'hb10, 12'hb11, 12'hb12, 12'hb13, 12'hb14, 12'hb15, 12'hb16, 12'hb17, 12'hb18, 12'hb19, 12'hb1a, 12'hb1b, 12'hb1c, 12'hb1d, 12'hb1e, 12'hb1f: csr_rdata_int = mhpmcounter[mhpmcounter_idx][31:0];
			12'hb80, 12'hb82, 12'hb83, 12'hb84, 12'hb85, 12'hb86, 12'hb87, 12'hb88, 12'hb89, 12'hb8a, 12'hb8b, 12'hb8c, 12'hb8d, 12'hb8e, 12'hb8f, 12'hb90, 12'hb91, 12'hb92, 12'hb93, 12'hb94, 12'hb95, 12'hb96, 12'hb97, 12'hb98, 12'hb99, 12'hb9a, 12'hb9b, 12'hb9c, 12'hb9d, 12'hb9e, 12'hb9f: csr_rdata_int = mhpmcounter[mhpmcounter_idx][63:32];
			12'h7a0: begin
				csr_rdata_int = tselect_rdata;
				illegal_csr = ~DbgTriggerEn;
			end
			12'h7a1: begin
				csr_rdata_int = tmatch_control_rdata;
				illegal_csr = ~DbgTriggerEn;
			end
			12'h7a2: begin
				csr_rdata_int = tmatch_value_rdata;
				illegal_csr = ~DbgTriggerEn;
			end
			12'h7a3: begin
				csr_rdata_int = 1'sb0;
				illegal_csr = ~DbgTriggerEn;
			end
			12'h7a8: begin
				csr_rdata_int = 1'sb0;
				illegal_csr = ~DbgTriggerEn;
			end
			12'h5a8: begin
				csr_rdata_int = 1'sb0;
				illegal_csr = ~DbgTriggerEn;
			end
			12'h7aa: begin
				csr_rdata_int = 1'sb0;
				illegal_csr = ~DbgTriggerEn;
			end
			12'h7c0: csr_rdata_int = {{23 {1'b0}}, cpuctrlsts_ic_scr_key_valid_q, cpuctrlsts_part_q};
			12'h7c1: csr_rdata_int = 1'sb0;
			default: illegal_csr = 1'b1;
		endcase
		if (!PMPEnable)
			if (|{csr_addr == 12'h3a0, csr_addr == 12'h3a1, csr_addr == 12'h3a2, csr_addr == 12'h3a3, csr_addr == 12'h3b0, csr_addr == 12'h3b1, csr_addr == 12'h3b2, csr_addr == 12'h3b3, csr_addr == 12'h3b4, csr_addr == 12'h3b5, csr_addr == 12'h3b6, csr_addr == 12'h3b7, csr_addr == 12'h3b8, csr_addr == 12'h3b9, csr_addr == 12'h3ba, csr_addr == 12'h3bb, csr_addr == 12'h3bc, csr_addr == 12'h3bd, csr_addr == 12'h3be, csr_addr == 12'h3bf})
				illegal_csr = 1'b1;
	end
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	always @(*) begin
		exception_pc = pc_id_i;
		priv_lvl_d = priv_lvl_q;
		mstatus_en = 1'b0;
		mstatus_d = mstatus_q;
		mie_en = 1'b0;
		mscratch_en = 1'b0;
		mepc_en = 1'b0;
		mepc_d = {csr_wdata_int[31:1], 1'b0};
		mcause_en = 1'b0;
		mcause_d = {csr_wdata_int[31:30] == 2'b11, csr_wdata_int[31:30] == 2'b10, csr_wdata_int[4:0]};
		mtval_en = 1'b0;
		mtval_d = csr_wdata_int;
		mtvec_en = csr_mtvec_init_i;
		mtvec_d = (csr_mtvec_init_i ? {boot_addr_i[31:8], 6'b000000, 2'b01} : {csr_wdata_int[31:8], 6'b000000, 2'b01});
		dcsr_en = 1'b0;
		dcsr_d = dcsr_q;
		depc_d = {csr_wdata_int[31:1], 1'b0};
		depc_en = 1'b0;
		dscratch0_en = 1'b0;
		dscratch1_en = 1'b0;
		mstack_en = 1'b0;
		mstack_d[2] = mstatus_q[4];
		mstack_d[1-:2] = mstatus_q[3-:2];
		mstack_epc_d = mepc_q;
		mstack_cause_d = mcause_q;
		mcountinhibit_we = 1'b0;
		mhpmcounter_we = 1'sb0;
		mhpmcounterh_we = 1'sb0;
		cpuctrlsts_part_we = 1'b0;
		cpuctrlsts_part_d = cpuctrlsts_part_q;
		double_fault_seen_o = 1'b0;
		if (csr_we_int)
			case (csr_addr_i)
				12'h300: begin
					mstatus_en = 1'b1;
					mstatus_d = {csr_wdata_int[ibex_pkg_CSR_MSTATUS_MIE_BIT], csr_wdata_int[ibex_pkg_CSR_MSTATUS_MPIE_BIT], sv2v_cast_2(csr_wdata_int[ibex_pkg_CSR_MSTATUS_MPP_BIT_HIGH:ibex_pkg_CSR_MSTATUS_MPP_BIT_LOW]), csr_wdata_int[ibex_pkg_CSR_MSTATUS_MPRV_BIT], csr_wdata_int[ibex_pkg_CSR_MSTATUS_TW_BIT]};
					if ((mstatus_d[3-:2] != 2'b11) && (mstatus_d[3-:2] != 2'b00))
						mstatus_d[3-:2] = 2'b00;
				end
				12'h304: mie_en = 1'b1;
				12'h340: mscratch_en = 1'b1;
				12'h341: mepc_en = 1'b1;
				12'h342: mcause_en = 1'b1;
				12'h343: mtval_en = 1'b1;
				12'h305: mtvec_en = 1'b1;
				12'h7b0: begin
					dcsr_d = csr_wdata_int;
					dcsr_d[31-:4] = 4'd4;
					if ((dcsr_d[1-:2] != 2'b11) && (dcsr_d[1-:2] != 2'b00))
						dcsr_d[1-:2] = 2'b00;
					dcsr_d[8-:3] = dcsr_q[8-:3];
					dcsr_d[11] = 1'b0;
					dcsr_d[3] = 1'b0;
					dcsr_d[4] = 1'b0;
					dcsr_d[10] = 1'b0;
					dcsr_d[9] = 1'b0;
					dcsr_d[5] = 1'b0;
					dcsr_d[14] = 1'b0;
					dcsr_d[27-:12] = 12'h000;
					dcsr_en = 1'b1;
				end
				12'h7b1: depc_en = 1'b1;
				12'h7b2: dscratch0_en = 1'b1;
				12'h7b3: dscratch1_en = 1'b1;
				12'h320: mcountinhibit_we = 1'b1;
				12'hb00, 12'hb02, 12'hb03, 12'hb04, 12'hb05, 12'hb06, 12'hb07, 12'hb08, 12'hb09, 12'hb0a, 12'hb0b, 12'hb0c, 12'hb0d, 12'hb0e, 12'hb0f, 12'hb10, 12'hb11, 12'hb12, 12'hb13, 12'hb14, 12'hb15, 12'hb16, 12'hb17, 12'hb18, 12'hb19, 12'hb1a, 12'hb1b, 12'hb1c, 12'hb1d, 12'hb1e, 12'hb1f: mhpmcounter_we[mhpmcounter_idx] = 1'b1;
				12'hb80, 12'hb82, 12'hb83, 12'hb84, 12'hb85, 12'hb86, 12'hb87, 12'hb88, 12'hb89, 12'hb8a, 12'hb8b, 12'hb8c, 12'hb8d, 12'hb8e, 12'hb8f, 12'hb90, 12'hb91, 12'hb92, 12'hb93, 12'hb94, 12'hb95, 12'hb96, 12'hb97, 12'hb98, 12'hb99, 12'hb9a, 12'hb9b, 12'hb9c, 12'hb9d, 12'hb9e, 12'hb9f: mhpmcounterh_we[mhpmcounter_idx] = 1'b1;
				12'h7c0: begin
					cpuctrlsts_part_d = cpuctrlsts_part_wdata;
					cpuctrlsts_part_we = 1'b1;
				end
				default:
					;
			endcase
		case (1'b1)
			csr_save_cause_i: begin
				case (1'b1)
					csr_save_if_i: exception_pc = pc_if_i;
					csr_save_id_i: exception_pc = pc_id_i;
					csr_save_wb_i: exception_pc = pc_wb_i;
					default:
						;
				endcase
				priv_lvl_d = 2'b11;
				if (debug_csr_save_i) begin
					dcsr_d[1-:2] = priv_lvl_q;
					dcsr_d[8-:3] = debug_cause_i;
					dcsr_en = 1'b1;
					depc_d = exception_pc;
					depc_en = 1'b1;
				end
				else if (!debug_mode_i) begin
					mtval_en = 1'b1;
					mtval_d = csr_mtval_i;
					mstatus_en = 1'b1;
					mstatus_d[5] = 1'b0;
					mstatus_d[4] = mstatus_q[5];
					mstatus_d[3-:2] = priv_lvl_q;
					mepc_en = 1'b1;
					mepc_d = exception_pc;
					mcause_en = 1'b1;
					mcause_d = csr_mcause_i;
					mstack_en = 1'b1;
					if (!(mcause_d[5] || mcause_d[6])) begin
						cpuctrlsts_part_we = 1'b1;
						cpuctrlsts_part_d[6] = 1'b1;
						if (cpuctrlsts_part_q[6]) begin
							double_fault_seen_o = 1'b1;
							cpuctrlsts_part_d[7] = 1'b1;
						end
					end
				end
			end
			csr_restore_dret_i: priv_lvl_d = dcsr_q[1-:2];
			csr_restore_mret_i: begin
				priv_lvl_d = mstatus_q[3-:2];
				mstatus_en = 1'b1;
				mstatus_d[5] = mstatus_q[4];
				if (mstatus_q[3-:2] != 2'b11)
					mstatus_d[1] = 1'b0;
				cpuctrlsts_part_we = 1'b1;
				cpuctrlsts_part_d[6] = 1'b0;
				if (nmi_mode_i) begin
					mstatus_d[4] = mstack_q[2];
					mstatus_d[3-:2] = mstack_q[1-:2];
					mepc_en = 1'b1;
					mepc_d = mstack_epc_q;
					mcause_en = 1'b1;
					mcause_d = mstack_cause_q;
				end
				else begin
					mstatus_d[4] = 1'b1;
					mstatus_d[3-:2] = 2'b00;
				end
			end
			default:
				;
		endcase
	end
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			priv_lvl_q <= 2'b11;
		else
			priv_lvl_q <= priv_lvl_d;
	assign priv_mode_id_o = priv_lvl_q;
	assign priv_mode_lsu_o = (mstatus_q[1] ? mstatus_q[3-:2] : priv_lvl_q);
	always @(*)
		case (csr_op_i)
			2'd1: csr_wdata_int = csr_wdata_i;
			2'd2: csr_wdata_int = csr_wdata_i | csr_rdata_o;
			2'd3: csr_wdata_int = ~csr_wdata_i & csr_rdata_o;
			2'd0: csr_wdata_int = csr_wdata_i;
			default: csr_wdata_int = csr_wdata_i;
		endcase
	assign csr_wr = |{csr_op_i == 2'd1, csr_op_i == 2'd2, csr_op_i == 2'd3};
	assign csr_we_int = (csr_wr & csr_op_en_i) & ~illegal_csr_insn_o;
	assign csr_rdata_o = csr_rdata_int;
	assign csr_mepc_o = mepc_q;
	assign csr_depc_o = depc_q;
	assign csr_mtvec_o = mtvec_q;
	assign csr_mtval_o = mtval_q;
	assign csr_mstatus_mie_o = mstatus_q[5];
	assign csr_mstatus_tw_o = mstatus_q[0];
	assign debug_single_step_o = dcsr_q[2];
	assign debug_ebreakm_o = dcsr_q[15];
	assign debug_ebreaku_o = dcsr_q[12];
	assign irqs_o = mip & mie_q;
	assign irq_pending_o = |irqs_o;
	localparam [5:0] MSTATUS_RST_VAL = 6'b010000;
	ibex_csr #(
		.Width(6),
		.ShadowCopy(ShadowCSR),
		.ResetValue({MSTATUS_RST_VAL})
	) u_mstatus_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i({mstatus_d}),
		.wr_en_i(mstatus_en),
		.rd_data_o(mstatus_q),
		.rd_error_o(mstatus_err)
	);
	ibex_csr #(
		.Width(32),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_mepc_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(mepc_d),
		.wr_en_i(mepc_en),
		.rd_data_o(mepc_q)
	);
	assign mie_d[17] = csr_wdata_int[ibex_pkg_CSR_MSIX_BIT];
	assign mie_d[16] = csr_wdata_int[ibex_pkg_CSR_MTIX_BIT];
	assign mie_d[15] = csr_wdata_int[ibex_pkg_CSR_MEIX_BIT];
	assign mie_d[14-:15] = csr_wdata_int[ibex_pkg_CSR_MFIX_BIT_HIGH:ibex_pkg_CSR_MFIX_BIT_LOW];
	ibex_csr #(
		.Width(18),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_mie_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i({mie_d}),
		.wr_en_i(mie_en),
		.rd_data_o(mie_q)
	);
	ibex_csr #(
		.Width(32),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_mscratch_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(csr_wdata_int),
		.wr_en_i(mscratch_en),
		.rd_data_o(mscratch_q)
	);
	ibex_csr #(
		.Width(7),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_mcause_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i({mcause_d}),
		.wr_en_i(mcause_en),
		.rd_data_o(mcause_q)
	);
	ibex_csr #(
		.Width(32),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_mtval_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(mtval_d),
		.wr_en_i(mtval_en),
		.rd_data_o(mtval_q)
	);
	ibex_csr #(
		.Width(32),
		.ShadowCopy(ShadowCSR),
		.ResetValue(32'd1)
	) u_mtvec_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(mtvec_d),
		.wr_en_i(mtvec_en),
		.rd_data_o(mtvec_q),
		.rd_error_o(mtvec_err)
	);
	localparam [31:0] DCSR_RESET_VAL = 32'b01000000000000000000000000000011;
	ibex_csr #(
		.Width(32),
		.ShadowCopy(1'b0),
		.ResetValue({DCSR_RESET_VAL})
	) u_dcsr_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i({dcsr_d}),
		.wr_en_i(dcsr_en),
		.rd_data_o(dcsr_q)
	);
	ibex_csr #(
		.Width(32),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_depc_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(depc_d),
		.wr_en_i(depc_en),
		.rd_data_o(depc_q)
	);
	ibex_csr #(
		.Width(32),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_dscratch0_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(csr_wdata_int),
		.wr_en_i(dscratch0_en),
		.rd_data_o(dscratch0_q)
	);
	ibex_csr #(
		.Width(32),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_dscratch1_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(csr_wdata_int),
		.wr_en_i(dscratch1_en),
		.rd_data_o(dscratch1_q)
	);
	localparam [2:0] MSTACK_RESET_VAL = 3'b100;
	ibex_csr #(
		.Width(3),
		.ShadowCopy(1'b0),
		.ResetValue({MSTACK_RESET_VAL})
	) u_mstack_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i({mstack_d}),
		.wr_en_i(mstack_en),
		.rd_data_o(mstack_q)
	);
	ibex_csr #(
		.Width(32),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_mstack_epc_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(mstack_epc_d),
		.wr_en_i(mstack_en),
		.rd_data_o(mstack_epc_q)
	);
	ibex_csr #(
		.Width(7),
		.ShadowCopy(1'b0),
		.ResetValue(1'sb0)
	) u_mstack_cause_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i(mstack_cause_d),
		.wr_en_i(mstack_en),
		.rd_data_o(mstack_cause_q)
	);
	localparam [11:0] ibex_pkg_CSR_OFF_PMP_ADDR = 12'h3b0;
	localparam [11:0] ibex_pkg_CSR_OFF_PMP_CFG = 12'h3a0;
	generate
		if (PMPEnable) begin : g_pmp_registers
			localparam [95:0] pmp_cfg_rst = 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			localparam [543:0] pmp_addr_rst = 544'h0;
			localparam [2:0] pmp_mseccfg_rst = 3'b000;
			wire [2:0] pmp_mseccfg_q;
			wire [2:0] pmp_mseccfg_d;
			wire pmp_mseccfg_we;
			wire pmp_mseccfg_err;
			wire [5:0] pmp_cfg [0:PMPNumRegions - 1];
			wire [PMPNumRegions - 1:0] pmp_cfg_locked;
			wire [PMPNumRegions - 1:0] pmp_cfg_wr_suppress;
			reg [5:0] pmp_cfg_wdata [0:PMPNumRegions - 1];
			wire [PMPAddrWidth - 1:0] pmp_addr [0:PMPNumRegions - 1];
			wire [PMPNumRegions - 1:0] pmp_cfg_we;
			wire [PMPNumRegions - 1:0] pmp_cfg_err;
			wire [PMPNumRegions - 1:0] pmp_addr_we;
			wire [PMPNumRegions - 1:0] pmp_addr_err;
			wire any_pmp_entry_locked;
			genvar i;
			for (i = 0; i < ibex_pkg_PMP_MAX_REGIONS; i = i + 1) begin : g_exp_rd_data
				if (i < PMPNumRegions) begin : g_implemented_regions
					assign pmp_cfg_rdata[i] = {pmp_cfg[i][5], 2'b00, pmp_cfg[i][4-:2], pmp_cfg[i][2], pmp_cfg[i][1], pmp_cfg[i][0]};
					if (PMPGranularity == 0) begin : g_pmp_g0
						wire [32:1] sv2v_tmp_646D9;
						assign sv2v_tmp_646D9 = pmp_addr[i];
						always @(*) pmp_addr_rdata[i] = sv2v_tmp_646D9;
					end
					else if (PMPGranularity == 1) begin : g_pmp_g1
						always @(*) begin
							pmp_addr_rdata[i] = pmp_addr[i];
							if ((pmp_cfg[i][4-:2] == 2'b00) || (pmp_cfg[i][4-:2] == 2'b01))
								pmp_addr_rdata[i][PMPGranularity - 1:0] = 1'sb0;
						end
					end
					else begin : g_pmp_g2
						always @(*) begin
							pmp_addr_rdata[i] = {pmp_addr[i], {PMPGranularity - 1 {1'b1}}};
							if ((pmp_cfg[i][4-:2] == 2'b00) || (pmp_cfg[i][4-:2] == 2'b01))
								pmp_addr_rdata[i][PMPGranularity - 1:0] = 1'sb0;
						end
					end
				end
				else begin : g_other_regions
					assign pmp_cfg_rdata[i] = 1'sb0;
					wire [32:1] sv2v_tmp_96282;
					assign sv2v_tmp_96282 = 1'sb0;
					always @(*) pmp_addr_rdata[i] = sv2v_tmp_96282;
				end
			end
			for (i = 0; i < PMPNumRegions; i = i + 1) begin : g_pmp_csrs
				assign pmp_cfg_we[i] = ((csr_we_int & ~pmp_cfg_locked[i]) & ~pmp_cfg_wr_suppress[i]) & (csr_addr == (ibex_pkg_CSR_OFF_PMP_CFG + (i[11:0] >> 2)));
				wire [1:1] sv2v_tmp_43D04;
				assign sv2v_tmp_43D04 = csr_wdata_int[((i % 4) * ibex_pkg_PMP_CFG_W) + 7];
				always @(*) pmp_cfg_wdata[i][5] = sv2v_tmp_43D04;
				always @(*)
					case (csr_wdata_int[((i % 4) * ibex_pkg_PMP_CFG_W) + 3+:2])
						2'b00: pmp_cfg_wdata[i][4-:2] = 2'b00;
						2'b01: pmp_cfg_wdata[i][4-:2] = 2'b01;
						2'b10: pmp_cfg_wdata[i][4-:2] = (PMPGranularity == 0 ? 2'b10 : 2'b00);
						2'b11: pmp_cfg_wdata[i][4-:2] = 2'b11;
						default: pmp_cfg_wdata[i][4-:2] = 2'b00;
					endcase
				wire [1:1] sv2v_tmp_B5F8A;
				assign sv2v_tmp_B5F8A = csr_wdata_int[((i % 4) * ibex_pkg_PMP_CFG_W) + 2];
				always @(*) pmp_cfg_wdata[i][2] = sv2v_tmp_B5F8A;
				wire [1:1] sv2v_tmp_DA81D;
				assign sv2v_tmp_DA81D = (pmp_mseccfg_q[0] ? csr_wdata_int[((i % 4) * ibex_pkg_PMP_CFG_W) + 1] : &csr_wdata_int[(i % 4) * ibex_pkg_PMP_CFG_W+:2]);
				always @(*) pmp_cfg_wdata[i][1] = sv2v_tmp_DA81D;
				wire [1:1] sv2v_tmp_92290;
				assign sv2v_tmp_92290 = csr_wdata_int[(i % 4) * ibex_pkg_PMP_CFG_W];
				always @(*) pmp_cfg_wdata[i][0] = sv2v_tmp_92290;
				ibex_csr #(
					.Width(6),
					.ShadowCopy(ShadowCSR),
					.ResetValue(pmp_cfg_rst[(15 - i) * 6+:6])
				) u_pmp_cfg_csr(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.wr_data_i({pmp_cfg_wdata[i]}),
					.wr_en_i(pmp_cfg_we[i]),
					.rd_data_o(pmp_cfg[i]),
					.rd_error_o(pmp_cfg_err[i])
				);
				assign pmp_cfg_locked[i] = pmp_cfg[i][5] & ~pmp_mseccfg_q[2];
				assign pmp_cfg_wr_suppress[i] = (pmp_mseccfg_q[0] & ~pmp_mseccfg[2]) & is_mml_m_exec_cfg(pmp_cfg_wdata[i]);
				if (i < (PMPNumRegions - 1)) begin : g_lower
					assign pmp_addr_we[i] = ((csr_we_int & ~pmp_cfg_locked[i]) & (~pmp_cfg_locked[i + 1] | (pmp_cfg[i + 1][4-:2] != 2'b01))) & (csr_addr == (ibex_pkg_CSR_OFF_PMP_ADDR + i[11:0]));
				end
				else begin : g_upper
					assign pmp_addr_we[i] = (csr_we_int & ~pmp_cfg_locked[i]) & (csr_addr == (ibex_pkg_CSR_OFF_PMP_ADDR + i[11:0]));
				end
				ibex_csr #(
					.Width(PMPAddrWidth),
					.ShadowCopy(ShadowCSR),
					.ResetValue(pmp_addr_rst[((15 - i) * 34) + 33-:PMPAddrWidth])
				) u_pmp_addr_csr(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.wr_data_i(csr_wdata_int[31-:PMPAddrWidth]),
					.wr_en_i(pmp_addr_we[i]),
					.rd_data_o(pmp_addr[i]),
					.rd_error_o(pmp_addr_err[i])
				);
				assign csr_pmp_cfg_o[((PMPNumRegions - 1) - i) * 6+:6] = pmp_cfg[i];
				assign csr_pmp_addr_o[((PMPNumRegions - 1) - i) * 34+:34] = {pmp_addr_rdata[i], 2'b00};
			end
			assign pmp_mseccfg_we = csr_we_int & (csr_addr == 12'h747);
			assign pmp_mseccfg_d[0] = (pmp_mseccfg_q[0] ? 1'b1 : csr_wdata_int[ibex_pkg_CSR_MSECCFG_MML_BIT]);
			assign pmp_mseccfg_d[1] = (pmp_mseccfg_q[1] ? 1'b1 : csr_wdata_int[ibex_pkg_CSR_MSECCFG_MMWP_BIT]);
			assign any_pmp_entry_locked = |pmp_cfg_locked;
			assign pmp_mseccfg_d[2] = (any_pmp_entry_locked ? 1'b0 : csr_wdata_int[ibex_pkg_CSR_MSECCFG_RLB_BIT]);
			ibex_csr #(
				.Width(3),
				.ShadowCopy(ShadowCSR),
				.ResetValue(pmp_mseccfg_rst)
			) u_pmp_mseccfg(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.wr_data_i(pmp_mseccfg_d),
				.wr_en_i(pmp_mseccfg_we),
				.rd_data_o(pmp_mseccfg_q),
				.rd_error_o(pmp_mseccfg_err)
			);
			assign pmp_csr_err = (|pmp_cfg_err | |pmp_addr_err) | pmp_mseccfg_err;
			assign pmp_mseccfg = pmp_mseccfg_q;
		end
		else begin : g_no_pmp_tieoffs
			genvar i;
			for (i = 0; i < ibex_pkg_PMP_MAX_REGIONS; i = i + 1) begin : g_rdata
				wire [32:1] sv2v_tmp_96282;
				assign sv2v_tmp_96282 = 1'sb0;
				always @(*) pmp_addr_rdata[i] = sv2v_tmp_96282;
				assign pmp_cfg_rdata[i] = 1'sb0;
			end
			for (i = 0; i < PMPNumRegions; i = i + 1) begin : g_outputs
				assign csr_pmp_cfg_o[((PMPNumRegions - 1) - i) * 6+:6] = 6'b000000;
				assign csr_pmp_addr_o[((PMPNumRegions - 1) - i) * 34+:34] = 1'sb0;
			end
			assign pmp_csr_err = 1'b0;
			assign pmp_mseccfg = 1'sb0;
		end
	endgenerate
	assign csr_pmp_mseccfg_o = pmp_mseccfg;
	always @(*) begin : mcountinhibit_update
		if (mcountinhibit_we == 1'b1)
			mcountinhibit_d = {csr_wdata_int[MHPMCounterNum + 2:2], 1'b0, csr_wdata_int[0]};
		else
			mcountinhibit_d = mcountinhibit_q;
	end
	always @(*) begin : gen_mhpmcounter_incr
		begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < 32; i = i + 1)
				begin : gen_mhpmcounter_incr_inactive
					mhpmcounter_incr[i] = 1'b0;
				end
		end
		mhpmcounter_incr[0] = 1'b1;
		mhpmcounter_incr[1] = 1'b0;
		mhpmcounter_incr[2] = instr_ret_i;
		mhpmcounter_incr[3] = dside_wait_i;
		mhpmcounter_incr[4] = iside_wait_i;
		mhpmcounter_incr[5] = mem_load_i;
		mhpmcounter_incr[6] = mem_store_i;
		mhpmcounter_incr[7] = jump_i;
		mhpmcounter_incr[8] = branch_i;
		mhpmcounter_incr[9] = branch_taken_i;
		mhpmcounter_incr[10] = instr_ret_compressed_i;
		mhpmcounter_incr[11] = mul_wait_i;
		mhpmcounter_incr[12] = div_wait_i;
	end
	always @(*) begin : gen_mhpmevent
		begin : sv2v_autoblock_2
			reg signed [31:0] i;
			for (i = 0; i < 32; i = i + 1)
				begin : gen_mhpmevent_active
					mhpmevent[i] = 1'sb0;
					if (i >= 3)
						mhpmevent[i][i - 3] = 1'b1;
				end
		end
		mhpmevent[1] = 1'sb0;
		begin : sv2v_autoblock_3
			reg [31:0] i;
			for (i = 3 + MHPMCounterNum; i < 32; i = i + 1)
				begin : gen_mhpmevent_inactive
					mhpmevent[i] = 1'sb0;
				end
		end
	end
	ibex_counter #(.CounterWidth(64)) mcycle_counter_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.counter_inc_i(mhpmcounter_incr[0] & ~mcountinhibit[0]),
		.counterh_we_i(mhpmcounterh_we[0]),
		.counter_we_i(mhpmcounter_we[0]),
		.counter_val_i(csr_wdata_int),
		.counter_val_o(mhpmcounter[0])
	);
	ibex_counter #(
		.CounterWidth(64),
		.ProvideValUpd(1)
	) minstret_counter_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.counter_inc_i(mhpmcounter_incr[2] & ~mcountinhibit[2]),
		.counterh_we_i(mhpmcounterh_we[2]),
		.counter_we_i(mhpmcounter_we[2]),
		.counter_val_i(csr_wdata_int),
		.counter_val_o(minstret_raw),
		.counter_val_upd_o(minstret_next)
	);
	assign mhpmcounter[2] = (instr_ret_spec_i & ~mcountinhibit[2] ? minstret_next : minstret_raw);
	assign mhpmcounter[1] = 1'sb0;
	assign unused_mhpmcounter_we_1 = mhpmcounter_we[1];
	assign unused_mhpmcounterh_we_1 = mhpmcounterh_we[1];
	assign unused_mhpmcounter_incr_1 = mhpmcounter_incr[1];
	genvar i;
	generate
		for (i = 0; i < 29; i = i + 1) begin : gen_cntrs
			localparam signed [31:0] Cnt = i + 3;
			if (i < MHPMCounterNum) begin : gen_imp
				wire [63:0] mhpmcounter_raw;
				wire [63:0] mhpmcounter_next;
				ibex_counter #(
					.CounterWidth(MHPMCounterWidth),
					.ProvideValUpd(Cnt == 10)
				) mcounters_variable_i(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.counter_inc_i(mhpmcounter_incr[Cnt] & ~mcountinhibit[Cnt]),
					.counterh_we_i(mhpmcounterh_we[Cnt]),
					.counter_we_i(mhpmcounter_we[Cnt]),
					.counter_val_i(csr_wdata_int),
					.counter_val_o(mhpmcounter_raw),
					.counter_val_upd_o(mhpmcounter_next)
				);
				if (Cnt == 10) begin : gen_compressed_instr_cnt
					assign mhpmcounter[Cnt] = (instr_ret_compressed_spec_i & ~mcountinhibit[Cnt] ? mhpmcounter_next : mhpmcounter_raw);
				end
				else begin : gen_other_cnts
					wire [63:0] unused_mhpmcounter_next;
					assign mhpmcounter[Cnt] = mhpmcounter_raw;
					assign unused_mhpmcounter_next = mhpmcounter_next;
				end
			end
			else begin : gen_unimp
				assign mhpmcounter[Cnt] = 1'sb0;
				if (Cnt == 10) begin : gen_no_compressed_instr_cnt
					wire unused_instr_ret_compressed_spec_i;
					assign unused_instr_ret_compressed_spec_i = instr_ret_compressed_spec_i;
				end
			end
		end
		if (MHPMCounterNum < 29) begin : g_mcountinhibit_reduced
			wire [(29 - MHPMCounterNum) - 1:0] unused_mhphcounter_we;
			wire [(29 - MHPMCounterNum) - 1:0] unused_mhphcounterh_we;
			wire [(29 - MHPMCounterNum) - 1:0] unused_mhphcounter_incr;
			assign mcountinhibit = {{29 - MHPMCounterNum {1'b0}}, mcountinhibit_q};
			assign unused_mhphcounter_we = mhpmcounter_we[31:MHPMCounterNum + 3];
			assign unused_mhphcounterh_we = mhpmcounterh_we[31:MHPMCounterNum + 3];
			assign unused_mhphcounter_incr = mhpmcounter_incr[31:MHPMCounterNum + 3];
		end
		else begin : g_mcountinhibit_full
			assign mcountinhibit = mcountinhibit_q;
		end
	endgenerate
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			mcountinhibit_q <= 1'sb0;
		else
			mcountinhibit_q <= mcountinhibit_d;
	generate
		if (DbgTriggerEn) begin : gen_trigger_regs
			localparam [31:0] DbgHwNumLen = (DbgHwBreakNum > 1 ? $clog2(DbgHwBreakNum) : 1);
			localparam [31:0] MaxTselect = DbgHwBreakNum - 1;
			wire [DbgHwNumLen - 1:0] tselect_d;
			wire [DbgHwNumLen - 1:0] tselect_q;
			wire tmatch_control_d;
			wire [DbgHwBreakNum - 1:0] tmatch_control_q;
			wire [31:0] tmatch_value_d;
			wire [31:0] tmatch_value_q [0:DbgHwBreakNum - 1];
			wire selected_tmatch_control;
			wire [31:0] selected_tmatch_value;
			wire tselect_we;
			wire [DbgHwBreakNum - 1:0] tmatch_control_we;
			wire [DbgHwBreakNum - 1:0] tmatch_value_we;
			wire [DbgHwBreakNum - 1:0] trigger_match;
			assign tselect_we = (csr_we_int & debug_mode_i) & (csr_addr_i == 12'h7a0);
			genvar i;
			for (i = 0; i < DbgHwBreakNum; i = i + 1) begin : g_dbg_tmatch_we
				assign tmatch_control_we[i] = (((i[DbgHwNumLen - 1:0] == tselect_q) & csr_we_int) & debug_mode_i) & (csr_addr_i == 12'h7a1);
				assign tmatch_value_we[i] = (((i[DbgHwNumLen - 1:0] == tselect_q) & csr_we_int) & debug_mode_i) & (csr_addr_i == 12'h7a2);
			end
			assign tselect_d = (csr_wdata_int < DbgHwBreakNum ? csr_wdata_int[DbgHwNumLen - 1:0] : MaxTselect[DbgHwNumLen - 1:0]);
			assign tmatch_control_d = csr_wdata_int[2];
			assign tmatch_value_d = csr_wdata_int[31:0];
			ibex_csr #(
				.Width(DbgHwNumLen),
				.ShadowCopy(1'b0),
				.ResetValue(1'sb0)
			) u_tselect_csr(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.wr_data_i(tselect_d),
				.wr_en_i(tselect_we),
				.rd_data_o(tselect_q)
			);
			for (i = 0; i < DbgHwBreakNum; i = i + 1) begin : g_dbg_tmatch_reg
				ibex_csr #(
					.Width(1),
					.ShadowCopy(1'b0),
					.ResetValue(1'sb0)
				) u_tmatch_control_csr(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.wr_data_i(tmatch_control_d),
					.wr_en_i(tmatch_control_we[i]),
					.rd_data_o(tmatch_control_q[i])
				);
				ibex_csr #(
					.Width(32),
					.ShadowCopy(1'b0),
					.ResetValue(1'sb0)
				) u_tmatch_value_csr(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.wr_data_i(tmatch_value_d),
					.wr_en_i(tmatch_value_we[i]),
					.rd_data_o(tmatch_value_q[i])
				);
			end
			localparam [31:0] TSelectRdataPadlen = (DbgHwNumLen >= 32 ? 0 : 32 - DbgHwNumLen);
			assign tselect_rdata = {{TSelectRdataPadlen {1'b0}}, tselect_q};
			if (DbgHwBreakNum > 1) begin : g_dbg_tmatch_multiple_select
				assign selected_tmatch_control = tmatch_control_q[tselect_q];
				assign selected_tmatch_value = tmatch_value_q[tselect_q];
			end
			else begin : g_dbg_tmatch_single_select
				assign selected_tmatch_control = tmatch_control_q[0];
				assign selected_tmatch_value = tmatch_value_q[0];
			end
			assign tmatch_control_rdata = {29'b00101000000000000001000001001, selected_tmatch_control, 1'b0, 1'b0};
			assign tmatch_value_rdata = selected_tmatch_value;
			for (i = 0; i < DbgHwBreakNum; i = i + 1) begin : g_dbg_trigger_match
				assign trigger_match[i] = tmatch_control_q[i] & (pc_if_i[31:0] == tmatch_value_q[i]);
			end
			assign trigger_match_o = |trigger_match;
		end
		else begin : gen_no_trigger_regs
			assign tselect_rdata = 'b0;
			assign tmatch_control_rdata = 'b0;
			assign tmatch_value_rdata = 'b0;
			assign trigger_match_o = 'b0;
		end
	endgenerate
	assign cpuctrlsts_part_wdata_raw = csr_wdata_int[7:0];
	generate
		if (DataIndTiming) begin : gen_dit
			assign cpuctrlsts_part_wdata[1] = cpuctrlsts_part_wdata_raw[1];
		end
		else begin : gen_no_dit
			wire unused_dit;
			assign unused_dit = cpuctrlsts_part_wdata_raw[1];
			assign cpuctrlsts_part_wdata[1] = 1'b0;
		end
	endgenerate
	assign data_ind_timing_o = cpuctrlsts_part_q[1];
	generate
		if (DummyInstructions) begin : gen_dummy
			assign cpuctrlsts_part_wdata[2] = cpuctrlsts_part_wdata_raw[2];
			assign cpuctrlsts_part_wdata[5-:3] = cpuctrlsts_part_wdata_raw[5-:3];
			assign dummy_instr_seed_en_o = csr_we_int && (csr_addr == 12'h7c1);
			assign dummy_instr_seed_o = csr_wdata_int;
		end
		else begin : gen_no_dummy
			wire unused_dummy_en;
			wire [2:0] unused_dummy_mask;
			assign unused_dummy_en = cpuctrlsts_part_wdata_raw[2];
			assign unused_dummy_mask = cpuctrlsts_part_wdata_raw[5-:3];
			assign cpuctrlsts_part_wdata[2] = 1'b0;
			assign cpuctrlsts_part_wdata[5-:3] = 3'b000;
			assign dummy_instr_seed_en_o = 1'b0;
			assign dummy_instr_seed_o = 1'sb0;
		end
	endgenerate
	assign dummy_instr_en_o = cpuctrlsts_part_q[2];
	assign dummy_instr_mask_o = cpuctrlsts_part_q[5-:3];
	generate
		if (ICache) begin : gen_icache_enable
			assign cpuctrlsts_part_wdata[0] = cpuctrlsts_part_wdata_raw[0];
			ibex_csr #(
				.Width(1),
				.ShadowCopy(ShadowCSR),
				.ResetValue(1'b0)
			) u_cpuctrlsts_ic_scr_key_valid_q_csr(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.wr_data_i(ic_scr_key_valid_i),
				.wr_en_i(1'b1),
				.rd_data_o(cpuctrlsts_ic_scr_key_valid_q),
				.rd_error_o(cpuctrlsts_ic_scr_key_err)
			);
		end
		else begin : gen_no_icache
			wire unused_icen;
			assign unused_icen = cpuctrlsts_part_wdata_raw[0];
			assign cpuctrlsts_part_wdata[0] = 1'b0;
			wire unused_ic_scr_key_valid;
			assign unused_ic_scr_key_valid = ic_scr_key_valid_i;
			assign cpuctrlsts_ic_scr_key_valid_q = 1'b0;
			assign cpuctrlsts_ic_scr_key_err = 1'b0;
		end
	endgenerate
	assign cpuctrlsts_part_wdata[7] = cpuctrlsts_part_wdata_raw[7];
	assign cpuctrlsts_part_wdata[6] = cpuctrlsts_part_wdata_raw[6];
	assign icache_enable_o = cpuctrlsts_part_q[0] & ~(debug_mode_i | debug_mode_entering_i);
	ibex_csr #(
		.Width(8),
		.ShadowCopy(ShadowCSR),
		.ResetValue(1'sb0)
	) u_cpuctrlsts_part_csr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.wr_data_i({cpuctrlsts_part_d}),
		.wr_en_i(cpuctrlsts_part_we),
		.rd_data_o(cpuctrlsts_part_q),
		.rd_error_o(cpuctrlsts_part_err)
	);
	assign csr_shadow_err_o = (((mstatus_err | mtvec_err) | pmp_csr_err) | cpuctrlsts_part_err) | cpuctrlsts_ic_scr_key_err;
endmodule
module ibex_csr (
	clk_i,
	rst_ni,
	wr_data_i,
	wr_en_i,
	rd_data_o,
	rd_error_o
);
	parameter [31:0] Width = 32;
	parameter [0:0] ShadowCopy = 1'b0;
	parameter [Width - 1:0] ResetValue = 1'sb0;
	input wire clk_i;
	input wire rst_ni;
	input wire [Width - 1:0] wr_data_i;
	input wire wr_en_i;
	output wire [Width - 1:0] rd_data_o;
	output wire rd_error_o;
	reg [Width - 1:0] rdata_q;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			rdata_q <= ResetValue;
		else if (wr_en_i)
			rdata_q <= wr_data_i;
	assign rd_data_o = rdata_q;
	generate
		if (ShadowCopy) begin : gen_shadow
			reg [Width - 1:0] shadow_q;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					shadow_q <= ~ResetValue;
				else if (wr_en_i)
					shadow_q <= ~wr_data_i;
			assign rd_error_o = rdata_q != ~shadow_q;
		end
		else begin : gen_no_shadow
			assign rd_error_o = 1'b0;
		end
	endgenerate
endmodule
module ibex_decoder (
	clk_i,
	rst_ni,
	illegal_insn_o,
	ebrk_insn_o,
	mret_insn_o,
	dret_insn_o,
	ecall_insn_o,
	wfi_insn_o,
	jump_set_o,
	branch_taken_i,
	icache_inval_o,
	instr_first_cycle_i,
	instr_rdata_i,
	instr_rdata_alu_i,
	illegal_c_insn_i,
	imm_a_mux_sel_o,
	imm_b_mux_sel_o,
	bt_a_mux_sel_o,
	bt_b_mux_sel_o,
	imm_i_type_o,
	imm_s_type_o,
	imm_b_type_o,
	imm_u_type_o,
	imm_j_type_o,
	zimm_rs1_type_o,
	rf_wdata_sel_o,
	rf_we_o,
	rf_raddr_a_o,
	rf_raddr_b_o,
	rf_waddr_o,
	rf_ren_a_o,
	rf_ren_b_o,
	alu_operator_o,
	alu_op_a_mux_sel_o,
	alu_op_b_mux_sel_o,
	alu_multicycle_o,
	mult_en_o,
	div_en_o,
	mult_sel_o,
	div_sel_o,
	multdiv_operator_o,
	multdiv_signed_mode_o,
	csr_access_o,
	csr_op_o,
	data_req_o,
	data_we_o,
	data_type_o,
	data_sign_extension_o,
	jump_in_dec_o,
	branch_in_dec_o
);
	parameter [0:0] RV32E = 0;
	parameter integer RV32M = 32'sd2;
	parameter integer RV32B = 32'sd0;
	parameter [0:0] BranchTargetALU = 0;
	input wire clk_i;
	input wire rst_ni;
	output wire illegal_insn_o;
	output reg ebrk_insn_o;
	output reg mret_insn_o;
	output reg dret_insn_o;
	output reg ecall_insn_o;
	output reg wfi_insn_o;
	output reg jump_set_o;
	input wire branch_taken_i;
	output reg icache_inval_o;
	input wire instr_first_cycle_i;
	input wire [31:0] instr_rdata_i;
	input wire [31:0] instr_rdata_alu_i;
	input wire illegal_c_insn_i;
	output reg imm_a_mux_sel_o;
	output reg [2:0] imm_b_mux_sel_o;
	output reg [1:0] bt_a_mux_sel_o;
	output reg [2:0] bt_b_mux_sel_o;
	output wire [31:0] imm_i_type_o;
	output wire [31:0] imm_s_type_o;
	output wire [31:0] imm_b_type_o;
	output wire [31:0] imm_u_type_o;
	output wire [31:0] imm_j_type_o;
	output wire [31:0] zimm_rs1_type_o;
	output reg rf_wdata_sel_o;
	output wire rf_we_o;
	output wire [4:0] rf_raddr_a_o;
	output wire [4:0] rf_raddr_b_o;
	output wire [4:0] rf_waddr_o;
	output reg rf_ren_a_o;
	output reg rf_ren_b_o;
	output reg [6:0] alu_operator_o;
	output reg [1:0] alu_op_a_mux_sel_o;
	output reg alu_op_b_mux_sel_o;
	output reg alu_multicycle_o;
	output wire mult_en_o;
	output wire div_en_o;
	output reg mult_sel_o;
	output reg div_sel_o;
	output reg [1:0] multdiv_operator_o;
	output reg [1:0] multdiv_signed_mode_o;
	output reg csr_access_o;
	output reg [1:0] csr_op_o;
	output reg data_req_o;
	output reg data_we_o;
	output reg [1:0] data_type_o;
	output reg data_sign_extension_o;
	output reg jump_in_dec_o;
	output reg branch_in_dec_o;
	reg illegal_insn;
	wire illegal_reg_rv32e;
	reg csr_illegal;
	reg rf_we;
	wire [31:0] instr;
	wire [31:0] instr_alu;
	wire [9:0] unused_instr_alu;
	wire [4:0] instr_rs1;
	wire [4:0] instr_rs2;
	wire [4:0] instr_rs3;
	wire [4:0] instr_rd;
	reg use_rs3_d;
	reg use_rs3_q;
	reg [1:0] csr_op;
	reg [6:0] opcode;
	reg [6:0] opcode_alu;
	assign instr = instr_rdata_i;
	assign instr_alu = instr_rdata_alu_i;
	assign imm_i_type_o = {{20 {instr[31]}}, instr[31:20]};
	assign imm_s_type_o = {{20 {instr[31]}}, instr[31:25], instr[11:7]};
	assign imm_b_type_o = {{19 {instr[31]}}, instr[31], instr[7], instr[30:25], instr[11:8], 1'b0};
	assign imm_u_type_o = {instr[31:12], 12'b000000000000};
	assign imm_j_type_o = {{12 {instr[31]}}, instr[19:12], instr[20], instr[30:21], 1'b0};
	assign zimm_rs1_type_o = {27'b000000000000000000000000000, instr_rs1};
	generate
		if (RV32B != 32'sd0) begin : gen_rs3_flop
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					use_rs3_q <= 1'b0;
				else
					use_rs3_q <= use_rs3_d;
		end
		else begin : gen_no_rs3_flop
			wire unused_clk;
			wire unused_rst_n;
			assign unused_clk = clk_i;
			assign unused_rst_n = rst_ni;
			wire [1:1] sv2v_tmp_44B6F;
			assign sv2v_tmp_44B6F = use_rs3_d;
			always @(*) use_rs3_q = sv2v_tmp_44B6F;
		end
	endgenerate
	assign instr_rs1 = instr[19:15];
	assign instr_rs2 = instr[24:20];
	assign instr_rs3 = instr[31:27];
	assign rf_raddr_a_o = (use_rs3_q & ~instr_first_cycle_i ? instr_rs3 : instr_rs1);
	assign rf_raddr_b_o = instr_rs2;
	assign instr_rd = instr[11:7];
	assign rf_waddr_o = instr_rd;
	generate
		if (RV32E) begin : gen_rv32e_reg_check_active
			assign illegal_reg_rv32e = ((rf_raddr_a_o[4] & (alu_op_a_mux_sel_o == 2'd0)) | (rf_raddr_b_o[4] & (alu_op_b_mux_sel_o == 1'd0))) | (rf_waddr_o[4] & rf_we);
		end
		else begin : gen_rv32e_reg_check_inactive
			assign illegal_reg_rv32e = 1'b0;
		end
	endgenerate
	always @(*) begin : csr_operand_check
		csr_op_o = csr_op;
		if (((csr_op == 2'd2) || (csr_op == 2'd3)) && (instr_rs1 == {5 {1'sb0}}))
			csr_op_o = 2'd0;
	end
	always @(*) begin
		jump_in_dec_o = 1'b0;
		jump_set_o = 1'b0;
		branch_in_dec_o = 1'b0;
		icache_inval_o = 1'b0;
		multdiv_operator_o = 2'd0;
		multdiv_signed_mode_o = 2'b00;
		rf_wdata_sel_o = 1'd0;
		rf_we = 1'b0;
		rf_ren_a_o = 1'b0;
		rf_ren_b_o = 1'b0;
		csr_access_o = 1'b0;
		csr_illegal = 1'b0;
		csr_op = 2'd0;
		data_we_o = 1'b0;
		data_type_o = 2'b00;
		data_sign_extension_o = 1'b0;
		data_req_o = 1'b0;
		illegal_insn = 1'b0;
		ebrk_insn_o = 1'b0;
		mret_insn_o = 1'b0;
		dret_insn_o = 1'b0;
		ecall_insn_o = 1'b0;
		wfi_insn_o = 1'b0;
		opcode = instr[6:0];
		case (opcode)
			7'h6f: begin
				jump_in_dec_o = 1'b1;
				if (instr_first_cycle_i) begin
					rf_we = BranchTargetALU;
					jump_set_o = 1'b1;
				end
				else
					rf_we = 1'b1;
			end
			7'h67: begin
				jump_in_dec_o = 1'b1;
				if (instr_first_cycle_i) begin
					rf_we = BranchTargetALU;
					jump_set_o = 1'b1;
				end
				else
					rf_we = 1'b1;
				if (instr[14:12] != 3'b000)
					illegal_insn = 1'b1;
				rf_ren_a_o = 1'b1;
			end
			7'h63: begin
				branch_in_dec_o = 1'b1;
				case (instr[14:12])
					3'b000, 3'b001, 3'b100, 3'b101, 3'b110, 3'b111: illegal_insn = 1'b0;
					default: illegal_insn = 1'b1;
				endcase
				rf_ren_a_o = 1'b1;
				rf_ren_b_o = 1'b1;
			end
			7'h23: begin
				rf_ren_a_o = 1'b1;
				rf_ren_b_o = 1'b1;
				data_req_o = 1'b1;
				data_we_o = 1'b1;
				if (instr[14])
					illegal_insn = 1'b1;
				case (instr[13:12])
					2'b00: data_type_o = 2'b10;
					2'b01: data_type_o = 2'b01;
					2'b10: data_type_o = 2'b00;
					default: illegal_insn = 1'b1;
				endcase
			end
			7'h03: begin
				rf_ren_a_o = 1'b1;
				data_req_o = 1'b1;
				data_type_o = 2'b00;
				data_sign_extension_o = ~instr[14];
				case (instr[13:12])
					2'b00: data_type_o = 2'b10;
					2'b01: data_type_o = 2'b01;
					2'b10: begin
						data_type_o = 2'b00;
						if (instr[14])
							illegal_insn = 1'b1;
					end
					default: illegal_insn = 1'b1;
				endcase
			end
			7'h37: rf_we = 1'b1;
			7'h17: rf_we = 1'b1;
			7'h13: begin
				rf_ren_a_o = 1'b1;
				rf_we = 1'b1;
				case (instr[14:12])
					3'b000, 3'b010, 3'b011, 3'b100, 3'b110, 3'b111: illegal_insn = 1'b0;
					3'b001:
						case (instr[31:27])
							5'b00000: illegal_insn = (instr[26:25] == 2'b00 ? 1'b0 : 1'b1);
							5'b00100: illegal_insn = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? 1'b0 : 1'b1);
							5'b01001, 5'b00101, 5'b01101: illegal_insn = (RV32B != 32'sd0 ? 1'b0 : 1'b1);
							5'b00001:
								if (instr[26] == 1'b0)
									illegal_insn = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? 1'b0 : 1'b1);
								else
									illegal_insn = 1'b1;
							5'b01100:
								case (instr[26:20])
									7'b0000000, 7'b0000001, 7'b0000010, 7'b0000100, 7'b0000101: illegal_insn = (RV32B != 32'sd0 ? 1'b0 : 1'b1);
									7'b0010000, 7'b0010001, 7'b0010010, 7'b0011000, 7'b0011001, 7'b0011010: illegal_insn = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? 1'b0 : 1'b1);
									default: illegal_insn = 1'b1;
								endcase
							default: illegal_insn = 1'b1;
						endcase
					3'b101:
						if (instr[26])
							illegal_insn = (RV32B != 32'sd0 ? 1'b0 : 1'b1);
						else
							case (instr[31:27])
								5'b00000, 5'b01000: illegal_insn = (instr[26:25] == 2'b00 ? 1'b0 : 1'b1);
								5'b00100: illegal_insn = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? 1'b0 : 1'b1);
								5'b01100, 5'b01001: illegal_insn = (RV32B != 32'sd0 ? 1'b0 : 1'b1);
								5'b01101:
									if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
										illegal_insn = 1'b0;
									else if (RV32B == 32'sd1)
										illegal_insn = (instr[24:20] == 5'b11000 ? 1'b0 : 1'b1);
									else
										illegal_insn = 1'b1;
								5'b00101:
									if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
										illegal_insn = 1'b0;
									else if (instr[24:20] == 5'b00111)
										illegal_insn = (RV32B == 32'sd1 ? 1'b0 : 1'b1);
									else
										illegal_insn = 1'b1;
								5'b00001:
									if (instr[26] == 1'b0)
										illegal_insn = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? 1'b0 : 1'b1);
									else
										illegal_insn = 1'b1;
								default: illegal_insn = 1'b1;
							endcase
					default: illegal_insn = 1'b1;
				endcase
			end
			7'h33: begin
				rf_ren_a_o = 1'b1;
				rf_ren_b_o = 1'b1;
				rf_we = 1'b1;
				if ({instr[26], instr[13:12]} == 3'b101)
					illegal_insn = (RV32B != 32'sd0 ? 1'b0 : 1'b1);
				else
					case ({instr[31:25], instr[14:12]})
						10'b0000000000, 10'b0100000000, 10'b0000000010, 10'b0000000011, 10'b0000000100, 10'b0000000110, 10'b0000000111, 10'b0000000001, 10'b0000000101, 10'b0100000101: illegal_insn = 1'b0;
						10'b0010000010, 10'b0010000100, 10'b0010000110, 10'b0100000111, 10'b0100000110, 10'b0100000100, 10'b0110000001, 10'b0110000101, 10'b0000101100, 10'b0000101110, 10'b0000101101, 10'b0000101111, 10'b0000100100, 10'b0100100100, 10'b0000100111, 10'b0100100001, 10'b0010100001, 10'b0110100001, 10'b0100100101, 10'b0100100111: illegal_insn = (RV32B != 32'sd0 ? 1'b0 : 1'b1);
						10'b0110100101, 10'b0010100101, 10'b0000100001, 10'b0000100101, 10'b0010100010, 10'b0010100100, 10'b0010100110, 10'b0010000001, 10'b0010000101, 10'b0000101001, 10'b0000101010, 10'b0000101011: illegal_insn = ((RV32B == 32'sd2) || (RV32B == 32'sd3) ? 1'b0 : 1'b1);
						10'b0100100110, 10'b0000100110: illegal_insn = (RV32B == 32'sd3 ? 1'b0 : 1'b1);
						10'b0000001000: begin
							multdiv_operator_o = 2'd0;
							multdiv_signed_mode_o = 2'b00;
							illegal_insn = (RV32M == 32'sd0 ? 1'b1 : 1'b0);
						end
						10'b0000001001: begin
							multdiv_operator_o = 2'd1;
							multdiv_signed_mode_o = 2'b11;
							illegal_insn = (RV32M == 32'sd0 ? 1'b1 : 1'b0);
						end
						10'b0000001010: begin
							multdiv_operator_o = 2'd1;
							multdiv_signed_mode_o = 2'b01;
							illegal_insn = (RV32M == 32'sd0 ? 1'b1 : 1'b0);
						end
						10'b0000001011: begin
							multdiv_operator_o = 2'd1;
							multdiv_signed_mode_o = 2'b00;
							illegal_insn = (RV32M == 32'sd0 ? 1'b1 : 1'b0);
						end
						10'b0000001100: begin
							multdiv_operator_o = 2'd2;
							multdiv_signed_mode_o = 2'b11;
							illegal_insn = (RV32M == 32'sd0 ? 1'b1 : 1'b0);
						end
						10'b0000001101: begin
							multdiv_operator_o = 2'd2;
							multdiv_signed_mode_o = 2'b00;
							illegal_insn = (RV32M == 32'sd0 ? 1'b1 : 1'b0);
						end
						10'b0000001110: begin
							multdiv_operator_o = 2'd3;
							multdiv_signed_mode_o = 2'b11;
							illegal_insn = (RV32M == 32'sd0 ? 1'b1 : 1'b0);
						end
						10'b0000001111: begin
							multdiv_operator_o = 2'd3;
							multdiv_signed_mode_o = 2'b00;
							illegal_insn = (RV32M == 32'sd0 ? 1'b1 : 1'b0);
						end
						default: illegal_insn = 1'b1;
					endcase
			end
			7'h0f:
				case (instr[14:12])
					3'b000: rf_we = 1'b0;
					3'b001: begin
						jump_in_dec_o = 1'b1;
						rf_we = 1'b0;
						if (instr_first_cycle_i) begin
							jump_set_o = 1'b1;
							icache_inval_o = 1'b1;
						end
					end
					default: illegal_insn = 1'b1;
				endcase
			7'h73:
				if (instr[14:12] == 3'b000) begin
					case (instr[31:20])
						12'h000: ecall_insn_o = 1'b1;
						12'h001: ebrk_insn_o = 1'b1;
						12'h302: mret_insn_o = 1'b1;
						12'h7b2: dret_insn_o = 1'b1;
						12'h105: wfi_insn_o = 1'b1;
						default: illegal_insn = 1'b1;
					endcase
					if ((instr_rs1 != 5'b00000) || (instr_rd != 5'b00000))
						illegal_insn = 1'b1;
				end
				else begin
					csr_access_o = 1'b1;
					rf_wdata_sel_o = 1'd1;
					rf_we = 1'b1;
					if (~instr[14])
						rf_ren_a_o = 1'b1;
					case (instr[13:12])
						2'b01: csr_op = 2'd1;
						2'b10: csr_op = 2'd2;
						2'b11: csr_op = 2'd3;
						default: csr_illegal = 1'b1;
					endcase
					illegal_insn = csr_illegal;
				end
			default: illegal_insn = 1'b1;
		endcase
		if (illegal_c_insn_i)
			illegal_insn = 1'b1;
		if (illegal_insn) begin
			rf_we = 1'b0;
			data_req_o = 1'b0;
			data_we_o = 1'b0;
			jump_in_dec_o = 1'b0;
			jump_set_o = 1'b0;
			branch_in_dec_o = 1'b0;
			csr_access_o = 1'b0;
		end
	end
	always @(*) begin
		alu_operator_o = 7'd44;
		alu_op_a_mux_sel_o = 2'd3;
		alu_op_b_mux_sel_o = 1'd1;
		imm_a_mux_sel_o = 1'd1;
		imm_b_mux_sel_o = 3'd0;
		bt_a_mux_sel_o = 2'd2;
		bt_b_mux_sel_o = 3'd0;
		opcode_alu = instr_alu[6:0];
		use_rs3_d = 1'b0;
		alu_multicycle_o = 1'b0;
		mult_sel_o = 1'b0;
		div_sel_o = 1'b0;
		case (opcode_alu)
			7'h6f: begin
				if (BranchTargetALU) begin
					bt_a_mux_sel_o = 2'd2;
					bt_b_mux_sel_o = 3'd4;
				end
				if (instr_first_cycle_i && !BranchTargetALU) begin
					alu_op_a_mux_sel_o = 2'd2;
					alu_op_b_mux_sel_o = 1'd1;
					imm_b_mux_sel_o = 3'd4;
					alu_operator_o = 7'd0;
				end
				else begin
					alu_op_a_mux_sel_o = 2'd2;
					alu_op_b_mux_sel_o = 1'd1;
					imm_b_mux_sel_o = 3'd5;
					alu_operator_o = 7'd0;
				end
			end
			7'h67: begin
				if (BranchTargetALU) begin
					bt_a_mux_sel_o = 2'd0;
					bt_b_mux_sel_o = 3'd0;
				end
				if (instr_first_cycle_i && !BranchTargetALU) begin
					alu_op_a_mux_sel_o = 2'd0;
					alu_op_b_mux_sel_o = 1'd1;
					imm_b_mux_sel_o = 3'd0;
					alu_operator_o = 7'd0;
				end
				else begin
					alu_op_a_mux_sel_o = 2'd2;
					alu_op_b_mux_sel_o = 1'd1;
					imm_b_mux_sel_o = 3'd5;
					alu_operator_o = 7'd0;
				end
			end
			7'h63: begin
				case (instr_alu[14:12])
					3'b000: alu_operator_o = 7'd29;
					3'b001: alu_operator_o = 7'd30;
					3'b100: alu_operator_o = 7'd25;
					3'b101: alu_operator_o = 7'd27;
					3'b110: alu_operator_o = 7'd26;
					3'b111: alu_operator_o = 7'd28;
					default:
						;
				endcase
				if (BranchTargetALU) begin
					bt_a_mux_sel_o = 2'd2;
					bt_b_mux_sel_o = (branch_taken_i ? 3'd2 : 3'd5);
				end
				if (instr_first_cycle_i) begin
					alu_op_a_mux_sel_o = 2'd0;
					alu_op_b_mux_sel_o = 1'd0;
				end
				else if (!BranchTargetALU) begin
					alu_op_a_mux_sel_o = 2'd2;
					alu_op_b_mux_sel_o = 1'd1;
					imm_b_mux_sel_o = (branch_taken_i ? 3'd2 : 3'd5);
					alu_operator_o = 7'd0;
				end
			end
			7'h23: begin
				alu_op_a_mux_sel_o = 2'd0;
				alu_op_b_mux_sel_o = 1'd0;
				alu_operator_o = 7'd0;
				if (!instr_alu[14]) begin
					imm_b_mux_sel_o = 3'd1;
					alu_op_b_mux_sel_o = 1'd1;
				end
			end
			7'h03: begin
				alu_op_a_mux_sel_o = 2'd0;
				alu_operator_o = 7'd0;
				alu_op_b_mux_sel_o = 1'd1;
				imm_b_mux_sel_o = 3'd0;
			end
			7'h37: begin
				alu_op_a_mux_sel_o = 2'd3;
				alu_op_b_mux_sel_o = 1'd1;
				imm_a_mux_sel_o = 1'd1;
				imm_b_mux_sel_o = 3'd3;
				alu_operator_o = 7'd0;
			end
			7'h17: begin
				alu_op_a_mux_sel_o = 2'd2;
				alu_op_b_mux_sel_o = 1'd1;
				imm_b_mux_sel_o = 3'd3;
				alu_operator_o = 7'd0;
			end
			7'h13: begin
				alu_op_a_mux_sel_o = 2'd0;
				alu_op_b_mux_sel_o = 1'd1;
				imm_b_mux_sel_o = 3'd0;
				case (instr_alu[14:12])
					3'b000: alu_operator_o = 7'd0;
					3'b010: alu_operator_o = 7'd43;
					3'b011: alu_operator_o = 7'd44;
					3'b100: alu_operator_o = 7'd2;
					3'b110: alu_operator_o = 7'd3;
					3'b111: alu_operator_o = 7'd4;
					3'b001:
						if (RV32B != 32'sd0)
							case (instr_alu[31:27])
								5'b00000: alu_operator_o = 7'd10;
								5'b00100:
									if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
										alu_operator_o = 7'd12;
								5'b01001: alu_operator_o = 7'd50;
								5'b00101: alu_operator_o = 7'd49;
								5'b01101: alu_operator_o = 7'd51;
								5'b00001:
									if (instr_alu[26] == 0)
										alu_operator_o = 7'd17;
								5'b01100:
									case (instr_alu[26:20])
										7'b0000000: alu_operator_o = 7'd40;
										7'b0000001: alu_operator_o = 7'd41;
										7'b0000010: alu_operator_o = 7'd42;
										7'b0000100: alu_operator_o = 7'd38;
										7'b0000101: alu_operator_o = 7'd39;
										7'b0010000:
											if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin
												alu_operator_o = 7'd59;
												alu_multicycle_o = 1'b1;
											end
										7'b0010001:
											if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin
												alu_operator_o = 7'd61;
												alu_multicycle_o = 1'b1;
											end
										7'b0010010:
											if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin
												alu_operator_o = 7'd63;
												alu_multicycle_o = 1'b1;
											end
										7'b0011000:
											if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin
												alu_operator_o = 7'd60;
												alu_multicycle_o = 1'b1;
											end
										7'b0011001:
											if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin
												alu_operator_o = 7'd62;
												alu_multicycle_o = 1'b1;
											end
										7'b0011010:
											if ((RV32B == 32'sd2) || (RV32B == 32'sd3)) begin
												alu_operator_o = 7'd64;
												alu_multicycle_o = 1'b1;
											end
										default:
											;
									endcase
								default:
									;
							endcase
						else
							alu_operator_o = 7'd10;
					3'b101:
						if (RV32B != 32'sd0) begin
							if (instr_alu[26] == 1'b1) begin
								alu_operator_o = 7'd48;
								alu_multicycle_o = 1'b1;
								if (instr_first_cycle_i)
									use_rs3_d = 1'b1;
								else
									use_rs3_d = 1'b0;
							end
							else
								case (instr_alu[31:27])
									5'b00000: alu_operator_o = 7'd9;
									5'b01000: alu_operator_o = 7'd8;
									5'b00100:
										if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
											alu_operator_o = 7'd11;
									5'b01001: alu_operator_o = 7'd52;
									5'b01100: begin
										alu_operator_o = 7'd13;
										alu_multicycle_o = 1'b1;
									end
									5'b01101: alu_operator_o = 7'd15;
									5'b00101: alu_operator_o = 7'd16;
									5'b00001:
										if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
											if (instr_alu[26] == 1'b0)
												alu_operator_o = 7'd18;
									default:
										;
								endcase
						end
						else if (instr_alu[31:27] == 5'b00000)
							alu_operator_o = 7'd9;
						else if (instr_alu[31:27] == 5'b01000)
							alu_operator_o = 7'd8;
					default:
						;
				endcase
			end
			7'h33: begin
				alu_op_a_mux_sel_o = 2'd0;
				alu_op_b_mux_sel_o = 1'd0;
				if (instr_alu[26]) begin
					if (RV32B != 32'sd0)
						case ({instr_alu[26:25], instr_alu[14:12]})
							5'b11001: begin
								alu_operator_o = 7'd46;
								alu_multicycle_o = 1'b1;
								if (instr_first_cycle_i)
									use_rs3_d = 1'b1;
								else
									use_rs3_d = 1'b0;
							end
							5'b11101: begin
								alu_operator_o = 7'd45;
								alu_multicycle_o = 1'b1;
								if (instr_first_cycle_i)
									use_rs3_d = 1'b1;
								else
									use_rs3_d = 1'b0;
							end
							5'b10001: begin
								alu_operator_o = 7'd47;
								alu_multicycle_o = 1'b1;
								if (instr_first_cycle_i)
									use_rs3_d = 1'b1;
								else
									use_rs3_d = 1'b0;
							end
							5'b10101: begin
								alu_operator_o = 7'd48;
								alu_multicycle_o = 1'b1;
								if (instr_first_cycle_i)
									use_rs3_d = 1'b1;
								else
									use_rs3_d = 1'b0;
							end
							default:
								;
						endcase
				end
				else
					case ({instr_alu[31:25], instr_alu[14:12]})
						10'b0000000000: alu_operator_o = 7'd0;
						10'b0100000000: alu_operator_o = 7'd1;
						10'b0000000010: alu_operator_o = 7'd43;
						10'b0000000011: alu_operator_o = 7'd44;
						10'b0000000100: alu_operator_o = 7'd2;
						10'b0000000110: alu_operator_o = 7'd3;
						10'b0000000111: alu_operator_o = 7'd4;
						10'b0000000001: alu_operator_o = 7'd10;
						10'b0000000101: alu_operator_o = 7'd9;
						10'b0100000101: alu_operator_o = 7'd8;
						10'b0110000001:
							if (RV32B != 32'sd0) begin
								alu_operator_o = 7'd14;
								alu_multicycle_o = 1'b1;
							end
						10'b0110000101:
							if (RV32B != 32'sd0) begin
								alu_operator_o = 7'd13;
								alu_multicycle_o = 1'b1;
							end
						10'b0000101100:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd31;
						10'b0000101110:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd33;
						10'b0000101101:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd32;
						10'b0000101111:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd34;
						10'b0000100100:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd35;
						10'b0100100100:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd36;
						10'b0000100111:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd37;
						10'b0100000100:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd5;
						10'b0100000110:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd6;
						10'b0100000111:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd7;
						10'b0010000010:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd22;
						10'b0010000100:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd23;
						10'b0010000110:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd24;
						10'b0100100001:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd50;
						10'b0010100001:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd49;
						10'b0110100001:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd51;
						10'b0100100101:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd52;
						10'b0100100111:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd55;
						10'b0110100101:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd15;
						10'b0010100101:
							if (RV32B != 32'sd0)
								alu_operator_o = 7'd16;
						10'b0000100001:
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								alu_operator_o = 7'd17;
						10'b0000100101:
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								alu_operator_o = 7'd18;
						10'b0010100010:
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								alu_operator_o = 7'd19;
						10'b0010100100:
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								alu_operator_o = 7'd20;
						10'b0010100110:
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								alu_operator_o = 7'd21;
						10'b0010000001:
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								alu_operator_o = 7'd12;
						10'b0010000101:
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								alu_operator_o = 7'd11;
						10'b0000101001:
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								alu_operator_o = 7'd56;
						10'b0000101010:
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								alu_operator_o = 7'd57;
						10'b0000101011:
							if ((RV32B == 32'sd2) || (RV32B == 32'sd3))
								alu_operator_o = 7'd58;
						10'b0100100110:
							if (RV32B == 32'sd3) begin
								alu_operator_o = 7'd54;
								alu_multicycle_o = 1'b1;
							end
						10'b0000100110:
							if (RV32B == 32'sd3) begin
								alu_operator_o = 7'd53;
								alu_multicycle_o = 1'b1;
							end
						10'b0000001000: begin
							alu_operator_o = 7'd0;
							mult_sel_o = (RV32M == 32'sd0 ? 1'b0 : 1'b1);
						end
						10'b0000001001: begin
							alu_operator_o = 7'd0;
							mult_sel_o = (RV32M == 32'sd0 ? 1'b0 : 1'b1);
						end
						10'b0000001010: begin
							alu_operator_o = 7'd0;
							mult_sel_o = (RV32M == 32'sd0 ? 1'b0 : 1'b1);
						end
						10'b0000001011: begin
							alu_operator_o = 7'd0;
							mult_sel_o = (RV32M == 32'sd0 ? 1'b0 : 1'b1);
						end
						10'b0000001100: begin
							alu_operator_o = 7'd0;
							div_sel_o = (RV32M == 32'sd0 ? 1'b0 : 1'b1);
						end
						10'b0000001101: begin
							alu_operator_o = 7'd0;
							div_sel_o = (RV32M == 32'sd0 ? 1'b0 : 1'b1);
						end
						10'b0000001110: begin
							alu_operator_o = 7'd0;
							div_sel_o = (RV32M == 32'sd0 ? 1'b0 : 1'b1);
						end
						10'b0000001111: begin
							alu_operator_o = 7'd0;
							div_sel_o = (RV32M == 32'sd0 ? 1'b0 : 1'b1);
						end
						default:
							;
					endcase
			end
			7'h0f:
				case (instr_alu[14:12])
					3'b000: begin
						alu_operator_o = 7'd0;
						alu_op_a_mux_sel_o = 2'd0;
						alu_op_b_mux_sel_o = 1'd1;
					end
					3'b001:
						if (BranchTargetALU) begin
							bt_a_mux_sel_o = 2'd2;
							bt_b_mux_sel_o = 3'd5;
						end
						else begin
							alu_op_a_mux_sel_o = 2'd2;
							alu_op_b_mux_sel_o = 1'd1;
							imm_b_mux_sel_o = 3'd5;
							alu_operator_o = 7'd0;
						end
					default:
						;
				endcase
			7'h73:
				if (instr_alu[14:12] == 3'b000) begin
					alu_op_a_mux_sel_o = 2'd0;
					alu_op_b_mux_sel_o = 1'd1;
				end
				else begin
					alu_op_b_mux_sel_o = 1'd1;
					imm_a_mux_sel_o = 1'd0;
					imm_b_mux_sel_o = 3'd0;
					if (instr_alu[14])
						alu_op_a_mux_sel_o = 2'd3;
					else
						alu_op_a_mux_sel_o = 2'd0;
				end
			default:
				;
		endcase
	end
	assign mult_en_o = (illegal_insn ? 1'b0 : mult_sel_o);
	assign div_en_o = (illegal_insn ? 1'b0 : div_sel_o);
	assign illegal_insn_o = illegal_insn | illegal_reg_rv32e;
	assign rf_we_o = rf_we & ~illegal_reg_rv32e;
	assign unused_instr_alu = {instr_alu[19:15], instr_alu[11:7]};
endmodule
module ibex_dummy_instr (
	clk_i,
	rst_ni,
	dummy_instr_en_i,
	dummy_instr_mask_i,
	dummy_instr_seed_en_i,
	dummy_instr_seed_i,
	fetch_valid_i,
	id_in_ready_i,
	insert_dummy_instr_o,
	dummy_instr_data_o
);
	localparam signed [31:0] ibex_pkg_LfsrWidth = 32;
	localparam [31:0] ibex_pkg_RndCnstLfsrSeedDefault = 32'hac533bf4;
	parameter [31:0] RndCnstLfsrSeed = ibex_pkg_RndCnstLfsrSeedDefault;
	localparam [159:0] ibex_pkg_RndCnstLfsrPermDefault = 160'h1e35ecba467fd1b12e958152c04fa43878a8daed;
	parameter [159:0] RndCnstLfsrPerm = ibex_pkg_RndCnstLfsrPermDefault;
	input wire clk_i;
	input wire rst_ni;
	input wire dummy_instr_en_i;
	input wire [2:0] dummy_instr_mask_i;
	input wire dummy_instr_seed_en_i;
	input wire [31:0] dummy_instr_seed_i;
	input wire fetch_valid_i;
	input wire id_in_ready_i;
	output wire insert_dummy_instr_o;
	output wire [31:0] dummy_instr_data_o;
	localparam [31:0] TIMEOUT_CNT_W = 5;
	localparam [31:0] OP_W = 5;
	localparam [31:0] LFSR_OUT_W = 17;
	wire [16:0] lfsr_data;
	wire [4:0] dummy_cnt_incr;
	wire [4:0] dummy_cnt_threshold;
	wire [4:0] dummy_cnt_d;
	reg [4:0] dummy_cnt_q;
	wire dummy_cnt_en;
	wire lfsr_en;
	wire [16:0] lfsr_state;
	wire insert_dummy_instr;
	reg [6:0] dummy_set;
	reg [2:0] dummy_opcode;
	wire [31:0] dummy_instr;
	reg [31:0] dummy_instr_seed_q;
	wire [31:0] dummy_instr_seed_d;
	assign lfsr_en = insert_dummy_instr & id_in_ready_i;
	assign dummy_instr_seed_d = dummy_instr_seed_q ^ dummy_instr_seed_i;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			dummy_instr_seed_q <= 1'sb0;
		else if (dummy_instr_seed_en_i)
			dummy_instr_seed_q <= dummy_instr_seed_d;
	prim_lfsr #(
		.LfsrDw(ibex_pkg_LfsrWidth),
		.StateOutDw(LFSR_OUT_W),
		.DefaultSeed(RndCnstLfsrSeed),
		.StatePermEn(1'b1),
		.StatePerm(RndCnstLfsrPerm)
	) lfsr_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.seed_en_i(dummy_instr_seed_en_i),
		.seed_i(dummy_instr_seed_d),
		.lfsr_en_i(lfsr_en),
		.entropy_i(1'sb0),
		.state_o(lfsr_state)
	);
	function automatic [16:0] sv2v_cast_B5B52;
		input reg [16:0] inp;
		sv2v_cast_B5B52 = inp;
	endfunction
	assign lfsr_data = sv2v_cast_B5B52(lfsr_state);
	assign dummy_cnt_threshold = lfsr_data[4-:TIMEOUT_CNT_W] & {dummy_instr_mask_i, {2 {1'b1}}};
	assign dummy_cnt_incr = dummy_cnt_q + {{4 {1'b0}}, 1'b1};
	assign dummy_cnt_d = (insert_dummy_instr ? {5 {1'sb0}} : dummy_cnt_incr);
	assign dummy_cnt_en = (dummy_instr_en_i & id_in_ready_i) & (fetch_valid_i | insert_dummy_instr);
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			dummy_cnt_q <= 1'sb0;
		else if (dummy_cnt_en)
			dummy_cnt_q <= dummy_cnt_d;
	assign insert_dummy_instr = dummy_instr_en_i & (dummy_cnt_q == dummy_cnt_threshold);
	always @(*)
		case (lfsr_data[16-:2])
			2'b00: begin
				dummy_set = 7'b0000000;
				dummy_opcode = 3'b000;
			end
			2'b01: begin
				dummy_set = 7'b0000001;
				dummy_opcode = 3'b000;
			end
			2'b10: begin
				dummy_set = 7'b0000001;
				dummy_opcode = 3'b100;
			end
			2'b11: begin
				dummy_set = 7'b0000000;
				dummy_opcode = 3'b111;
			end
			default: begin
				dummy_set = 7'b0000000;
				dummy_opcode = 3'b000;
			end
		endcase
	assign dummy_instr = {dummy_set, lfsr_data[14-:5], lfsr_data[9-:5], dummy_opcode, 5'h00, 7'h33};
	assign insert_dummy_instr_o = insert_dummy_instr;
	assign dummy_instr_data_o = dummy_instr;
endmodule
module ibex_ex_block (
	clk_i,
	rst_ni,
	alu_operator_i,
	alu_operand_a_i,
	alu_operand_b_i,
	alu_instr_first_cycle_i,
	bt_a_operand_i,
	bt_b_operand_i,
	multdiv_operator_i,
	mult_en_i,
	div_en_i,
	mult_sel_i,
	div_sel_i,
	multdiv_signed_mode_i,
	multdiv_operand_a_i,
	multdiv_operand_b_i,
	multdiv_ready_id_i,
	data_ind_timing_i,
	imd_val_we_o,
	imd_val_d_o,
	imd_val_q_i,
	alu_adder_result_ex_o,
	result_ex_o,
	branch_target_o,
	branch_decision_o,
	ex_valid_o
);
	parameter integer RV32M = 32'sd2;
	parameter integer RV32B = 32'sd0;
	parameter [0:0] BranchTargetALU = 0;
	input wire clk_i;
	input wire rst_ni;
	input wire [6:0] alu_operator_i;
	input wire [31:0] alu_operand_a_i;
	input wire [31:0] alu_operand_b_i;
	input wire alu_instr_first_cycle_i;
	input wire [31:0] bt_a_operand_i;
	input wire [31:0] bt_b_operand_i;
	input wire [1:0] multdiv_operator_i;
	input wire mult_en_i;
	input wire div_en_i;
	input wire mult_sel_i;
	input wire div_sel_i;
	input wire [1:0] multdiv_signed_mode_i;
	input wire [31:0] multdiv_operand_a_i;
	input wire [31:0] multdiv_operand_b_i;
	input wire multdiv_ready_id_i;
	input wire data_ind_timing_i;
	output wire [1:0] imd_val_we_o;
	output wire [67:0] imd_val_d_o;
	input wire [67:0] imd_val_q_i;
	output wire [31:0] alu_adder_result_ex_o;
	output wire [31:0] result_ex_o;
	output wire [31:0] branch_target_o;
	output wire branch_decision_o;
	output wire ex_valid_o;
	wire [31:0] alu_result;
	wire [31:0] multdiv_result;
	wire [32:0] multdiv_alu_operand_b;
	wire [32:0] multdiv_alu_operand_a;
	wire [33:0] alu_adder_result_ext;
	wire alu_cmp_result;
	wire alu_is_equal_result;
	wire multdiv_valid;
	wire multdiv_sel;
	wire [63:0] alu_imd_val_q;
	wire [63:0] alu_imd_val_d;
	wire [1:0] alu_imd_val_we;
	wire [67:0] multdiv_imd_val_d;
	wire [1:0] multdiv_imd_val_we;
	generate
		if (RV32M != 32'sd0) begin : gen_multdiv_m
			assign multdiv_sel = mult_sel_i | div_sel_i;
		end
		else begin : gen_multdiv_no_m
			assign multdiv_sel = 1'b0;
		end
	endgenerate
	assign imd_val_d_o[34+:34] = (multdiv_sel ? multdiv_imd_val_d[34+:34] : {2'b00, alu_imd_val_d[32+:32]});
	assign imd_val_d_o[0+:34] = (multdiv_sel ? multdiv_imd_val_d[0+:34] : {2'b00, alu_imd_val_d[0+:32]});
	assign imd_val_we_o = (multdiv_sel ? multdiv_imd_val_we : alu_imd_val_we);
	assign alu_imd_val_q = {imd_val_q_i[65-:32], imd_val_q_i[31-:32]};
	assign result_ex_o = (multdiv_sel ? multdiv_result : alu_result);
	assign branch_decision_o = alu_cmp_result;
	generate
		if (BranchTargetALU) begin : g_branch_target_alu
			wire [32:0] bt_alu_result;
			wire unused_bt_carry;
			assign bt_alu_result = bt_a_operand_i + bt_b_operand_i;
			assign unused_bt_carry = bt_alu_result[32];
			assign branch_target_o = bt_alu_result[31:0];
		end
		else begin : g_no_branch_target_alu
			wire [31:0] unused_bt_a_operand;
			wire [31:0] unused_bt_b_operand;
			assign unused_bt_a_operand = bt_a_operand_i;
			assign unused_bt_b_operand = bt_b_operand_i;
			assign branch_target_o = alu_adder_result_ex_o;
		end
	endgenerate
	ibex_alu #(.RV32B(RV32B)) alu_i(
		.operator_i(alu_operator_i),
		.operand_a_i(alu_operand_a_i),
		.operand_b_i(alu_operand_b_i),
		.instr_first_cycle_i(alu_instr_first_cycle_i),
		.imd_val_q_i(alu_imd_val_q),
		.imd_val_we_o(alu_imd_val_we),
		.imd_val_d_o(alu_imd_val_d),
		.multdiv_operand_a_i(multdiv_alu_operand_a),
		.multdiv_operand_b_i(multdiv_alu_operand_b),
		.multdiv_sel_i(multdiv_sel),
		.adder_result_o(alu_adder_result_ex_o),
		.adder_result_ext_o(alu_adder_result_ext),
		.result_o(alu_result),
		.comparison_result_o(alu_cmp_result),
		.is_equal_result_o(alu_is_equal_result)
	);
	generate
		if (RV32M == 32'sd1) begin : gen_multdiv_slow
			ibex_multdiv_slow multdiv_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.mult_en_i(mult_en_i),
				.div_en_i(div_en_i),
				.mult_sel_i(mult_sel_i),
				.div_sel_i(div_sel_i),
				.operator_i(multdiv_operator_i),
				.signed_mode_i(multdiv_signed_mode_i),
				.op_a_i(multdiv_operand_a_i),
				.op_b_i(multdiv_operand_b_i),
				.alu_adder_ext_i(alu_adder_result_ext),
				.alu_adder_i(alu_adder_result_ex_o),
				.equal_to_zero_i(alu_is_equal_result),
				.data_ind_timing_i(data_ind_timing_i),
				.valid_o(multdiv_valid),
				.alu_operand_a_o(multdiv_alu_operand_a),
				.alu_operand_b_o(multdiv_alu_operand_b),
				.imd_val_q_i(imd_val_q_i),
				.imd_val_d_o(multdiv_imd_val_d),
				.imd_val_we_o(multdiv_imd_val_we),
				.multdiv_ready_id_i(multdiv_ready_id_i),
				.multdiv_result_o(multdiv_result)
			);
		end
		else if ((RV32M == 32'sd2) || (RV32M == 32'sd3)) begin : gen_multdiv_fast
			ibex_multdiv_fast #(.RV32M(RV32M)) multdiv_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.mult_en_i(mult_en_i),
				.div_en_i(div_en_i),
				.mult_sel_i(mult_sel_i),
				.div_sel_i(div_sel_i),
				.operator_i(multdiv_operator_i),
				.signed_mode_i(multdiv_signed_mode_i),
				.op_a_i(multdiv_operand_a_i),
				.op_b_i(multdiv_operand_b_i),
				.alu_operand_a_o(multdiv_alu_operand_a),
				.alu_operand_b_o(multdiv_alu_operand_b),
				.alu_adder_ext_i(alu_adder_result_ext),
				.alu_adder_i(alu_adder_result_ex_o),
				.equal_to_zero_i(alu_is_equal_result),
				.data_ind_timing_i(data_ind_timing_i),
				.imd_val_q_i(imd_val_q_i),
				.imd_val_d_o(multdiv_imd_val_d),
				.imd_val_we_o(multdiv_imd_val_we),
				.multdiv_ready_id_i(multdiv_ready_id_i),
				.valid_o(multdiv_valid),
				.multdiv_result_o(multdiv_result)
			);
		end
	endgenerate
	assign ex_valid_o = (multdiv_sel ? multdiv_valid : ~(|alu_imd_val_we));
endmodule
module ibex_fetch_fifo (
	clk_i,
	rst_ni,
	clear_i,
	busy_o,
	in_valid_i,
	in_addr_i,
	in_rdata_i,
	in_err_i,
	out_valid_o,
	out_ready_i,
	out_addr_o,
	out_rdata_o,
	out_err_o,
	out_err_plus2_o
);
	parameter [31:0] NUM_REQS = 2;
	parameter [0:0] ResetAll = 1'b0;
	input wire clk_i;
	input wire rst_ni;
	input wire clear_i;
	output wire [NUM_REQS - 1:0] busy_o;
	input wire in_valid_i;
	input wire [31:0] in_addr_i;
	input wire [31:0] in_rdata_i;
	input wire in_err_i;
	output reg out_valid_o;
	input wire out_ready_i;
	output wire [31:0] out_addr_o;
	output reg [31:0] out_rdata_o;
	output reg out_err_o;
	output reg out_err_plus2_o;
	localparam [31:0] DEPTH = NUM_REQS + 1;
	wire [(DEPTH * 32) - 1:0] rdata_d;
	reg [(DEPTH * 32) - 1:0] rdata_q;
	wire [DEPTH - 1:0] err_d;
	reg [DEPTH - 1:0] err_q;
	wire [DEPTH - 1:0] valid_d;
	reg [DEPTH - 1:0] valid_q;
	wire [DEPTH - 1:0] lowest_free_entry;
	wire [DEPTH - 1:0] valid_pushed;
	wire [DEPTH - 1:0] valid_popped;
	wire [DEPTH - 1:0] entry_en;
	wire pop_fifo;
	wire [31:0] rdata;
	wire [31:0] rdata_unaligned;
	wire err;
	wire err_unaligned;
	wire err_plus2;
	wire valid;
	wire valid_unaligned;
	wire aligned_is_compressed;
	wire unaligned_is_compressed;
	wire addr_incr_two;
	wire [31:1] instr_addr_next;
	wire [31:1] instr_addr_d;
	reg [31:1] instr_addr_q;
	wire instr_addr_en;
	wire unused_addr_in;
	assign rdata = (valid_q[0] ? rdata_q[0+:32] : in_rdata_i);
	assign err = (valid_q[0] ? err_q[0] : in_err_i);
	assign valid = valid_q[0] | in_valid_i;
	assign rdata_unaligned = (valid_q[1] ? {rdata_q[47-:16], rdata[31:16]} : {in_rdata_i[15:0], rdata[31:16]});
	assign err_unaligned = (valid_q[1] ? (err_q[1] & ~unaligned_is_compressed) | err_q[0] : (valid_q[0] & err_q[0]) | (in_err_i & (~valid_q[0] | ~unaligned_is_compressed)));
	assign err_plus2 = (valid_q[1] ? err_q[1] & ~err_q[0] : (in_err_i & valid_q[0]) & ~err_q[0]);
	assign valid_unaligned = (valid_q[1] ? 1'b1 : valid_q[0] & in_valid_i);
	assign unaligned_is_compressed = (rdata[17:16] != 2'b11) & ~err;
	assign aligned_is_compressed = (rdata[1:0] != 2'b11) & ~err;
	always @(*)
		if (out_addr_o[1]) begin
			out_rdata_o = rdata_unaligned;
			out_err_o = err_unaligned;
			out_err_plus2_o = err_plus2;
			if (unaligned_is_compressed)
				out_valid_o = valid;
			else
				out_valid_o = valid_unaligned;
		end
		else begin
			out_rdata_o = rdata;
			out_err_o = err;
			out_err_plus2_o = 1'b0;
			out_valid_o = valid;
		end
	assign instr_addr_en = clear_i | (out_ready_i & out_valid_o);
	assign addr_incr_two = (instr_addr_q[1] ? unaligned_is_compressed : aligned_is_compressed);
	assign instr_addr_next = instr_addr_q[31:1] + {29'd0, ~addr_incr_two, addr_incr_two};
	assign instr_addr_d = (clear_i ? in_addr_i[31:1] : instr_addr_next);
	generate
		if (ResetAll) begin : g_instr_addr_ra
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					instr_addr_q <= 1'sb0;
				else if (instr_addr_en)
					instr_addr_q <= instr_addr_d;
		end
		else begin : g_instr_addr_nr
			always @(posedge clk_i)
				if (instr_addr_en)
					instr_addr_q <= instr_addr_d;
		end
	endgenerate
	assign out_addr_o = {instr_addr_q, 1'b0};
	assign unused_addr_in = in_addr_i[0];
	assign busy_o = valid_q[DEPTH - 1:DEPTH - NUM_REQS];
	assign pop_fifo = (out_ready_i & out_valid_o) & (~aligned_is_compressed | out_addr_o[1]);
	genvar i;
	generate
		for (i = 0; i < (DEPTH - 1); i = i + 1) begin : g_fifo_next
			if (i == 0) begin : g_ent0
				assign lowest_free_entry[i] = ~valid_q[i];
			end
			else begin : g_ent_others
				assign lowest_free_entry[i] = ~valid_q[i] & valid_q[i - 1];
			end
			assign valid_pushed[i] = (in_valid_i & lowest_free_entry[i]) | valid_q[i];
			assign valid_popped[i] = (pop_fifo ? valid_pushed[i + 1] : valid_pushed[i]);
			assign valid_d[i] = valid_popped[i] & ~clear_i;
			assign entry_en[i] = (valid_pushed[i + 1] & pop_fifo) | ((in_valid_i & lowest_free_entry[i]) & ~pop_fifo);
			assign rdata_d[i * 32+:32] = (valid_q[i + 1] ? rdata_q[(i + 1) * 32+:32] : in_rdata_i);
			assign err_d[i] = (valid_q[i + 1] ? err_q[i + 1] : in_err_i);
		end
	endgenerate
	assign lowest_free_entry[DEPTH - 1] = ~valid_q[DEPTH - 1] & valid_q[DEPTH - 2];
	assign valid_pushed[DEPTH - 1] = valid_q[DEPTH - 1] | (in_valid_i & lowest_free_entry[DEPTH - 1]);
	assign valid_popped[DEPTH - 1] = (pop_fifo ? 1'b0 : valid_pushed[DEPTH - 1]);
	assign valid_d[DEPTH - 1] = valid_popped[DEPTH - 1] & ~clear_i;
	assign entry_en[DEPTH - 1] = in_valid_i & lowest_free_entry[DEPTH - 1];
	assign rdata_d[(DEPTH - 1) * 32+:32] = in_rdata_i;
	assign err_d[DEPTH - 1] = in_err_i;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			valid_q <= 1'sb0;
		else
			valid_q <= valid_d;
	generate
		for (i = 0; i < DEPTH; i = i + 1) begin : g_fifo_regs
			if (ResetAll) begin : g_rdata_ra
				always @(posedge clk_i or negedge rst_ni)
					if (!rst_ni) begin
						rdata_q[i * 32+:32] <= 1'sb0;
						err_q[i] <= 1'sb0;
					end
					else if (entry_en[i]) begin
						rdata_q[i * 32+:32] <= rdata_d[i * 32+:32];
						err_q[i] <= err_d[i];
					end
			end
			else begin : g_rdata_nr
				always @(posedge clk_i)
					if (entry_en[i]) begin
						rdata_q[i * 32+:32] <= rdata_d[i * 32+:32];
						err_q[i] <= err_d[i];
					end
			end
		end
	endgenerate
endmodule
module ibex_icache (
	clk_i,
	rst_ni,
	req_i,
	branch_i,
	addr_i,
	ready_i,
	valid_o,
	rdata_o,
	addr_o,
	err_o,
	err_plus2_o,
	instr_req_o,
	instr_gnt_i,
	instr_addr_o,
	instr_rdata_i,
	instr_err_i,
	instr_rvalid_i,
	ic_tag_req_o,
	ic_tag_write_o,
	ic_tag_addr_o,
	ic_tag_wdata_o,
	ic_tag_rdata_i,
	ic_data_req_o,
	ic_data_write_o,
	ic_data_addr_o,
	ic_data_wdata_o,
	ic_data_rdata_i,
	ic_scr_key_valid_i,
	ic_scr_key_req_o,
	icache_enable_i,
	icache_inval_i,
	busy_o,
	ecc_error_o
);
	parameter [0:0] ICacheECC = 1'b0;
	parameter [0:0] ResetAll = 1'b0;
	localparam [31:0] ibex_pkg_BUS_SIZE = 32;
	parameter [31:0] BusSizeECC = ibex_pkg_BUS_SIZE;
	localparam [31:0] ibex_pkg_ADDR_W = 32;
	localparam [31:0] ibex_pkg_IC_LINE_SIZE = 64;
	localparam [31:0] ibex_pkg_IC_LINE_BYTES = 8;
	localparam [31:0] ibex_pkg_IC_NUM_WAYS = 2;
	localparam [31:0] ibex_pkg_IC_SIZE_BYTES = 4096;
	localparam [31:0] ibex_pkg_IC_NUM_LINES = (ibex_pkg_IC_SIZE_BYTES / ibex_pkg_IC_NUM_WAYS) / ibex_pkg_IC_LINE_BYTES;
	localparam [31:0] ibex_pkg_IC_INDEX_W = $clog2(ibex_pkg_IC_NUM_LINES);
	localparam [31:0] ibex_pkg_IC_LINE_W = 3;
	localparam [31:0] ibex_pkg_IC_TAG_SIZE = ((ibex_pkg_ADDR_W - ibex_pkg_IC_INDEX_W) - ibex_pkg_IC_LINE_W) + 1;
	parameter [31:0] TagSizeECC = ibex_pkg_IC_TAG_SIZE;
	parameter [31:0] LineSizeECC = ibex_pkg_IC_LINE_SIZE;
	parameter [0:0] BranchCache = 1'b0;
	input wire clk_i;
	input wire rst_ni;
	input wire req_i;
	input wire branch_i;
	input wire [31:0] addr_i;
	input wire ready_i;
	output wire valid_o;
	output wire [31:0] rdata_o;
	output wire [31:0] addr_o;
	output wire err_o;
	output wire err_plus2_o;
	output wire instr_req_o;
	input wire instr_gnt_i;
	output wire [31:0] instr_addr_o;
	input wire [31:0] instr_rdata_i;
	input wire instr_err_i;
	input wire instr_rvalid_i;
	output wire [1:0] ic_tag_req_o;
	output wire ic_tag_write_o;
	output wire [ibex_pkg_IC_INDEX_W - 1:0] ic_tag_addr_o;
	output wire [TagSizeECC - 1:0] ic_tag_wdata_o;
	input wire [(ibex_pkg_IC_NUM_WAYS * TagSizeECC) - 1:0] ic_tag_rdata_i;
	output wire [1:0] ic_data_req_o;
	output wire ic_data_write_o;
	output wire [ibex_pkg_IC_INDEX_W - 1:0] ic_data_addr_o;
	output wire [LineSizeECC - 1:0] ic_data_wdata_o;
	input wire [(ibex_pkg_IC_NUM_WAYS * LineSizeECC) - 1:0] ic_data_rdata_i;
	input wire ic_scr_key_valid_i;
	output reg ic_scr_key_req_o;
	input wire icache_enable_i;
	input wire icache_inval_i;
	output wire busy_o;
	output wire ecc_error_o;
	localparam [31:0] NUM_FB = 4;
	localparam [31:0] FB_THRESHOLD = 2;
	wire [31:0] lookup_addr_aligned;
	wire [31:0] prefetch_addr_d;
	reg [31:0] prefetch_addr_q;
	wire prefetch_addr_en;
	wire lookup_throttle;
	wire lookup_req_ic0;
	wire [31:0] lookup_addr_ic0;
	wire [ibex_pkg_IC_INDEX_W - 1:0] lookup_index_ic0;
	wire fill_req_ic0;
	wire [ibex_pkg_IC_INDEX_W - 1:0] fill_index_ic0;
	wire [ibex_pkg_IC_TAG_SIZE - 1:0] fill_tag_ic0;
	wire [63:0] fill_wdata_ic0;
	wire lookup_grant_ic0;
	wire lookup_actual_ic0;
	wire fill_grant_ic0;
	wire tag_req_ic0;
	wire [ibex_pkg_IC_INDEX_W - 1:0] tag_index_ic0;
	wire [1:0] tag_banks_ic0;
	wire tag_write_ic0;
	wire [TagSizeECC - 1:0] tag_wdata_ic0;
	wire data_req_ic0;
	wire [ibex_pkg_IC_INDEX_W - 1:0] data_index_ic0;
	wire [1:0] data_banks_ic0;
	wire data_write_ic0;
	wire [LineSizeECC - 1:0] data_wdata_ic0;
	wire [(ibex_pkg_IC_NUM_WAYS * TagSizeECC) - 1:0] tag_rdata_ic1;
	wire [(ibex_pkg_IC_NUM_WAYS * LineSizeECC) - 1:0] data_rdata_ic1;
	reg [LineSizeECC - 1:0] hit_data_ecc_ic1;
	wire [63:0] hit_data_ic1;
	reg lookup_valid_ic1;
	localparam [31:0] ibex_pkg_IC_INDEX_HI = (ibex_pkg_IC_INDEX_W + ibex_pkg_IC_LINE_W) - 1;
	reg [31:ibex_pkg_IC_INDEX_HI + 1] lookup_addr_ic1;
	wire [1:0] tag_match_ic1;
	wire tag_hit_ic1;
	wire [1:0] tag_invalid_ic1;
	wire [1:0] lowest_invalid_way_ic1;
	wire [1:0] round_robin_way_ic1;
	reg [1:0] round_robin_way_q;
	wire [1:0] sel_way_ic1;
	wire ecc_err_ic1;
	wire ecc_write_req;
	wire [1:0] ecc_write_ways;
	wire [ibex_pkg_IC_INDEX_W - 1:0] ecc_write_index;
	reg [1:0] fb_fill_level;
	wire fill_cache_new;
	wire fill_new_alloc;
	wire fill_spec_req;
	wire fill_spec_done;
	wire fill_spec_hold;
	wire [(NUM_FB * NUM_FB) - 1:0] fill_older_d;
	reg [(NUM_FB * NUM_FB) - 1:0] fill_older_q;
	wire [3:0] fill_alloc_sel;
	wire [3:0] fill_alloc;
	wire [3:0] fill_busy_d;
	reg [3:0] fill_busy_q;
	wire [3:0] fill_done;
	reg [3:0] fill_in_ic1;
	wire [3:0] fill_stale_d;
	reg [3:0] fill_stale_q;
	wire [3:0] fill_cache_d;
	reg [3:0] fill_cache_q;
	wire [3:0] fill_hit_ic1;
	wire [3:0] fill_hit_d;
	reg [3:0] fill_hit_q;
	localparam [31:0] ibex_pkg_BUS_BYTES = 4;
	localparam [31:0] ibex_pkg_IC_LINE_BEATS = ibex_pkg_IC_LINE_BYTES / ibex_pkg_BUS_BYTES;
	localparam [31:0] ibex_pkg_IC_LINE_BEATS_W = $clog2(ibex_pkg_IC_LINE_BEATS);
	wire [(ibex_pkg_IC_LINE_BEATS_W >= 0 ? (NUM_FB * (ibex_pkg_IC_LINE_BEATS_W + 1)) - 1 : (NUM_FB * (1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W - 1)):(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W + 0)] fill_ext_cnt_d;
	reg [(ibex_pkg_IC_LINE_BEATS_W >= 0 ? (NUM_FB * (ibex_pkg_IC_LINE_BEATS_W + 1)) - 1 : (NUM_FB * (1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W - 1)):(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W + 0)] fill_ext_cnt_q;
	wire [3:0] fill_ext_hold_d;
	reg [3:0] fill_ext_hold_q;
	wire [3:0] fill_ext_done_d;
	reg [3:0] fill_ext_done_q;
	wire [(ibex_pkg_IC_LINE_BEATS_W >= 0 ? (NUM_FB * (ibex_pkg_IC_LINE_BEATS_W + 1)) - 1 : (NUM_FB * (1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W - 1)):(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W + 0)] fill_rvd_cnt_d;
	reg [(ibex_pkg_IC_LINE_BEATS_W >= 0 ? (NUM_FB * (ibex_pkg_IC_LINE_BEATS_W + 1)) - 1 : (NUM_FB * (1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W - 1)):(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W + 0)] fill_rvd_cnt_q;
	wire [3:0] fill_rvd_done;
	wire [3:0] fill_ram_done_d;
	reg [3:0] fill_ram_done_q;
	wire [3:0] fill_out_grant;
	wire [(ibex_pkg_IC_LINE_BEATS_W >= 0 ? (NUM_FB * (ibex_pkg_IC_LINE_BEATS_W + 1)) - 1 : (NUM_FB * (1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W - 1)):(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W + 0)] fill_out_cnt_d;
	reg [(ibex_pkg_IC_LINE_BEATS_W >= 0 ? (NUM_FB * (ibex_pkg_IC_LINE_BEATS_W + 1)) - 1 : (NUM_FB * (1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W - 1)):(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W + 0)] fill_out_cnt_q;
	wire [3:0] fill_out_done;
	wire [3:0] fill_ext_req;
	wire [3:0] fill_rvd_exp;
	wire [3:0] fill_ram_req;
	wire [3:0] fill_out_req;
	wire [3:0] fill_data_sel;
	wire [3:0] fill_data_reg;
	wire [3:0] fill_data_hit;
	wire [3:0] fill_data_rvd;
	wire [(NUM_FB * ibex_pkg_IC_LINE_BEATS_W) - 1:0] fill_ext_off;
	wire [(NUM_FB * ibex_pkg_IC_LINE_BEATS_W) - 1:0] fill_rvd_off;
	wire [(ibex_pkg_IC_LINE_BEATS_W >= 0 ? (NUM_FB * (ibex_pkg_IC_LINE_BEATS_W + 1)) - 1 : (NUM_FB * (1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W - 1)):(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W + 0)] fill_ext_beat;
	wire [(ibex_pkg_IC_LINE_BEATS_W >= 0 ? (NUM_FB * (ibex_pkg_IC_LINE_BEATS_W + 1)) - 1 : (NUM_FB * (1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W - 1)):(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W + 0)] fill_rvd_beat;
	wire [3:0] fill_ext_arb;
	wire [3:0] fill_ram_arb;
	wire [3:0] fill_out_arb;
	wire [3:0] fill_rvd_arb;
	wire [3:0] fill_entry_en;
	wire [3:0] fill_addr_en;
	wire [3:0] fill_way_en;
	wire [(NUM_FB * ibex_pkg_IC_LINE_BEATS) - 1:0] fill_data_en;
	wire [(NUM_FB * ibex_pkg_IC_LINE_BEATS) - 1:0] fill_err_d;
	reg [(NUM_FB * ibex_pkg_IC_LINE_BEATS) - 1:0] fill_err_q;
	reg [31:0] fill_addr_q [0:3];
	reg [1:0] fill_way_q [0:3];
	wire [63:0] fill_data_d [0:3];
	reg [63:0] fill_data_q [0:3];
	localparam [31:0] ibex_pkg_BUS_W = 2;
	reg [31:ibex_pkg_BUS_W] fill_ext_req_addr;
	reg [31:0] fill_ram_req_addr;
	reg [1:0] fill_ram_req_way;
	reg [63:0] fill_ram_req_data;
	reg [63:0] fill_out_data;
	reg [ibex_pkg_IC_LINE_BEATS - 1:0] fill_out_err;
	wire instr_req;
	wire [31:ibex_pkg_BUS_W] instr_addr;
	wire skid_complete_instr;
	wire skid_ready;
	wire output_compressed;
	wire skid_valid_d;
	reg skid_valid_q;
	wire skid_en;
	wire [15:0] skid_data_d;
	reg [15:0] skid_data_q;
	reg skid_err_q;
	wire output_valid;
	wire addr_incr_two;
	wire output_addr_en;
	wire [31:1] output_addr_incr;
	wire [31:1] output_addr_d;
	reg [31:1] output_addr_q;
	reg [15:0] output_data_lo;
	reg [15:0] output_data_hi;
	wire data_valid;
	wire output_ready;
	wire [63:0] line_data;
	wire [ibex_pkg_IC_LINE_BEATS - 1:0] line_err;
	reg [31:0] line_data_muxed;
	reg line_err_muxed;
	wire [31:0] output_data;
	wire output_err;
	reg [1:0] inval_state_q;
	reg [1:0] inval_state_d;
	reg inval_write_req;
	reg inval_block_cache;
	reg [ibex_pkg_IC_INDEX_W - 1:0] inval_index_d;
	reg [ibex_pkg_IC_INDEX_W - 1:0] inval_index_q;
	reg inval_index_en;
	wire inval_active;
	assign lookup_addr_aligned = {lookup_addr_ic0[31:ibex_pkg_IC_LINE_W], {ibex_pkg_IC_LINE_W {1'b0}}};
	assign prefetch_addr_d = (lookup_grant_ic0 ? lookup_addr_aligned + {{(ibex_pkg_ADDR_W - ibex_pkg_IC_LINE_W) - 1 {1'b0}}, 1'b1, {ibex_pkg_IC_LINE_W {1'b0}}} : addr_i);
	assign prefetch_addr_en = branch_i | lookup_grant_ic0;
	generate
		if (ResetAll) begin : g_prefetch_addr_ra
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					prefetch_addr_q <= 1'sb0;
				else if (prefetch_addr_en)
					prefetch_addr_q <= prefetch_addr_d;
		end
		else begin : g_prefetch_addr_nr
			always @(posedge clk_i)
				if (prefetch_addr_en)
					prefetch_addr_q <= prefetch_addr_d;
		end
	endgenerate
	assign lookup_throttle = fb_fill_level > FB_THRESHOLD[1:0];
	assign lookup_req_ic0 = ((req_i & ~&fill_busy_q) & (branch_i | ~lookup_throttle)) & ~ecc_write_req;
	assign lookup_addr_ic0 = (branch_i ? addr_i : prefetch_addr_q);
	assign lookup_index_ic0 = lookup_addr_ic0[ibex_pkg_IC_INDEX_HI:ibex_pkg_IC_LINE_W];
	assign fill_req_ic0 = |fill_ram_req;
	assign fill_index_ic0 = fill_ram_req_addr[ibex_pkg_IC_INDEX_HI:ibex_pkg_IC_LINE_W];
	assign fill_tag_ic0 = {~inval_write_req & ~ecc_write_req, fill_ram_req_addr[31:ibex_pkg_IC_INDEX_HI + 1]};
	assign fill_wdata_ic0 = fill_ram_req_data;
	assign lookup_grant_ic0 = lookup_req_ic0;
	assign fill_grant_ic0 = ((fill_req_ic0 & ~lookup_req_ic0) & ~inval_write_req) & ~ecc_write_req;
	assign lookup_actual_ic0 = (lookup_grant_ic0 & icache_enable_i) & ~inval_block_cache;
	assign tag_req_ic0 = ((lookup_req_ic0 | fill_req_ic0) | inval_write_req) | ecc_write_req;
	assign tag_index_ic0 = (inval_write_req ? inval_index_q : (ecc_write_req ? ecc_write_index : (fill_grant_ic0 ? fill_index_ic0 : lookup_index_ic0)));
	assign tag_banks_ic0 = (ecc_write_req ? ecc_write_ways : (fill_grant_ic0 ? fill_ram_req_way : {ibex_pkg_IC_NUM_WAYS {1'b1}}));
	assign tag_write_ic0 = (fill_grant_ic0 | inval_write_req) | ecc_write_req;
	assign data_req_ic0 = lookup_req_ic0 | fill_req_ic0;
	assign data_index_ic0 = tag_index_ic0;
	assign data_banks_ic0 = tag_banks_ic0;
	assign data_write_ic0 = tag_write_ic0;
	generate
		if (ICacheECC) begin : gen_ecc_wdata
			wire [21:0] tag_ecc_input_padded;
			wire [27:0] tag_ecc_output_padded;
			wire [22 - ibex_pkg_IC_TAG_SIZE:0] unused_tag_ecc_output;
			assign tag_ecc_input_padded = {{22 - ibex_pkg_IC_TAG_SIZE {1'b0}}, fill_tag_ic0};
			assign unused_tag_ecc_output = tag_ecc_output_padded[21:ibex_pkg_IC_TAG_SIZE - 1];
			prim_secded_inv_28_22_enc tag_ecc_enc(
				.data_i(tag_ecc_input_padded),
				.data_o(tag_ecc_output_padded)
			);
			assign tag_wdata_ic0 = {tag_ecc_output_padded[27:22], tag_ecc_output_padded[ibex_pkg_IC_TAG_SIZE - 1:0]};
			genvar bank;
			for (bank = 0; bank < ibex_pkg_IC_LINE_BEATS; bank = bank + 1) begin : gen_ecc_banks
				prim_secded_inv_39_32_enc data_ecc_enc(
					.data_i(fill_wdata_ic0[bank * ibex_pkg_BUS_SIZE+:ibex_pkg_BUS_SIZE]),
					.data_o(data_wdata_ic0[bank * BusSizeECC+:BusSizeECC])
				);
			end
		end
		else begin : gen_noecc_wdata
			assign tag_wdata_ic0 = fill_tag_ic0;
			assign data_wdata_ic0 = fill_wdata_ic0;
		end
	endgenerate
	assign ic_tag_req_o = {ibex_pkg_IC_NUM_WAYS {tag_req_ic0}} & tag_banks_ic0;
	assign ic_tag_write_o = tag_write_ic0;
	assign ic_tag_addr_o = tag_index_ic0;
	assign ic_tag_wdata_o = tag_wdata_ic0;
	assign tag_rdata_ic1 = ic_tag_rdata_i;
	assign ic_data_req_o = {ibex_pkg_IC_NUM_WAYS {data_req_ic0}} & data_banks_ic0;
	assign ic_data_write_o = data_write_ic0;
	assign ic_data_addr_o = data_index_ic0;
	assign ic_data_wdata_o = data_wdata_ic0;
	assign data_rdata_ic1 = ic_data_rdata_i;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			lookup_valid_ic1 <= 1'b0;
		else
			lookup_valid_ic1 <= lookup_actual_ic0;
	generate
		if (ResetAll) begin : g_lookup_addr_ra
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni) begin
					lookup_addr_ic1 <= 1'sb0;
					fill_in_ic1 <= 1'sb0;
				end
				else if (lookup_grant_ic0) begin
					lookup_addr_ic1 <= lookup_addr_ic0[31:ibex_pkg_IC_INDEX_HI + 1];
					fill_in_ic1 <= fill_alloc_sel;
				end
		end
		else begin : g_lookup_addr_nr
			always @(posedge clk_i)
				if (lookup_grant_ic0) begin
					lookup_addr_ic1 <= lookup_addr_ic0[31:ibex_pkg_IC_INDEX_HI + 1];
					fill_in_ic1 <= fill_alloc_sel;
				end
		end
	endgenerate
	genvar way;
	generate
		for (way = 0; way < ibex_pkg_IC_NUM_WAYS; way = way + 1) begin : gen_tag_match
			assign tag_match_ic1[way] = tag_rdata_ic1[((1 - way) * TagSizeECC) + (ibex_pkg_IC_TAG_SIZE - 1)-:ibex_pkg_IC_TAG_SIZE] == {1'b1, lookup_addr_ic1[31:ibex_pkg_IC_INDEX_HI + 1]};
			assign tag_invalid_ic1[way] = ~tag_rdata_ic1[((1 - way) * TagSizeECC) + (ibex_pkg_IC_TAG_SIZE - 1)];
		end
	endgenerate
	assign tag_hit_ic1 = |tag_match_ic1;
	always @(*) begin
		hit_data_ecc_ic1 = 'b0;
		begin : sv2v_autoblock_1
			reg signed [31:0] way;
			for (way = 0; way < ibex_pkg_IC_NUM_WAYS; way = way + 1)
				if (tag_match_ic1[way])
					hit_data_ecc_ic1 = hit_data_ecc_ic1 | data_rdata_ic1[(1 - way) * LineSizeECC+:LineSizeECC];
		end
	end
	assign lowest_invalid_way_ic1[0] = tag_invalid_ic1[0];
	assign round_robin_way_ic1[0] = round_robin_way_q[1];
	generate
		for (way = 1; way < ibex_pkg_IC_NUM_WAYS; way = way + 1) begin : gen_lowest_way
			assign lowest_invalid_way_ic1[way] = tag_invalid_ic1[way] & ~|tag_invalid_ic1[way - 1:0];
			assign round_robin_way_ic1[way] = round_robin_way_q[way - 1];
		end
	endgenerate
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			round_robin_way_q <= 2'b01;
		else if (lookup_valid_ic1)
			round_robin_way_q <= round_robin_way_ic1;
	assign sel_way_ic1 = (|tag_invalid_ic1 ? lowest_invalid_way_ic1 : round_robin_way_q);
	generate
		if (ICacheECC) begin : gen_data_ecc_checking
			wire [1:0] tag_err_ic1;
			wire [(ibex_pkg_IC_LINE_BEATS * 2) - 1:0] data_err_ic1;
			wire ecc_correction_write_d;
			reg ecc_correction_write_q;
			wire [1:0] ecc_correction_ways_d;
			reg [1:0] ecc_correction_ways_q;
			reg [ibex_pkg_IC_INDEX_W - 1:0] lookup_index_ic1;
			reg [ibex_pkg_IC_INDEX_W - 1:0] ecc_correction_index_q;
			genvar way;
			for (way = 0; way < ibex_pkg_IC_NUM_WAYS; way = way + 1) begin : gen_tag_ecc
				wire [1:0] tag_err_bank_ic1;
				wire [27:0] tag_rdata_padded_ic1;
				assign tag_rdata_padded_ic1 = {tag_rdata_ic1[((1 - way) * TagSizeECC) + (TagSizeECC - 1)-:6], {22 - ibex_pkg_IC_TAG_SIZE {1'b0}}, tag_rdata_ic1[((1 - way) * TagSizeECC) + (ibex_pkg_IC_TAG_SIZE - 1)-:ibex_pkg_IC_TAG_SIZE]};
				prim_secded_inv_28_22_dec data_ecc_dec(
					.data_i(tag_rdata_padded_ic1),
					.err_o(tag_err_bank_ic1)
				);
				assign tag_err_ic1[way] = |tag_err_bank_ic1;
			end
			genvar bank;
			for (bank = 0; bank < ibex_pkg_IC_LINE_BEATS; bank = bank + 1) begin : gen_ecc_banks
				prim_secded_inv_39_32_dec data_ecc_dec(
					.data_i(hit_data_ecc_ic1[bank * BusSizeECC+:BusSizeECC]),
					.err_o(data_err_ic1[bank * 2+:2])
				);
				assign hit_data_ic1[bank * ibex_pkg_BUS_SIZE+:ibex_pkg_BUS_SIZE] = hit_data_ecc_ic1[bank * BusSizeECC+:ibex_pkg_BUS_SIZE];
			end
			assign ecc_err_ic1 = lookup_valid_ic1 & ((|data_err_ic1 & tag_hit_ic1) | |tag_err_ic1);
			assign ecc_correction_ways_d = {ibex_pkg_IC_NUM_WAYS {|tag_err_ic1}} | (tag_match_ic1 & {ibex_pkg_IC_NUM_WAYS {|data_err_ic1}});
			assign ecc_correction_write_d = ecc_err_ic1;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					ecc_correction_write_q <= 1'b0;
				else
					ecc_correction_write_q <= ecc_correction_write_d;
			if (ResetAll) begin : g_lookup_ind_ra
				always @(posedge clk_i or negedge rst_ni)
					if (!rst_ni)
						lookup_index_ic1 <= 1'sb0;
					else if (lookup_grant_ic0)
						lookup_index_ic1 <= lookup_addr_ic0[ibex_pkg_IC_INDEX_HI-:ibex_pkg_IC_INDEX_W];
			end
			else begin : g_lookup_ind_nr
				always @(posedge clk_i)
					if (lookup_grant_ic0)
						lookup_index_ic1 <= lookup_addr_ic0[ibex_pkg_IC_INDEX_HI-:ibex_pkg_IC_INDEX_W];
			end
			if (ResetAll) begin : g_ecc_correction_ra
				always @(posedge clk_i or negedge rst_ni)
					if (!rst_ni) begin
						ecc_correction_ways_q <= 1'sb0;
						ecc_correction_index_q <= 1'sb0;
					end
					else if (ecc_err_ic1) begin
						ecc_correction_ways_q <= ecc_correction_ways_d;
						ecc_correction_index_q <= lookup_index_ic1;
					end
			end
			else begin : g_ecc_correction_nr
				always @(posedge clk_i)
					if (ecc_err_ic1) begin
						ecc_correction_ways_q <= ecc_correction_ways_d;
						ecc_correction_index_q <= lookup_index_ic1;
					end
			end
			assign ecc_write_req = ecc_correction_write_q;
			assign ecc_write_ways = ecc_correction_ways_q;
			assign ecc_write_index = ecc_correction_index_q;
			assign ecc_error_o = ecc_err_ic1;
		end
		else begin : gen_no_data_ecc
			assign ecc_err_ic1 = 1'b0;
			assign ecc_write_req = 1'b0;
			assign ecc_write_ways = 1'sb0;
			assign ecc_write_index = 1'sb0;
			assign hit_data_ic1 = hit_data_ecc_ic1;
			assign ecc_error_o = 1'b0;
		end
		if (BranchCache) begin : gen_caching_logic
			localparam [31:0] CACHE_AHEAD = 2;
			localparam [31:0] CACHE_CNT_W = 2;
			wire cache_cnt_dec;
			wire [1:0] cache_cnt_d;
			reg [1:0] cache_cnt_q;
			assign cache_cnt_dec = lookup_grant_ic0 & |cache_cnt_q;
			assign cache_cnt_d = (branch_i ? CACHE_AHEAD[1:0] : cache_cnt_q - {1'b0, cache_cnt_dec});
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					cache_cnt_q <= 1'sb0;
				else
					cache_cnt_q <= cache_cnt_d;
			assign fill_cache_new = ((branch_i | |cache_cnt_q) & icache_enable_i) & ~inval_block_cache;
		end
		else begin : gen_cache_all
			assign fill_cache_new = icache_enable_i & ~inval_block_cache;
		end
	endgenerate
	always @(*) begin
		fb_fill_level = 1'sb0;
		begin : sv2v_autoblock_2
			reg signed [31:0] i;
			for (i = 0; i < NUM_FB; i = i + 1)
				if (fill_busy_q[i] & ~fill_stale_q[i])
					fb_fill_level = fb_fill_level + 2'b01;
		end
	end
	assign fill_new_alloc = lookup_grant_ic0;
	assign fill_spec_req = (~icache_enable_i | branch_i) & ~|fill_ext_req;
	assign fill_spec_done = fill_spec_req & instr_gnt_i;
	assign fill_spec_hold = fill_spec_req & ~instr_gnt_i;
	genvar fb;
	generate
		for (fb = 0; fb < NUM_FB; fb = fb + 1) begin : gen_fbs
			if (fb == 0) begin : gen_fb_zero
				assign fill_alloc_sel[fb] = ~fill_busy_q[fb];
			end
			else begin : gen_fb_rest
				assign fill_alloc_sel[fb] = ~fill_busy_q[fb] & &fill_busy_q[fb - 1:0];
			end
			assign fill_alloc[fb] = fill_alloc_sel[fb] & fill_new_alloc;
			assign fill_busy_d[fb] = fill_alloc[fb] | (fill_busy_q[fb] & ~fill_done[fb]);
			assign fill_older_d[fb * NUM_FB+:NUM_FB] = (fill_alloc[fb] ? fill_busy_q : fill_older_q[fb * NUM_FB+:NUM_FB]) & ~fill_done;
			assign fill_done[fb] = ((((fill_ram_done_q[fb] | fill_hit_q[fb]) | ~fill_cache_q[fb]) | |fill_err_q[fb * ibex_pkg_IC_LINE_BEATS+:ibex_pkg_IC_LINE_BEATS]) & ((fill_out_done[fb] | fill_stale_q[fb]) | branch_i)) & fill_rvd_done[fb];
			assign fill_stale_d[fb] = fill_busy_q[fb] & (branch_i | fill_stale_q[fb]);
			assign fill_cache_d[fb] = (fill_alloc[fb] & fill_cache_new) | (((fill_cache_q[fb] & fill_busy_q[fb]) & icache_enable_i) & ~icache_inval_i);
			assign fill_hit_ic1[fb] = ((lookup_valid_ic1 & fill_in_ic1[fb]) & tag_hit_ic1) & ~ecc_err_ic1;
			assign fill_hit_d[fb] = fill_hit_ic1[fb] | (fill_hit_q[fb] & fill_busy_q[fb]);
			assign fill_ext_req[fb] = fill_busy_q[fb] & ~fill_ext_done_d[fb];
			assign fill_ext_cnt_d[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] = (fill_alloc[fb] ? {{ibex_pkg_IC_LINE_BEATS_W {1'b0}}, fill_spec_done} : fill_ext_cnt_q[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] + {{ibex_pkg_IC_LINE_BEATS_W {1'b0}}, fill_ext_arb[fb] & instr_gnt_i});
			assign fill_ext_hold_d[fb] = (fill_alloc[fb] & fill_spec_hold) | (fill_ext_arb[fb] & ~instr_gnt_i);
			assign fill_ext_done_d[fb] = ((((fill_ext_cnt_q[(fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W : ibex_pkg_IC_LINE_BEATS_W - ibex_pkg_IC_LINE_BEATS_W)] | fill_hit_ic1[fb]) | fill_hit_q[fb]) | (~fill_cache_q[fb] & ((branch_i | fill_stale_q[fb]) | fill_ext_beat[(fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W : ibex_pkg_IC_LINE_BEATS_W - ibex_pkg_IC_LINE_BEATS_W)]))) & ~fill_ext_hold_q[fb]) & fill_busy_q[fb];
			assign fill_rvd_exp[fb] = fill_busy_q[fb] & ~fill_rvd_done[fb];
			assign fill_rvd_cnt_d[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] = (fill_alloc[fb] ? {(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W) * 1 {1'sb0}} : fill_rvd_cnt_q[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] + {{ibex_pkg_IC_LINE_BEATS_W {1'b0}}, fill_rvd_arb[fb]});
			assign fill_rvd_done[fb] = (fill_ext_done_q[fb] & ~fill_ext_hold_q[fb]) & (fill_rvd_cnt_q[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] == fill_ext_cnt_q[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)]);
			assign fill_out_req[fb] = ((fill_busy_q[fb] & ~fill_stale_q[fb]) & ~fill_out_done[fb]) & (((fill_hit_ic1[fb] | fill_hit_q[fb]) | (fill_rvd_beat[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] > fill_out_cnt_q[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)])) | fill_rvd_arb[fb]);
			assign fill_out_grant[fb] = fill_out_arb[fb] & output_ready;
			assign fill_out_cnt_d[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] = (fill_alloc[fb] ? {1'b0, lookup_addr_ic0[2:ibex_pkg_BUS_W]} : fill_out_cnt_q[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] + {{ibex_pkg_IC_LINE_BEATS_W {1'b0}}, fill_out_grant[fb]});
			assign fill_out_done[fb] = fill_out_cnt_q[(fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W : ibex_pkg_IC_LINE_BEATS_W - ibex_pkg_IC_LINE_BEATS_W)];
			assign fill_ram_req[fb] = ((((fill_busy_q[fb] & fill_rvd_cnt_q[(fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W : ibex_pkg_IC_LINE_BEATS_W - ibex_pkg_IC_LINE_BEATS_W)]) & ~fill_hit_q[fb]) & fill_cache_q[fb]) & ~|fill_err_q[fb * ibex_pkg_IC_LINE_BEATS+:ibex_pkg_IC_LINE_BEATS]) & ~fill_ram_done_q[fb];
			assign fill_ram_done_d[fb] = fill_ram_arb[fb] | (fill_ram_done_q[fb] & fill_busy_q[fb]);
			assign fill_ext_beat[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] = {1'b0, fill_addr_q[fb][2:ibex_pkg_BUS_W]} + fill_ext_cnt_q[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W : (ibex_pkg_IC_LINE_BEATS_W + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) - 1) : ibex_pkg_IC_LINE_BEATS_W - (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W : (ibex_pkg_IC_LINE_BEATS_W + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) - 1)) : (((fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W : (ibex_pkg_IC_LINE_BEATS_W + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) - 1) : ibex_pkg_IC_LINE_BEATS_W - (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W : (ibex_pkg_IC_LINE_BEATS_W + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) - 1))) + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) - 1)-:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)];
			assign fill_ext_off[fb * ibex_pkg_IC_LINE_BEATS_W+:ibex_pkg_IC_LINE_BEATS_W] = fill_ext_beat[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W - 1 : ibex_pkg_IC_LINE_BEATS_W - (ibex_pkg_IC_LINE_BEATS_W - 1)) : (((fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W - 1 : ibex_pkg_IC_LINE_BEATS_W - (ibex_pkg_IC_LINE_BEATS_W - 1))) + ibex_pkg_IC_LINE_BEATS_W) - 1)-:ibex_pkg_IC_LINE_BEATS_W];
			assign fill_rvd_beat[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] = {1'b0, fill_addr_q[fb][2:ibex_pkg_BUS_W]} + fill_rvd_cnt_q[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W : (ibex_pkg_IC_LINE_BEATS_W + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) - 1) : ibex_pkg_IC_LINE_BEATS_W - (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W : (ibex_pkg_IC_LINE_BEATS_W + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) - 1)) : (((fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W : (ibex_pkg_IC_LINE_BEATS_W + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) - 1) : ibex_pkg_IC_LINE_BEATS_W - (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W : (ibex_pkg_IC_LINE_BEATS_W + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) - 1))) + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) - 1)-:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)];
			assign fill_rvd_off[fb * ibex_pkg_IC_LINE_BEATS_W+:ibex_pkg_IC_LINE_BEATS_W] = fill_rvd_beat[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W - 1 : ibex_pkg_IC_LINE_BEATS_W - (ibex_pkg_IC_LINE_BEATS_W - 1)) : (((fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)) + (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W - 1 : ibex_pkg_IC_LINE_BEATS_W - (ibex_pkg_IC_LINE_BEATS_W - 1))) + ibex_pkg_IC_LINE_BEATS_W) - 1)-:ibex_pkg_IC_LINE_BEATS_W];
			assign fill_ext_arb[fb] = fill_ext_req[fb] & ~|(fill_ext_req & fill_older_q[fb * NUM_FB+:NUM_FB]);
			assign fill_ram_arb[fb] = (fill_ram_req[fb] & fill_grant_ic0) & ~|(fill_ram_req & fill_older_q[fb * NUM_FB+:NUM_FB]);
			assign fill_data_sel[fb] = ~|(((fill_busy_q & ~fill_out_done) & ~fill_stale_q) & fill_older_q[fb * NUM_FB+:NUM_FB]);
			assign fill_out_arb[fb] = fill_out_req[fb] & fill_data_sel[fb];
			assign fill_rvd_arb[fb] = (instr_rvalid_i & fill_rvd_exp[fb]) & ~|(fill_rvd_exp & fill_older_q[fb * NUM_FB+:NUM_FB]);
			assign fill_data_reg[fb] = (((fill_busy_q[fb] & ~fill_stale_q[fb]) & ~fill_out_done[fb]) & fill_data_sel[fb]) & (((fill_rvd_beat[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] > fill_out_cnt_q[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)]) | fill_hit_q[fb]) | |fill_err_q[fb * ibex_pkg_IC_LINE_BEATS+:ibex_pkg_IC_LINE_BEATS]);
			assign fill_data_hit[fb] = (fill_busy_q[fb] & fill_hit_ic1[fb]) & fill_data_sel[fb];
			assign fill_data_rvd[fb] = ((((((fill_busy_q[fb] & fill_rvd_arb[fb]) & ~fill_hit_q[fb]) & ~fill_hit_ic1[fb]) & ~fill_stale_q[fb]) & ~fill_out_done[fb]) & (fill_rvd_beat[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] == fill_out_cnt_q[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)])) & fill_data_sel[fb];
			assign fill_entry_en[fb] = fill_alloc[fb] | fill_busy_q[fb];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni) begin
					fill_busy_q[fb] <= 1'b0;
					fill_older_q[fb * NUM_FB+:NUM_FB] <= 1'sb0;
					fill_stale_q[fb] <= 1'b0;
					fill_cache_q[fb] <= 1'b0;
					fill_hit_q[fb] <= 1'b0;
					fill_ext_cnt_q[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] <= 1'sb0;
					fill_ext_hold_q[fb] <= 1'b0;
					fill_ext_done_q[fb] <= 1'b0;
					fill_rvd_cnt_q[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] <= 1'sb0;
					fill_ram_done_q[fb] <= 1'b0;
					fill_out_cnt_q[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] <= 1'sb0;
				end
				else if (fill_entry_en[fb]) begin
					fill_busy_q[fb] <= fill_busy_d[fb];
					fill_older_q[fb * NUM_FB+:NUM_FB] <= fill_older_d[fb * NUM_FB+:NUM_FB];
					fill_stale_q[fb] <= fill_stale_d[fb];
					fill_cache_q[fb] <= fill_cache_d[fb];
					fill_hit_q[fb] <= fill_hit_d[fb];
					fill_ext_cnt_q[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] <= fill_ext_cnt_d[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)];
					fill_ext_hold_q[fb] <= fill_ext_hold_d[fb];
					fill_ext_done_q[fb] <= fill_ext_done_d[fb];
					fill_rvd_cnt_q[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] <= fill_rvd_cnt_d[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)];
					fill_ram_done_q[fb] <= fill_ram_done_d[fb];
					fill_out_cnt_q[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)] <= fill_out_cnt_d[(ibex_pkg_IC_LINE_BEATS_W >= 0 ? 0 : ibex_pkg_IC_LINE_BEATS_W) + (fb * (ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W))+:(ibex_pkg_IC_LINE_BEATS_W >= 0 ? ibex_pkg_IC_LINE_BEATS_W + 1 : 1 - ibex_pkg_IC_LINE_BEATS_W)];
				end
			assign fill_addr_en[fb] = fill_alloc[fb];
			assign fill_way_en[fb] = lookup_valid_ic1 & fill_in_ic1[fb];
			if (ResetAll) begin : g_fill_addr_ra
				always @(posedge clk_i or negedge rst_ni)
					if (!rst_ni)
						fill_addr_q[fb] <= 1'sb0;
					else if (fill_addr_en[fb])
						fill_addr_q[fb] <= lookup_addr_ic0;
			end
			else begin : g_fill_addr_nr
				always @(posedge clk_i)
					if (fill_addr_en[fb])
						fill_addr_q[fb] <= lookup_addr_ic0;
			end
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					fill_way_q[fb] <= 1'sb0;
				else if (fill_way_en[fb])
					fill_way_q[fb] <= sel_way_ic1;
			assign fill_data_d[fb] = (fill_hit_ic1[fb] ? hit_data_ic1 : {ibex_pkg_IC_LINE_BEATS {instr_rdata_i}});
			genvar b;
			for (b = 0; b < ibex_pkg_IC_LINE_BEATS; b = b + 1) begin : gen_data_buf
				assign fill_err_d[(fb * ibex_pkg_IC_LINE_BEATS) + b] = ((fill_rvd_arb[fb] & instr_err_i) & (fill_rvd_off[fb * ibex_pkg_IC_LINE_BEATS_W+:ibex_pkg_IC_LINE_BEATS_W] == b[ibex_pkg_IC_LINE_BEATS_W - 1:0])) | (fill_busy_q[fb] & fill_err_q[(fb * ibex_pkg_IC_LINE_BEATS) + b]);
				always @(posedge clk_i or negedge rst_ni)
					if (!rst_ni)
						fill_err_q[(fb * ibex_pkg_IC_LINE_BEATS) + b] <= 1'sb0;
					else if (fill_entry_en[fb])
						fill_err_q[(fb * ibex_pkg_IC_LINE_BEATS) + b] <= fill_err_d[(fb * ibex_pkg_IC_LINE_BEATS) + b];
				assign fill_data_en[(fb * ibex_pkg_IC_LINE_BEATS) + b] = fill_hit_ic1[fb] | ((fill_rvd_arb[fb] & ~fill_hit_q[fb]) & (fill_rvd_off[fb * ibex_pkg_IC_LINE_BEATS_W+:ibex_pkg_IC_LINE_BEATS_W] == b[ibex_pkg_IC_LINE_BEATS_W - 1:0]));
				if (ResetAll) begin : g_fill_data_ra
					always @(posedge clk_i or negedge rst_ni)
						if (!rst_ni)
							fill_data_q[fb][b * ibex_pkg_BUS_SIZE+:ibex_pkg_BUS_SIZE] <= 1'sb0;
						else if (fill_data_en[(fb * ibex_pkg_IC_LINE_BEATS) + b])
							fill_data_q[fb][b * ibex_pkg_BUS_SIZE+:ibex_pkg_BUS_SIZE] <= fill_data_d[fb][b * ibex_pkg_BUS_SIZE+:ibex_pkg_BUS_SIZE];
				end
				else begin : g_fill_data_nr
					always @(posedge clk_i)
						if (fill_data_en[(fb * ibex_pkg_IC_LINE_BEATS) + b])
							fill_data_q[fb][b * ibex_pkg_BUS_SIZE+:ibex_pkg_BUS_SIZE] <= fill_data_d[fb][b * ibex_pkg_BUS_SIZE+:ibex_pkg_BUS_SIZE];
				end
			end
		end
	endgenerate
	always @(*) begin
		fill_ext_req_addr = 1'sb0;
		begin : sv2v_autoblock_3
			reg signed [31:0] i;
			for (i = 0; i < NUM_FB; i = i + 1)
				if (fill_ext_arb[i])
					fill_ext_req_addr = fill_ext_req_addr | {fill_addr_q[i][31:ibex_pkg_IC_LINE_W], fill_ext_off[i * ibex_pkg_IC_LINE_BEATS_W+:ibex_pkg_IC_LINE_BEATS_W]};
		end
	end
	always @(*) begin
		fill_ram_req_addr = 1'sb0;
		fill_ram_req_way = 1'sb0;
		fill_ram_req_data = 1'sb0;
		begin : sv2v_autoblock_4
			reg signed [31:0] i;
			for (i = 0; i < NUM_FB; i = i + 1)
				if (fill_ram_arb[i]) begin
					fill_ram_req_addr = fill_ram_req_addr | fill_addr_q[i];
					fill_ram_req_way = fill_ram_req_way | fill_way_q[i];
					fill_ram_req_data = fill_ram_req_data | fill_data_q[i];
				end
		end
	end
	always @(*) begin
		fill_out_data = 1'sb0;
		fill_out_err = 1'sb0;
		begin : sv2v_autoblock_5
			reg signed [31:0] i;
			for (i = 0; i < NUM_FB; i = i + 1)
				if (fill_data_reg[i]) begin
					fill_out_data = fill_out_data | fill_data_q[i];
					fill_out_err = fill_out_err | (fill_err_q[i * ibex_pkg_IC_LINE_BEATS+:ibex_pkg_IC_LINE_BEATS] & ~{ibex_pkg_IC_LINE_BEATS {fill_hit_q[i]}});
				end
		end
	end
	assign instr_req = ((~icache_enable_i | branch_i) & lookup_grant_ic0) | |fill_ext_req;
	assign instr_addr = (|fill_ext_req ? fill_ext_req_addr : lookup_addr_ic0[31:ibex_pkg_BUS_W]);
	assign instr_req_o = instr_req;
	assign instr_addr_o = {instr_addr[31:ibex_pkg_BUS_W], {ibex_pkg_BUS_W {1'b0}}};
	assign line_data = (|fill_data_hit ? hit_data_ic1 : fill_out_data);
	assign line_err = (|fill_data_hit ? {ibex_pkg_IC_LINE_BEATS {1'b0}} : fill_out_err);
	always @(*) begin
		line_data_muxed = 1'sb0;
		line_err_muxed = 1'b0;
		begin : sv2v_autoblock_6
			reg [31:0] i;
			for (i = 0; i < ibex_pkg_IC_LINE_BEATS; i = i + 1)
				if ((output_addr_q[2:ibex_pkg_BUS_W] + {{ibex_pkg_IC_LINE_BEATS_W - 1 {1'b0}}, skid_valid_q}) == i[ibex_pkg_IC_LINE_BEATS_W - 1:0]) begin
					line_data_muxed = line_data_muxed | line_data[i * 32+:32];
					line_err_muxed = line_err_muxed | line_err[i];
				end
		end
	end
	assign output_data = (|fill_data_rvd ? instr_rdata_i : line_data_muxed);
	assign output_err = (|fill_data_rvd ? instr_err_i : line_err_muxed);
	assign data_valid = |fill_out_arb;
	assign skid_data_d = output_data[31:16];
	assign skid_en = data_valid & (ready_i | skid_ready);
	generate
		if (ResetAll) begin : g_skid_data_ra
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni) begin
					skid_data_q <= 1'sb0;
					skid_err_q <= 1'sb0;
				end
				else if (skid_en) begin
					skid_data_q <= skid_data_d;
					skid_err_q <= output_err;
				end
		end
		else begin : g_skid_data_nr
			always @(posedge clk_i)
				if (skid_en) begin
					skid_data_q <= skid_data_d;
					skid_err_q <= output_err;
				end
		end
	endgenerate
	assign skid_complete_instr = skid_valid_q & ((skid_data_q[1:0] != 2'b11) | skid_err_q);
	assign skid_ready = (output_addr_q[1] & ~skid_valid_q) & (~output_compressed | output_err);
	assign output_ready = (ready_i | skid_ready) & ~skid_complete_instr;
	assign output_compressed = rdata_o[1:0] != 2'b11;
	assign skid_valid_d = (branch_i ? 1'b0 : (skid_valid_q ? ~(ready_i & ((skid_data_q[1:0] != 2'b11) | skid_err_q)) : data_valid & ((output_addr_q[1] & (~output_compressed | output_err)) | (((~output_addr_q[1] & output_compressed) & ~output_err) & ready_i))));
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			skid_valid_q <= 1'b0;
		else
			skid_valid_q <= skid_valid_d;
	assign output_valid = skid_complete_instr | (data_valid & (((~output_addr_q[1] | skid_valid_q) | output_err) | (output_data[17:16] != 2'b11)));
	assign output_addr_en = branch_i | (ready_i & valid_o);
	assign addr_incr_two = output_compressed & ~err_o;
	assign output_addr_incr = output_addr_q[31:1] + {29'd0, ~addr_incr_two, addr_incr_two};
	assign output_addr_d = (branch_i ? addr_i[31:1] : output_addr_incr);
	generate
		if (ResetAll) begin : g_output_addr_ra
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					output_addr_q <= 1'sb0;
				else if (output_addr_en)
					output_addr_q <= output_addr_d;
		end
		else begin : g_output_addr_nr
			always @(posedge clk_i)
				if (output_addr_en)
					output_addr_q <= output_addr_d;
		end
	endgenerate
	localparam [31:0] ibex_pkg_IC_OUTPUT_BEATS = 2;
	always @(*) begin
		output_data_lo = 1'sb0;
		begin : sv2v_autoblock_7
			reg [31:0] i;
			for (i = 0; i < ibex_pkg_IC_OUTPUT_BEATS; i = i + 1)
				if (output_addr_q[1:1] == i[0:0])
					output_data_lo = output_data_lo | output_data[i * 16+:16];
		end
	end
	always @(*) begin
		output_data_hi = 1'sb0;
		begin : sv2v_autoblock_8
			reg [31:0] i;
			for (i = 0; i < 1; i = i + 1)
				if (output_addr_q[1:1] == i[0:0])
					output_data_hi = output_data_hi | output_data[(i + 1) * 16+:16];
		end
		if (&output_addr_q[1:1])
			output_data_hi = output_data_hi | output_data[15:0];
	end
	assign valid_o = output_valid;
	assign rdata_o = {output_data_hi, (skid_valid_q ? skid_data_q : output_data_lo)};
	assign addr_o = {output_addr_q, 1'b0};
	assign err_o = (skid_valid_q & skid_err_q) | (~skid_complete_instr & output_err);
	assign err_plus2_o = skid_valid_q & ~skid_err_q;
	always @(*) begin
		inval_state_d = inval_state_q;
		inval_index_d = inval_index_q;
		inval_index_en = 1'b0;
		inval_write_req = 1'b0;
		ic_scr_key_req_o = 1'b0;
		inval_block_cache = 1'b1;
		case (inval_state_q)
			2'd0: begin
				inval_state_d = 2'd1;
				if (~ic_scr_key_valid_i)
					ic_scr_key_req_o = 1'b1;
			end
			2'd1:
				if (ic_scr_key_valid_i) begin
					inval_state_d = 2'd2;
					inval_index_d = 1'sb0;
					inval_index_en = 1'b1;
				end
			2'd2: begin
				inval_write_req = 1'b1;
				inval_index_d = inval_index_q + {{ibex_pkg_IC_INDEX_W - 1 {1'b0}}, 1'b1};
				inval_index_en = 1'b1;
				if (icache_inval_i) begin
					ic_scr_key_req_o = 1'b1;
					inval_state_d = 2'd1;
				end
				else if (&inval_index_q)
					inval_state_d = 2'd3;
			end
			2'd3:
				if (icache_inval_i) begin
					ic_scr_key_req_o = 1'b1;
					inval_state_d = 2'd1;
				end
				else
					inval_block_cache = 1'b0;
			default:
				;
		endcase
	end
	assign inval_active = inval_state_q != 2'd3;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			inval_state_q <= 2'd0;
		else
			inval_state_q <= inval_state_d;
	generate
		if (ResetAll) begin : g_inval_index_ra
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inval_index_q <= 1'sb0;
				else if (inval_index_en)
					inval_index_q <= inval_index_d;
		end
		else begin : g_inval_index_nr
			always @(posedge clk_i)
				if (inval_index_en)
					inval_index_q <= inval_index_d;
		end
	endgenerate
	assign busy_o = inval_active | |(fill_busy_q & ~fill_rvd_done);
endmodule
module ibex_id_stage (
	clk_i,
	rst_ni,
	ctrl_busy_o,
	illegal_insn_o,
	instr_valid_i,
	instr_rdata_i,
	instr_rdata_alu_i,
	instr_rdata_c_i,
	instr_is_compressed_i,
	instr_bp_taken_i,
	instr_req_o,
	instr_first_cycle_id_o,
	instr_valid_clear_o,
	id_in_ready_o,
	instr_exec_i,
	icache_inval_o,
	branch_decision_i,
	pc_set_o,
	pc_mux_o,
	nt_branch_mispredict_o,
	nt_branch_addr_o,
	exc_pc_mux_o,
	exc_cause_o,
	illegal_c_insn_i,
	instr_fetch_err_i,
	instr_fetch_err_plus2_i,
	pc_id_i,
	ex_valid_i,
	lsu_resp_valid_i,
	alu_operator_ex_o,
	alu_operand_a_ex_o,
	alu_operand_b_ex_o,
	imd_val_we_ex_i,
	imd_val_d_ex_i,
	imd_val_q_ex_o,
	bt_a_operand_o,
	bt_b_operand_o,
	mult_en_ex_o,
	div_en_ex_o,
	mult_sel_ex_o,
	div_sel_ex_o,
	multdiv_operator_ex_o,
	multdiv_signed_mode_ex_o,
	multdiv_operand_a_ex_o,
	multdiv_operand_b_ex_o,
	multdiv_ready_id_o,
	csr_access_o,
	csr_op_o,
	csr_op_en_o,
	csr_save_if_o,
	csr_save_id_o,
	csr_save_wb_o,
	csr_restore_mret_id_o,
	csr_restore_dret_id_o,
	csr_save_cause_o,
	csr_mtval_o,
	priv_mode_i,
	csr_mstatus_tw_i,
	illegal_csr_insn_i,
	data_ind_timing_i,
	lsu_req_o,
	lsu_we_o,
	lsu_type_o,
	lsu_sign_ext_o,
	lsu_wdata_o,
	lsu_req_done_i,
	lsu_addr_incr_req_i,
	lsu_addr_last_i,
	csr_mstatus_mie_i,
	irq_pending_i,
	irqs_i,
	irq_nm_i,
	nmi_mode_o,
	lsu_load_err_i,
	lsu_load_resp_intg_err_i,
	lsu_store_err_i,
	lsu_store_resp_intg_err_i,
	debug_mode_o,
	debug_mode_entering_o,
	debug_cause_o,
	debug_csr_save_o,
	debug_req_i,
	debug_single_step_i,
	debug_ebreakm_i,
	debug_ebreaku_i,
	trigger_match_i,
	result_ex_i,
	csr_rdata_i,
	rf_raddr_a_o,
	rf_rdata_a_i,
	rf_raddr_b_o,
	rf_rdata_b_i,
	rf_ren_a_o,
	rf_ren_b_o,
	rf_waddr_id_o,
	rf_wdata_id_o,
	rf_we_id_o,
	rf_rd_a_wb_match_o,
	rf_rd_b_wb_match_o,
	rf_waddr_wb_i,
	rf_wdata_fwd_wb_i,
	rf_write_wb_i,
	en_wb_o,
	instr_type_wb_o,
	instr_perf_count_id_o,
	ready_wb_i,
	outstanding_load_wb_i,
	outstanding_store_wb_i,
	perf_jump_o,
	perf_branch_o,
	perf_tbranch_o,
	perf_dside_wait_o,
	perf_mul_wait_o,
	perf_div_wait_o,
	instr_id_done_o
);
	parameter [0:0] RV32E = 0;
	parameter integer RV32M = 32'sd2;
	parameter integer RV32B = 32'sd0;
	parameter [0:0] DataIndTiming = 1'b0;
	parameter [0:0] BranchTargetALU = 0;
	parameter [0:0] WritebackStage = 0;
	parameter [0:0] BranchPredictor = 0;
	parameter [0:0] MemECC = 1'b0;
	input wire clk_i;
	input wire rst_ni;
	output wire ctrl_busy_o;
	output wire illegal_insn_o;
	input wire instr_valid_i;
	input wire [31:0] instr_rdata_i;
	input wire [31:0] instr_rdata_alu_i;
	input wire [15:0] instr_rdata_c_i;
	input wire instr_is_compressed_i;
	input wire instr_bp_taken_i;
	output wire instr_req_o;
	output wire instr_first_cycle_id_o;
	output wire instr_valid_clear_o;
	output wire id_in_ready_o;
	input wire instr_exec_i;
	output wire icache_inval_o;
	input wire branch_decision_i;
	output wire pc_set_o;
	output wire [2:0] pc_mux_o;
	output wire nt_branch_mispredict_o;
	output wire [31:0] nt_branch_addr_o;
	output wire [1:0] exc_pc_mux_o;
	output wire [6:0] exc_cause_o;
	input wire illegal_c_insn_i;
	input wire instr_fetch_err_i;
	input wire instr_fetch_err_plus2_i;
	input wire [31:0] pc_id_i;
	input wire ex_valid_i;
	input wire lsu_resp_valid_i;
	output wire [6:0] alu_operator_ex_o;
	output wire [31:0] alu_operand_a_ex_o;
	output wire [31:0] alu_operand_b_ex_o;
	input wire [1:0] imd_val_we_ex_i;
	input wire [67:0] imd_val_d_ex_i;
	output wire [67:0] imd_val_q_ex_o;
	output reg [31:0] bt_a_operand_o;
	output reg [31:0] bt_b_operand_o;
	output wire mult_en_ex_o;
	output wire div_en_ex_o;
	output wire mult_sel_ex_o;
	output wire div_sel_ex_o;
	output wire [1:0] multdiv_operator_ex_o;
	output wire [1:0] multdiv_signed_mode_ex_o;
	output wire [31:0] multdiv_operand_a_ex_o;
	output wire [31:0] multdiv_operand_b_ex_o;
	output wire multdiv_ready_id_o;
	output wire csr_access_o;
	output wire [1:0] csr_op_o;
	output wire csr_op_en_o;
	output wire csr_save_if_o;
	output wire csr_save_id_o;
	output wire csr_save_wb_o;
	output wire csr_restore_mret_id_o;
	output wire csr_restore_dret_id_o;
	output wire csr_save_cause_o;
	output wire [31:0] csr_mtval_o;
	input wire [1:0] priv_mode_i;
	input wire csr_mstatus_tw_i;
	input wire illegal_csr_insn_i;
	input wire data_ind_timing_i;
	output wire lsu_req_o;
	output wire lsu_we_o;
	output wire [1:0] lsu_type_o;
	output wire lsu_sign_ext_o;
	output wire [31:0] lsu_wdata_o;
	input wire lsu_req_done_i;
	input wire lsu_addr_incr_req_i;
	input wire [31:0] lsu_addr_last_i;
	input wire csr_mstatus_mie_i;
	input wire irq_pending_i;
	input wire [17:0] irqs_i;
	input wire irq_nm_i;
	output wire nmi_mode_o;
	input wire lsu_load_err_i;
	input wire lsu_load_resp_intg_err_i;
	input wire lsu_store_err_i;
	input wire lsu_store_resp_intg_err_i;
	output wire debug_mode_o;
	output wire debug_mode_entering_o;
	output wire [2:0] debug_cause_o;
	output wire debug_csr_save_o;
	input wire debug_req_i;
	input wire debug_single_step_i;
	input wire debug_ebreakm_i;
	input wire debug_ebreaku_i;
	input wire trigger_match_i;
	input wire [31:0] result_ex_i;
	input wire [31:0] csr_rdata_i;
	output wire [4:0] rf_raddr_a_o;
	input wire [31:0] rf_rdata_a_i;
	output wire [4:0] rf_raddr_b_o;
	input wire [31:0] rf_rdata_b_i;
	output wire rf_ren_a_o;
	output wire rf_ren_b_o;
	output wire [4:0] rf_waddr_id_o;
	output reg [31:0] rf_wdata_id_o;
	output wire rf_we_id_o;
	output wire rf_rd_a_wb_match_o;
	output wire rf_rd_b_wb_match_o;
	input wire [4:0] rf_waddr_wb_i;
	input wire [31:0] rf_wdata_fwd_wb_i;
	input wire rf_write_wb_i;
	output wire en_wb_o;
	output wire [1:0] instr_type_wb_o;
	output wire instr_perf_count_id_o;
	input wire ready_wb_i;
	input wire outstanding_load_wb_i;
	input wire outstanding_store_wb_i;
	output wire perf_jump_o;
	output reg perf_branch_o;
	output wire perf_tbranch_o;
	output wire perf_dside_wait_o;
	output wire perf_mul_wait_o;
	output wire perf_div_wait_o;
	output wire instr_id_done_o;
	wire illegal_insn_dec;
	wire illegal_dret_insn;
	wire illegal_umode_insn;
	wire ebrk_insn;
	wire mret_insn_dec;
	wire dret_insn_dec;
	wire ecall_insn_dec;
	wire wfi_insn_dec;
	wire wb_exception;
	wire id_exception;
	wire branch_in_dec;
	wire branch_set;
	wire branch_set_raw;
	reg branch_set_raw_d;
	reg branch_jump_set_done_q;
	wire branch_jump_set_done_d;
	reg branch_not_set;
	wire branch_taken;
	wire jump_in_dec;
	wire jump_set_dec;
	wire jump_set;
	reg jump_set_raw;
	wire instr_first_cycle;
	wire instr_executing_spec;
	wire instr_executing;
	wire instr_done;
	wire controller_run;
	wire stall_ld_hz;
	wire stall_mem;
	reg stall_multdiv;
	reg stall_branch;
	reg stall_jump;
	wire stall_id;
	wire stall_wb;
	wire flush_id;
	wire multicycle_done;
	wire mem_resp_intg_err;
	wire [31:0] imm_i_type;
	wire [31:0] imm_s_type;
	wire [31:0] imm_b_type;
	wire [31:0] imm_u_type;
	wire [31:0] imm_j_type;
	wire [31:0] zimm_rs1_type;
	wire [31:0] imm_a;
	reg [31:0] imm_b;
	wire rf_wdata_sel;
	wire rf_we_dec;
	reg rf_we_raw;
	wire rf_ren_a;
	wire rf_ren_b;
	wire rf_ren_a_dec;
	wire rf_ren_b_dec;
	assign rf_ren_a = ((instr_valid_i & ~instr_fetch_err_i) & ~illegal_insn_o) & rf_ren_a_dec;
	assign rf_ren_b = ((instr_valid_i & ~instr_fetch_err_i) & ~illegal_insn_o) & rf_ren_b_dec;
	assign rf_ren_a_o = rf_ren_a;
	assign rf_ren_b_o = rf_ren_b;
	wire [31:0] rf_rdata_a_fwd;
	wire [31:0] rf_rdata_b_fwd;
	wire [6:0] alu_operator;
	wire [1:0] alu_op_a_mux_sel;
	wire [1:0] alu_op_a_mux_sel_dec;
	wire alu_op_b_mux_sel;
	wire alu_op_b_mux_sel_dec;
	wire alu_multicycle_dec;
	reg stall_alu;
	reg [67:0] imd_val_q;
	wire [1:0] bt_a_mux_sel;
	wire [2:0] bt_b_mux_sel;
	wire imm_a_mux_sel;
	wire [2:0] imm_b_mux_sel;
	wire [2:0] imm_b_mux_sel_dec;
	wire mult_en_id;
	wire mult_en_dec;
	wire div_en_id;
	wire div_en_dec;
	wire multdiv_en_dec;
	wire [1:0] multdiv_operator;
	wire [1:0] multdiv_signed_mode;
	wire lsu_we;
	wire [1:0] lsu_type;
	wire lsu_sign_ext;
	wire lsu_req;
	wire lsu_req_dec;
	wire data_req_allowed;
	reg csr_pipe_flush;
	reg [31:0] alu_operand_a;
	wire [31:0] alu_operand_b;
	assign alu_op_a_mux_sel = (lsu_addr_incr_req_i ? 2'd1 : alu_op_a_mux_sel_dec);
	assign alu_op_b_mux_sel = (lsu_addr_incr_req_i ? 1'd1 : alu_op_b_mux_sel_dec);
	assign imm_b_mux_sel = (lsu_addr_incr_req_i ? 3'd6 : imm_b_mux_sel_dec);
	assign imm_a = (imm_a_mux_sel == 1'd0 ? zimm_rs1_type : {32 {1'sb0}});
	always @(*) begin : alu_operand_a_mux
		case (alu_op_a_mux_sel)
			2'd0: alu_operand_a = rf_rdata_a_fwd;
			2'd1: alu_operand_a = lsu_addr_last_i;
			2'd2: alu_operand_a = pc_id_i;
			2'd3: alu_operand_a = imm_a;
			default: alu_operand_a = pc_id_i;
		endcase
	end
	generate
		if (BranchTargetALU) begin : g_btalu_muxes
			always @(*) begin : bt_operand_a_mux
				case (bt_a_mux_sel)
					2'd0: bt_a_operand_o = rf_rdata_a_fwd;
					2'd2: bt_a_operand_o = pc_id_i;
					default: bt_a_operand_o = pc_id_i;
				endcase
			end
			always @(*) begin : bt_immediate_b_mux
				case (bt_b_mux_sel)
					3'd0: bt_b_operand_o = imm_i_type;
					3'd2: bt_b_operand_o = imm_b_type;
					3'd4: bt_b_operand_o = imm_j_type;
					3'd5: bt_b_operand_o = (instr_is_compressed_i ? 32'h00000002 : 32'h00000004);
					default: bt_b_operand_o = (instr_is_compressed_i ? 32'h00000002 : 32'h00000004);
				endcase
			end
			always @(*) begin : immediate_b_mux
				case (imm_b_mux_sel)
					3'd0: imm_b = imm_i_type;
					3'd1: imm_b = imm_s_type;
					3'd3: imm_b = imm_u_type;
					3'd5: imm_b = (instr_is_compressed_i ? 32'h00000002 : 32'h00000004);
					3'd6: imm_b = 32'h00000004;
					default: imm_b = 32'h00000004;
				endcase
			end
		end
		else begin : g_nobtalu
			wire [1:0] unused_a_mux_sel;
			wire [2:0] unused_b_mux_sel;
			assign unused_a_mux_sel = bt_a_mux_sel;
			assign unused_b_mux_sel = bt_b_mux_sel;
			wire [32:1] sv2v_tmp_FACAA;
			assign sv2v_tmp_FACAA = 1'sb0;
			always @(*) bt_a_operand_o = sv2v_tmp_FACAA;
			wire [32:1] sv2v_tmp_A4AF9;
			assign sv2v_tmp_A4AF9 = 1'sb0;
			always @(*) bt_b_operand_o = sv2v_tmp_A4AF9;
			always @(*) begin : immediate_b_mux
				case (imm_b_mux_sel)
					3'd0: imm_b = imm_i_type;
					3'd1: imm_b = imm_s_type;
					3'd2: imm_b = imm_b_type;
					3'd3: imm_b = imm_u_type;
					3'd4: imm_b = imm_j_type;
					3'd5: imm_b = (instr_is_compressed_i ? 32'h00000002 : 32'h00000004);
					3'd6: imm_b = 32'h00000004;
					default: imm_b = 32'h00000004;
				endcase
			end
		end
	endgenerate
	assign alu_operand_b = (alu_op_b_mux_sel == 1'd1 ? imm_b : rf_rdata_b_fwd);
	genvar i;
	generate
		for (i = 0; i < 2; i = i + 1) begin : gen_intermediate_val_reg
			always @(posedge clk_i or negedge rst_ni) begin : intermediate_val_reg
				if (!rst_ni)
					imd_val_q[(1 - i) * 34+:34] <= 1'sb0;
				else if (imd_val_we_ex_i[i])
					imd_val_q[(1 - i) * 34+:34] <= imd_val_d_ex_i[(1 - i) * 34+:34];
			end
		end
	endgenerate
	assign imd_val_q_ex_o = imd_val_q;
	assign rf_we_id_o = (rf_we_raw & instr_executing) & ~illegal_csr_insn_i;
	always @(*) begin : rf_wdata_id_mux
		case (rf_wdata_sel)
			1'd0: rf_wdata_id_o = result_ex_i;
			1'd1: rf_wdata_id_o = csr_rdata_i;
			default: rf_wdata_id_o = result_ex_i;
		endcase
	end
	ibex_decoder #(
		.RV32E(RV32E),
		.RV32M(RV32M),
		.RV32B(RV32B),
		.BranchTargetALU(BranchTargetALU)
	) decoder_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.illegal_insn_o(illegal_insn_dec),
		.ebrk_insn_o(ebrk_insn),
		.mret_insn_o(mret_insn_dec),
		.dret_insn_o(dret_insn_dec),
		.ecall_insn_o(ecall_insn_dec),
		.wfi_insn_o(wfi_insn_dec),
		.jump_set_o(jump_set_dec),
		.branch_taken_i(branch_taken),
		.icache_inval_o(icache_inval_o),
		.instr_first_cycle_i(instr_first_cycle),
		.instr_rdata_i(instr_rdata_i),
		.instr_rdata_alu_i(instr_rdata_alu_i),
		.illegal_c_insn_i(illegal_c_insn_i),
		.imm_a_mux_sel_o(imm_a_mux_sel),
		.imm_b_mux_sel_o(imm_b_mux_sel_dec),
		.bt_a_mux_sel_o(bt_a_mux_sel),
		.bt_b_mux_sel_o(bt_b_mux_sel),
		.imm_i_type_o(imm_i_type),
		.imm_s_type_o(imm_s_type),
		.imm_b_type_o(imm_b_type),
		.imm_u_type_o(imm_u_type),
		.imm_j_type_o(imm_j_type),
		.zimm_rs1_type_o(zimm_rs1_type),
		.rf_wdata_sel_o(rf_wdata_sel),
		.rf_we_o(rf_we_dec),
		.rf_raddr_a_o(rf_raddr_a_o),
		.rf_raddr_b_o(rf_raddr_b_o),
		.rf_waddr_o(rf_waddr_id_o),
		.rf_ren_a_o(rf_ren_a_dec),
		.rf_ren_b_o(rf_ren_b_dec),
		.alu_operator_o(alu_operator),
		.alu_op_a_mux_sel_o(alu_op_a_mux_sel_dec),
		.alu_op_b_mux_sel_o(alu_op_b_mux_sel_dec),
		.alu_multicycle_o(alu_multicycle_dec),
		.mult_en_o(mult_en_dec),
		.div_en_o(div_en_dec),
		.mult_sel_o(mult_sel_ex_o),
		.div_sel_o(div_sel_ex_o),
		.multdiv_operator_o(multdiv_operator),
		.multdiv_signed_mode_o(multdiv_signed_mode),
		.csr_access_o(csr_access_o),
		.csr_op_o(csr_op_o),
		.data_req_o(lsu_req_dec),
		.data_we_o(lsu_we),
		.data_type_o(lsu_type),
		.data_sign_extension_o(lsu_sign_ext),
		.jump_in_dec_o(jump_in_dec),
		.branch_in_dec_o(branch_in_dec)
	);
	always @(*) begin : csr_pipeline_flushes
		csr_pipe_flush = 1'b0;
		if ((csr_op_en_o == 1'b1) && ((csr_op_o == 2'd1) || (csr_op_o == 2'd2))) begin
			if ((((instr_rdata_i[31:20] == 12'h300) || (instr_rdata_i[31:20] == 12'h304)) || (instr_rdata_i[31:20] == 12'h747)) || (instr_rdata_i[31:25] == 7'h1d))
				csr_pipe_flush = 1'b1;
		end
		else if ((csr_op_en_o == 1'b1) && (csr_op_o != 2'd0))
			if ((((instr_rdata_i[31:20] == 12'h7b0) || (instr_rdata_i[31:20] == 12'h7b1)) || (instr_rdata_i[31:20] == 12'h7b2)) || (instr_rdata_i[31:20] == 12'h7b3))
				csr_pipe_flush = 1'b1;
	end
	assign illegal_dret_insn = dret_insn_dec & ~debug_mode_o;
	assign illegal_umode_insn = (priv_mode_i != 2'b11) & (mret_insn_dec | (csr_mstatus_tw_i & wfi_insn_dec));
	assign illegal_insn_o = instr_valid_i & (((illegal_insn_dec | illegal_csr_insn_i) | illegal_dret_insn) | illegal_umode_insn);
	assign mem_resp_intg_err = lsu_load_resp_intg_err_i | lsu_store_resp_intg_err_i;
	ibex_controller #(
		.WritebackStage(WritebackStage),
		.BranchPredictor(BranchPredictor),
		.MemECC(MemECC)
	) controller_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.ctrl_busy_o(ctrl_busy_o),
		.illegal_insn_i(illegal_insn_o),
		.ecall_insn_i(ecall_insn_dec),
		.mret_insn_i(mret_insn_dec),
		.dret_insn_i(dret_insn_dec),
		.wfi_insn_i(wfi_insn_dec),
		.ebrk_insn_i(ebrk_insn),
		.csr_pipe_flush_i(csr_pipe_flush),
		.instr_valid_i(instr_valid_i),
		.instr_i(instr_rdata_i),
		.instr_compressed_i(instr_rdata_c_i),
		.instr_is_compressed_i(instr_is_compressed_i),
		.instr_bp_taken_i(instr_bp_taken_i),
		.instr_fetch_err_i(instr_fetch_err_i),
		.instr_fetch_err_plus2_i(instr_fetch_err_plus2_i),
		.pc_id_i(pc_id_i),
		.instr_valid_clear_o(instr_valid_clear_o),
		.id_in_ready_o(id_in_ready_o),
		.controller_run_o(controller_run),
		.instr_exec_i(instr_exec_i),
		.instr_req_o(instr_req_o),
		.pc_set_o(pc_set_o),
		.pc_mux_o(pc_mux_o),
		.nt_branch_mispredict_o(nt_branch_mispredict_o),
		.exc_pc_mux_o(exc_pc_mux_o),
		.exc_cause_o(exc_cause_o),
		.lsu_addr_last_i(lsu_addr_last_i),
		.load_err_i(lsu_load_err_i),
		.mem_resp_intg_err_i(mem_resp_intg_err),
		.store_err_i(lsu_store_err_i),
		.wb_exception_o(wb_exception),
		.id_exception_o(id_exception),
		.branch_set_i(branch_set),
		.branch_not_set_i(branch_not_set),
		.jump_set_i(jump_set),
		.csr_mstatus_mie_i(csr_mstatus_mie_i),
		.irq_pending_i(irq_pending_i),
		.irqs_i(irqs_i),
		.irq_nm_ext_i(irq_nm_i),
		.nmi_mode_o(nmi_mode_o),
		.csr_save_if_o(csr_save_if_o),
		.csr_save_id_o(csr_save_id_o),
		.csr_save_wb_o(csr_save_wb_o),
		.csr_restore_mret_id_o(csr_restore_mret_id_o),
		.csr_restore_dret_id_o(csr_restore_dret_id_o),
		.csr_save_cause_o(csr_save_cause_o),
		.csr_mtval_o(csr_mtval_o),
		.priv_mode_i(priv_mode_i),
		.debug_mode_o(debug_mode_o),
		.debug_mode_entering_o(debug_mode_entering_o),
		.debug_cause_o(debug_cause_o),
		.debug_csr_save_o(debug_csr_save_o),
		.debug_req_i(debug_req_i),
		.debug_single_step_i(debug_single_step_i),
		.debug_ebreakm_i(debug_ebreakm_i),
		.debug_ebreaku_i(debug_ebreaku_i),
		.trigger_match_i(trigger_match_i),
		.stall_id_i(stall_id),
		.stall_wb_i(stall_wb),
		.flush_id_o(flush_id),
		.ready_wb_i(ready_wb_i),
		.perf_jump_o(perf_jump_o),
		.perf_tbranch_o(perf_tbranch_o)
	);
	assign multdiv_en_dec = mult_en_dec | div_en_dec;
	assign lsu_req = (instr_executing ? data_req_allowed & lsu_req_dec : 1'b0);
	assign mult_en_id = (instr_executing ? mult_en_dec : 1'b0);
	assign div_en_id = (instr_executing ? div_en_dec : 1'b0);
	assign lsu_req_o = lsu_req;
	assign lsu_we_o = lsu_we;
	assign lsu_type_o = lsu_type;
	assign lsu_sign_ext_o = lsu_sign_ext;
	assign lsu_wdata_o = rf_rdata_b_fwd;
	assign csr_op_en_o = (csr_access_o & instr_executing) & instr_id_done_o;
	assign alu_operator_ex_o = alu_operator;
	assign alu_operand_a_ex_o = alu_operand_a;
	assign alu_operand_b_ex_o = alu_operand_b;
	assign mult_en_ex_o = mult_en_id;
	assign div_en_ex_o = div_en_id;
	assign multdiv_operator_ex_o = multdiv_operator;
	assign multdiv_signed_mode_ex_o = multdiv_signed_mode;
	assign multdiv_operand_a_ex_o = rf_rdata_a_fwd;
	assign multdiv_operand_b_ex_o = rf_rdata_b_fwd;
	generate
		if (BranchTargetALU && !DataIndTiming) begin : g_branch_set_direct
			assign branch_set_raw = branch_set_raw_d;
		end
		else begin : g_branch_set_flop
			reg branch_set_raw_q;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					branch_set_raw_q <= 1'b0;
				else
					branch_set_raw_q <= branch_set_raw_d;
			assign branch_set_raw = (BranchTargetALU && !data_ind_timing_i ? branch_set_raw_d : branch_set_raw_q);
		end
	endgenerate
	assign branch_jump_set_done_d = ((branch_set_raw | jump_set_raw) | branch_jump_set_done_q) & ~instr_valid_clear_o;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			branch_jump_set_done_q <= 1'b0;
		else
			branch_jump_set_done_q <= branch_jump_set_done_d;
	assign jump_set = jump_set_raw & ~branch_jump_set_done_q;
	assign branch_set = branch_set_raw & ~branch_jump_set_done_q;
	generate
		if (DataIndTiming) begin : g_sec_branch_taken
			reg branch_taken_q;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					branch_taken_q <= 1'b0;
				else
					branch_taken_q <= branch_decision_i;
			assign branch_taken = ~data_ind_timing_i | branch_taken_q;
		end
		else begin : g_nosec_branch_taken
			assign branch_taken = 1'b1;
		end
		if (BranchPredictor) begin : g_calc_nt_addr
			assign nt_branch_addr_o = pc_id_i + (instr_is_compressed_i ? 32'd2 : 32'd4);
		end
		else begin : g_n_calc_nt_addr
			assign nt_branch_addr_o = 32'd0;
		end
	endgenerate
	reg id_fsm_q;
	reg id_fsm_d;
	always @(posedge clk_i or negedge rst_ni) begin : id_pipeline_reg
		if (!rst_ni)
			id_fsm_q <= 1'd0;
		else if (instr_executing)
			id_fsm_q <= id_fsm_d;
	end
	always @(*) begin
		id_fsm_d = id_fsm_q;
		rf_we_raw = rf_we_dec;
		stall_multdiv = 1'b0;
		stall_jump = 1'b0;
		stall_branch = 1'b0;
		stall_alu = 1'b0;
		branch_set_raw_d = 1'b0;
		branch_not_set = 1'b0;
		jump_set_raw = 1'b0;
		perf_branch_o = 1'b0;
		if (instr_executing_spec)
			case (id_fsm_q)
				1'd0:
					case (1'b1)
						lsu_req_dec:
							if (!WritebackStage)
								id_fsm_d = 1'd1;
							else if (~lsu_req_done_i)
								id_fsm_d = 1'd1;
						multdiv_en_dec:
							if (~ex_valid_i) begin
								id_fsm_d = 1'd1;
								rf_we_raw = 1'b0;
								stall_multdiv = 1'b1;
							end
						branch_in_dec: begin
							id_fsm_d = (data_ind_timing_i || (!BranchTargetALU && branch_decision_i) ? 1'd1 : 1'd0);
							stall_branch = (~BranchTargetALU & branch_decision_i) | data_ind_timing_i;
							branch_set_raw_d = branch_decision_i | data_ind_timing_i;
							if (BranchPredictor)
								branch_not_set = ~branch_decision_i;
							perf_branch_o = 1'b1;
						end
						jump_in_dec: begin
							id_fsm_d = (BranchTargetALU ? 1'd0 : 1'd1);
							stall_jump = ~BranchTargetALU;
							jump_set_raw = jump_set_dec;
						end
						alu_multicycle_dec: begin
							stall_alu = 1'b1;
							id_fsm_d = 1'd1;
							rf_we_raw = 1'b0;
						end
						default: id_fsm_d = 1'd0;
					endcase
				1'd1: begin
					if (multdiv_en_dec)
						rf_we_raw = rf_we_dec & ex_valid_i;
					if (multicycle_done & ready_wb_i)
						id_fsm_d = 1'd0;
					else begin
						stall_multdiv = multdiv_en_dec;
						stall_branch = branch_in_dec;
						stall_jump = jump_in_dec;
					end
				end
				default: id_fsm_d = 1'd0;
			endcase
	end
	assign multdiv_ready_id_o = ready_wb_i;
	assign stall_id = ((((stall_ld_hz | stall_mem) | stall_multdiv) | stall_jump) | stall_branch) | stall_alu;
	assign instr_done = (~stall_id & ~flush_id) & instr_executing;
	assign instr_first_cycle = instr_valid_i & (id_fsm_q == 1'd0);
	assign instr_first_cycle_id_o = instr_first_cycle;
	generate
		if (WritebackStage) begin : gen_stall_mem
			wire rf_rd_a_wb_match;
			wire rf_rd_b_wb_match;
			wire rf_rd_a_hz;
			wire rf_rd_b_hz;
			wire outstanding_memory_access;
			wire instr_kill;
			assign multicycle_done = (lsu_req_dec ? ~stall_mem : ex_valid_i);
			assign outstanding_memory_access = (outstanding_load_wb_i | outstanding_store_wb_i) & ~lsu_resp_valid_i;
			assign data_req_allowed = ~outstanding_memory_access;
			assign instr_kill = ((instr_fetch_err_i | wb_exception) | id_exception) | ~controller_run;
			assign instr_executing_spec = ((instr_valid_i & ~instr_fetch_err_i) & controller_run) & ~stall_ld_hz;
			assign instr_executing = ((instr_valid_i & ~instr_kill) & ~stall_ld_hz) & ~outstanding_memory_access;
			assign stall_mem = instr_valid_i & (outstanding_memory_access | (lsu_req_dec & ~lsu_req_done_i));
			assign rf_rd_a_wb_match = (rf_waddr_wb_i == rf_raddr_a_o) & |rf_raddr_a_o;
			assign rf_rd_b_wb_match = (rf_waddr_wb_i == rf_raddr_b_o) & |rf_raddr_b_o;
			assign rf_rd_a_wb_match_o = rf_rd_a_wb_match;
			assign rf_rd_b_wb_match_o = rf_rd_b_wb_match;
			assign rf_rd_a_hz = rf_rd_a_wb_match & rf_ren_a;
			assign rf_rd_b_hz = rf_rd_b_wb_match & rf_ren_b;
			assign rf_rdata_a_fwd = (rf_rd_a_wb_match & rf_write_wb_i ? rf_wdata_fwd_wb_i : rf_rdata_a_i);
			assign rf_rdata_b_fwd = (rf_rd_b_wb_match & rf_write_wb_i ? rf_wdata_fwd_wb_i : rf_rdata_b_i);
			assign stall_ld_hz = outstanding_load_wb_i & (rf_rd_a_hz | rf_rd_b_hz);
			assign instr_type_wb_o = (~lsu_req_dec ? 2'd2 : (lsu_we ? 2'd1 : 2'd0));
			assign instr_id_done_o = en_wb_o & ready_wb_i;
			assign stall_wb = en_wb_o & ~ready_wb_i;
			assign perf_dside_wait_o = (instr_valid_i & ~instr_kill) & (outstanding_memory_access | stall_ld_hz);
		end
		else begin : gen_no_stall_mem
			assign multicycle_done = (lsu_req_dec ? lsu_resp_valid_i : ex_valid_i);
			assign data_req_allowed = instr_first_cycle;
			assign stall_mem = instr_valid_i & (lsu_req_dec & (~lsu_resp_valid_i | instr_first_cycle));
			assign stall_ld_hz = 1'b0;
			assign instr_executing_spec = (instr_valid_i & ~instr_fetch_err_i) & controller_run;
			assign instr_executing = instr_executing_spec;
			assign rf_rdata_a_fwd = rf_rdata_a_i;
			assign rf_rdata_b_fwd = rf_rdata_b_i;
			assign rf_rd_a_wb_match_o = 1'b0;
			assign rf_rd_b_wb_match_o = 1'b0;
			wire unused_data_req_done_ex;
			wire [4:0] unused_rf_waddr_wb;
			wire unused_rf_write_wb;
			wire unused_outstanding_load_wb;
			wire unused_outstanding_store_wb;
			wire unused_wb_exception;
			wire [31:0] unused_rf_wdata_fwd_wb;
			wire unused_id_exception;
			assign unused_data_req_done_ex = lsu_req_done_i;
			assign unused_rf_waddr_wb = rf_waddr_wb_i;
			assign unused_rf_write_wb = rf_write_wb_i;
			assign unused_outstanding_load_wb = outstanding_load_wb_i;
			assign unused_outstanding_store_wb = outstanding_store_wb_i;
			assign unused_wb_exception = wb_exception;
			assign unused_rf_wdata_fwd_wb = rf_wdata_fwd_wb_i;
			assign unused_id_exception = id_exception;
			assign instr_type_wb_o = 2'd2;
			assign stall_wb = 1'b0;
			assign perf_dside_wait_o = (instr_executing & lsu_req_dec) & ~lsu_resp_valid_i;
			assign instr_id_done_o = instr_done;
		end
	endgenerate
	assign instr_perf_count_id_o = (((~ebrk_insn & ~ecall_insn_dec) & ~illegal_insn_dec) & ~illegal_csr_insn_i) & ~instr_fetch_err_i;
	assign en_wb_o = instr_done;
	assign perf_mul_wait_o = stall_multdiv & mult_en_dec;
	assign perf_div_wait_o = stall_multdiv & div_en_dec;
endmodule
module ibex_if_stage (
	clk_i,
	rst_ni,
	boot_addr_i,
	req_i,
	instr_req_o,
	instr_addr_o,
	instr_gnt_i,
	instr_rvalid_i,
	instr_rdata_i,
	instr_bus_err_i,
	instr_intg_err_o,
	ic_tag_req_o,
	ic_tag_write_o,
	ic_tag_addr_o,
	ic_tag_wdata_o,
	ic_tag_rdata_i,
	ic_data_req_o,
	ic_data_write_o,
	ic_data_addr_o,
	ic_data_wdata_o,
	ic_data_rdata_i,
	ic_scr_key_valid_i,
	ic_scr_key_req_o,
	instr_valid_id_o,
	instr_new_id_o,
	instr_rdata_id_o,
	instr_rdata_alu_id_o,
	instr_rdata_c_id_o,
	instr_is_compressed_id_o,
	instr_bp_taken_o,
	instr_fetch_err_o,
	instr_fetch_err_plus2_o,
	illegal_c_insn_id_o,
	dummy_instr_id_o,
	pc_if_o,
	pc_id_o,
	pmp_err_if_i,
	pmp_err_if_plus2_i,
	instr_valid_clear_i,
	pc_set_i,
	pc_mux_i,
	nt_branch_mispredict_i,
	nt_branch_addr_i,
	exc_pc_mux_i,
	exc_cause,
	dummy_instr_en_i,
	dummy_instr_mask_i,
	dummy_instr_seed_en_i,
	dummy_instr_seed_i,
	icache_enable_i,
	icache_inval_i,
	icache_ecc_error_o,
	branch_target_ex_i,
	csr_mepc_i,
	csr_depc_i,
	csr_mtvec_i,
	csr_mtvec_init_o,
	id_in_ready_i,
	pc_mismatch_alert_o,
	if_busy_o
);
	parameter [31:0] DmHaltAddr = 32'h1a110800;
	parameter [31:0] DmExceptionAddr = 32'h1a110808;
	parameter [0:0] DummyInstructions = 1'b0;
	parameter [0:0] ICache = 1'b0;
	parameter [0:0] ICacheECC = 1'b0;
	localparam [31:0] ibex_pkg_BUS_SIZE = 32;
	parameter [31:0] BusSizeECC = ibex_pkg_BUS_SIZE;
	localparam [31:0] ibex_pkg_ADDR_W = 32;
	localparam [31:0] ibex_pkg_IC_LINE_SIZE = 64;
	localparam [31:0] ibex_pkg_IC_LINE_BYTES = 8;
	localparam [31:0] ibex_pkg_IC_NUM_WAYS = 2;
	localparam [31:0] ibex_pkg_IC_SIZE_BYTES = 4096;
	localparam [31:0] ibex_pkg_IC_NUM_LINES = (ibex_pkg_IC_SIZE_BYTES / ibex_pkg_IC_NUM_WAYS) / ibex_pkg_IC_LINE_BYTES;
	localparam [31:0] ibex_pkg_IC_INDEX_W = $clog2(ibex_pkg_IC_NUM_LINES);
	localparam [31:0] ibex_pkg_IC_LINE_W = 3;
	localparam [31:0] ibex_pkg_IC_TAG_SIZE = ((ibex_pkg_ADDR_W - ibex_pkg_IC_INDEX_W) - ibex_pkg_IC_LINE_W) + 1;
	parameter [31:0] TagSizeECC = ibex_pkg_IC_TAG_SIZE;
	parameter [31:0] LineSizeECC = ibex_pkg_IC_LINE_SIZE;
	parameter [0:0] PCIncrCheck = 1'b0;
	parameter [0:0] ResetAll = 1'b0;
	localparam signed [31:0] ibex_pkg_LfsrWidth = 32;
	localparam [31:0] ibex_pkg_RndCnstLfsrSeedDefault = 32'hac533bf4;
	parameter [31:0] RndCnstLfsrSeed = ibex_pkg_RndCnstLfsrSeedDefault;
	localparam [159:0] ibex_pkg_RndCnstLfsrPermDefault = 160'h1e35ecba467fd1b12e958152c04fa43878a8daed;
	parameter [159:0] RndCnstLfsrPerm = ibex_pkg_RndCnstLfsrPermDefault;
	parameter [0:0] BranchPredictor = 1'b0;
	parameter [0:0] MemECC = 1'b0;
	parameter [31:0] MemDataWidth = (MemECC ? 39 : 32);
	input wire clk_i;
	input wire rst_ni;
	input wire [31:0] boot_addr_i;
	input wire req_i;
	output wire instr_req_o;
	output wire [31:0] instr_addr_o;
	input wire instr_gnt_i;
	input wire instr_rvalid_i;
	input wire [MemDataWidth - 1:0] instr_rdata_i;
	input wire instr_bus_err_i;
	output wire instr_intg_err_o;
	output wire [1:0] ic_tag_req_o;
	output wire ic_tag_write_o;
	output wire [ibex_pkg_IC_INDEX_W - 1:0] ic_tag_addr_o;
	output wire [TagSizeECC - 1:0] ic_tag_wdata_o;
	input wire [(ibex_pkg_IC_NUM_WAYS * TagSizeECC) - 1:0] ic_tag_rdata_i;
	output wire [1:0] ic_data_req_o;
	output wire ic_data_write_o;
	output wire [ibex_pkg_IC_INDEX_W - 1:0] ic_data_addr_o;
	output wire [LineSizeECC - 1:0] ic_data_wdata_o;
	input wire [(ibex_pkg_IC_NUM_WAYS * LineSizeECC) - 1:0] ic_data_rdata_i;
	input wire ic_scr_key_valid_i;
	output wire ic_scr_key_req_o;
	output wire instr_valid_id_o;
	output wire instr_new_id_o;
	output reg [31:0] instr_rdata_id_o;
	output reg [31:0] instr_rdata_alu_id_o;
	output reg [15:0] instr_rdata_c_id_o;
	output reg instr_is_compressed_id_o;
	output wire instr_bp_taken_o;
	output reg instr_fetch_err_o;
	output reg instr_fetch_err_plus2_o;
	output reg illegal_c_insn_id_o;
	output reg dummy_instr_id_o;
	output wire [31:0] pc_if_o;
	output reg [31:0] pc_id_o;
	input wire pmp_err_if_i;
	input wire pmp_err_if_plus2_i;
	input wire instr_valid_clear_i;
	input wire pc_set_i;
	input wire [2:0] pc_mux_i;
	input wire nt_branch_mispredict_i;
	input wire [31:0] nt_branch_addr_i;
	input wire [1:0] exc_pc_mux_i;
	input wire [6:0] exc_cause;
	input wire dummy_instr_en_i;
	input wire [2:0] dummy_instr_mask_i;
	input wire dummy_instr_seed_en_i;
	input wire [31:0] dummy_instr_seed_i;
	input wire icache_enable_i;
	input wire icache_inval_i;
	output wire icache_ecc_error_o;
	input wire [31:0] branch_target_ex_i;
	input wire [31:0] csr_mepc_i;
	input wire [31:0] csr_depc_i;
	input wire [31:0] csr_mtvec_i;
	output wire csr_mtvec_init_o;
	input wire id_in_ready_i;
	output wire pc_mismatch_alert_o;
	output wire if_busy_o;
	wire instr_valid_id_d;
	reg instr_valid_id_q;
	wire instr_new_id_d;
	reg instr_new_id_q;
	wire instr_err;
	wire instr_intg_err;
	wire prefetch_busy;
	wire branch_req;
	reg [31:0] fetch_addr_n;
	wire unused_fetch_addr_n0;
	wire prefetch_branch;
	wire [31:0] prefetch_addr;
	wire fetch_valid_raw;
	wire fetch_valid;
	wire fetch_ready;
	wire [31:0] fetch_rdata;
	wire [31:0] fetch_addr;
	wire fetch_err;
	wire fetch_err_plus2;
	wire [31:0] instr_decompressed;
	wire illegal_c_insn;
	wire instr_is_compressed;
	wire if_instr_valid;
	wire [31:0] if_instr_rdata;
	wire [31:0] if_instr_addr;
	wire if_instr_bus_err;
	wire if_instr_pmp_err;
	wire if_instr_err;
	wire if_instr_err_plus2;
	reg [31:0] exc_pc;
	wire if_id_pipe_reg_we;
	wire stall_dummy_instr;
	wire [31:0] instr_out;
	wire instr_is_compressed_out;
	wire illegal_c_instr_out;
	wire instr_err_out;
	wire predict_branch_taken;
	wire [31:0] predict_branch_pc;
	reg [4:0] irq_vec;
	wire [2:0] pc_mux_internal;
	wire [7:0] unused_boot_addr;
	wire [7:0] unused_csr_mtvec;
	wire unused_exc_cause;
	assign unused_boot_addr = boot_addr_i[7:0];
	assign unused_csr_mtvec = csr_mtvec_i[7:0];
	assign unused_exc_cause = |{exc_cause[5], exc_cause[6]};
	localparam [6:0] ibex_pkg_ExcCauseIrqNm = 7'b0111111;
	always @(*) begin : exc_pc_mux
		irq_vec = exc_cause[4-:5];
		if (exc_cause[6])
			irq_vec = ibex_pkg_ExcCauseIrqNm[4-:5];
		case (exc_pc_mux_i)
			2'd0: exc_pc = {csr_mtvec_i[31:8], 8'h00};
			2'd1: exc_pc = {csr_mtvec_i[31:8], 1'b0, irq_vec, 2'b00};
			2'd2: exc_pc = DmHaltAddr;
			2'd3: exc_pc = DmExceptionAddr;
			default: exc_pc = {csr_mtvec_i[31:8], 8'h00};
		endcase
	end
	assign pc_mux_internal = ((BranchPredictor && predict_branch_taken) && !pc_set_i ? 3'd5 : pc_mux_i);
	always @(*) begin : fetch_addr_mux
		case (pc_mux_internal)
			3'd0: fetch_addr_n = {boot_addr_i[31:8], 8'h80};
			3'd1: fetch_addr_n = branch_target_ex_i;
			3'd2: fetch_addr_n = exc_pc;
			3'd3: fetch_addr_n = csr_mepc_i;
			3'd4: fetch_addr_n = csr_depc_i;
			3'd5: fetch_addr_n = (BranchPredictor ? predict_branch_pc : {boot_addr_i[31:8], 8'h80});
			default: fetch_addr_n = {boot_addr_i[31:8], 8'h80};
		endcase
	end
	assign csr_mtvec_init_o = (pc_mux_i == 3'd0) & pc_set_i;
	generate
		if (MemECC) begin : g_mem_ecc
			wire [1:0] ecc_err;
			wire [MemDataWidth - 1:0] instr_rdata_buf;
			prim_buf #(.Width(MemDataWidth)) u_prim_buf_instr_rdata(
				.in_i(instr_rdata_i),
				.out_o(instr_rdata_buf)
			);
			prim_secded_inv_39_32_dec u_instr_intg_dec(
				.data_i(instr_rdata_buf),
				.err_o(ecc_err)
			);
			assign instr_intg_err = |ecc_err;
		end
		else begin : g_no_mem_ecc
			assign instr_intg_err = 1'b0;
		end
	endgenerate
	assign instr_err = instr_intg_err | instr_bus_err_i;
	assign instr_intg_err_o = instr_intg_err & instr_rvalid_i;
	assign prefetch_branch = branch_req | nt_branch_mispredict_i;
	assign prefetch_addr = (branch_req ? {fetch_addr_n[31:1], 1'b0} : nt_branch_addr_i);
	assign fetch_valid = fetch_valid_raw & ~nt_branch_mispredict_i;
	generate
		if (ICache) begin : gen_icache
			ibex_icache #(
				.ICacheECC(ICacheECC),
				.ResetAll(ResetAll),
				.BusSizeECC(BusSizeECC),
				.TagSizeECC(TagSizeECC),
				.LineSizeECC(LineSizeECC)
			) icache_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_i(req_i),
				.branch_i(prefetch_branch),
				.addr_i(prefetch_addr),
				.ready_i(fetch_ready),
				.valid_o(fetch_valid_raw),
				.rdata_o(fetch_rdata),
				.addr_o(fetch_addr),
				.err_o(fetch_err),
				.err_plus2_o(fetch_err_plus2),
				.instr_req_o(instr_req_o),
				.instr_addr_o(instr_addr_o),
				.instr_gnt_i(instr_gnt_i),
				.instr_rvalid_i(instr_rvalid_i),
				.instr_rdata_i(instr_rdata_i[31:0]),
				.instr_err_i(instr_err),
				.ic_tag_req_o(ic_tag_req_o),
				.ic_tag_write_o(ic_tag_write_o),
				.ic_tag_addr_o(ic_tag_addr_o),
				.ic_tag_wdata_o(ic_tag_wdata_o),
				.ic_tag_rdata_i(ic_tag_rdata_i),
				.ic_data_req_o(ic_data_req_o),
				.ic_data_write_o(ic_data_write_o),
				.ic_data_addr_o(ic_data_addr_o),
				.ic_data_wdata_o(ic_data_wdata_o),
				.ic_data_rdata_i(ic_data_rdata_i),
				.ic_scr_key_valid_i(ic_scr_key_valid_i),
				.ic_scr_key_req_o(ic_scr_key_req_o),
				.icache_enable_i(icache_enable_i),
				.icache_inval_i(icache_inval_i),
				.busy_o(prefetch_busy),
				.ecc_error_o(icache_ecc_error_o)
			);
		end
		else begin : gen_prefetch_buffer
			ibex_prefetch_buffer #(.ResetAll(ResetAll)) prefetch_buffer_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_i(req_i),
				.branch_i(prefetch_branch),
				.addr_i(prefetch_addr),
				.ready_i(fetch_ready),
				.valid_o(fetch_valid_raw),
				.rdata_o(fetch_rdata),
				.addr_o(fetch_addr),
				.err_o(fetch_err),
				.err_plus2_o(fetch_err_plus2),
				.instr_req_o(instr_req_o),
				.instr_addr_o(instr_addr_o),
				.instr_gnt_i(instr_gnt_i),
				.instr_rvalid_i(instr_rvalid_i),
				.instr_rdata_i(instr_rdata_i[31:0]),
				.instr_err_i(instr_err),
				.busy_o(prefetch_busy)
			);
			wire unused_icen;
			wire unused_icinv;
			wire unused_scr_key_valid;
			wire [(ibex_pkg_IC_NUM_WAYS * TagSizeECC) - 1:0] unused_tag_ram_input;
			wire [(ibex_pkg_IC_NUM_WAYS * LineSizeECC) - 1:0] unused_data_ram_input;
			assign unused_icen = icache_enable_i;
			assign unused_icinv = icache_inval_i;
			assign unused_tag_ram_input = ic_tag_rdata_i;
			assign unused_data_ram_input = ic_data_rdata_i;
			assign unused_scr_key_valid = ic_scr_key_valid_i;
			assign ic_tag_req_o = 'b0;
			assign ic_tag_write_o = 'b0;
			assign ic_tag_addr_o = 'b0;
			assign ic_tag_wdata_o = 'b0;
			assign ic_data_req_o = 'b0;
			assign ic_data_write_o = 'b0;
			assign ic_data_addr_o = 'b0;
			assign ic_data_wdata_o = 'b0;
			assign ic_scr_key_req_o = 'b0;
			assign icache_ecc_error_o = 'b0;
		end
	endgenerate
	assign unused_fetch_addr_n0 = fetch_addr_n[0];
	assign branch_req = pc_set_i | predict_branch_taken;
	assign pc_if_o = if_instr_addr;
	assign if_busy_o = prefetch_busy;
	assign if_instr_pmp_err = pmp_err_if_i | ((if_instr_addr[1] & ~instr_is_compressed) & pmp_err_if_plus2_i);
	assign if_instr_err = if_instr_bus_err | if_instr_pmp_err;
	assign if_instr_err_plus2 = (((if_instr_addr[1] & ~instr_is_compressed) & pmp_err_if_plus2_i) | fetch_err_plus2) & ~pmp_err_if_i;
	ibex_compressed_decoder compressed_decoder_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.valid_i(fetch_valid & ~fetch_err),
		.instr_i(if_instr_rdata),
		.instr_o(instr_decompressed),
		.is_compressed_o(instr_is_compressed),
		.illegal_instr_o(illegal_c_insn)
	);
	generate
		if (DummyInstructions) begin : gen_dummy_instr
			wire insert_dummy_instr;
			wire [31:0] dummy_instr_data;
			ibex_dummy_instr #(
				.RndCnstLfsrSeed(RndCnstLfsrSeed),
				.RndCnstLfsrPerm(RndCnstLfsrPerm)
			) dummy_instr_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.dummy_instr_en_i(dummy_instr_en_i),
				.dummy_instr_mask_i(dummy_instr_mask_i),
				.dummy_instr_seed_en_i(dummy_instr_seed_en_i),
				.dummy_instr_seed_i(dummy_instr_seed_i),
				.fetch_valid_i(fetch_valid),
				.id_in_ready_i(id_in_ready_i),
				.insert_dummy_instr_o(insert_dummy_instr),
				.dummy_instr_data_o(dummy_instr_data)
			);
			assign instr_out = (insert_dummy_instr ? dummy_instr_data : instr_decompressed);
			assign instr_is_compressed_out = (insert_dummy_instr ? 1'b0 : instr_is_compressed);
			assign illegal_c_instr_out = (insert_dummy_instr ? 1'b0 : illegal_c_insn);
			assign instr_err_out = (insert_dummy_instr ? 1'b0 : if_instr_err);
			assign stall_dummy_instr = insert_dummy_instr;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					dummy_instr_id_o <= 1'b0;
				else if (if_id_pipe_reg_we)
					dummy_instr_id_o <= insert_dummy_instr;
		end
		else begin : gen_no_dummy_instr
			wire unused_dummy_en;
			wire [2:0] unused_dummy_mask;
			wire unused_dummy_seed_en;
			wire [31:0] unused_dummy_seed;
			assign unused_dummy_en = dummy_instr_en_i;
			assign unused_dummy_mask = dummy_instr_mask_i;
			assign unused_dummy_seed_en = dummy_instr_seed_en_i;
			assign unused_dummy_seed = dummy_instr_seed_i;
			assign instr_out = instr_decompressed;
			assign instr_is_compressed_out = instr_is_compressed;
			assign illegal_c_instr_out = illegal_c_insn;
			assign instr_err_out = if_instr_err;
			assign stall_dummy_instr = 1'b0;
			wire [1:1] sv2v_tmp_A80D7;
			assign sv2v_tmp_A80D7 = 1'b0;
			always @(*) dummy_instr_id_o = sv2v_tmp_A80D7;
		end
	endgenerate
	assign instr_valid_id_d = ((if_instr_valid & id_in_ready_i) & ~pc_set_i) | (instr_valid_id_q & ~instr_valid_clear_i);
	assign instr_new_id_d = if_instr_valid & id_in_ready_i;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			instr_valid_id_q <= 1'b0;
			instr_new_id_q <= 1'b0;
		end
		else begin
			instr_valid_id_q <= instr_valid_id_d;
			instr_new_id_q <= instr_new_id_d;
		end
	assign instr_valid_id_o = instr_valid_id_q;
	assign instr_new_id_o = instr_new_id_q;
	assign if_id_pipe_reg_we = instr_new_id_d;
	generate
		if (ResetAll) begin : g_instr_rdata_ra
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni) begin
					instr_rdata_id_o <= 1'sb0;
					instr_rdata_alu_id_o <= 1'sb0;
					instr_fetch_err_o <= 1'sb0;
					instr_fetch_err_plus2_o <= 1'sb0;
					instr_rdata_c_id_o <= 1'sb0;
					instr_is_compressed_id_o <= 1'sb0;
					illegal_c_insn_id_o <= 1'sb0;
					pc_id_o <= 1'sb0;
				end
				else if (if_id_pipe_reg_we) begin
					instr_rdata_id_o <= instr_out;
					instr_rdata_alu_id_o <= instr_out;
					instr_fetch_err_o <= instr_err_out;
					instr_fetch_err_plus2_o <= if_instr_err_plus2;
					instr_rdata_c_id_o <= if_instr_rdata[15:0];
					instr_is_compressed_id_o <= instr_is_compressed_out;
					illegal_c_insn_id_o <= illegal_c_instr_out;
					pc_id_o <= pc_if_o;
				end
		end
		else begin : g_instr_rdata_nr
			always @(posedge clk_i)
				if (if_id_pipe_reg_we) begin
					instr_rdata_id_o <= instr_out;
					instr_rdata_alu_id_o <= instr_out;
					instr_fetch_err_o <= instr_err_out;
					instr_fetch_err_plus2_o <= if_instr_err_plus2;
					instr_rdata_c_id_o <= if_instr_rdata[15:0];
					instr_is_compressed_id_o <= instr_is_compressed_out;
					illegal_c_insn_id_o <= illegal_c_instr_out;
					pc_id_o <= pc_if_o;
				end
		end
		if (PCIncrCheck) begin : g_secure_pc
			wire [31:0] prev_instr_addr_incr;
			wire [31:0] prev_instr_addr_incr_buf;
			reg prev_instr_seq_q;
			wire prev_instr_seq_d;
			assign prev_instr_seq_d = (((prev_instr_seq_q | instr_new_id_d) & ~branch_req) & ~if_instr_err) & ~stall_dummy_instr;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					prev_instr_seq_q <= 1'b0;
				else
					prev_instr_seq_q <= prev_instr_seq_d;
			assign prev_instr_addr_incr = pc_id_o + (instr_is_compressed_id_o ? 32'd2 : 32'd4);
			prim_buf #(.Width(32)) u_prev_instr_addr_incr_buf(
				.in_i(prev_instr_addr_incr),
				.out_o(prev_instr_addr_incr_buf)
			);
			assign pc_mismatch_alert_o = prev_instr_seq_q & (pc_if_o != prev_instr_addr_incr_buf);
		end
		else begin : g_no_secure_pc
			assign pc_mismatch_alert_o = 1'b0;
		end
		if (BranchPredictor) begin : g_branch_predictor
			reg [31:0] instr_skid_data_q;
			reg [31:0] instr_skid_addr_q;
			reg instr_skid_bp_taken_q;
			reg instr_skid_valid_q;
			wire instr_skid_valid_d;
			wire instr_skid_en;
			reg instr_bp_taken_q;
			wire instr_bp_taken_d;
			wire predict_branch_taken_raw;
			if (ResetAll) begin : g_bp_taken_ra
				always @(posedge clk_i or negedge rst_ni)
					if (!rst_ni)
						instr_bp_taken_q <= 1'sb0;
					else if (if_id_pipe_reg_we)
						instr_bp_taken_q <= instr_bp_taken_d;
			end
			else begin : g_bp_taken_nr
				always @(posedge clk_i)
					if (if_id_pipe_reg_we)
						instr_bp_taken_q <= instr_bp_taken_d;
			end
			assign instr_skid_en = ((predict_branch_taken & ~pc_set_i) & ~id_in_ready_i) & ~instr_skid_valid_q;
			assign instr_skid_valid_d = ((instr_skid_valid_q & ~id_in_ready_i) & ~stall_dummy_instr) | instr_skid_en;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					instr_skid_valid_q <= 1'b0;
				else
					instr_skid_valid_q <= instr_skid_valid_d;
			if (ResetAll) begin : g_instr_skid_ra
				always @(posedge clk_i or negedge rst_ni)
					if (!rst_ni) begin
						instr_skid_bp_taken_q <= 1'sb0;
						instr_skid_data_q <= 1'sb0;
						instr_skid_addr_q <= 1'sb0;
					end
					else if (instr_skid_en) begin
						instr_skid_bp_taken_q <= predict_branch_taken;
						instr_skid_data_q <= fetch_rdata;
						instr_skid_addr_q <= fetch_addr;
					end
			end
			else begin : g_instr_skid_nr
				always @(posedge clk_i)
					if (instr_skid_en) begin
						instr_skid_bp_taken_q <= predict_branch_taken;
						instr_skid_data_q <= fetch_rdata;
						instr_skid_addr_q <= fetch_addr;
					end
			end
			ibex_branch_predict branch_predict_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.fetch_rdata_i(fetch_rdata),
				.fetch_pc_i(fetch_addr),
				.fetch_valid_i(fetch_valid),
				.predict_branch_taken_o(predict_branch_taken_raw),
				.predict_branch_pc_o(predict_branch_pc)
			);
			assign predict_branch_taken = (predict_branch_taken_raw & ~instr_skid_valid_q) & ~fetch_err;
			assign if_instr_valid = fetch_valid | (instr_skid_valid_q & ~nt_branch_mispredict_i);
			assign if_instr_rdata = (instr_skid_valid_q ? instr_skid_data_q : fetch_rdata);
			assign if_instr_addr = (instr_skid_valid_q ? instr_skid_addr_q : fetch_addr);
			assign if_instr_bus_err = ~instr_skid_valid_q & fetch_err;
			assign instr_bp_taken_d = (instr_skid_valid_q ? instr_skid_bp_taken_q : predict_branch_taken);
			assign fetch_ready = (id_in_ready_i & ~stall_dummy_instr) & ~instr_skid_valid_q;
			assign instr_bp_taken_o = instr_bp_taken_q;
		end
		else begin : g_no_branch_predictor
			assign instr_bp_taken_o = 1'b0;
			assign predict_branch_taken = 1'b0;
			assign predict_branch_pc = 32'b00000000000000000000000000000000;
			assign if_instr_valid = fetch_valid;
			assign if_instr_rdata = fetch_rdata;
			assign if_instr_addr = fetch_addr;
			assign if_instr_bus_err = fetch_err;
			assign fetch_ready = id_in_ready_i & ~stall_dummy_instr;
		end
	endgenerate
endmodule
module ibex_load_store_unit (
	clk_i,
	rst_ni,
	data_req_o,
	data_gnt_i,
	data_rvalid_i,
	data_bus_err_i,
	data_pmp_err_i,
	data_addr_o,
	data_we_o,
	data_be_o,
	data_wdata_o,
	data_rdata_i,
	lsu_we_i,
	lsu_type_i,
	lsu_wdata_i,
	lsu_sign_ext_i,
	lsu_rdata_o,
	lsu_rdata_valid_o,
	lsu_req_i,
	adder_result_ex_i,
	addr_incr_req_o,
	addr_last_o,
	lsu_req_done_o,
	lsu_resp_valid_o,
	load_err_o,
	load_resp_intg_err_o,
	store_err_o,
	store_resp_intg_err_o,
	busy_o,
	perf_load_o,
	perf_store_o
);
	parameter [0:0] MemECC = 1'b0;
	parameter [31:0] MemDataWidth = (MemECC ? 39 : 32);
	input wire clk_i;
	input wire rst_ni;
	output reg data_req_o;
	input wire data_gnt_i;
	input wire data_rvalid_i;
	input wire data_bus_err_i;
	input wire data_pmp_err_i;
	output wire [31:0] data_addr_o;
	output wire data_we_o;
	output wire [3:0] data_be_o;
	output wire [MemDataWidth - 1:0] data_wdata_o;
	input wire [MemDataWidth - 1:0] data_rdata_i;
	input wire lsu_we_i;
	input wire [1:0] lsu_type_i;
	input wire [31:0] lsu_wdata_i;
	input wire lsu_sign_ext_i;
	output wire [31:0] lsu_rdata_o;
	output wire lsu_rdata_valid_o;
	input wire lsu_req_i;
	input wire [31:0] adder_result_ex_i;
	output reg addr_incr_req_o;
	output wire [31:0] addr_last_o;
	output wire lsu_req_done_o;
	output wire lsu_resp_valid_o;
	output wire load_err_o;
	output wire load_resp_intg_err_o;
	output wire store_err_o;
	output wire store_resp_intg_err_o;
	output wire busy_o;
	output reg perf_load_o;
	output reg perf_store_o;
	wire [31:0] data_addr;
	wire [31:0] data_addr_w_aligned;
	reg [31:0] addr_last_q;
	wire [31:0] addr_last_d;
	reg addr_update;
	reg ctrl_update;
	reg rdata_update;
	reg [31:8] rdata_q;
	reg [1:0] rdata_offset_q;
	reg [1:0] data_type_q;
	reg data_sign_ext_q;
	reg data_we_q;
	wire [1:0] data_offset;
	reg [3:0] data_be;
	reg [31:0] data_wdata;
	reg [31:0] data_rdata_ext;
	reg [31:0] rdata_w_ext;
	reg [31:0] rdata_h_ext;
	reg [31:0] rdata_b_ext;
	wire split_misaligned_access;
	reg handle_misaligned_q;
	reg handle_misaligned_d;
	reg pmp_err_q;
	reg pmp_err_d;
	reg lsu_err_q;
	reg lsu_err_d;
	wire data_intg_err;
	wire data_or_pmp_err;
	reg [2:0] ls_fsm_cs;
	reg [2:0] ls_fsm_ns;
	assign data_addr = adder_result_ex_i;
	assign data_offset = data_addr[1:0];
	always @(*)
		case (lsu_type_i)
			2'b00:
				if (!handle_misaligned_q)
					case (data_offset)
						2'b00: data_be = 4'b1111;
						2'b01: data_be = 4'b1110;
						2'b10: data_be = 4'b1100;
						2'b11: data_be = 4'b1000;
						default: data_be = 4'b1111;
					endcase
				else
					case (data_offset)
						2'b00: data_be = 4'b0000;
						2'b01: data_be = 4'b0001;
						2'b10: data_be = 4'b0011;
						2'b11: data_be = 4'b0111;
						default: data_be = 4'b1111;
					endcase
			2'b01:
				if (!handle_misaligned_q)
					case (data_offset)
						2'b00: data_be = 4'b0011;
						2'b01: data_be = 4'b0110;
						2'b10: data_be = 4'b1100;
						2'b11: data_be = 4'b1000;
						default: data_be = 4'b1111;
					endcase
				else
					data_be = 4'b0001;
			2'b10, 2'b11:
				case (data_offset)
					2'b00: data_be = 4'b0001;
					2'b01: data_be = 4'b0010;
					2'b10: data_be = 4'b0100;
					2'b11: data_be = 4'b1000;
					default: data_be = 4'b1111;
				endcase
			default: data_be = 4'b1111;
		endcase
	always @(*)
		case (data_offset)
			2'b00: data_wdata = lsu_wdata_i[31:0];
			2'b01: data_wdata = {lsu_wdata_i[23:0], lsu_wdata_i[31:24]};
			2'b10: data_wdata = {lsu_wdata_i[15:0], lsu_wdata_i[31:16]};
			2'b11: data_wdata = {lsu_wdata_i[7:0], lsu_wdata_i[31:8]};
			default: data_wdata = lsu_wdata_i[31:0];
		endcase
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			rdata_q <= 1'sb0;
		else if (rdata_update)
			rdata_q <= data_rdata_i[31:8];
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			rdata_offset_q <= 2'h0;
			data_type_q <= 2'h0;
			data_sign_ext_q <= 1'b0;
			data_we_q <= 1'b0;
		end
		else if (ctrl_update) begin
			rdata_offset_q <= data_offset;
			data_type_q <= lsu_type_i;
			data_sign_ext_q <= lsu_sign_ext_i;
			data_we_q <= lsu_we_i;
		end
	assign addr_last_d = (addr_incr_req_o ? data_addr_w_aligned : data_addr);
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			addr_last_q <= 1'sb0;
		else if (addr_update)
			addr_last_q <= addr_last_d;
	always @(*)
		case (rdata_offset_q)
			2'b00: rdata_w_ext = data_rdata_i[31:0];
			2'b01: rdata_w_ext = {data_rdata_i[7:0], rdata_q[31:8]};
			2'b10: rdata_w_ext = {data_rdata_i[15:0], rdata_q[31:16]};
			2'b11: rdata_w_ext = {data_rdata_i[23:0], rdata_q[31:24]};
			default: rdata_w_ext = data_rdata_i[31:0];
		endcase
	always @(*)
		case (rdata_offset_q)
			2'b00:
				if (!data_sign_ext_q)
					rdata_h_ext = {16'h0000, data_rdata_i[15:0]};
				else
					rdata_h_ext = {{16 {data_rdata_i[15]}}, data_rdata_i[15:0]};
			2'b01:
				if (!data_sign_ext_q)
					rdata_h_ext = {16'h0000, data_rdata_i[23:8]};
				else
					rdata_h_ext = {{16 {data_rdata_i[23]}}, data_rdata_i[23:8]};
			2'b10:
				if (!data_sign_ext_q)
					rdata_h_ext = {16'h0000, data_rdata_i[31:16]};
				else
					rdata_h_ext = {{16 {data_rdata_i[31]}}, data_rdata_i[31:16]};
			2'b11:
				if (!data_sign_ext_q)
					rdata_h_ext = {16'h0000, data_rdata_i[7:0], rdata_q[31:24]};
				else
					rdata_h_ext = {{16 {data_rdata_i[7]}}, data_rdata_i[7:0], rdata_q[31:24]};
			default: rdata_h_ext = {16'h0000, data_rdata_i[15:0]};
		endcase
	always @(*)
		case (rdata_offset_q)
			2'b00:
				if (!data_sign_ext_q)
					rdata_b_ext = {24'h000000, data_rdata_i[7:0]};
				else
					rdata_b_ext = {{24 {data_rdata_i[7]}}, data_rdata_i[7:0]};
			2'b01:
				if (!data_sign_ext_q)
					rdata_b_ext = {24'h000000, data_rdata_i[15:8]};
				else
					rdata_b_ext = {{24 {data_rdata_i[15]}}, data_rdata_i[15:8]};
			2'b10:
				if (!data_sign_ext_q)
					rdata_b_ext = {24'h000000, data_rdata_i[23:16]};
				else
					rdata_b_ext = {{24 {data_rdata_i[23]}}, data_rdata_i[23:16]};
			2'b11:
				if (!data_sign_ext_q)
					rdata_b_ext = {24'h000000, data_rdata_i[31:24]};
				else
					rdata_b_ext = {{24 {data_rdata_i[31]}}, data_rdata_i[31:24]};
			default: rdata_b_ext = {24'h000000, data_rdata_i[7:0]};
		endcase
	always @(*)
		case (data_type_q)
			2'b00: data_rdata_ext = rdata_w_ext;
			2'b01: data_rdata_ext = rdata_h_ext;
			2'b10, 2'b11: data_rdata_ext = rdata_b_ext;
			default: data_rdata_ext = rdata_w_ext;
		endcase
	generate
		if (MemECC) begin : g_mem_rdata_ecc
			wire [1:0] ecc_err;
			wire [MemDataWidth - 1:0] data_rdata_buf;
			prim_buf #(.Width(MemDataWidth)) u_prim_buf_instr_rdata(
				.in_i(data_rdata_i),
				.out_o(data_rdata_buf)
			);
			prim_secded_inv_39_32_dec u_data_intg_dec(
				.data_i(data_rdata_buf),
				.err_o(ecc_err)
			);
			assign data_intg_err = |ecc_err;
		end
		else begin : g_no_mem_data_ecc
			assign data_intg_err = 1'b0;
		end
	endgenerate
	assign split_misaligned_access = ((lsu_type_i == 2'b00) && (data_offset != 2'b00)) || ((lsu_type_i == 2'b01) && (data_offset == 2'b11));
	always @(*) begin
		ls_fsm_ns = ls_fsm_cs;
		data_req_o = 1'b0;
		addr_incr_req_o = 1'b0;
		handle_misaligned_d = handle_misaligned_q;
		pmp_err_d = pmp_err_q;
		lsu_err_d = lsu_err_q;
		addr_update = 1'b0;
		ctrl_update = 1'b0;
		rdata_update = 1'b0;
		perf_load_o = 1'b0;
		perf_store_o = 1'b0;
		case (ls_fsm_cs)
			3'd0: begin
				pmp_err_d = 1'b0;
				if (lsu_req_i) begin
					data_req_o = 1'b1;
					pmp_err_d = data_pmp_err_i;
					lsu_err_d = 1'b0;
					perf_load_o = ~lsu_we_i;
					perf_store_o = lsu_we_i;
					if (data_gnt_i) begin
						ctrl_update = 1'b1;
						addr_update = 1'b1;
						handle_misaligned_d = split_misaligned_access;
						ls_fsm_ns = (split_misaligned_access ? 3'd2 : 3'd0);
					end
					else
						ls_fsm_ns = (split_misaligned_access ? 3'd1 : 3'd3);
				end
			end
			3'd1: begin
				data_req_o = 1'b1;
				if (data_gnt_i || pmp_err_q) begin
					addr_update = 1'b1;
					ctrl_update = 1'b1;
					handle_misaligned_d = 1'b1;
					ls_fsm_ns = 3'd2;
				end
			end
			3'd2: begin
				data_req_o = 1'b1;
				addr_incr_req_o = 1'b1;
				if (data_rvalid_i || pmp_err_q) begin
					pmp_err_d = data_pmp_err_i;
					lsu_err_d = data_bus_err_i | pmp_err_q;
					rdata_update = ~data_we_q;
					ls_fsm_ns = (data_gnt_i ? 3'd0 : 3'd3);
					addr_update = data_gnt_i & ~(data_bus_err_i | pmp_err_q);
					handle_misaligned_d = ~data_gnt_i;
				end
				else if (data_gnt_i) begin
					ls_fsm_ns = 3'd4;
					handle_misaligned_d = 1'b0;
				end
			end
			3'd3: begin
				addr_incr_req_o = handle_misaligned_q;
				data_req_o = 1'b1;
				if (data_gnt_i || pmp_err_q) begin
					ctrl_update = 1'b1;
					addr_update = ~lsu_err_q;
					ls_fsm_ns = 3'd0;
					handle_misaligned_d = 1'b0;
				end
			end
			3'd4: begin
				addr_incr_req_o = 1'b1;
				if (data_rvalid_i) begin
					pmp_err_d = data_pmp_err_i;
					lsu_err_d = data_bus_err_i;
					addr_update = ~data_bus_err_i;
					rdata_update = ~data_we_q;
					ls_fsm_ns = 3'd0;
				end
			end
			default: ls_fsm_ns = 3'd0;
		endcase
	end
	assign lsu_req_done_o = (lsu_req_i | (ls_fsm_cs != 3'd0)) & (ls_fsm_ns == 3'd0);
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			ls_fsm_cs <= 3'd0;
			handle_misaligned_q <= 1'sb0;
			pmp_err_q <= 1'sb0;
			lsu_err_q <= 1'sb0;
		end
		else begin
			ls_fsm_cs <= ls_fsm_ns;
			handle_misaligned_q <= handle_misaligned_d;
			pmp_err_q <= pmp_err_d;
			lsu_err_q <= lsu_err_d;
		end
	assign data_or_pmp_err = (lsu_err_q | data_bus_err_i) | pmp_err_q;
	assign lsu_resp_valid_o = (data_rvalid_i | pmp_err_q) & (ls_fsm_cs == 3'd0);
	assign lsu_rdata_valid_o = ((((ls_fsm_cs == 3'd0) & data_rvalid_i) & ~data_or_pmp_err) & ~data_we_q) & ~data_intg_err;
	assign lsu_rdata_o = data_rdata_ext;
	assign data_addr_w_aligned = {data_addr[31:2], 2'b00};
	assign data_addr_o = data_addr_w_aligned;
	assign data_we_o = lsu_we_i;
	assign data_be_o = data_be;
	generate
		if (MemECC) begin : g_mem_wdata_ecc
			prim_secded_inv_39_32_enc u_data_gen(
				.data_i(data_wdata),
				.data_o(data_wdata_o)
			);
		end
		else begin : g_no_mem_wdata_ecc
			assign data_wdata_o = data_wdata;
		end
	endgenerate
	assign addr_last_o = addr_last_q;
	assign load_err_o = (data_or_pmp_err & ~data_we_q) & lsu_resp_valid_o;
	assign store_err_o = (data_or_pmp_err & data_we_q) & lsu_resp_valid_o;
	assign load_resp_intg_err_o = (data_intg_err & data_rvalid_i) & ~data_we_q;
	assign store_resp_intg_err_o = (data_intg_err & data_rvalid_i) & data_we_q;
	assign busy_o = ls_fsm_cs != 3'd0;
endmodule
module ibex_lockstep (
	clk_i,
	rst_ni,
	hart_id_i,
	boot_addr_i,
	instr_req_i,
	instr_gnt_i,
	instr_rvalid_i,
	instr_addr_i,
	instr_rdata_i,
	instr_err_i,
	data_req_i,
	data_gnt_i,
	data_rvalid_i,
	data_we_i,
	data_be_i,
	data_addr_i,
	data_wdata_i,
	data_rdata_i,
	data_err_i,
	dummy_instr_id_i,
	dummy_instr_wb_i,
	rf_raddr_a_i,
	rf_raddr_b_i,
	rf_waddr_wb_i,
	rf_we_wb_i,
	rf_wdata_wb_ecc_i,
	rf_rdata_a_ecc_i,
	rf_rdata_b_ecc_i,
	ic_tag_req_i,
	ic_tag_write_i,
	ic_tag_addr_i,
	ic_tag_wdata_i,
	ic_tag_rdata_i,
	ic_data_req_i,
	ic_data_write_i,
	ic_data_addr_i,
	ic_data_wdata_i,
	ic_data_rdata_i,
	ic_scr_key_valid_i,
	ic_scr_key_req_i,
	irq_software_i,
	irq_timer_i,
	irq_external_i,
	irq_fast_i,
	irq_nm_i,
	irq_pending_i,
	debug_req_i,
	crash_dump_i,
	double_fault_seen_i,
	fetch_enable_i,
	alert_minor_o,
	alert_major_internal_o,
	alert_major_bus_o,
	core_busy_i,
	test_en_i,
	scan_rst_ni
);
	parameter [31:0] LockstepOffset = 2;
	parameter [0:0] PMPEnable = 1'b0;
	parameter [31:0] PMPGranularity = 0;
	parameter [31:0] PMPNumRegions = 4;
	parameter [31:0] MHPMCounterNum = 0;
	parameter [31:0] MHPMCounterWidth = 40;
	parameter [0:0] RV32E = 1'b0;
	parameter integer RV32M = 32'sd2;
	parameter integer RV32B = 32'sd0;
	parameter [0:0] BranchTargetALU = 1'b0;
	parameter [0:0] WritebackStage = 1'b0;
	parameter [0:0] ICache = 1'b0;
	parameter [0:0] ICacheECC = 1'b0;
	localparam [31:0] ibex_pkg_BUS_SIZE = 32;
	parameter [31:0] BusSizeECC = ibex_pkg_BUS_SIZE;
	localparam [31:0] ibex_pkg_ADDR_W = 32;
	localparam [31:0] ibex_pkg_IC_LINE_SIZE = 64;
	localparam [31:0] ibex_pkg_IC_LINE_BYTES = 8;
	localparam [31:0] ibex_pkg_IC_NUM_WAYS = 2;
	localparam [31:0] ibex_pkg_IC_SIZE_BYTES = 4096;
	localparam [31:0] ibex_pkg_IC_NUM_LINES = (ibex_pkg_IC_SIZE_BYTES / ibex_pkg_IC_NUM_WAYS) / ibex_pkg_IC_LINE_BYTES;
	localparam [31:0] ibex_pkg_IC_INDEX_W = $clog2(ibex_pkg_IC_NUM_LINES);
	localparam [31:0] ibex_pkg_IC_LINE_W = 3;
	localparam [31:0] ibex_pkg_IC_TAG_SIZE = ((ibex_pkg_ADDR_W - ibex_pkg_IC_INDEX_W) - ibex_pkg_IC_LINE_W) + 1;
	parameter [31:0] TagSizeECC = ibex_pkg_IC_TAG_SIZE;
	parameter [31:0] LineSizeECC = ibex_pkg_IC_LINE_SIZE;
	parameter [0:0] BranchPredictor = 1'b0;
	parameter [0:0] DbgTriggerEn = 1'b0;
	parameter [31:0] DbgHwBreakNum = 1;
	parameter [0:0] ResetAll = 1'b0;
	localparam signed [31:0] ibex_pkg_LfsrWidth = 32;
	localparam [31:0] ibex_pkg_RndCnstLfsrSeedDefault = 32'hac533bf4;
	parameter [31:0] RndCnstLfsrSeed = ibex_pkg_RndCnstLfsrSeedDefault;
	localparam [159:0] ibex_pkg_RndCnstLfsrPermDefault = 160'h1e35ecba467fd1b12e958152c04fa43878a8daed;
	parameter [159:0] RndCnstLfsrPerm = ibex_pkg_RndCnstLfsrPermDefault;
	parameter [0:0] SecureIbex = 1'b0;
	parameter [0:0] DummyInstructions = 1'b0;
	parameter [0:0] RegFileECC = 1'b0;
	parameter [31:0] RegFileDataWidth = 32;
	parameter [0:0] MemECC = 1'b0;
	parameter [31:0] MemDataWidth = (MemECC ? 39 : 32);
	parameter [31:0] DmHaltAddr = 32'h1a110800;
	parameter [31:0] DmExceptionAddr = 32'h1a110808;
	input wire clk_i;
	input wire rst_ni;
	input wire [31:0] hart_id_i;
	input wire [31:0] boot_addr_i;
	input wire instr_req_i;
	input wire instr_gnt_i;
	input wire instr_rvalid_i;
	input wire [31:0] instr_addr_i;
	input wire [MemDataWidth - 1:0] instr_rdata_i;
	input wire instr_err_i;
	input wire data_req_i;
	input wire data_gnt_i;
	input wire data_rvalid_i;
	input wire data_we_i;
	input wire [3:0] data_be_i;
	input wire [31:0] data_addr_i;
	input wire [MemDataWidth - 1:0] data_wdata_i;
	input wire [MemDataWidth - 1:0] data_rdata_i;
	input wire data_err_i;
	input wire dummy_instr_id_i;
	input wire dummy_instr_wb_i;
	input wire [4:0] rf_raddr_a_i;
	input wire [4:0] rf_raddr_b_i;
	input wire [4:0] rf_waddr_wb_i;
	input wire rf_we_wb_i;
	input wire [RegFileDataWidth - 1:0] rf_wdata_wb_ecc_i;
	input wire [RegFileDataWidth - 1:0] rf_rdata_a_ecc_i;
	input wire [RegFileDataWidth - 1:0] rf_rdata_b_ecc_i;
	input wire [1:0] ic_tag_req_i;
	input wire ic_tag_write_i;
	input wire [ibex_pkg_IC_INDEX_W - 1:0] ic_tag_addr_i;
	input wire [TagSizeECC - 1:0] ic_tag_wdata_i;
	input wire [(ibex_pkg_IC_NUM_WAYS * TagSizeECC) - 1:0] ic_tag_rdata_i;
	input wire [1:0] ic_data_req_i;
	input wire ic_data_write_i;
	input wire [ibex_pkg_IC_INDEX_W - 1:0] ic_data_addr_i;
	input wire [LineSizeECC - 1:0] ic_data_wdata_i;
	input wire [(ibex_pkg_IC_NUM_WAYS * LineSizeECC) - 1:0] ic_data_rdata_i;
	input wire ic_scr_key_valid_i;
	input wire ic_scr_key_req_i;
	input wire irq_software_i;
	input wire irq_timer_i;
	input wire irq_external_i;
	input wire [14:0] irq_fast_i;
	input wire irq_nm_i;
	input wire irq_pending_i;
	input wire debug_req_i;
	input wire [159:0] crash_dump_i;
	input wire double_fault_seen_i;
	input wire [3:0] fetch_enable_i;
	output wire alert_minor_o;
	output wire alert_major_internal_o;
	output wire alert_major_bus_o;
	input wire [3:0] core_busy_i;
	input wire test_en_i;
	input wire scan_rst_ni;
	localparam [31:0] LockstepOffsetW = $clog2(LockstepOffset);
	localparam [31:0] OutputsOffset = LockstepOffset + 1;
	wire [LockstepOffsetW - 1:0] rst_shadow_cnt_d;
	reg [LockstepOffsetW - 1:0] rst_shadow_cnt_q;
	wire [LockstepOffsetW - 1:0] rst_shadow_cnt_incr;
	wire rst_shadow_set_d;
	wire rst_shadow_set_q;
	wire rst_shadow_n;
	reg enable_cmp_q;
	assign rst_shadow_cnt_incr = rst_shadow_cnt_q + 1'b1;
	function automatic [LockstepOffsetW - 1:0] sv2v_cast_3B624;
		input reg [LockstepOffsetW - 1:0] inp;
		sv2v_cast_3B624 = inp;
	endfunction
	assign rst_shadow_set_d = rst_shadow_cnt_q == sv2v_cast_3B624(LockstepOffset - 1);
	assign rst_shadow_cnt_d = (rst_shadow_set_d ? rst_shadow_cnt_q : rst_shadow_cnt_incr);
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			rst_shadow_cnt_q <= 1'sb0;
			enable_cmp_q <= 1'sb0;
		end
		else begin
			rst_shadow_cnt_q <= rst_shadow_cnt_d;
			enable_cmp_q <= rst_shadow_set_q;
		end
	prim_flop #(
		.Width(1),
		.ResetValue(1'b0)
	) u_prim_rst_shadow_set_flop(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(rst_shadow_set_d),
		.q_o(rst_shadow_set_q)
	);
	prim_clock_mux2 #(.NoFpgaBufG(1'b1)) u_prim_rst_shadow_n_mux2(
		.clk0_i(rst_shadow_set_q),
		.clk1_i(scan_rst_ni),
		.sel_i(test_en_i),
		.clk_o(rst_shadow_n)
	);
	reg [((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? (LockstepOffset * (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 25)) - 1 : (LockstepOffset * (1 - (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24))) + (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 23)):((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 0 : ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24)] shadow_inputs_q;
	wire [((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24:0] shadow_inputs_in;
	reg [(LockstepOffset * TagSizeECC) - 1:0] shadow_tag_rdata_q [0:1];
	reg [(LockstepOffset * LineSizeECC) - 1:0] shadow_data_rdata_q [0:1];
	assign shadow_inputs_in[2 + (MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))))] = instr_gnt_i;
	assign shadow_inputs_in[1 + (MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))))] = instr_rvalid_i;
	assign shadow_inputs_in[MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))))-:((MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))))) >= (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 25))))) ? ((MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))))) - (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 25)))))) + 1 : ((3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 25))))) - (MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))))) + 1)] = instr_rdata_i;
	assign shadow_inputs_in[3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))] = instr_err_i;
	assign shadow_inputs_in[2 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))] = data_gnt_i;
	assign shadow_inputs_in[1 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))] = data_rvalid_i;
	assign shadow_inputs_in[MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))-:((MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))) >= (1 + (RegFileDataWidth + (RegFileDataWidth + 25))) ? ((MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))) - (1 + (RegFileDataWidth + (RegFileDataWidth + 25)))) + 1 : ((1 + (RegFileDataWidth + (RegFileDataWidth + 25))) - (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))) + 1)] = data_rdata_i;
	assign shadow_inputs_in[1 + (RegFileDataWidth + (RegFileDataWidth + 24))] = data_err_i;
	assign shadow_inputs_in[RegFileDataWidth + (RegFileDataWidth + 24)-:((RegFileDataWidth + (RegFileDataWidth + 24)) >= (RegFileDataWidth + 25) ? ((RegFileDataWidth + (RegFileDataWidth + 24)) - (RegFileDataWidth + 25)) + 1 : ((RegFileDataWidth + 25) - (RegFileDataWidth + (RegFileDataWidth + 24))) + 1)] = rf_rdata_a_ecc_i;
	assign shadow_inputs_in[RegFileDataWidth + 24-:((RegFileDataWidth + 24) >= 25 ? RegFileDataWidth + 0 : 26 - (RegFileDataWidth + 24))] = rf_rdata_b_ecc_i;
	assign shadow_inputs_in[24] = irq_software_i;
	assign shadow_inputs_in[23] = irq_timer_i;
	assign shadow_inputs_in[22] = irq_external_i;
	assign shadow_inputs_in[21-:15] = irq_fast_i;
	assign shadow_inputs_in[6] = irq_nm_i;
	assign shadow_inputs_in[5] = debug_req_i;
	assign shadow_inputs_in[4-:4] = fetch_enable_i;
	assign shadow_inputs_in[0] = ic_scr_key_valid_i;
	function automatic [((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 25 : 1 - (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24)) - 1:0] sv2v_cast_6AC9E;
		input reg [((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 25 : 1 - (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24)) - 1:0] inp;
		sv2v_cast_6AC9E = inp;
	endfunction
	function automatic [TagSizeECC - 1:0] sv2v_cast_CA15E;
		input reg [TagSizeECC - 1:0] inp;
		sv2v_cast_CA15E = inp;
	endfunction
	function automatic [LineSizeECC - 1:0] sv2v_cast_B1C65;
		input reg [LineSizeECC - 1:0] inp;
		sv2v_cast_B1C65 = inp;
	endfunction
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < LockstepOffset; i = i + 1)
				begin
					shadow_inputs_q[((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 0 : ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) + (i * ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 25 : 1 - (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24)))+:((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 25 : 1 - (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24))] <= sv2v_cast_6AC9E(1'sb0);
					shadow_tag_rdata_q[i] <= {LockstepOffset {sv2v_cast_CA15E(0)}};
					shadow_data_rdata_q[i] <= {LockstepOffset {sv2v_cast_B1C65(0)}};
				end
		end
		else begin
			begin : sv2v_autoblock_2
				reg [31:0] i;
				for (i = 0; i < (LockstepOffset - 1); i = i + 1)
					begin
						shadow_inputs_q[((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 0 : ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) + (i * ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 25 : 1 - (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24)))+:((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 25 : 1 - (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24))] <= shadow_inputs_q[((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 0 : ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) + ((i + 1) * ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 25 : 1 - (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24)))+:((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 25 : 1 - (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24))];
						shadow_tag_rdata_q[i] <= shadow_tag_rdata_q[i + 1];
						shadow_data_rdata_q[i] <= shadow_data_rdata_q[i + 1];
					end
			end
			shadow_inputs_q[((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 0 : ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) + ((LockstepOffset - 1) * ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 25 : 1 - (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24)))+:((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 25 : 1 - (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24))] <= shadow_inputs_in;
			shadow_tag_rdata_q[LockstepOffset - 1] <= ic_tag_rdata_i;
			shadow_data_rdata_q[LockstepOffset - 1] <= ic_data_rdata_i;
		end
	reg [(((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + 3) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + 3) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) >= 0 ? (OutputsOffset * ((((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 167)) - 1 : (OutputsOffset * (1 - ((((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166))) + ((((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 165)):(((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + 3) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + 3) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) >= 0 ? 0 : (((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166)] core_outputs_q;
	wire [(((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166:0] core_outputs_in;
	wire [(((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166:0] shadow_outputs_d;
	reg [(((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166:0] shadow_outputs_q;
	assign core_outputs_in[71 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))] = instr_req_i;
	assign core_outputs_in[70 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))-:((70 + (MemDataWidth + (18 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))) >= (38 + (MemDataWidth + (18 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))) ? ((70 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))) - (38 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))))))) + 1 : ((38 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))))) - (70 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))))))) + 1)] = instr_addr_i;
	assign core_outputs_in[38 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))] = data_req_i;
	assign core_outputs_in[37 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))] = data_we_i;
	assign core_outputs_in[36 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))-:((36 + (MemDataWidth + (18 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))) >= (32 + (MemDataWidth + (18 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))) ? ((36 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))) - (32 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))))))) + 1 : ((32 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))))) - (36 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))))))) + 1)] = data_be_i;
	assign core_outputs_in[32 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))-:((32 + (MemDataWidth + (18 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))) >= (MemDataWidth + (18 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))) ? ((32 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))) - (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))))) + 1 : ((MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))))) - (32 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))))))) + 1)] = data_addr_i;
	assign core_outputs_in[MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))))-:((MemDataWidth + (18 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))) >= (18 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))) ? ((MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))))) - (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))))) + 1 : ((18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))) - (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))) + 1)] = data_wdata_i;
	assign core_outputs_in[18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))] = dummy_instr_id_i;
	assign core_outputs_in[17 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))] = dummy_instr_wb_i;
	assign core_outputs_in[16 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))-:((16 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))) >= (11 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))) ? ((16 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))) - (11 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))))) + 1 : ((11 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))) - (16 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))))) + 1)] = rf_raddr_a_i;
	assign core_outputs_in[11 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))-:((11 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))) >= (6 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))) ? ((11 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))) - (6 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))))) + 1 : ((6 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))) - (11 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))))) + 1)] = rf_raddr_b_i;
	assign core_outputs_in[6 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))-:((6 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))) >= (1 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))) ? ((6 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))) - (1 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))))) + 1 : ((1 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))) - (6 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))))) + 1)] = rf_waddr_wb_i;
	assign core_outputs_in[1 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))] = rf_we_wb_i;
	assign core_outputs_in[RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))-:((RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))) >= (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))) ? ((RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))) - (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))) + 1 : ((ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))) - (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))) + 1)] = rf_wdata_wb_ecc_i;
	assign core_outputs_in[ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))-:((3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))) >= (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))) ? ((ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))) - (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))) + 1 : ((1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))) - (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))) + 1)] = ic_tag_req_i;
	assign core_outputs_in[1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))] = ic_tag_write_i;
	assign core_outputs_in[ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))-:((ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))) >= (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))) ? ((ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))) - (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))) + 1 : ((TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))) - (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))) + 1)] = ic_tag_addr_i;
	assign core_outputs_in[TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))-:((TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))) >= (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))) ? ((TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))) - (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))) + 1 : ((ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))) - (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))) + 1)] = ic_tag_wdata_i;
	assign core_outputs_in[ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))-:((3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))) >= (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))) ? ((ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))) - (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))) + 1 : ((1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))) - (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))) + 1)] = ic_data_req_i;
	assign core_outputs_in[1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))] = ic_data_write_i;
	assign core_outputs_in[ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)-:((ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)) >= (LineSizeECC + 167) ? ((ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)) - (LineSizeECC + 167)) + 1 : ((LineSizeECC + 167) - (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))) + 1)] = ic_data_addr_i;
	assign core_outputs_in[LineSizeECC + 166-:((LineSizeECC + 166) >= 167 ? LineSizeECC + 0 : 168 - (LineSizeECC + 166))] = ic_data_wdata_i;
	assign core_outputs_in[166] = ic_scr_key_req_i;
	assign core_outputs_in[165] = irq_pending_i;
	assign core_outputs_in[164-:160] = crash_dump_i;
	assign core_outputs_in[4] = double_fault_seen_i;
	assign core_outputs_in[3-:4] = core_busy_i;
	always @(posedge clk_i) begin
		begin : sv2v_autoblock_3
			reg [31:0] i;
			for (i = 0; i < (OutputsOffset - 1); i = i + 1)
				core_outputs_q[(((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + 3) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + 3) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) >= 0 ? 0 : (((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) + (i * (((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + 3) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + 3) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) >= 0 ? (((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 167 : 1 - ((((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166)))+:(((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + 3) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + 3) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) >= 0 ? (((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 167 : 1 - ((((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166))] <= core_outputs_q[(((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + 3) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + 3) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) >= 0 ? 0 : (((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) + ((i + 1) * (((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + 3) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + 3) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) >= 0 ? (((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 167 : 1 - ((((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166)))+:(((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + 3) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + 3) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) >= 0 ? (((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 167 : 1 - ((((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166))];
		end
		core_outputs_q[(((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + 3) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + 3) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) >= 0 ? 0 : (((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) + ((OutputsOffset - 1) * (((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + 3) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + 3) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) >= 0 ? (((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 167 : 1 - ((((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166)))+:(((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + 3) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + 3) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) >= 0 ? (((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 167 : 1 - ((((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166))] <= core_outputs_in;
	end
	wire shadow_alert_minor;
	wire shadow_alert_major_internal;
	wire shadow_alert_major_bus;
	ibex_core #(
		.PMPEnable(PMPEnable),
		.PMPGranularity(PMPGranularity),
		.PMPNumRegions(PMPNumRegions),
		.MHPMCounterNum(MHPMCounterNum),
		.MHPMCounterWidth(MHPMCounterWidth),
		.RV32E(RV32E),
		.RV32M(RV32M),
		.RV32B(RV32B),
		.BranchTargetALU(BranchTargetALU),
		.ICache(ICache),
		.ICacheECC(ICacheECC),
		.BusSizeECC(BusSizeECC),
		.TagSizeECC(TagSizeECC),
		.LineSizeECC(LineSizeECC),
		.BranchPredictor(BranchPredictor),
		.DbgTriggerEn(DbgTriggerEn),
		.DbgHwBreakNum(DbgHwBreakNum),
		.WritebackStage(WritebackStage),
		.ResetAll(ResetAll),
		.RndCnstLfsrSeed(RndCnstLfsrSeed),
		.RndCnstLfsrPerm(RndCnstLfsrPerm),
		.SecureIbex(SecureIbex),
		.DummyInstructions(DummyInstructions),
		.RegFileECC(RegFileECC),
		.RegFileDataWidth(RegFileDataWidth),
		.MemECC(MemECC),
		.MemDataWidth(MemDataWidth),
		.DmHaltAddr(DmHaltAddr),
		.DmExceptionAddr(DmExceptionAddr)
	) u_shadow_core(
		.clk_i(clk_i),
		.rst_ni(rst_shadow_n),
		.hart_id_i(hart_id_i),
		.boot_addr_i(boot_addr_i),
		.instr_req_o(shadow_outputs_d[71 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))]),
		.instr_gnt_i(shadow_inputs_q[0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 2 + (MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))))) : (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) - (2 + (MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))))))]),
		.instr_rvalid_i(shadow_inputs_q[0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 1 + (MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))))) : (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) - (1 + (MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))))))]),
		.instr_addr_o(shadow_outputs_d[70 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))-:((70 + (MemDataWidth + (18 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))) >= (38 + (MemDataWidth + (18 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))) ? ((70 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))) - (38 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))))))) + 1 : ((38 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))))) - (70 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))))))) + 1)]),
		.instr_rdata_i(shadow_inputs_q[((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))) : (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) - (MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))))) : ((0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))) : (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) - (MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))))))) + ((MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))))) >= (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 25))))) ? ((MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))))) - (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 25)))))) + 1 : ((3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 25))))) - (MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))))) + 1)) - 1)-:((MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))))) >= (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 25))))) ? ((MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))))) - (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 25)))))) + 1 : ((3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 25))))) - (MemDataWidth + (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))))) + 1)]),
		.instr_err_i(shadow_inputs_q[0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))) : (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) - (3 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))))]),
		.data_req_o(shadow_outputs_d[38 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))]),
		.data_gnt_i(shadow_inputs_q[0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 2 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))) : (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) - (2 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))))]),
		.data_rvalid_i(shadow_inputs_q[0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 1 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))) : (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) - (1 + (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))))]),
		.data_we_o(shadow_outputs_d[37 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))]),
		.data_be_o(shadow_outputs_d[36 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))-:((36 + (MemDataWidth + (18 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))) >= (32 + (MemDataWidth + (18 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))) ? ((36 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))) - (32 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))))))) + 1 : ((32 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))))) - (36 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))))))) + 1)]),
		.data_addr_o(shadow_outputs_d[32 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))-:((32 + (MemDataWidth + (18 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))) >= (MemDataWidth + (18 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))) ? ((32 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))) - (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))))) + 1 : ((MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))))) - (32 + (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))))))) + 1)]),
		.data_wdata_o(shadow_outputs_d[MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))))-:((MemDataWidth + (18 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))) >= (18 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))) ? ((MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))))) - (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))))) + 1 : ((18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))) - (MemDataWidth + (18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))))) + 1)]),
		.data_rdata_i(shadow_inputs_q[((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))) : (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) - (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))) : ((0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))) : (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) - (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))))) + ((MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))) >= (1 + (RegFileDataWidth + (RegFileDataWidth + 25))) ? ((MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))) - (1 + (RegFileDataWidth + (RegFileDataWidth + 25)))) + 1 : ((1 + (RegFileDataWidth + (RegFileDataWidth + 25))) - (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))) + 1)) - 1)-:((MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))) >= (1 + (RegFileDataWidth + (RegFileDataWidth + 25))) ? ((MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24)))) - (1 + (RegFileDataWidth + (RegFileDataWidth + 25)))) + 1 : ((1 + (RegFileDataWidth + (RegFileDataWidth + 25))) - (MemDataWidth + (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))) + 1)]),
		.data_err_i(shadow_inputs_q[0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 1 + (RegFileDataWidth + (RegFileDataWidth + 24)) : (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) - (1 + (RegFileDataWidth + (RegFileDataWidth + 24))))]),
		.dummy_instr_id_o(shadow_outputs_d[18 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))]),
		.dummy_instr_wb_o(shadow_outputs_d[17 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))]),
		.rf_raddr_a_o(shadow_outputs_d[16 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))-:((16 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))) >= (11 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))) ? ((16 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))) - (11 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))))) + 1 : ((11 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))) - (16 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))))) + 1)]),
		.rf_raddr_b_o(shadow_outputs_d[11 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))-:((11 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))) >= (6 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))) ? ((11 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))) - (6 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))))) + 1 : ((6 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))) - (11 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))))) + 1)]),
		.rf_waddr_wb_o(shadow_outputs_d[6 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))-:((6 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))) >= (1 + (RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))) ? ((6 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))) - (1 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))))) + 1 : ((1 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))))) - (6 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))))) + 1)]),
		.rf_we_wb_o(shadow_outputs_d[1 + (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))]),
		.rf_wdata_wb_ecc_o(shadow_outputs_d[RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))-:((RegFileDataWidth + (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))) >= (3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))) ? ((RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))) - (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))))) + 1 : ((ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))) - (RegFileDataWidth + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))))) + 1)]),
		.rf_rdata_a_ecc_i(shadow_inputs_q[((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? RegFileDataWidth + (RegFileDataWidth + 24) : (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) - (RegFileDataWidth + (RegFileDataWidth + 24))) : ((0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? RegFileDataWidth + (RegFileDataWidth + 24) : (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) - (RegFileDataWidth + (RegFileDataWidth + 24)))) + ((RegFileDataWidth + (RegFileDataWidth + 24)) >= (RegFileDataWidth + 25) ? ((RegFileDataWidth + (RegFileDataWidth + 24)) - (RegFileDataWidth + 25)) + 1 : ((RegFileDataWidth + 25) - (RegFileDataWidth + (RegFileDataWidth + 24))) + 1)) - 1)-:((RegFileDataWidth + (RegFileDataWidth + 24)) >= (RegFileDataWidth + 25) ? ((RegFileDataWidth + (RegFileDataWidth + 24)) - (RegFileDataWidth + 25)) + 1 : ((RegFileDataWidth + 25) - (RegFileDataWidth + (RegFileDataWidth + 24))) + 1)]),
		.rf_rdata_b_ecc_i(shadow_inputs_q[((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? RegFileDataWidth + 24 : (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) - (RegFileDataWidth + 24)) : ((0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? RegFileDataWidth + 24 : (((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) - (RegFileDataWidth + 24))) + ((RegFileDataWidth + 24) >= 25 ? RegFileDataWidth + 0 : 26 - (RegFileDataWidth + 24))) - 1)-:((RegFileDataWidth + 24) >= 25 ? RegFileDataWidth + 0 : 26 - (RegFileDataWidth + 24))]),
		.ic_tag_req_o(shadow_outputs_d[ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))-:((3 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))) >= (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))) ? ((ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))))) - (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))))) + 1 : ((1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))))) - (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))))) + 1)]),
		.ic_tag_write_o(shadow_outputs_d[1 + (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))]),
		.ic_tag_addr_o(shadow_outputs_d[ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))-:((ibex_pkg_IC_INDEX_W + (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))) >= (TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))) ? ((ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))) - (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))))) + 1 : ((TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))) - (ibex_pkg_IC_INDEX_W + (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))))) + 1)]),
		.ic_tag_wdata_o(shadow_outputs_d[TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))-:((TagSizeECC + (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))) >= (3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))) ? ((TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))) - (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))))) + 1 : ((ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))) - (TagSizeECC + (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))))) + 1)]),
		.ic_tag_rdata_i(shadow_tag_rdata_q[0]),
		.ic_data_req_o(shadow_outputs_d[ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))-:((3 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))) >= (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))) ? ((ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)))) - (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167)))) + 1 : ((1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 167))) - (ibex_pkg_IC_NUM_WAYS + (1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))))) + 1)]),
		.ic_data_write_o(shadow_outputs_d[1 + (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))]),
		.ic_data_addr_o(shadow_outputs_d[ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)-:((ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)) >= (LineSizeECC + 167) ? ((ibex_pkg_IC_INDEX_W + (LineSizeECC + 166)) - (LineSizeECC + 167)) + 1 : ((LineSizeECC + 167) - (ibex_pkg_IC_INDEX_W + (LineSizeECC + 166))) + 1)]),
		.ic_data_wdata_o(shadow_outputs_d[LineSizeECC + 166-:((LineSizeECC + 166) >= 167 ? LineSizeECC + 0 : 168 - (LineSizeECC + 166))]),
		.ic_data_rdata_i(shadow_data_rdata_q[0]),
		.ic_scr_key_valid_i(shadow_inputs_q[0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 0 : ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24)]),
		.ic_scr_key_req_o(shadow_outputs_d[166]),
		.irq_software_i(shadow_inputs_q[0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 24 : ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 0)]),
		.irq_timer_i(shadow_inputs_q[0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 23 : ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 1)]),
		.irq_external_i(shadow_inputs_q[0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 22 : ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 2)]),
		.irq_fast_i(shadow_inputs_q[((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 21 : ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 3) : (0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 21 : ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 3)) + 14)-:15]),
		.irq_nm_i(shadow_inputs_q[0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 6 : ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 18)]),
		.irq_pending_o(shadow_outputs_d[165]),
		.debug_req_i(shadow_inputs_q[0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 5 : ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 19)]),
		.crash_dump_o(shadow_outputs_d[164-:160]),
		.double_fault_seen_o(shadow_outputs_d[4]),
		.fetch_enable_i(shadow_inputs_q[((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 4 : ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 20) : (0 + ((((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 24) >= 0 ? 4 : ((((((2 + MemDataWidth) + 3) + MemDataWidth) + 1) + RegFileDataWidth) + RegFileDataWidth) + 20)) + 3)-:4]),
		.alert_minor_o(shadow_alert_minor),
		.alert_major_internal_o(shadow_alert_major_internal),
		.alert_major_bus_o(shadow_alert_major_bus),
		.core_busy_o(shadow_outputs_d[3-:4])
	);
	always @(posedge clk_i) shadow_outputs_q <= shadow_outputs_d;
	wire outputs_mismatch;
	assign outputs_mismatch = enable_cmp_q & (shadow_outputs_q != core_outputs_q[(((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + 3) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + 3) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) >= 0 ? 0 : (((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) + 0+:(((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + 3) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + 3) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166) >= 0 ? (((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 167 : 1 - ((((((((((((71 + MemDataWidth) + 18) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 166))]);
	assign alert_major_internal_o = outputs_mismatch | shadow_alert_major_internal;
	assign alert_major_bus_o = shadow_alert_major_bus;
	assign alert_minor_o = shadow_alert_minor;
endmodule
module ibex_multdiv_fast (
	clk_i,
	rst_ni,
	mult_en_i,
	div_en_i,
	mult_sel_i,
	div_sel_i,
	operator_i,
	signed_mode_i,
	op_a_i,
	op_b_i,
	alu_adder_ext_i,
	alu_adder_i,
	equal_to_zero_i,
	data_ind_timing_i,
	alu_operand_a_o,
	alu_operand_b_o,
	imd_val_q_i,
	imd_val_d_o,
	imd_val_we_o,
	multdiv_ready_id_i,
	multdiv_result_o,
	valid_o
);
	parameter integer RV32M = 32'sd2;
	input wire clk_i;
	input wire rst_ni;
	input wire mult_en_i;
	input wire div_en_i;
	input wire mult_sel_i;
	input wire div_sel_i;
	input wire [1:0] operator_i;
	input wire [1:0] signed_mode_i;
	input wire [31:0] op_a_i;
	input wire [31:0] op_b_i;
	input wire [33:0] alu_adder_ext_i;
	input wire [31:0] alu_adder_i;
	input wire equal_to_zero_i;
	input wire data_ind_timing_i;
	output reg [32:0] alu_operand_a_o;
	output reg [32:0] alu_operand_b_o;
	input wire [67:0] imd_val_q_i;
	output wire [67:0] imd_val_d_o;
	output wire [1:0] imd_val_we_o;
	input wire multdiv_ready_id_i;
	output wire [31:0] multdiv_result_o;
	output wire valid_o;
	wire signed [34:0] mac_res_signed;
	wire [34:0] mac_res_ext;
	reg [33:0] accum;
	reg sign_a;
	reg sign_b;
	reg mult_valid;
	wire signed_mult;
	reg [33:0] mac_res_d;
	reg [33:0] op_remainder_d;
	wire [33:0] mac_res;
	wire div_sign_a;
	wire div_sign_b;
	reg is_greater_equal;
	wire div_change_sign;
	wire rem_change_sign;
	wire [31:0] one_shift;
	wire [31:0] op_denominator_q;
	reg [31:0] op_numerator_q;
	reg [31:0] op_quotient_q;
	reg [31:0] op_denominator_d;
	reg [31:0] op_numerator_d;
	reg [31:0] op_quotient_d;
	wire [31:0] next_remainder;
	wire [32:0] next_quotient;
	wire [31:0] res_adder_h;
	reg div_valid;
	reg [4:0] div_counter_q;
	reg [4:0] div_counter_d;
	wire multdiv_en;
	reg mult_hold;
	reg div_hold;
	reg div_by_zero_d;
	reg div_by_zero_q;
	wire mult_en_internal;
	wire div_en_internal;
	reg [2:0] md_state_q;
	reg [2:0] md_state_d;
	wire unused_mult_sel_i;
	assign unused_mult_sel_i = mult_sel_i;
	assign mult_en_internal = mult_en_i & ~mult_hold;
	assign div_en_internal = div_en_i & ~div_hold;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			div_counter_q <= 1'sb0;
			md_state_q <= 3'd0;
			op_numerator_q <= 1'sb0;
			op_quotient_q <= 1'sb0;
			div_by_zero_q <= 1'sb0;
		end
		else if (div_en_internal) begin
			div_counter_q <= div_counter_d;
			op_numerator_q <= op_numerator_d;
			op_quotient_q <= op_quotient_d;
			md_state_q <= md_state_d;
			div_by_zero_q <= div_by_zero_d;
		end
	assign multdiv_en = mult_en_internal | div_en_internal;
	assign imd_val_d_o[34+:34] = (div_sel_i ? op_remainder_d : mac_res_d);
	assign imd_val_we_o[0] = multdiv_en;
	assign imd_val_d_o[0+:34] = {2'b00, op_denominator_d};
	assign imd_val_we_o[1] = div_en_internal;
	assign op_denominator_q = imd_val_q_i[31-:32];
	wire [1:0] unused_imd_val;
	assign unused_imd_val = imd_val_q_i[33-:2];
	wire unused_mac_res_ext;
	assign unused_mac_res_ext = mac_res_ext[34];
	assign signed_mult = signed_mode_i != 2'b00;
	assign multdiv_result_o = (div_sel_i ? imd_val_q_i[65-:32] : mac_res_d[31:0]);
	generate
		if (RV32M == 32'sd3) begin : gen_mult_single_cycle
			reg mult_state_q;
			reg mult_state_d;
			wire signed [33:0] mult1_res;
			wire signed [33:0] mult2_res;
			wire signed [33:0] mult3_res;
			wire [33:0] mult1_res_uns;
			wire [33:32] unused_mult1_res_uns;
			wire [15:0] mult1_op_a;
			wire [15:0] mult1_op_b;
			wire [15:0] mult2_op_a;
			wire [15:0] mult2_op_b;
			reg [15:0] mult3_op_a;
			reg [15:0] mult3_op_b;
			wire mult1_sign_a;
			wire mult1_sign_b;
			wire mult2_sign_a;
			wire mult2_sign_b;
			reg mult3_sign_a;
			reg mult3_sign_b;
			reg [33:0] summand1;
			reg [33:0] summand2;
			reg [33:0] summand3;
			assign mult1_res = $signed({mult1_sign_a, mult1_op_a}) * $signed({mult1_sign_b, mult1_op_b});
			assign mult2_res = $signed({mult2_sign_a, mult2_op_a}) * $signed({mult2_sign_b, mult2_op_b});
			assign mult3_res = $signed({mult3_sign_a, mult3_op_a}) * $signed({mult3_sign_b, mult3_op_b});
			assign mac_res_signed = ($signed(summand1) + $signed(summand2)) + $signed(summand3);
			assign mult1_res_uns = $unsigned(mult1_res);
			assign mac_res_ext = $unsigned(mac_res_signed);
			assign mac_res = mac_res_ext[33:0];
			wire [1:1] sv2v_tmp_822BD;
			assign sv2v_tmp_822BD = signed_mode_i[0] & op_a_i[31];
			always @(*) sign_a = sv2v_tmp_822BD;
			wire [1:1] sv2v_tmp_4DE54;
			assign sv2v_tmp_4DE54 = signed_mode_i[1] & op_b_i[31];
			always @(*) sign_b = sv2v_tmp_4DE54;
			assign mult1_sign_a = 1'b0;
			assign mult1_sign_b = 1'b0;
			assign mult1_op_a = op_a_i[15:0];
			assign mult1_op_b = op_b_i[15:0];
			assign mult2_sign_a = 1'b0;
			assign mult2_sign_b = sign_b;
			assign mult2_op_a = op_a_i[15:0];
			assign mult2_op_b = op_b_i[31:16];
			wire [18:1] sv2v_tmp_915C6;
			assign sv2v_tmp_915C6 = imd_val_q_i[67-:18];
			always @(*) accum[17:0] = sv2v_tmp_915C6;
			wire [16:1] sv2v_tmp_2094F;
			assign sv2v_tmp_2094F = {16 {signed_mult & imd_val_q_i[67]}};
			always @(*) accum[33:18] = sv2v_tmp_2094F;
			always @(*) begin
				mult3_sign_a = sign_a;
				mult3_sign_b = 1'b0;
				mult3_op_a = op_a_i[31:16];
				mult3_op_b = op_b_i[15:0];
				summand1 = {18'h00000, mult1_res_uns[31:16]};
				summand2 = $unsigned(mult2_res);
				summand3 = $unsigned(mult3_res);
				mac_res_d = {2'b00, mac_res[15:0], mult1_res_uns[15:0]};
				mult_valid = mult_en_i;
				mult_state_d = 1'd0;
				mult_hold = 1'b0;
				case (mult_state_q)
					1'd0:
						if (operator_i != 2'd0) begin
							mac_res_d = mac_res;
							mult_valid = 1'b0;
							mult_state_d = 1'd1;
						end
						else
							mult_hold = ~multdiv_ready_id_i;
					1'd1: begin
						mult3_sign_a = sign_a;
						mult3_sign_b = sign_b;
						mult3_op_a = op_a_i[31:16];
						mult3_op_b = op_b_i[31:16];
						mac_res_d = mac_res;
						summand1 = 1'sb0;
						summand2 = accum;
						summand3 = $unsigned(mult3_res);
						mult_state_d = 1'd0;
						mult_valid = 1'b1;
						mult_hold = ~multdiv_ready_id_i;
					end
					default: mult_state_d = 1'd0;
				endcase
			end
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mult_state_q <= 1'd0;
				else if (mult_en_internal)
					mult_state_q <= mult_state_d;
			assign unused_mult1_res_uns = mult1_res_uns[33:32];
		end
		else begin : gen_mult_fast
			reg [15:0] mult_op_a;
			reg [15:0] mult_op_b;
			reg [1:0] mult_state_q;
			reg [1:0] mult_state_d;
			assign mac_res_signed = ($signed({sign_a, mult_op_a}) * $signed({sign_b, mult_op_b})) + $signed(accum);
			assign mac_res_ext = $unsigned(mac_res_signed);
			assign mac_res = mac_res_ext[33:0];
			always @(*) begin
				mult_op_a = op_a_i[15:0];
				mult_op_b = op_b_i[15:0];
				sign_a = 1'b0;
				sign_b = 1'b0;
				accum = imd_val_q_i[34+:34];
				mac_res_d = mac_res;
				mult_state_d = mult_state_q;
				mult_valid = 1'b0;
				mult_hold = 1'b0;
				case (mult_state_q)
					2'd0: begin
						mult_op_a = op_a_i[15:0];
						mult_op_b = op_b_i[15:0];
						sign_a = 1'b0;
						sign_b = 1'b0;
						accum = 1'sb0;
						mac_res_d = mac_res;
						mult_state_d = 2'd1;
					end
					2'd1: begin
						mult_op_a = op_a_i[15:0];
						mult_op_b = op_b_i[31:16];
						sign_a = 1'b0;
						sign_b = signed_mode_i[1] & op_b_i[31];
						accum = {18'b000000000000000000, imd_val_q_i[65-:16]};
						if (operator_i == 2'd0)
							mac_res_d = {2'b00, mac_res[15:0], imd_val_q_i[49-:16]};
						else
							mac_res_d = mac_res;
						mult_state_d = 2'd2;
					end
					2'd2: begin
						mult_op_a = op_a_i[31:16];
						mult_op_b = op_b_i[15:0];
						sign_a = signed_mode_i[0] & op_a_i[31];
						sign_b = 1'b0;
						if (operator_i == 2'd0) begin
							accum = {18'b000000000000000000, imd_val_q_i[65-:16]};
							mac_res_d = {2'b00, mac_res[15:0], imd_val_q_i[49-:16]};
							mult_valid = 1'b1;
							mult_state_d = 2'd0;
							mult_hold = ~multdiv_ready_id_i;
						end
						else begin
							accum = imd_val_q_i[34+:34];
							mac_res_d = mac_res;
							mult_state_d = 2'd3;
						end
					end
					2'd3: begin
						mult_op_a = op_a_i[31:16];
						mult_op_b = op_b_i[31:16];
						sign_a = signed_mode_i[0] & op_a_i[31];
						sign_b = signed_mode_i[1] & op_b_i[31];
						accum[17:0] = imd_val_q_i[67-:18];
						accum[33:18] = {16 {signed_mult & imd_val_q_i[67]}};
						mac_res_d = mac_res;
						mult_valid = 1'b1;
						mult_state_d = 2'd0;
						mult_hold = ~multdiv_ready_id_i;
					end
					default: mult_state_d = 2'd0;
				endcase
			end
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mult_state_q <= 2'd0;
				else if (mult_en_internal)
					mult_state_q <= mult_state_d;
		end
	endgenerate
	assign res_adder_h = alu_adder_ext_i[32:1];
	wire [1:0] unused_alu_adder_ext;
	assign unused_alu_adder_ext = {alu_adder_ext_i[33], alu_adder_ext_i[0]};
	assign next_remainder = (is_greater_equal ? res_adder_h[31:0] : imd_val_q_i[65-:32]);
	assign next_quotient = (is_greater_equal ? {1'b0, op_quotient_q} | {1'b0, one_shift} : {1'b0, op_quotient_q});
	assign one_shift = 32'b00000000000000000000000000000001 << div_counter_q;
	always @(*)
		if ((imd_val_q_i[65] ^ op_denominator_q[31]) == 1'b0)
			is_greater_equal = res_adder_h[31] == 1'b0;
		else
			is_greater_equal = imd_val_q_i[65];
	assign div_sign_a = op_a_i[31] & signed_mode_i[0];
	assign div_sign_b = op_b_i[31] & signed_mode_i[1];
	assign div_change_sign = (div_sign_a ^ div_sign_b) & ~div_by_zero_q;
	assign rem_change_sign = div_sign_a;
	always @(*) begin
		div_counter_d = div_counter_q - 5'h01;
		op_remainder_d = imd_val_q_i[34+:34];
		op_quotient_d = op_quotient_q;
		md_state_d = md_state_q;
		op_numerator_d = op_numerator_q;
		op_denominator_d = op_denominator_q;
		alu_operand_a_o = 33'b000000000000000000000000000000001;
		alu_operand_b_o = {~op_b_i, 1'b1};
		div_valid = 1'b0;
		div_hold = 1'b0;
		div_by_zero_d = div_by_zero_q;
		case (md_state_q)
			3'd0: begin
				if (operator_i == 2'd2) begin
					op_remainder_d = 1'sb1;
					md_state_d = (!data_ind_timing_i && equal_to_zero_i ? 3'd6 : 3'd1);
					div_by_zero_d = equal_to_zero_i;
				end
				else begin
					op_remainder_d = {2'b00, op_a_i};
					md_state_d = (!data_ind_timing_i && equal_to_zero_i ? 3'd6 : 3'd1);
				end
				alu_operand_a_o = 33'b000000000000000000000000000000001;
				alu_operand_b_o = {~op_b_i, 1'b1};
				div_counter_d = 5'd31;
			end
			3'd1: begin
				op_quotient_d = 1'sb0;
				op_numerator_d = (div_sign_a ? alu_adder_i : op_a_i);
				md_state_d = 3'd2;
				div_counter_d = 5'd31;
				alu_operand_a_o = 33'b000000000000000000000000000000001;
				alu_operand_b_o = {~op_a_i, 1'b1};
			end
			3'd2: begin
				op_remainder_d = {33'h000000000, op_numerator_q[31]};
				op_denominator_d = (div_sign_b ? alu_adder_i : op_b_i);
				md_state_d = 3'd3;
				div_counter_d = 5'd31;
				alu_operand_a_o = 33'b000000000000000000000000000000001;
				alu_operand_b_o = {~op_b_i, 1'b1};
			end
			3'd3: begin
				op_remainder_d = {1'b0, next_remainder[31:0], op_numerator_q[div_counter_d]};
				op_quotient_d = next_quotient[31:0];
				md_state_d = (div_counter_q == 5'd1 ? 3'd4 : 3'd3);
				alu_operand_a_o = {imd_val_q_i[65-:32], 1'b1};
				alu_operand_b_o = {~op_denominator_q[31:0], 1'b1};
			end
			3'd4: begin
				if (operator_i == 2'd2)
					op_remainder_d = {1'b0, next_quotient};
				else
					op_remainder_d = {2'b00, next_remainder[31:0]};
				alu_operand_a_o = {imd_val_q_i[65-:32], 1'b1};
				alu_operand_b_o = {~op_denominator_q[31:0], 1'b1};
				md_state_d = 3'd5;
			end
			3'd5: begin
				md_state_d = 3'd6;
				if (operator_i == 2'd2)
					op_remainder_d = (div_change_sign ? {2'h0, alu_adder_i} : imd_val_q_i[34+:34]);
				else
					op_remainder_d = (rem_change_sign ? {2'h0, alu_adder_i} : imd_val_q_i[34+:34]);
				alu_operand_a_o = 33'b000000000000000000000000000000001;
				alu_operand_b_o = {~imd_val_q_i[65-:32], 1'b1};
			end
			3'd6: begin
				md_state_d = 3'd0;
				div_hold = ~multdiv_ready_id_i;
				div_valid = 1'b1;
			end
			default: md_state_d = 3'd0;
		endcase
	end
	assign valid_o = mult_valid | div_valid;
endmodule
module ibex_multdiv_slow (
	clk_i,
	rst_ni,
	mult_en_i,
	div_en_i,
	mult_sel_i,
	div_sel_i,
	operator_i,
	signed_mode_i,
	op_a_i,
	op_b_i,
	alu_adder_ext_i,
	alu_adder_i,
	equal_to_zero_i,
	data_ind_timing_i,
	alu_operand_a_o,
	alu_operand_b_o,
	imd_val_q_i,
	imd_val_d_o,
	imd_val_we_o,
	multdiv_ready_id_i,
	multdiv_result_o,
	valid_o
);
	input wire clk_i;
	input wire rst_ni;
	input wire mult_en_i;
	input wire div_en_i;
	input wire mult_sel_i;
	input wire div_sel_i;
	input wire [1:0] operator_i;
	input wire [1:0] signed_mode_i;
	input wire [31:0] op_a_i;
	input wire [31:0] op_b_i;
	input wire [33:0] alu_adder_ext_i;
	input wire [31:0] alu_adder_i;
	input wire equal_to_zero_i;
	input wire data_ind_timing_i;
	output reg [32:0] alu_operand_a_o;
	output reg [32:0] alu_operand_b_o;
	input wire [67:0] imd_val_q_i;
	output wire [67:0] imd_val_d_o;
	output wire [1:0] imd_val_we_o;
	input wire multdiv_ready_id_i;
	output wire [31:0] multdiv_result_o;
	output wire valid_o;
	reg [2:0] md_state_q;
	reg [2:0] md_state_d;
	wire [32:0] accum_window_q;
	reg [32:0] accum_window_d;
	wire unused_imd_val0;
	wire [1:0] unused_imd_val1;
	wire [32:0] res_adder_l;
	wire [32:0] res_adder_h;
	reg [4:0] multdiv_count_q;
	reg [4:0] multdiv_count_d;
	reg [32:0] op_b_shift_q;
	reg [32:0] op_b_shift_d;
	reg [32:0] op_a_shift_q;
	reg [32:0] op_a_shift_d;
	wire [32:0] op_a_ext;
	wire [32:0] op_b_ext;
	wire [32:0] one_shift;
	wire [32:0] op_a_bw_pp;
	wire [32:0] op_a_bw_last_pp;
	wire [31:0] b_0;
	wire sign_a;
	wire sign_b;
	wire [32:0] next_quotient;
	wire [31:0] next_remainder;
	wire [31:0] op_numerator_q;
	reg [31:0] op_numerator_d;
	wire is_greater_equal;
	wire div_change_sign;
	wire rem_change_sign;
	reg div_by_zero_d;
	reg div_by_zero_q;
	reg multdiv_hold;
	wire multdiv_en;
	assign res_adder_l = alu_adder_ext_i[32:0];
	assign res_adder_h = alu_adder_ext_i[33:1];
	assign imd_val_d_o[34+:34] = {1'b0, accum_window_d};
	assign imd_val_we_o[0] = ~multdiv_hold;
	assign accum_window_q = imd_val_q_i[66-:33];
	assign unused_imd_val0 = imd_val_q_i[67];
	assign imd_val_d_o[0+:34] = {2'b00, op_numerator_d};
	assign imd_val_we_o[1] = multdiv_en;
	assign op_numerator_q = imd_val_q_i[31-:32];
	assign unused_imd_val1 = imd_val_q_i[33-:2];
	always @(*) begin
		alu_operand_a_o = accum_window_q;
		case (operator_i)
			2'd0: alu_operand_b_o = op_a_bw_pp;
			2'd1: alu_operand_b_o = (md_state_q == 3'd4 ? op_a_bw_last_pp : op_a_bw_pp);
			2'd2, 2'd3:
				case (md_state_q)
					3'd0: begin
						alu_operand_a_o = 33'b000000000000000000000000000000001;
						alu_operand_b_o = {~op_b_i, 1'b1};
					end
					3'd1: begin
						alu_operand_a_o = 33'b000000000000000000000000000000001;
						alu_operand_b_o = {~op_a_i, 1'b1};
					end
					3'd2: begin
						alu_operand_a_o = 33'b000000000000000000000000000000001;
						alu_operand_b_o = {~op_b_i, 1'b1};
					end
					3'd5: begin
						alu_operand_a_o = 33'b000000000000000000000000000000001;
						alu_operand_b_o = {~accum_window_q[31:0], 1'b1};
					end
					default: begin
						alu_operand_a_o = {accum_window_q[31:0], 1'b1};
						alu_operand_b_o = {~op_b_shift_q[31:0], 1'b1};
					end
				endcase
			default: begin
				alu_operand_a_o = accum_window_q;
				alu_operand_b_o = {~op_b_shift_q[31:0], 1'b1};
			end
		endcase
	end
	assign b_0 = {32 {op_b_shift_q[0]}};
	assign op_a_bw_pp = {~(op_a_shift_q[32] & op_b_shift_q[0]), op_a_shift_q[31:0] & b_0};
	assign op_a_bw_last_pp = {op_a_shift_q[32] & op_b_shift_q[0], ~(op_a_shift_q[31:0] & b_0)};
	assign sign_a = op_a_i[31] & signed_mode_i[0];
	assign sign_b = op_b_i[31] & signed_mode_i[1];
	assign op_a_ext = {sign_a, op_a_i};
	assign op_b_ext = {sign_b, op_b_i};
	assign is_greater_equal = (accum_window_q[31] == op_b_shift_q[31] ? ~res_adder_h[31] : accum_window_q[31]);
	assign one_shift = 33'b000000000000000000000000000000001 << multdiv_count_q;
	assign next_remainder = (is_greater_equal ? res_adder_h[31:0] : accum_window_q[31:0]);
	assign next_quotient = (is_greater_equal ? op_a_shift_q | one_shift : op_a_shift_q);
	assign div_change_sign = (sign_a ^ sign_b) & ~div_by_zero_q;
	assign rem_change_sign = sign_a;
	always @(*) begin
		multdiv_count_d = multdiv_count_q;
		accum_window_d = accum_window_q;
		op_b_shift_d = op_b_shift_q;
		op_a_shift_d = op_a_shift_q;
		op_numerator_d = op_numerator_q;
		md_state_d = md_state_q;
		multdiv_hold = 1'b0;
		div_by_zero_d = div_by_zero_q;
		if (mult_sel_i || div_sel_i)
			case (md_state_q)
				3'd0: begin
					case (operator_i)
						2'd0: begin
							op_a_shift_d = op_a_ext << 1;
							accum_window_d = {~(op_a_ext[32] & op_b_i[0]), op_a_ext[31:0] & {32 {op_b_i[0]}}};
							op_b_shift_d = op_b_ext >> 1;
							md_state_d = (!data_ind_timing_i && ((op_b_ext >> 1) == 0) ? 3'd4 : 3'd3);
						end
						2'd1: begin
							op_a_shift_d = op_a_ext;
							accum_window_d = {1'b1, ~(op_a_ext[32] & op_b_i[0]), op_a_ext[31:1] & {31 {op_b_i[0]}}};
							op_b_shift_d = op_b_ext >> 1;
							md_state_d = 3'd3;
						end
						2'd2: begin
							accum_window_d = {33 {1'b1}};
							md_state_d = (!data_ind_timing_i && equal_to_zero_i ? 3'd6 : 3'd1);
							div_by_zero_d = equal_to_zero_i;
						end
						2'd3: begin
							accum_window_d = op_a_ext;
							md_state_d = (!data_ind_timing_i && equal_to_zero_i ? 3'd6 : 3'd1);
						end
						default:
							;
					endcase
					multdiv_count_d = 5'd31;
				end
				3'd1: begin
					op_a_shift_d = 1'sb0;
					op_numerator_d = (sign_a ? alu_adder_i : op_a_i);
					md_state_d = 3'd2;
				end
				3'd2: begin
					accum_window_d = {32'h00000000, op_numerator_q[31]};
					op_b_shift_d = (sign_b ? {1'b0, alu_adder_i} : {1'b0, op_b_i});
					md_state_d = 3'd3;
				end
				3'd3: begin
					multdiv_count_d = multdiv_count_q - 5'h01;
					case (operator_i)
						2'd0: begin
							accum_window_d = res_adder_l;
							op_a_shift_d = op_a_shift_q << 1;
							op_b_shift_d = op_b_shift_q >> 1;
							md_state_d = ((!data_ind_timing_i && (op_b_shift_d == 0)) || (multdiv_count_q == 5'd1) ? 3'd4 : 3'd3);
						end
						2'd1: begin
							accum_window_d = res_adder_h;
							op_a_shift_d = op_a_shift_q;
							op_b_shift_d = op_b_shift_q >> 1;
							md_state_d = (multdiv_count_q == 5'd1 ? 3'd4 : 3'd3);
						end
						2'd2, 2'd3: begin
							accum_window_d = {next_remainder[31:0], op_numerator_q[multdiv_count_d]};
							op_a_shift_d = next_quotient;
							md_state_d = (multdiv_count_q == 5'd1 ? 3'd4 : 3'd3);
						end
						default:
							;
					endcase
				end
				3'd4:
					case (operator_i)
						2'd0: begin
							accum_window_d = res_adder_l;
							md_state_d = 3'd0;
							multdiv_hold = ~multdiv_ready_id_i;
						end
						2'd1: begin
							accum_window_d = res_adder_l;
							md_state_d = 3'd0;
							md_state_d = 3'd0;
							multdiv_hold = ~multdiv_ready_id_i;
						end
						2'd2: begin
							accum_window_d = next_quotient;
							md_state_d = 3'd5;
						end
						2'd3: begin
							accum_window_d = {1'b0, next_remainder[31:0]};
							md_state_d = 3'd5;
						end
						default:
							;
					endcase
				3'd5: begin
					md_state_d = 3'd6;
					case (operator_i)
						2'd2: accum_window_d = (div_change_sign ? {1'b0, alu_adder_i} : accum_window_q);
						2'd3: accum_window_d = (rem_change_sign ? {1'b0, alu_adder_i} : accum_window_q);
						default:
							;
					endcase
				end
				3'd6: begin
					md_state_d = 3'd0;
					multdiv_hold = ~multdiv_ready_id_i;
				end
				default: md_state_d = 3'd0;
			endcase
	end
	assign multdiv_en = (mult_en_i | div_en_i) & ~multdiv_hold;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			multdiv_count_q <= 5'h00;
			op_b_shift_q <= 33'h000000000;
			op_a_shift_q <= 33'h000000000;
			md_state_q <= 3'd0;
			div_by_zero_q <= 1'b0;
		end
		else if (multdiv_en) begin
			multdiv_count_q <= multdiv_count_d;
			op_b_shift_q <= op_b_shift_d;
			op_a_shift_q <= op_a_shift_d;
			md_state_q <= md_state_d;
			div_by_zero_q <= div_by_zero_d;
		end
	assign valid_o = (md_state_q == 3'd6) | ((md_state_q == 3'd4) & ((operator_i == 2'd0) | (operator_i == 2'd1)));
	assign multdiv_result_o = (div_en_i ? accum_window_q[31:0] : res_adder_l[31:0]);
endmodule
module ibex_pmp (
	csr_pmp_cfg_i,
	csr_pmp_addr_i,
	csr_pmp_mseccfg_i,
	priv_mode_i,
	pmp_req_addr_i,
	pmp_req_type_i,
	pmp_req_err_o
);
	parameter [31:0] PMPGranularity = 0;
	parameter [31:0] PMPNumChan = 2;
	parameter [31:0] PMPNumRegions = 4;
	input wire [(PMPNumRegions * 6) - 1:0] csr_pmp_cfg_i;
	input wire [(PMPNumRegions * 34) - 1:0] csr_pmp_addr_i;
	input wire [2:0] csr_pmp_mseccfg_i;
	input wire [(PMPNumChan * 2) - 1:0] priv_mode_i;
	input wire [(PMPNumChan * 34) - 1:0] pmp_req_addr_i;
	input wire [(PMPNumChan * 2) - 1:0] pmp_req_type_i;
	output wire [0:PMPNumChan - 1] pmp_req_err_o;
	wire [33:0] region_start_addr [0:PMPNumRegions - 1];
	wire [33:PMPGranularity + 2] region_addr_mask [0:PMPNumRegions - 1];
	wire [(PMPNumChan * PMPNumRegions) - 1:0] region_match_gt;
	wire [(PMPNumChan * PMPNumRegions) - 1:0] region_match_lt;
	wire [(PMPNumChan * PMPNumRegions) - 1:0] region_match_eq;
	reg [(PMPNumChan * PMPNumRegions) - 1:0] region_match_all;
	wire [(PMPNumChan * PMPNumRegions) - 1:0] region_basic_perm_check;
	wire [(PMPNumChan * PMPNumRegions) - 1:0] region_perm_check;
	function automatic mml_perm_check;
		input reg [5:0] csr_pmp_cfg;
		input reg [1:0] pmp_req_type;
		input reg [1:0] priv_mode;
		input reg permission_check;
		reg result;
		reg unused_cfg;
		begin
			result = 1'b0;
			unused_cfg = |csr_pmp_cfg[4-:2];
			if (!csr_pmp_cfg[0] && csr_pmp_cfg[1])
				case ({csr_pmp_cfg[5], csr_pmp_cfg[2]})
					2'b00: result = (pmp_req_type == 2'b10) | ((pmp_req_type == 2'b01) & (priv_mode == 2'b11));
					2'b01: result = (pmp_req_type == 2'b10) | (pmp_req_type == 2'b01);
					2'b10: result = pmp_req_type == 2'b00;
					2'b11: result = (pmp_req_type == 2'b00) | ((pmp_req_type == 2'b10) & (priv_mode == 2'b11));
					default:
						;
				endcase
			else if (((csr_pmp_cfg[0] & csr_pmp_cfg[1]) & csr_pmp_cfg[2]) & csr_pmp_cfg[5])
				result = pmp_req_type == 2'b10;
			else
				result = permission_check & (priv_mode == 2'b11 ? csr_pmp_cfg[5] : ~csr_pmp_cfg[5]);
			mml_perm_check = result;
		end
	endfunction
	function automatic orig_perm_check;
		input reg pmp_cfg_lock;
		input reg [1:0] priv_mode;
		input reg permission_check;
		orig_perm_check = (priv_mode == 2'b11 ? ~pmp_cfg_lock | permission_check : permission_check);
	endfunction
	function automatic perm_check_wrapper;
		input reg csr_pmp_mseccfg_mml;
		input reg [5:0] csr_pmp_cfg;
		input reg [1:0] pmp_req_type;
		input reg [1:0] priv_mode;
		input reg permission_check;
		perm_check_wrapper = (csr_pmp_mseccfg_mml ? mml_perm_check(csr_pmp_cfg, pmp_req_type, priv_mode, permission_check) : orig_perm_check(csr_pmp_cfg[5], priv_mode, permission_check));
	endfunction
	function automatic access_fault_check;
		input reg csr_pmp_mseccfg_mmwp;
		input reg csr_pmp_mseccfg_mml;
		input reg [1:0] pmp_req_type;
		input reg [PMPNumRegions - 1:0] match_all;
		input reg [1:0] priv_mode;
		input reg [PMPNumRegions - 1:0] final_perm_check;
		reg access_fail;
		reg matched;
		begin
			access_fail = (csr_pmp_mseccfg_mmwp | (priv_mode != 2'b11)) | (csr_pmp_mseccfg_mml && (pmp_req_type == 2'b00));
			matched = 1'b0;
			begin : sv2v_autoblock_1
				reg signed [31:0] r;
				for (r = 0; r < PMPNumRegions; r = r + 1)
					if (!matched && match_all[r]) begin
						access_fail = ~final_perm_check[r];
						matched = 1'b1;
					end
			end
			access_fault_check = access_fail;
		end
	endfunction
	genvar r;
	generate
		for (r = 0; r < PMPNumRegions; r = r + 1) begin : g_addr_exp
			if (r == 0) begin : g_entry0
				assign region_start_addr[r] = (csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 4-:2] == 2'b01 ? 34'h000000000 : csr_pmp_addr_i[((PMPNumRegions - 1) - r) * 34+:34]);
			end
			else begin : g_oth
				assign region_start_addr[r] = (csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 4-:2] == 2'b01 ? csr_pmp_addr_i[((PMPNumRegions - 1) - (r - 1)) * 34+:34] : csr_pmp_addr_i[((PMPNumRegions - 1) - r) * 34+:34]);
			end
			genvar b;
			for (b = PMPGranularity + 2; b < 34; b = b + 1) begin : g_bitmask
				if (b == 2) begin : g_bit0
					assign region_addr_mask[r][b] = csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 4-:2] != 2'b11;
				end
				else begin : g_others
					if (PMPGranularity == 0) begin : g_region_addr_mask_zero_granularity
						assign region_addr_mask[r][b] = (csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 4-:2] != 2'b11) | ~&csr_pmp_addr_i[(((PMPNumRegions - 1) - r) * 34) + ((b - 1) >= 2 ? b - 1 : ((b - 1) + ((b - 1) >= 2 ? b - 2 : 4 - b)) - 1)-:((b - 1) >= 2 ? b - 2 : 4 - b)];
					end
					else begin : g_region_addr_mask_other_granularity
						assign region_addr_mask[r][b] = (csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 4-:2] != 2'b11) | ~&csr_pmp_addr_i[(((PMPNumRegions - 1) - r) * 34) + ((b - 1) >= (PMPGranularity + 1) ? b - 1 : ((b - 1) + ((b - 1) >= (PMPGranularity + 1) ? ((b - 1) - (PMPGranularity + 1)) + 1 : ((PMPGranularity + 1) - (b - 1)) + 1)) - 1)-:((b - 1) >= (PMPGranularity + 1) ? ((b - 1) - (PMPGranularity + 1)) + 1 : ((PMPGranularity + 1) - (b - 1)) + 1)];
					end
				end
			end
		end
	endgenerate
	genvar c;
	generate
		for (c = 0; c < PMPNumChan; c = c + 1) begin : g_access_check
			genvar r;
			for (r = 0; r < PMPNumRegions; r = r + 1) begin : g_regions
				assign region_match_eq[(c * PMPNumRegions) + r] = (pmp_req_addr_i[(((PMPNumChan - 1) - c) * 34) + (33 >= (PMPGranularity + 2) ? 33 : (33 + (33 >= (PMPGranularity + 2) ? 34 - (PMPGranularity + 2) : PMPGranularity - 30)) - 1)-:(33 >= (PMPGranularity + 2) ? 34 - (PMPGranularity + 2) : PMPGranularity - 30)] & region_addr_mask[r]) == (region_start_addr[r][33:PMPGranularity + 2] & region_addr_mask[r]);
				assign region_match_gt[(c * PMPNumRegions) + r] = pmp_req_addr_i[(((PMPNumChan - 1) - c) * 34) + (33 >= (PMPGranularity + 2) ? 33 : (33 + (33 >= (PMPGranularity + 2) ? 34 - (PMPGranularity + 2) : PMPGranularity - 30)) - 1)-:(33 >= (PMPGranularity + 2) ? 34 - (PMPGranularity + 2) : PMPGranularity - 30)] > region_start_addr[r][33:PMPGranularity + 2];
				assign region_match_lt[(c * PMPNumRegions) + r] = pmp_req_addr_i[(((PMPNumChan - 1) - c) * 34) + (33 >= (PMPGranularity + 2) ? 33 : (33 + (33 >= (PMPGranularity + 2) ? 34 - (PMPGranularity + 2) : PMPGranularity - 30)) - 1)-:(33 >= (PMPGranularity + 2) ? 34 - (PMPGranularity + 2) : PMPGranularity - 30)] < csr_pmp_addr_i[(((PMPNumRegions - 1) - r) * 34) + (33 >= (PMPGranularity + 2) ? 33 : (33 + (33 >= (PMPGranularity + 2) ? 34 - (PMPGranularity + 2) : PMPGranularity - 30)) - 1)-:(33 >= (PMPGranularity + 2) ? 34 - (PMPGranularity + 2) : PMPGranularity - 30)];
				always @(*) begin
					region_match_all[(c * PMPNumRegions) + r] = 1'b0;
					case (csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 4-:2])
						2'b00: region_match_all[(c * PMPNumRegions) + r] = 1'b0;
						2'b10: region_match_all[(c * PMPNumRegions) + r] = region_match_eq[(c * PMPNumRegions) + r];
						2'b11: region_match_all[(c * PMPNumRegions) + r] = region_match_eq[(c * PMPNumRegions) + r];
						2'b01: region_match_all[(c * PMPNumRegions) + r] = (region_match_eq[(c * PMPNumRegions) + r] | region_match_gt[(c * PMPNumRegions) + r]) & region_match_lt[(c * PMPNumRegions) + r];
						default: region_match_all[(c * PMPNumRegions) + r] = 1'b0;
					endcase
				end
				assign region_basic_perm_check[(c * PMPNumRegions) + r] = (((pmp_req_type_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b00) & csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 2]) | ((pmp_req_type_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b01) & csr_pmp_cfg_i[(((PMPNumRegions - 1) - r) * 6) + 1])) | ((pmp_req_type_i[((PMPNumChan - 1) - c) * 2+:2] == 2'b10) & csr_pmp_cfg_i[((PMPNumRegions - 1) - r) * 6]);
				assign region_perm_check[(c * PMPNumRegions) + r] = perm_check_wrapper(csr_pmp_mseccfg_i[0], csr_pmp_cfg_i[((PMPNumRegions - 1) - r) * 6+:6], pmp_req_type_i[((PMPNumChan - 1) - c) * 2+:2], priv_mode_i[((PMPNumChan - 1) - c) * 2+:2], region_basic_perm_check[(c * PMPNumRegions) + r]);
				wire unused_sigs;
				assign unused_sigs = ^{region_start_addr[r][PMPGranularity + 1:0], pmp_req_addr_i[(((PMPNumChan - 1) - c) * 34) + ((PMPGranularity + 1) >= 0 ? PMPGranularity + 1 : ((PMPGranularity + 1) + ((PMPGranularity + 1) >= 0 ? PMPGranularity + 2 : 1 - (PMPGranularity + 1))) - 1)-:((PMPGranularity + 1) >= 0 ? PMPGranularity + 2 : 1 - (PMPGranularity + 1))]};
			end
			assign pmp_req_err_o[c] = access_fault_check(csr_pmp_mseccfg_i[1], csr_pmp_mseccfg_i[0], pmp_req_type_i[((PMPNumChan - 1) - c) * 2+:2], region_match_all[c * PMPNumRegions+:PMPNumRegions], priv_mode_i[((PMPNumChan - 1) - c) * 2+:2], region_perm_check[c * PMPNumRegions+:PMPNumRegions]);
		end
	endgenerate
	wire unused_csr_pmp_mseccfg_rlb;
	assign unused_csr_pmp_mseccfg_rlb = csr_pmp_mseccfg_i[2];
endmodule
module ibex_prefetch_buffer (
	clk_i,
	rst_ni,
	req_i,
	branch_i,
	addr_i,
	ready_i,
	valid_o,
	rdata_o,
	addr_o,
	err_o,
	err_plus2_o,
	instr_req_o,
	instr_gnt_i,
	instr_addr_o,
	instr_rdata_i,
	instr_err_i,
	instr_rvalid_i,
	busy_o
);
	parameter [0:0] ResetAll = 1'b0;
	input wire clk_i;
	input wire rst_ni;
	input wire req_i;
	input wire branch_i;
	input wire [31:0] addr_i;
	input wire ready_i;
	output wire valid_o;
	output wire [31:0] rdata_o;
	output wire [31:0] addr_o;
	output wire err_o;
	output wire err_plus2_o;
	output wire instr_req_o;
	input wire instr_gnt_i;
	output wire [31:0] instr_addr_o;
	input wire [31:0] instr_rdata_i;
	input wire instr_err_i;
	input wire instr_rvalid_i;
	output wire busy_o;
	localparam [31:0] NUM_REQS = 2;
	wire valid_new_req;
	wire valid_req;
	wire valid_req_d;
	reg valid_req_q;
	wire discard_req_d;
	reg discard_req_q;
	wire [1:0] rdata_outstanding_n;
	wire [1:0] rdata_outstanding_s;
	reg [1:0] rdata_outstanding_q;
	wire [1:0] branch_discard_n;
	wire [1:0] branch_discard_s;
	reg [1:0] branch_discard_q;
	wire [1:0] rdata_outstanding_rev;
	wire [31:0] stored_addr_d;
	reg [31:0] stored_addr_q;
	wire stored_addr_en;
	wire [31:0] fetch_addr_d;
	reg [31:0] fetch_addr_q;
	wire fetch_addr_en;
	wire [31:0] instr_addr;
	wire [31:0] instr_addr_w_aligned;
	wire fifo_valid;
	wire [31:0] fifo_addr;
	wire fifo_ready;
	wire fifo_clear;
	wire [1:0] fifo_busy;
	assign busy_o = |rdata_outstanding_q | instr_req_o;
	assign fifo_clear = branch_i;
	genvar i;
	generate
		for (i = 0; i < NUM_REQS; i = i + 1) begin : gen_rd_rev
			assign rdata_outstanding_rev[i] = rdata_outstanding_q[1 - i];
		end
	endgenerate
	assign fifo_ready = ~&(fifo_busy | rdata_outstanding_rev);
	ibex_fetch_fifo #(
		.NUM_REQS(NUM_REQS),
		.ResetAll(ResetAll)
	) fifo_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clear_i(fifo_clear),
		.busy_o(fifo_busy),
		.in_valid_i(fifo_valid),
		.in_addr_i(fifo_addr),
		.in_rdata_i(instr_rdata_i),
		.in_err_i(instr_err_i),
		.out_valid_o(valid_o),
		.out_ready_i(ready_i),
		.out_rdata_o(rdata_o),
		.out_addr_o(addr_o),
		.out_err_o(err_o),
		.out_err_plus2_o(err_plus2_o)
	);
	assign valid_new_req = (req_i & (fifo_ready | branch_i)) & ~rdata_outstanding_q[1];
	assign valid_req = valid_req_q | valid_new_req;
	assign valid_req_d = valid_req & ~instr_gnt_i;
	assign discard_req_d = valid_req_q & (branch_i | discard_req_q);
	assign stored_addr_en = (valid_new_req & ~valid_req_q) & ~instr_gnt_i;
	assign stored_addr_d = instr_addr;
	generate
		if (ResetAll) begin : g_stored_addr_ra
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					stored_addr_q <= 1'sb0;
				else if (stored_addr_en)
					stored_addr_q <= stored_addr_d;
		end
		else begin : g_stored_addr_nr
			always @(posedge clk_i)
				if (stored_addr_en)
					stored_addr_q <= stored_addr_d;
		end
	endgenerate
	assign fetch_addr_en = branch_i | (valid_new_req & ~valid_req_q);
	assign fetch_addr_d = (branch_i ? addr_i : {fetch_addr_q[31:2], 2'b00}) + {{29 {1'b0}}, valid_new_req & ~valid_req_q, 2'b00};
	generate
		if (ResetAll) begin : g_fetch_addr_ra
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					fetch_addr_q <= 1'sb0;
				else if (fetch_addr_en)
					fetch_addr_q <= fetch_addr_d;
		end
		else begin : g_fetch_addr_nr
			always @(posedge clk_i)
				if (fetch_addr_en)
					fetch_addr_q <= fetch_addr_d;
		end
	endgenerate
	assign instr_addr = (valid_req_q ? stored_addr_q : (branch_i ? addr_i : fetch_addr_q));
	assign instr_addr_w_aligned = {instr_addr[31:2], 2'b00};
	generate
		for (i = 0; i < NUM_REQS; i = i + 1) begin : g_outstanding_reqs
			if (i == 0) begin : g_req0
				assign rdata_outstanding_n[i] = (valid_req & instr_gnt_i) | rdata_outstanding_q[i];
				assign branch_discard_n[i] = (((valid_req & instr_gnt_i) & discard_req_d) | (branch_i & rdata_outstanding_q[i])) | branch_discard_q[i];
			end
			else begin : g_reqtop
				assign rdata_outstanding_n[i] = ((valid_req & instr_gnt_i) & rdata_outstanding_q[i - 1]) | rdata_outstanding_q[i];
				assign branch_discard_n[i] = ((((valid_req & instr_gnt_i) & discard_req_d) & rdata_outstanding_q[i - 1]) | (branch_i & rdata_outstanding_q[i])) | branch_discard_q[i];
			end
		end
	endgenerate
	assign rdata_outstanding_s = (instr_rvalid_i ? {1'b0, rdata_outstanding_n[1:1]} : rdata_outstanding_n);
	assign branch_discard_s = (instr_rvalid_i ? {1'b0, branch_discard_n[1:1]} : branch_discard_n);
	assign fifo_valid = instr_rvalid_i & ~branch_discard_q[0];
	assign fifo_addr = addr_i;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			valid_req_q <= 1'b0;
			discard_req_q <= 1'b0;
			rdata_outstanding_q <= 'b0;
			branch_discard_q <= 'b0;
		end
		else begin
			valid_req_q <= valid_req_d;
			discard_req_q <= discard_req_d;
			rdata_outstanding_q <= rdata_outstanding_s;
			branch_discard_q <= branch_discard_s;
		end
	assign instr_req_o = valid_req;
	assign instr_addr_o = instr_addr_w_aligned;
endmodule
module ibex_register_file_ff (
	clk_i,
	rst_ni,
	test_en_i,
	dummy_instr_id_i,
	dummy_instr_wb_i,
	raddr_a_i,
	rdata_a_o,
	raddr_b_i,
	rdata_b_o,
	waddr_a_i,
	wdata_a_i,
	we_a_i,
	err_o
);
	parameter [0:0] RV32E = 0;
	parameter [31:0] DataWidth = 32;
	parameter [0:0] DummyInstructions = 0;
	parameter [0:0] WrenCheck = 0;
	parameter [DataWidth - 1:0] WordZeroVal = 1'sb0;
	input wire clk_i;
	input wire rst_ni;
	input wire test_en_i;
	input wire dummy_instr_id_i;
	input wire dummy_instr_wb_i;
	input wire [4:0] raddr_a_i;
	output wire [DataWidth - 1:0] rdata_a_o;
	input wire [4:0] raddr_b_i;
	output wire [DataWidth - 1:0] rdata_b_o;
	input wire [4:0] waddr_a_i;
	input wire [DataWidth - 1:0] wdata_a_i;
	input wire we_a_i;
	output wire err_o;
	localparam [31:0] ADDR_WIDTH = (RV32E ? 4 : 5);
	localparam [31:0] NUM_WORDS = 2 ** ADDR_WIDTH;
	wire [DataWidth - 1:0] rf_reg [0:NUM_WORDS - 1];
	reg [NUM_WORDS - 1:0] we_a_dec;
	function automatic [4:0] sv2v_cast_5;
		input reg [4:0] inp;
		sv2v_cast_5 = inp;
	endfunction
	always @(*) begin : we_a_decoder
		begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < NUM_WORDS; i = i + 1)
				we_a_dec[i] = (waddr_a_i == sv2v_cast_5(i) ? we_a_i : 1'b0);
		end
	end
	generate
		if (WrenCheck) begin : gen_wren_check
			wire [NUM_WORDS - 1:0] we_a_dec_buf;
			prim_buf #(.Width(NUM_WORDS)) u_prim_buf(
				.in_i(we_a_dec),
				.out_o(we_a_dec_buf)
			);
			prim_onehot_check #(
				.AddrWidth(ADDR_WIDTH),
				.AddrCheck(1),
				.EnableCheck(1)
			) u_prim_onehot_check(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.oh_i(we_a_dec_buf),
				.addr_i(waddr_a_i),
				.en_i(we_a_i),
				.err_o(err_o)
			);
		end
		else begin : gen_no_wren_check
			wire unused_strobe;
			assign unused_strobe = we_a_dec[0];
			assign err_o = 1'b0;
		end
	endgenerate
	genvar i;
	generate
		for (i = 1; i < NUM_WORDS; i = i + 1) begin : g_rf_flops
			reg [DataWidth - 1:0] rf_reg_q;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					rf_reg_q <= WordZeroVal;
				else if (we_a_dec[i])
					rf_reg_q <= wdata_a_i;
			assign rf_reg[i] = rf_reg_q;
		end
		if (DummyInstructions) begin : g_dummy_r0
			wire we_r0_dummy;
			reg [DataWidth - 1:0] rf_r0_q;
			assign we_r0_dummy = we_a_i & dummy_instr_wb_i;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					rf_r0_q <= WordZeroVal;
				else if (we_r0_dummy)
					rf_r0_q <= wdata_a_i;
			assign rf_reg[0] = (dummy_instr_id_i ? rf_r0_q : WordZeroVal);
		end
		else begin : g_normal_r0
			wire unused_dummy_instr;
			assign unused_dummy_instr = dummy_instr_id_i ^ dummy_instr_wb_i;
			assign rf_reg[0] = WordZeroVal;
		end
	endgenerate
	assign rdata_a_o = rf_reg[raddr_a_i];
	assign rdata_b_o = rf_reg[raddr_b_i];
	wire unused_test_en;
	assign unused_test_en = test_en_i;
endmodule
module ibex_top (
	clk_i,
	rst_ni,
	test_en_i,
	ram_cfg_i,
	hart_id_i,
	boot_addr_i,
	instr_req_o,
	instr_gnt_i,
	instr_rvalid_i,
	instr_addr_o,
	instr_rdata_i,
	instr_rdata_intg_i,
	instr_err_i,
	data_req_o,
	data_gnt_i,
	data_rvalid_i,
	data_we_o,
	data_be_o,
	data_addr_o,
	data_wdata_o,
	data_wdata_intg_o,
	data_rdata_i,
	data_rdata_intg_i,
	data_err_i,
	irq_software_i,
	irq_timer_i,
	irq_external_i,
	irq_fast_i,
	irq_nm_i,
	scramble_key_valid_i,
	scramble_key_i,
	scramble_nonce_i,
	scramble_req_o,
	debug_req_i,
	crash_dump_o,
	double_fault_seen_o,
	fetch_enable_i,
	alert_minor_o,
	alert_major_internal_o,
	alert_major_bus_o,
	core_sleep_o,
	scan_rst_ni
);
	parameter [0:0] PMPEnable = 1'b0;
	parameter [31:0] PMPGranularity = 0;
	parameter [31:0] PMPNumRegions = 4;
	parameter [31:0] MHPMCounterNum = 0;
	parameter [31:0] MHPMCounterWidth = 40;
	parameter [0:0] RV32E = 1'b0;
	parameter integer RV32M = 32'sd1;
	parameter integer RV32B = 32'sd0;
	parameter integer RegFile = 32'sd0;
	parameter [0:0] BranchTargetALU = 1'b0;
	parameter [0:0] WritebackStage = 1'b0;
	parameter [0:0] ICache = 1'b0;
	parameter [0:0] ICacheECC = 1'b0;
	parameter [0:0] BranchPredictor = 1'b0;
	parameter [0:0] DbgTriggerEn = 1'b0;
	parameter [31:0] DbgHwBreakNum = 1;
	parameter [0:0] SecureIbex = 1'b1;
	parameter [0:0] ICacheScramble = 1'b0;
	localparam signed [31:0] ibex_pkg_LfsrWidth = 32;
	localparam [31:0] ibex_pkg_RndCnstLfsrSeedDefault = 32'hac533bf4;
	parameter [31:0] RndCnstLfsrSeed = ibex_pkg_RndCnstLfsrSeedDefault;
	localparam [159:0] ibex_pkg_RndCnstLfsrPermDefault = 160'h1e35ecba467fd1b12e958152c04fa43878a8daed;
	parameter [159:0] RndCnstLfsrPerm = ibex_pkg_RndCnstLfsrPermDefault;
	parameter [31:0] DmHaltAddr = 32'h1a110800;
	parameter [31:0] DmExceptionAddr = 32'h1a110808;
	localparam [31:0] ibex_pkg_SCRAMBLE_KEY_W = 128;
	localparam [127:0] ibex_pkg_RndCnstIbexKeyDefault = 128'h14e8cecae3040d5e12286bb3cc113298;
	parameter [127:0] RndCnstIbexKey = ibex_pkg_RndCnstIbexKeyDefault;
	localparam [31:0] ibex_pkg_SCRAMBLE_NONCE_W = 64;
	localparam [63:0] ibex_pkg_RndCnstIbexNonceDefault = 64'hf79780bc735f3843;
	parameter [63:0] RndCnstIbexNonce = ibex_pkg_RndCnstIbexNonceDefault;
	input wire clk_i;
	input wire rst_ni;
	input wire test_en_i;
	input wire [9:0] ram_cfg_i;
	input wire [31:0] hart_id_i;
	input wire [31:0] boot_addr_i;
	output wire instr_req_o;
	input wire instr_gnt_i;
	input wire instr_rvalid_i;
	output wire [31:0] instr_addr_o;
	input wire [31:0] instr_rdata_i;
	input wire [6:0] instr_rdata_intg_i;
	input wire instr_err_i;
	output wire data_req_o;
	input wire data_gnt_i;
	input wire data_rvalid_i;
	output wire data_we_o;
	output wire [3:0] data_be_o;
	output wire [31:0] data_addr_o;
	output wire [31:0] data_wdata_o;
	output wire [6:0] data_wdata_intg_o;
	input wire [31:0] data_rdata_i;
	input wire [6:0] data_rdata_intg_i;
	input wire data_err_i;
	input wire irq_software_i;
	input wire irq_timer_i;
	input wire irq_external_i;
	input wire [14:0] irq_fast_i;
	input wire irq_nm_i;
	input wire scramble_key_valid_i;
	input wire [127:0] scramble_key_i;
	input wire [63:0] scramble_nonce_i;
	output wire scramble_req_o;
	input wire debug_req_i;
	output wire [159:0] crash_dump_o;
	output wire double_fault_seen_o;
	input wire [3:0] fetch_enable_i;
	output wire alert_minor_o;
	output wire alert_major_internal_o;
	output wire alert_major_bus_o;
	output wire core_sleep_o;
	input wire scan_rst_ni;
	localparam [0:0] Lockstep = 1'b0;
	localparam [0:0] ResetAll = 1'b1;
	localparam [0:0] DummyInstructions = SecureIbex;
	localparam [0:0] RegFileECC = SecureIbex;
	localparam [0:0] RegFileWrenCheck = SecureIbex;
	localparam [31:0] RegFileDataWidth = (RegFileECC ? 39 : 32);
	localparam [0:0] MemECC = SecureIbex;
	localparam [31:0] MemDataWidth = (MemECC ? 39 : 32);
	localparam [31:0] ibex_pkg_BUS_SIZE = 32;
	localparam [31:0] BusSizeECC = (ICacheECC ? 39 : ibex_pkg_BUS_SIZE);
	localparam [31:0] ibex_pkg_BUS_BYTES = 4;
	localparam [31:0] ibex_pkg_IC_LINE_SIZE = 64;
	localparam [31:0] ibex_pkg_IC_LINE_BYTES = 8;
	localparam [31:0] ibex_pkg_IC_LINE_BEATS = ibex_pkg_IC_LINE_BYTES / ibex_pkg_BUS_BYTES;
	localparam [31:0] LineSizeECC = BusSizeECC * ibex_pkg_IC_LINE_BEATS;
	localparam [31:0] ibex_pkg_ADDR_W = 32;
	localparam [31:0] ibex_pkg_IC_NUM_WAYS = 2;
	localparam [31:0] ibex_pkg_IC_SIZE_BYTES = 4096;
	localparam [31:0] ibex_pkg_IC_NUM_LINES = (ibex_pkg_IC_SIZE_BYTES / ibex_pkg_IC_NUM_WAYS) / ibex_pkg_IC_LINE_BYTES;
	localparam [31:0] ibex_pkg_IC_INDEX_W = $clog2(ibex_pkg_IC_NUM_LINES);
	localparam [31:0] ibex_pkg_IC_LINE_W = 3;
	localparam [31:0] ibex_pkg_IC_TAG_SIZE = ((ibex_pkg_ADDR_W - ibex_pkg_IC_INDEX_W) - ibex_pkg_IC_LINE_W) + 1;
	localparam [31:0] TagSizeECC = (ICacheECC ? ibex_pkg_IC_TAG_SIZE + 6 : ibex_pkg_IC_TAG_SIZE);
	localparam [31:0] NumAddrScrRounds = (ICacheScramble ? 2 : 0);
	localparam [31:0] NumDiffRounds = NumAddrScrRounds;
	wire clk;
	wire [3:0] core_busy_d;
	reg [3:0] core_busy_q;
	wire clock_en;
	wire irq_pending;
	wire dummy_instr_id;
	wire dummy_instr_wb;
	wire [4:0] rf_raddr_a;
	wire [4:0] rf_raddr_b;
	wire [4:0] rf_waddr_wb;
	wire rf_we_wb;
	wire [RegFileDataWidth - 1:0] rf_wdata_wb_ecc;
	wire [RegFileDataWidth - 1:0] rf_rdata_a_ecc;
	wire [RegFileDataWidth - 1:0] rf_rdata_a_ecc_buf;
	wire [RegFileDataWidth - 1:0] rf_rdata_b_ecc;
	wire [RegFileDataWidth - 1:0] rf_rdata_b_ecc_buf;
	wire [MemDataWidth - 1:0] data_wdata_core;
	wire [MemDataWidth - 1:0] data_rdata_core;
	wire [MemDataWidth - 1:0] instr_rdata_core;
	wire [1:0] ic_tag_req;
	wire ic_tag_write;
	wire [ibex_pkg_IC_INDEX_W - 1:0] ic_tag_addr;
	wire [TagSizeECC - 1:0] ic_tag_wdata;
	wire [(ibex_pkg_IC_NUM_WAYS * TagSizeECC) - 1:0] ic_tag_rdata;
	wire [1:0] ic_data_req;
	wire ic_data_write;
	wire [ibex_pkg_IC_INDEX_W - 1:0] ic_data_addr;
	wire [LineSizeECC - 1:0] ic_data_wdata;
	wire [(ibex_pkg_IC_NUM_WAYS * LineSizeECC) - 1:0] ic_data_rdata;
	wire ic_scr_key_req;
	wire core_alert_major_internal;
	wire core_alert_major_bus;
	wire core_alert_minor;
	wire lockstep_alert_major_internal;
	wire lockstep_alert_major_bus;
	wire lockstep_alert_minor;
	reg [127:0] scramble_key_q;
	reg [63:0] scramble_nonce_q;
	wire scramble_key_valid_d;
	reg scramble_key_valid_q;
	wire scramble_req_d;
	reg scramble_req_q;
	wire [3:0] fetch_enable_buf;
	localparam [3:0] ibex_pkg_IbexMuBiOff = 4'b1010;
	generate
		if (SecureIbex) begin : g_clock_en_secure
			wire [4:1] sv2v_tmp_u_prim_core_busy_flop_q_o;
			always @(*) core_busy_q = sv2v_tmp_u_prim_core_busy_flop_q_o;
			prim_flop #(
				.Width(4),
				.ResetValue(ibex_pkg_IbexMuBiOff)
			) u_prim_core_busy_flop(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(core_busy_d),
				.q_o(sv2v_tmp_u_prim_core_busy_flop_q_o)
			);
			assign clock_en = (((core_busy_q != ibex_pkg_IbexMuBiOff) | debug_req_i) | irq_pending) | irq_nm_i;
		end
		else begin : g_clock_en_non_secure
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					core_busy_q <= ibex_pkg_IbexMuBiOff;
				else
					core_busy_q <= core_busy_d;
			assign clock_en = ((core_busy_q[0] | debug_req_i) | irq_pending) | irq_nm_i;
			wire unused_core_busy;
			assign unused_core_busy = ^core_busy_q[3:1];
		end
	endgenerate
	assign core_sleep_o = ~clock_en;
	prim_clock_gating core_clock_gate_i(
		.clk_i(clk_i),
		.en_i(clock_en),
		.test_en_i(test_en_i),
		.clk_o(clk)
	);
	prim_buf #(.Width(4)) u_fetch_enable_buf(
		.in_i(fetch_enable_i),
		.out_o(fetch_enable_buf)
	);
	prim_buf #(.Width(RegFileDataWidth)) u_rf_rdata_a_ecc_buf(
		.in_i(rf_rdata_a_ecc),
		.out_o(rf_rdata_a_ecc_buf)
	);
	prim_buf #(.Width(RegFileDataWidth)) u_rf_rdata_b_ecc_buf(
		.in_i(rf_rdata_b_ecc),
		.out_o(rf_rdata_b_ecc_buf)
	);
	assign data_rdata_core[31:0] = data_rdata_i;
	assign instr_rdata_core[31:0] = instr_rdata_i;
	generate
		if (MemECC) begin : gen_mem_rdata_ecc
			assign data_rdata_core[38:32] = data_rdata_intg_i;
			assign instr_rdata_core[38:32] = instr_rdata_intg_i;
		end
		else begin : gen_non_mem_rdata_ecc
			wire unused_intg;
			assign unused_intg = ^{instr_rdata_intg_i, data_rdata_intg_i};
		end
	endgenerate
	ibex_core #(
		.PMPEnable(PMPEnable),
		.PMPGranularity(PMPGranularity),
		.PMPNumRegions(PMPNumRegions),
		.MHPMCounterNum(MHPMCounterNum),
		.MHPMCounterWidth(MHPMCounterWidth),
		.RV32E(RV32E),
		.RV32M(RV32M),
		.RV32B(RV32B),
		.BranchTargetALU(BranchTargetALU),
		.ICache(ICache),
		.ICacheECC(ICacheECC),
		.BusSizeECC(BusSizeECC),
		.TagSizeECC(TagSizeECC),
		.LineSizeECC(LineSizeECC),
		.BranchPredictor(BranchPredictor),
		.DbgTriggerEn(DbgTriggerEn),
		.DbgHwBreakNum(DbgHwBreakNum),
		.WritebackStage(WritebackStage),
		.ResetAll(ResetAll),
		.RndCnstLfsrSeed(RndCnstLfsrSeed),
		.RndCnstLfsrPerm(RndCnstLfsrPerm),
		.SecureIbex(SecureIbex),
		.DummyInstructions(DummyInstructions),
		.RegFileECC(RegFileECC),
		.RegFileDataWidth(RegFileDataWidth),
		.MemECC(MemECC),
		.MemDataWidth(MemDataWidth),
		.DmHaltAddr(DmHaltAddr),
		.DmExceptionAddr(DmExceptionAddr)
	) u_ibex_core(
		.clk_i(clk),
		.rst_ni(rst_ni),
		.hart_id_i(hart_id_i),
		.boot_addr_i(boot_addr_i),
		.instr_req_o(instr_req_o),
		.instr_gnt_i(instr_gnt_i),
		.instr_rvalid_i(instr_rvalid_i),
		.instr_addr_o(instr_addr_o),
		.instr_rdata_i(instr_rdata_core),
		.instr_err_i(instr_err_i),
		.data_req_o(data_req_o),
		.data_gnt_i(data_gnt_i),
		.data_rvalid_i(data_rvalid_i),
		.data_we_o(data_we_o),
		.data_be_o(data_be_o),
		.data_addr_o(data_addr_o),
		.data_wdata_o(data_wdata_core),
		.data_rdata_i(data_rdata_core),
		.data_err_i(data_err_i),
		.dummy_instr_id_o(dummy_instr_id),
		.dummy_instr_wb_o(dummy_instr_wb),
		.rf_raddr_a_o(rf_raddr_a),
		.rf_raddr_b_o(rf_raddr_b),
		.rf_waddr_wb_o(rf_waddr_wb),
		.rf_we_wb_o(rf_we_wb),
		.rf_wdata_wb_ecc_o(rf_wdata_wb_ecc),
		.rf_rdata_a_ecc_i(rf_rdata_a_ecc_buf),
		.rf_rdata_b_ecc_i(rf_rdata_b_ecc_buf),
		.ic_tag_req_o(ic_tag_req),
		.ic_tag_write_o(ic_tag_write),
		.ic_tag_addr_o(ic_tag_addr),
		.ic_tag_wdata_o(ic_tag_wdata),
		.ic_tag_rdata_i(ic_tag_rdata),
		.ic_data_req_o(ic_data_req),
		.ic_data_write_o(ic_data_write),
		.ic_data_addr_o(ic_data_addr),
		.ic_data_wdata_o(ic_data_wdata),
		.ic_data_rdata_i(ic_data_rdata),
		.ic_scr_key_valid_i(scramble_key_valid_q),
		.ic_scr_key_req_o(ic_scr_key_req),
		.irq_software_i(irq_software_i),
		.irq_timer_i(irq_timer_i),
		.irq_external_i(irq_external_i),
		.irq_fast_i(irq_fast_i),
		.irq_nm_i(irq_nm_i),
		.irq_pending_o(irq_pending),
		.debug_req_i(debug_req_i),
		.crash_dump_o(crash_dump_o),
		.double_fault_seen_o(double_fault_seen_o),
		.fetch_enable_i(fetch_enable_buf),
		.alert_minor_o(core_alert_minor),
		.alert_major_internal_o(core_alert_major_internal),
		.alert_major_bus_o(core_alert_major_bus),
		.core_busy_o(core_busy_d)
	);
	wire rf_alert_major_internal;
	localparam [38:0] prim_secded_pkg_SecdedInv3932ZeroWord = 39'h2a00000000;
	function automatic [RegFileDataWidth - 1:0] sv2v_cast_E67BC;
		input reg [RegFileDataWidth - 1:0] inp;
		sv2v_cast_E67BC = inp;
	endfunction
	generate
		if (RegFile == 32'sd0) begin : gen_regfile_ff
			ibex_register_file_ff #(
				.RV32E(RV32E),
				.DataWidth(RegFileDataWidth),
				.DummyInstructions(DummyInstructions),
				.WrenCheck(RegFileWrenCheck),
				.WordZeroVal(sv2v_cast_E67BC(prim_secded_pkg_SecdedInv3932ZeroWord))
			) register_file_i(
				.clk_i(clk),
				.rst_ni(rst_ni),
				.test_en_i(test_en_i),
				.dummy_instr_id_i(dummy_instr_id),
				.dummy_instr_wb_i(dummy_instr_wb),
				.raddr_a_i(rf_raddr_a),
				.rdata_a_o(rf_rdata_a_ecc),
				.raddr_b_i(rf_raddr_b),
				.rdata_b_o(rf_rdata_b_ecc),
				.waddr_a_i(rf_waddr_wb),
				.wdata_a_i(rf_wdata_wb_ecc),
				.we_a_i(rf_we_wb),
				.err_o(rf_alert_major_internal)
			);
		end
		else if (RegFile == 32'sd1) begin : gen_regfile_fpga
			ibex_register_file_fpga #(
				.RV32E(RV32E),
				.DataWidth(RegFileDataWidth),
				.DummyInstructions(DummyInstructions),
				.WrenCheck(RegFileWrenCheck),
				.WordZeroVal(sv2v_cast_E67BC(prim_secded_pkg_SecdedInv3932ZeroWord))
			) register_file_i(
				.clk_i(clk),
				.rst_ni(rst_ni),
				.test_en_i(test_en_i),
				.dummy_instr_id_i(dummy_instr_id),
				.dummy_instr_wb_i(dummy_instr_wb),
				.raddr_a_i(rf_raddr_a),
				.rdata_a_o(rf_rdata_a_ecc),
				.raddr_b_i(rf_raddr_b),
				.rdata_b_o(rf_rdata_b_ecc),
				.waddr_a_i(rf_waddr_wb),
				.wdata_a_i(rf_wdata_wb_ecc),
				.we_a_i(rf_we_wb),
				.err_o(rf_alert_major_internal)
			);
		end
		else if (RegFile == 32'sd2) begin : gen_regfile_latch
			ibex_register_file_latch #(
				.RV32E(RV32E),
				.DataWidth(RegFileDataWidth),
				.DummyInstructions(DummyInstructions),
				.WrenCheck(RegFileWrenCheck),
				.WordZeroVal(sv2v_cast_E67BC(prim_secded_pkg_SecdedInv3932ZeroWord))
			) register_file_i(
				.clk_i(clk),
				.rst_ni(rst_ni),
				.test_en_i(test_en_i),
				.dummy_instr_id_i(dummy_instr_id),
				.dummy_instr_wb_i(dummy_instr_wb),
				.raddr_a_i(rf_raddr_a),
				.rdata_a_o(rf_rdata_a_ecc),
				.raddr_b_i(rf_raddr_b),
				.rdata_b_o(rf_rdata_b_ecc),
				.waddr_a_i(rf_waddr_wb),
				.wdata_a_i(rf_wdata_wb_ecc),
				.we_a_i(rf_we_wb),
				.err_o(rf_alert_major_internal)
			);
		end
		if (ICacheScramble) begin : gen_scramble
			assign scramble_key_valid_d = (scramble_req_q ? scramble_key_valid_i : (ic_scr_key_req ? 1'b0 : scramble_key_valid_q));
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni) begin
					scramble_key_q <= RndCnstIbexKey;
					scramble_nonce_q <= RndCnstIbexNonce;
				end
				else if (scramble_key_valid_i) begin
					scramble_key_q <= scramble_key_i;
					scramble_nonce_q <= scramble_nonce_i;
				end
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni) begin
					scramble_key_valid_q <= 1'b1;
					scramble_req_q <= 1'sb0;
				end
				else begin
					scramble_key_valid_q <= scramble_key_valid_d;
					scramble_req_q <= scramble_req_d;
				end
			assign scramble_req_d = (scramble_req_q ? ~scramble_key_valid_i : ic_scr_key_req);
			assign scramble_req_o = scramble_req_q;
		end
		else begin : gen_noscramble
			reg unused_scramble_inputs = (((((((scramble_key_valid_i & |scramble_key_i) & |RndCnstIbexKey) & |scramble_nonce_i) & |RndCnstIbexNonce) & scramble_req_q) & ic_scr_key_req) & scramble_key_valid_d) & scramble_req_d;
			assign scramble_req_d = 1'b0;
			wire [1:1] sv2v_tmp_AE3A4;
			assign sv2v_tmp_AE3A4 = 1'b0;
			always @(*) scramble_req_q = sv2v_tmp_AE3A4;
			assign scramble_req_o = 1'b0;
			wire [128:1] sv2v_tmp_A2325;
			assign sv2v_tmp_A2325 = 1'sb0;
			always @(*) scramble_key_q = sv2v_tmp_A2325;
			wire [64:1] sv2v_tmp_70913;
			assign sv2v_tmp_70913 = 1'sb0;
			always @(*) scramble_nonce_q = sv2v_tmp_70913;
			wire [1:1] sv2v_tmp_92821;
			assign sv2v_tmp_92821 = 1'b1;
			always @(*) scramble_key_valid_q = sv2v_tmp_92821;
			assign scramble_key_valid_d = 1'b1;
		end
	endgenerate
	function automatic [TagSizeECC - 1:0] sv2v_cast_CFEC9;
		input reg [TagSizeECC - 1:0] inp;
		sv2v_cast_CFEC9 = inp;
	endfunction
	function automatic [LineSizeECC - 1:0] sv2v_cast_80844;
		input reg [LineSizeECC - 1:0] inp;
		sv2v_cast_80844 = inp;
	endfunction
	generate
		if (ICache) begin : gen_rams
			genvar way;
			for (way = 0; way < ibex_pkg_IC_NUM_WAYS; way = way + 1) begin : gen_rams_inner
				if (ICacheScramble) begin : gen_scramble_rams
					prim_ram_1p_scr #(
						.Width(TagSizeECC),
						.Depth(ibex_pkg_IC_NUM_LINES),
						.DataBitsPerMask(TagSizeECC),
						.EnableParity(0),
						.DiffWidth(TagSizeECC),
						.NumAddrScrRounds(NumAddrScrRounds),
						.NumDiffRounds(NumDiffRounds)
					) tag_bank(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.key_valid_i(scramble_key_valid_q),
						.key_i(scramble_key_q),
						.nonce_i(scramble_nonce_q),
						.req_i(ic_tag_req[way]),
						.write_i(ic_tag_write),
						.addr_i(ic_tag_addr),
						.wdata_i(ic_tag_wdata),
						.wmask_i({TagSizeECC {1'b1}}),
						.intg_error_i(1'b0),
						.rdata_o(ic_tag_rdata[(1 - way) * TagSizeECC+:TagSizeECC]),
						.cfg_i(ram_cfg_i)
					);
					prim_ram_1p_scr #(
						.Width(LineSizeECC),
						.Depth(ibex_pkg_IC_NUM_LINES),
						.DataBitsPerMask(LineSizeECC),
						.ReplicateKeyStream(1),
						.EnableParity(0),
						.DiffWidth(LineSizeECC),
						.NumAddrScrRounds(NumAddrScrRounds),
						.NumDiffRounds(NumDiffRounds)
					) data_bank(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.key_valid_i(scramble_key_valid_q),
						.key_i(scramble_key_q),
						.nonce_i(scramble_nonce_q),
						.req_i(ic_data_req[way]),
						.write_i(ic_data_write),
						.addr_i(ic_data_addr),
						.wdata_i(ic_data_wdata),
						.wmask_i({LineSizeECC {1'b1}}),
						.intg_error_i(1'b0),
						.rdata_o(ic_data_rdata[(1 - way) * LineSizeECC+:LineSizeECC]),
						.cfg_i(ram_cfg_i)
					);
				end
				else begin : gen_noscramble_rams
					prim_ram_1p #(
						.Width(TagSizeECC),
						.Depth(ibex_pkg_IC_NUM_LINES),
						.DataBitsPerMask(TagSizeECC)
					) tag_bank(
						.clk_i(clk_i),
						.req_i(ic_tag_req[way]),
						.write_i(ic_tag_write),
						.addr_i(ic_tag_addr),
						.wdata_i(ic_tag_wdata),
						.wmask_i({TagSizeECC {1'b1}}),
						.rdata_o(ic_tag_rdata[(1 - way) * TagSizeECC+:TagSizeECC]),
						.cfg_i(ram_cfg_i)
					);
					prim_ram_1p #(
						.Width(LineSizeECC),
						.Depth(ibex_pkg_IC_NUM_LINES),
						.DataBitsPerMask(LineSizeECC)
					) data_bank(
						.clk_i(clk_i),
						.req_i(ic_data_req[way]),
						.write_i(ic_data_write),
						.addr_i(ic_data_addr),
						.wdata_i(ic_data_wdata),
						.wmask_i({LineSizeECC {1'b1}}),
						.rdata_o(ic_data_rdata[(1 - way) * LineSizeECC+:LineSizeECC]),
						.cfg_i(ram_cfg_i)
					);
				end
			end
		end
		else begin : gen_norams
			wire [9:0] unused_ram_cfg;
			wire unused_ram_inputs;
			assign unused_ram_cfg = ram_cfg_i;
			assign unused_ram_inputs = ((((((((((((|ic_tag_req & ic_tag_write) & |ic_tag_addr) & |ic_tag_wdata) & |ic_data_req) & ic_data_write) & |ic_data_addr) & |ic_data_wdata) & |scramble_key_q) & |scramble_nonce_q) & scramble_key_valid_q) & scramble_key_valid_d) & |scramble_nonce_q) & |NumAddrScrRounds;
			assign ic_tag_rdata = {ibex_pkg_IC_NUM_WAYS {sv2v_cast_CFEC9('b0)}};
			assign ic_data_rdata = {ibex_pkg_IC_NUM_WAYS {sv2v_cast_80844('b0)}};
		end
	endgenerate
	assign data_wdata_o = data_wdata_core[31:0];
	generate
		if (MemECC) begin : gen_mem_wdata_ecc
			prim_buf #(.Width(7)) u_prim_buf_data_wdata_intg(
				.in_i(data_wdata_core[38:32]),
				.out_o(data_wdata_intg_o)
			);
		end
		else begin : gen_no_mem_ecc
			assign data_wdata_intg_o = 1'sb0;
		end
		if (Lockstep) begin : gen_lockstep
			localparam signed [31:0] NumBufferBits = ((((((((((((((((99 + MemDataWidth) + 41) + MemDataWidth) + MemDataWidth) + 19) + RegFileDataWidth) + RegFileDataWidth) + RegFileDataWidth) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + TagSizeECC) + ibex_pkg_IC_NUM_WAYS) + 1) + ibex_pkg_IC_INDEX_W) + LineSizeECC) + 192;
			wire [NumBufferBits - 1:0] buf_in;
			wire [NumBufferBits - 1:0] buf_out;
			wire [31:0] hart_id_local;
			wire [31:0] boot_addr_local;
			wire instr_req_local;
			wire instr_gnt_local;
			wire instr_rvalid_local;
			wire [31:0] instr_addr_local;
			wire [MemDataWidth - 1:0] instr_rdata_local;
			wire instr_err_local;
			wire data_req_local;
			wire data_gnt_local;
			wire data_rvalid_local;
			wire data_we_local;
			wire [3:0] data_be_local;
			wire [31:0] data_addr_local;
			wire [MemDataWidth - 1:0] data_wdata_local;
			wire [MemDataWidth - 1:0] data_rdata_local;
			wire data_err_local;
			wire dummy_instr_id_local;
			wire dummy_instr_wb_local;
			wire [4:0] rf_raddr_a_local;
			wire [4:0] rf_raddr_b_local;
			wire [4:0] rf_waddr_wb_local;
			wire rf_we_wb_local;
			wire [RegFileDataWidth - 1:0] rf_wdata_wb_ecc_local;
			wire [RegFileDataWidth - 1:0] rf_rdata_a_ecc_local;
			wire [RegFileDataWidth - 1:0] rf_rdata_b_ecc_local;
			wire [1:0] ic_tag_req_local;
			wire ic_tag_write_local;
			wire [ibex_pkg_IC_INDEX_W - 1:0] ic_tag_addr_local;
			wire [TagSizeECC - 1:0] ic_tag_wdata_local;
			wire [1:0] ic_data_req_local;
			wire ic_data_write_local;
			wire [ibex_pkg_IC_INDEX_W - 1:0] ic_data_addr_local;
			wire [LineSizeECC - 1:0] ic_data_wdata_local;
			wire scramble_key_valid_local;
			wire ic_scr_key_req_local;
			wire irq_software_local;
			wire irq_timer_local;
			wire irq_external_local;
			wire [14:0] irq_fast_local;
			wire irq_nm_local;
			wire irq_pending_local;
			wire debug_req_local;
			wire [159:0] crash_dump_local;
			wire double_fault_seen_local;
			wire [3:0] fetch_enable_local;
			wire [3:0] core_busy_local;
			assign buf_in = {hart_id_i, boot_addr_i, instr_req_o, instr_gnt_i, instr_rvalid_i, instr_addr_o, instr_rdata_core, instr_err_i, data_req_o, data_gnt_i, data_rvalid_i, data_we_o, data_be_o, data_addr_o, data_wdata_core, data_rdata_core, data_err_i, dummy_instr_id, dummy_instr_wb, rf_raddr_a, rf_raddr_b, rf_waddr_wb, rf_we_wb, rf_wdata_wb_ecc, rf_rdata_a_ecc, rf_rdata_b_ecc, ic_tag_req, ic_tag_write, ic_tag_addr, ic_tag_wdata, ic_data_req, ic_data_write, ic_data_addr, ic_data_wdata, scramble_key_valid_q, ic_scr_key_req, irq_software_i, irq_timer_i, irq_external_i, irq_fast_i, irq_nm_i, irq_pending, debug_req_i, crash_dump_o, double_fault_seen_o, fetch_enable_i, core_busy_d};
			assign {hart_id_local, boot_addr_local, instr_req_local, instr_gnt_local, instr_rvalid_local, instr_addr_local, instr_rdata_local, instr_err_local, data_req_local, data_gnt_local, data_rvalid_local, data_we_local, data_be_local, data_addr_local, data_wdata_local, data_rdata_local, data_err_local, dummy_instr_id_local, dummy_instr_wb_local, rf_raddr_a_local, rf_raddr_b_local, rf_waddr_wb_local, rf_we_wb_local, rf_wdata_wb_ecc_local, rf_rdata_a_ecc_local, rf_rdata_b_ecc_local, ic_tag_req_local, ic_tag_write_local, ic_tag_addr_local, ic_tag_wdata_local, ic_data_req_local, ic_data_write_local, ic_data_addr_local, ic_data_wdata_local, scramble_key_valid_local, ic_scr_key_req_local, irq_software_local, irq_timer_local, irq_external_local, irq_fast_local, irq_nm_local, irq_pending_local, debug_req_local, crash_dump_local, double_fault_seen_local, fetch_enable_local, core_busy_local} = buf_out;
			prim_buf #(.Width(NumBufferBits)) u_signals_prim_buf(
				.in_i(buf_in),
				.out_o(buf_out)
			);
			wire [(ibex_pkg_IC_NUM_WAYS * TagSizeECC) - 1:0] ic_tag_rdata_local;
			wire [(ibex_pkg_IC_NUM_WAYS * LineSizeECC) - 1:0] ic_data_rdata_local;
			genvar k;
			for (k = 0; k < ibex_pkg_IC_NUM_WAYS; k = k + 1) begin : gen_ways
				prim_buf #(.Width(TagSizeECC)) u_tag_prim_buf(
					.in_i(ic_tag_rdata[(1 - k) * TagSizeECC+:TagSizeECC]),
					.out_o(ic_tag_rdata_local[(1 - k) * TagSizeECC+:TagSizeECC])
				);
				prim_buf #(.Width(LineSizeECC)) u_data_prim_buf(
					.in_i(ic_data_rdata[(1 - k) * LineSizeECC+:LineSizeECC]),
					.out_o(ic_data_rdata_local[(1 - k) * LineSizeECC+:LineSizeECC])
				);
			end
			wire lockstep_alert_minor_local;
			wire lockstep_alert_major_internal_local;
			wire lockstep_alert_major_bus_local;
			ibex_lockstep #(
				.PMPEnable(PMPEnable),
				.PMPGranularity(PMPGranularity),
				.PMPNumRegions(PMPNumRegions),
				.MHPMCounterNum(MHPMCounterNum),
				.MHPMCounterWidth(MHPMCounterWidth),
				.RV32E(RV32E),
				.RV32M(RV32M),
				.RV32B(RV32B),
				.BranchTargetALU(BranchTargetALU),
				.ICache(ICache),
				.ICacheECC(ICacheECC),
				.BusSizeECC(BusSizeECC),
				.TagSizeECC(TagSizeECC),
				.LineSizeECC(LineSizeECC),
				.BranchPredictor(BranchPredictor),
				.DbgTriggerEn(DbgTriggerEn),
				.DbgHwBreakNum(DbgHwBreakNum),
				.WritebackStage(WritebackStage),
				.ResetAll(ResetAll),
				.RndCnstLfsrSeed(RndCnstLfsrSeed),
				.RndCnstLfsrPerm(RndCnstLfsrPerm),
				.SecureIbex(SecureIbex),
				.DummyInstructions(DummyInstructions),
				.RegFileECC(RegFileECC),
				.RegFileDataWidth(RegFileDataWidth),
				.MemECC(MemECC),
				.DmHaltAddr(DmHaltAddr),
				.DmExceptionAddr(DmExceptionAddr)
			) u_ibex_lockstep(
				.clk_i(clk),
				.rst_ni(rst_ni),
				.hart_id_i(hart_id_local),
				.boot_addr_i(boot_addr_local),
				.instr_req_i(instr_req_local),
				.instr_gnt_i(instr_gnt_local),
				.instr_rvalid_i(instr_rvalid_local),
				.instr_addr_i(instr_addr_local),
				.instr_rdata_i(instr_rdata_local),
				.instr_err_i(instr_err_local),
				.data_req_i(data_req_local),
				.data_gnt_i(data_gnt_local),
				.data_rvalid_i(data_rvalid_local),
				.data_we_i(data_we_local),
				.data_be_i(data_be_local),
				.data_addr_i(data_addr_local),
				.data_wdata_i(data_wdata_local),
				.data_rdata_i(data_rdata_local),
				.data_err_i(data_err_local),
				.dummy_instr_id_i(dummy_instr_id_local),
				.dummy_instr_wb_i(dummy_instr_wb_local),
				.rf_raddr_a_i(rf_raddr_a_local),
				.rf_raddr_b_i(rf_raddr_b_local),
				.rf_waddr_wb_i(rf_waddr_wb_local),
				.rf_we_wb_i(rf_we_wb_local),
				.rf_wdata_wb_ecc_i(rf_wdata_wb_ecc_local),
				.rf_rdata_a_ecc_i(rf_rdata_a_ecc_local),
				.rf_rdata_b_ecc_i(rf_rdata_b_ecc_local),
				.ic_tag_req_i(ic_tag_req_local),
				.ic_tag_write_i(ic_tag_write_local),
				.ic_tag_addr_i(ic_tag_addr_local),
				.ic_tag_wdata_i(ic_tag_wdata_local),
				.ic_tag_rdata_i(ic_tag_rdata_local),
				.ic_data_req_i(ic_data_req_local),
				.ic_data_write_i(ic_data_write_local),
				.ic_data_addr_i(ic_data_addr_local),
				.ic_data_wdata_i(ic_data_wdata_local),
				.ic_data_rdata_i(ic_data_rdata_local),
				.ic_scr_key_valid_i(scramble_key_valid_local),
				.ic_scr_key_req_i(ic_scr_key_req_local),
				.irq_software_i(irq_software_local),
				.irq_timer_i(irq_timer_local),
				.irq_external_i(irq_external_local),
				.irq_fast_i(irq_fast_local),
				.irq_nm_i(irq_nm_local),
				.irq_pending_i(irq_pending_local),
				.debug_req_i(debug_req_local),
				.crash_dump_i(crash_dump_local),
				.double_fault_seen_i(double_fault_seen_local),
				.fetch_enable_i(fetch_enable_local),
				.alert_minor_o(lockstep_alert_minor_local),
				.alert_major_internal_o(lockstep_alert_major_internal_local),
				.alert_major_bus_o(lockstep_alert_major_bus_local),
				.core_busy_i(core_busy_local),
				.test_en_i(test_en_i),
				.scan_rst_ni(scan_rst_ni)
			);
			prim_buf u_prim_buf_alert_minor(
				.in_i(lockstep_alert_minor_local),
				.out_o(lockstep_alert_minor)
			);
			prim_buf u_prim_buf_alert_major_internal(
				.in_i(lockstep_alert_major_internal_local),
				.out_o(lockstep_alert_major_internal)
			);
			prim_buf u_prim_buf_alert_major_bus(
				.in_i(lockstep_alert_major_bus_local),
				.out_o(lockstep_alert_major_bus)
			);
		end
		else begin : gen_no_lockstep
			assign lockstep_alert_major_internal = 1'b0;
			assign lockstep_alert_major_bus = 1'b0;
			assign lockstep_alert_minor = 1'b0;
			wire unused_scan;
			assign unused_scan = scan_rst_ni;
		end
	endgenerate
	assign alert_major_internal_o = (core_alert_major_internal | lockstep_alert_major_internal) | rf_alert_major_internal;
	assign alert_major_bus_o = core_alert_major_bus | lockstep_alert_major_bus;
	assign alert_minor_o = core_alert_minor | lockstep_alert_minor;
endmodule
module ibex_wb_stage (
	clk_i,
	rst_ni,
	en_wb_i,
	instr_type_wb_i,
	pc_id_i,
	instr_is_compressed_id_i,
	instr_perf_count_id_i,
	ready_wb_o,
	rf_write_wb_o,
	outstanding_load_wb_o,
	outstanding_store_wb_o,
	pc_wb_o,
	perf_instr_ret_wb_o,
	perf_instr_ret_compressed_wb_o,
	perf_instr_ret_wb_spec_o,
	perf_instr_ret_compressed_wb_spec_o,
	rf_waddr_id_i,
	rf_wdata_id_i,
	rf_we_id_i,
	dummy_instr_id_i,
	rf_wdata_lsu_i,
	rf_we_lsu_i,
	rf_wdata_fwd_wb_o,
	rf_waddr_wb_o,
	rf_wdata_wb_o,
	rf_we_wb_o,
	dummy_instr_wb_o,
	lsu_resp_valid_i,
	lsu_resp_err_i,
	instr_done_wb_o
);
	parameter [0:0] ResetAll = 1'b0;
	parameter [0:0] WritebackStage = 1'b0;
	parameter [0:0] DummyInstructions = 1'b0;
	input wire clk_i;
	input wire rst_ni;
	input wire en_wb_i;
	input wire [1:0] instr_type_wb_i;
	input wire [31:0] pc_id_i;
	input wire instr_is_compressed_id_i;
	input wire instr_perf_count_id_i;
	output wire ready_wb_o;
	output wire rf_write_wb_o;
	output wire outstanding_load_wb_o;
	output wire outstanding_store_wb_o;
	output wire [31:0] pc_wb_o;
	output wire perf_instr_ret_wb_o;
	output wire perf_instr_ret_compressed_wb_o;
	output wire perf_instr_ret_wb_spec_o;
	output wire perf_instr_ret_compressed_wb_spec_o;
	input wire [4:0] rf_waddr_id_i;
	input wire [31:0] rf_wdata_id_i;
	input wire rf_we_id_i;
	input wire dummy_instr_id_i;
	input wire [31:0] rf_wdata_lsu_i;
	input wire rf_we_lsu_i;
	output wire [31:0] rf_wdata_fwd_wb_o;
	output wire [4:0] rf_waddr_wb_o;
	output wire [31:0] rf_wdata_wb_o;
	output wire rf_we_wb_o;
	output wire dummy_instr_wb_o;
	input wire lsu_resp_valid_i;
	input wire lsu_resp_err_i;
	output wire instr_done_wb_o;
	wire [31:0] rf_wdata_wb_mux [0:1];
	wire [1:0] rf_wdata_wb_mux_we;
	generate
		if (WritebackStage) begin : g_writeback_stage
			reg [31:0] rf_wdata_wb_q;
			reg rf_we_wb_q;
			reg [4:0] rf_waddr_wb_q;
			wire wb_done;
			reg wb_valid_q;
			reg [31:0] wb_pc_q;
			reg wb_compressed_q;
			reg wb_count_q;
			reg [1:0] wb_instr_type_q;
			wire wb_valid_d;
			assign wb_valid_d = (en_wb_i & ready_wb_o) | (wb_valid_q & ~wb_done);
			assign wb_done = (wb_instr_type_q == 2'd2) | lsu_resp_valid_i;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					wb_valid_q <= 1'b0;
				else
					wb_valid_q <= wb_valid_d;
			if (ResetAll) begin : g_wb_regs_ra
				always @(posedge clk_i or negedge rst_ni)
					if (!rst_ni) begin
						rf_we_wb_q <= 1'sb0;
						rf_waddr_wb_q <= 1'sb0;
						rf_wdata_wb_q <= 1'sb0;
						wb_instr_type_q <= 2'd0;
						wb_pc_q <= 1'sb0;
						wb_compressed_q <= 1'sb0;
						wb_count_q <= 1'sb0;
					end
					else if (en_wb_i) begin
						rf_we_wb_q <= rf_we_id_i;
						rf_waddr_wb_q <= rf_waddr_id_i;
						rf_wdata_wb_q <= rf_wdata_id_i;
						wb_instr_type_q <= instr_type_wb_i;
						wb_pc_q <= pc_id_i;
						wb_compressed_q <= instr_is_compressed_id_i;
						wb_count_q <= instr_perf_count_id_i;
					end
			end
			else begin : g_wb_regs_nr
				always @(posedge clk_i)
					if (en_wb_i) begin
						rf_we_wb_q <= rf_we_id_i;
						rf_waddr_wb_q <= rf_waddr_id_i;
						rf_wdata_wb_q <= rf_wdata_id_i;
						wb_instr_type_q <= instr_type_wb_i;
						wb_pc_q <= pc_id_i;
						wb_compressed_q <= instr_is_compressed_id_i;
						wb_count_q <= instr_perf_count_id_i;
					end
			end
			assign rf_waddr_wb_o = rf_waddr_wb_q;
			assign rf_wdata_wb_mux[0] = rf_wdata_wb_q;
			assign rf_wdata_wb_mux_we[0] = rf_we_wb_q & wb_valid_q;
			assign ready_wb_o = ~wb_valid_q | wb_done;
			assign rf_write_wb_o = wb_valid_q & (rf_we_wb_q | (wb_instr_type_q == 2'd0));
			assign outstanding_load_wb_o = wb_valid_q & (wb_instr_type_q == 2'd0);
			assign outstanding_store_wb_o = wb_valid_q & (wb_instr_type_q == 2'd1);
			assign pc_wb_o = wb_pc_q;
			assign instr_done_wb_o = wb_valid_q & wb_done;
			assign perf_instr_ret_wb_spec_o = wb_count_q;
			assign perf_instr_ret_compressed_wb_spec_o = perf_instr_ret_wb_spec_o & wb_compressed_q;
			assign perf_instr_ret_wb_o = (instr_done_wb_o & wb_count_q) & ~(lsu_resp_valid_i & lsu_resp_err_i);
			assign perf_instr_ret_compressed_wb_o = perf_instr_ret_wb_o & wb_compressed_q;
			assign rf_wdata_fwd_wb_o = rf_wdata_wb_q;
			assign rf_wdata_wb_mux_we[1] = outstanding_load_wb_o & rf_we_lsu_i;
			if (DummyInstructions) begin : g_dummy_instr_wb
				reg dummy_instr_wb_q;
				if (ResetAll) begin : g_dummy_instr_wb_regs_ra
					always @(posedge clk_i or negedge rst_ni)
						if (!rst_ni)
							dummy_instr_wb_q <= 1'b0;
						else if (en_wb_i)
							dummy_instr_wb_q <= dummy_instr_id_i;
				end
				else begin : g_dummy_instr_wb_regs_nr
					always @(posedge clk_i)
						if (en_wb_i)
							dummy_instr_wb_q <= dummy_instr_id_i;
				end
				assign dummy_instr_wb_o = dummy_instr_wb_q;
			end
			else begin : g_no_dummy_instr_wb
				wire unused_dummy_instr_id;
				assign unused_dummy_instr_id = dummy_instr_id_i;
				assign dummy_instr_wb_o = 1'b0;
			end
		end
		else begin : g_bypass_wb
			assign rf_waddr_wb_o = rf_waddr_id_i;
			assign rf_wdata_wb_mux[0] = rf_wdata_id_i;
			assign rf_wdata_wb_mux_we[0] = rf_we_id_i;
			assign rf_wdata_wb_mux_we[1] = rf_we_lsu_i;
			assign dummy_instr_wb_o = dummy_instr_id_i;
			assign perf_instr_ret_wb_spec_o = 1'b0;
			assign perf_instr_ret_compressed_wb_spec_o = 1'b0;
			assign perf_instr_ret_wb_o = (instr_perf_count_id_i & en_wb_i) & ~(lsu_resp_valid_i & lsu_resp_err_i);
			assign perf_instr_ret_compressed_wb_o = perf_instr_ret_wb_o & instr_is_compressed_id_i;
			assign ready_wb_o = 1'b1;
			wire unused_clk;
			wire unused_rst;
			wire [1:0] unused_instr_type_wb;
			wire [31:0] unused_pc_id;
			wire unused_dummy_instr_id;
			assign unused_clk = clk_i;
			assign unused_rst = rst_ni;
			assign unused_instr_type_wb = instr_type_wb_i;
			assign unused_pc_id = pc_id_i;
			assign unused_dummy_instr_id = dummy_instr_id_i;
			assign outstanding_load_wb_o = 1'b0;
			assign outstanding_store_wb_o = 1'b0;
			assign pc_wb_o = 1'sb0;
			assign rf_write_wb_o = 1'b0;
			assign rf_wdata_fwd_wb_o = 32'b00000000000000000000000000000000;
			assign instr_done_wb_o = 1'b0;
		end
	endgenerate
	assign rf_wdata_wb_mux[1] = rf_wdata_lsu_i;
	assign rf_wdata_wb_o = ({32 {rf_wdata_wb_mux_we[0]}} & rf_wdata_wb_mux[0]) | ({32 {rf_wdata_wb_mux_we[1]}} & rf_wdata_wb_mux[1]);
	assign rf_we_wb_o = |rf_wdata_wb_mux_we;
endmodule
module noerr_rv_core_ibex (
	clk_i,
	rst_ni,
	clk_edn_i,
	rst_edn_ni,
	clk_esc_i,
	rst_esc_ni,
	rst_cpu_n_o,
	ram_cfg_i,
	hart_id_i,
	boot_addr_i,
	corei_tl_h_o,
	corei_tl_h_i,
	cored_tl_h_o,
	cored_tl_h_i,
	irq_software_i,
	irq_timer_i,
	irq_external_i,
	esc_tx_i,
	esc_rx_o,
	nmi_wdog_i,
	debug_req_i,
	crash_dump_o,
	lc_cpu_en_i,
	pwrmgr_cpu_en_i,
	pwrmgr_o,
	scan_rst_ni,
	scanmode_i,
	cfg_tl_d_i,
	cfg_tl_d_o,
	edn_o,
	edn_i,
	clk_otp_i,
	rst_otp_ni,
	icache_otp_key_o,
	icache_otp_key_i,
	fpga_info_i,
	alert_rx_i,
	alert_tx_o
);
	localparam signed [31:0] rv_core_ibex_reg_pkg_NumAlerts = 4;
	parameter [3:0] AlertAsyncOn = {rv_core_ibex_reg_pkg_NumAlerts {1'b1}};
	parameter [0:0] PMPEnable = 1'b1;
	parameter [31:0] PMPGranularity = 0;
	parameter [31:0] PMPNumRegions = 16;
	parameter [31:0] MHPMCounterNum = 10;
	parameter [31:0] MHPMCounterWidth = 32;
	parameter [0:0] RV32E = 0;
	parameter integer RV32M = 32'sd3;
	parameter integer RV32B = 32'sd2;
	parameter integer RegFile = 32'sd0;
	parameter [0:0] BranchTargetALU = 1'b1;
	parameter [0:0] WritebackStage = 1'b1;
	parameter [0:0] ICache = 1'b1;
	parameter [0:0] ICacheECC = 1'b1;
	parameter [0:0] ICacheScramble = 1'b1;
	parameter [0:0] BranchPredictor = 1'b0;
	parameter [0:0] DbgTriggerEn = 1'b1;
	parameter [31:0] DbgHwBreakNum = 4;
	parameter [0:0] SecureIbex = 1'b1;
	localparam signed [31:0] ibex_pkg_LfsrWidth = 32;
	localparam [31:0] ibex_pkg_RndCnstLfsrSeedDefault = 32'hac533bf4;
	parameter [31:0] RndCnstLfsrSeed = ibex_pkg_RndCnstLfsrSeedDefault;
	localparam [159:0] ibex_pkg_RndCnstLfsrPermDefault = 160'h1e35ecba467fd1b12e958152c04fa43878a8daed;
	parameter [159:0] RndCnstLfsrPerm = ibex_pkg_RndCnstLfsrPermDefault;
	parameter [31:0] DmHaltAddr = 32'h1a110800;
	parameter [31:0] DmExceptionAddr = 32'h1a110808;
	parameter [0:0] PipeLine = 1'b0;
	localparam [31:0] ibex_pkg_SCRAMBLE_KEY_W = 128;
	localparam [127:0] ibex_pkg_RndCnstIbexKeyDefault = 128'h14e8cecae3040d5e12286bb3cc113298;
	parameter [127:0] RndCnstIbexKeyDefault = ibex_pkg_RndCnstIbexKeyDefault;
	localparam [31:0] ibex_pkg_SCRAMBLE_NONCE_W = 64;
	localparam [63:0] ibex_pkg_RndCnstIbexNonceDefault = 64'hf79780bc735f3843;
	parameter [63:0] RndCnstIbexNonceDefault = ibex_pkg_RndCnstIbexNonceDefault;
	input wire clk_i;
	input wire rst_ni;
	input wire clk_edn_i;
	input wire rst_edn_ni;
	input wire clk_esc_i;
	input wire rst_esc_ni;
	output wire rst_cpu_n_o;
	input wire [9:0] ram_cfg_i;
	input wire [31:0] hart_id_i;
	input wire [31:0] boot_addr_i;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] corei_tl_h_o;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] corei_tl_h_i;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] cored_tl_h_o;
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] cored_tl_h_i;
	input wire irq_software_i;
	input wire irq_timer_i;
	input wire irq_external_i;
	input wire [1:0] esc_tx_i;
	output wire [1:0] esc_rx_o;
	input wire nmi_wdog_i;
	input wire debug_req_i;
	output wire [224:0] crash_dump_o;
	localparam signed [31:0] lc_ctrl_pkg_TxWidth = 4;
	input wire [3:0] lc_cpu_en_i;
	input wire [3:0] pwrmgr_cpu_en_i;
	output wire [0:0] pwrmgr_o;
	input scan_rst_ni;
	input wire [3:0] scanmode_i;
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] cfg_tl_d_i;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] cfg_tl_d_o;
	output wire [0:0] edn_o;
	localparam [31:0] edn_pkg_ENDPOINT_BUS_WIDTH = 32;
	input wire [33:0] edn_i;
	input clk_otp_i;
	input rst_otp_ni;
	output wire [0:0] icache_otp_key_o;
	localparam signed [31:0] otp_ctrl_pkg_SramKeyWidth = 128;
	localparam signed [31:0] otp_ctrl_pkg_SramNonceWidth = 128;
	input wire [257:0] icache_otp_key_i;
	input [31:0] fpga_info_i;
	input wire [15:0] alert_rx_i;
	output wire [7:0] alert_tx_o;
	wire [312:0] reg2hw;
	wire [82:0] hw2reg;
	localparam [0:0] FifoPass = (PipeLine ? 1'b0 : 1'b1);
	localparam [31:0] FifoDepth = (PipeLine ? 2 : 0);
	localparam signed [31:0] NumOutstandingReqs = (ICache ? 8 : 2);
	wire instr_req;
	wire instr_gnt;
	wire instr_rvalid;
	wire [31:0] instr_addr;
	wire [31:0] instr_rdata;
	wire [6:0] instr_rdata_intg;
	wire instr_err;
	wire data_req;
	wire data_gnt;
	wire data_rvalid;
	wire data_we;
	wire [3:0] data_be;
	wire [31:0] data_addr;
	wire [31:0] data_wdata;
	wire [6:0] data_wdata_intg;
	wire [31:0] data_rdata;
	wire [6:0] data_rdata_intg;
	wire data_err;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_i_ibex2fifo;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_i_fifo2ibex;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_d_ibex2fifo;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_d_fifo2ibex;
	wire core_sleep;
	wire ibex_top_clk_i;
	wire addr_trans_rst_ni;
	assign ibex_top_clk_i = clk_i;
	assign addr_trans_rst_ni = rst_ni;
	wire ibus_intg_err;
	wire dbus_intg_err;
	wire alert_minor;
	wire alert_major_internal;
	wire alert_major_bus;
	wire double_fault;
	wire fatal_intg_err;
	wire fatal_core_err;
	wire recov_core_err;
	wire fatal_intg_event;
	wire fatal_core_event;
	wire recov_core_event;
	assign fatal_intg_event = (ibus_intg_err | dbus_intg_err) | alert_major_bus;
	assign fatal_core_event = alert_major_internal | double_fault;
	assign recov_core_event = alert_minor;
	localparam signed [31:0] rv_core_ibex_reg_pkg_NumRegions = 2;
	wire [129:0] ibus_region_cfg;
	wire [129:0] dbus_region_cfg;
	assign rst_cpu_n_o = rst_ni;
	wire esc_irq_nm;
	localparam signed [31:0] alert_handler_reg_pkg_N_ESC_SEV = 4;
	localparam signed [31:0] alert_handler_reg_pkg_PING_CNT_DW = 16;
	prim_esc_receiver #(
		.N_ESC_SEV(alert_handler_reg_pkg_N_ESC_SEV),
		.PING_CNT_DW(alert_handler_reg_pkg_PING_CNT_DW)
	) u_prim_esc_receiver(
		.clk_i(clk_esc_i),
		.rst_ni(rst_esc_ni),
		.esc_req_o(esc_irq_nm),
		.esc_rx_o(esc_rx_o),
		.esc_tx_i(esc_tx_i)
	);
	wire alert_irq_nm;
	prim_flop_2sync #(.Width(1)) u_alert_nmi_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(esc_irq_nm),
		.q_o(alert_irq_nm)
	);
	wire wdog_irq_nm;
	prim_flop_2sync #(.Width(1)) u_wdog_nmi_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(nmi_wdog_i),
		.q_o(wdog_irq_nm)
	);
	assign hw2reg[77] = 1'b1;
	assign hw2reg[76] = alert_irq_nm;
	assign hw2reg[75] = 1'b1;
	assign hw2reg[74] = wdog_irq_nm;
	wire irq_nm;
	assign irq_nm = |(reg2hw[34-:2] & reg2hw[36-:2]);
	wire [3:0] lc_cpu_en;
	prim_lc_sync u_lc_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.lc_en_i(lc_cpu_en_i),
		.lc_en_o(lc_cpu_en)
	);
	wire [3:0] pwrmgr_cpu_en;
	prim_lc_sync u_pwrmgr_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.lc_en_i(pwrmgr_cpu_en_i),
		.lc_en_o(pwrmgr_cpu_en)
	);
	wire irq_timer_sync;
	prim_flop_2sync #(.Width(1)) u_intr_timer_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(irq_timer_i),
		.q_o(irq_timer_sync)
	);
	wire irq_software;
	wire irq_timer;
	wire irq_external;
	prim_sec_anchor_buf #(.Width(3)) u_prim_buf_irq(
		.in_i({irq_software_i, irq_timer_sync, irq_external_i}),
		.out_o({irq_software, irq_timer, irq_external})
	);
	wire key_req;
	wire key_ack;
	wire [127:0] key;
	wire [63:0] nonce;
	wire unused_seed_valid;
	localparam signed [31:0] PayLoadW = (ibex_pkg_SCRAMBLE_KEY_W + ibex_pkg_SCRAMBLE_NONCE_W) + 1;
	prim_sync_reqack_data #(
		.Width(PayLoadW),
		.DataSrc2Dst(1'b0)
	) u_prim_sync_reqack_data(
		.clk_src_i(clk_i),
		.rst_src_ni(rst_ni),
		.clk_dst_i(clk_otp_i),
		.rst_dst_ni(rst_otp_ni),
		.req_chk_i(1'b1),
		.src_req_i(key_req),
		.src_ack_o(key_ack),
		.dst_req_o(icache_otp_key_o[0]),
		.dst_ack_i(icache_otp_key_i[257]),
		.data_i({icache_otp_key_i[256-:128], icache_otp_key_i[64:1], icache_otp_key_i[0]}),
		.data_o({key, nonce, unused_seed_valid})
	);
	wire unused_nonce;
	assign unused_nonce = |icache_otp_key_i[128-:128];
	wire [3:0] local_fetch_enable_d;
	wire [3:0] local_fetch_enable_q;
	function automatic [3:0] sv2v_cast_A1913;
		input reg [3:0] inp;
		sv2v_cast_A1913 = inp;
	endfunction
	assign local_fetch_enable_d = (fatal_core_err ? sv2v_cast_A1913(4'b1010) : local_fetch_enable_q);
	prim_lc_sender #(
		.AsyncOn(1),
		.ResetValueIsOn(1)
	) u_prim_lc_sender(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.lc_en_i(local_fetch_enable_d),
		.lc_en_o(local_fetch_enable_q)
	);
	wire [3:0] fetch_enable;
	function automatic [3:0] lc_ctrl_pkg_lc_tx_and;
		input reg [3:0] a;
		input reg [3:0] b;
		input reg [3:0] act;
		reg [3:0] a_in;
		reg [3:0] b_in;
		reg [3:0] act_in;
		reg [3:0] out;
		begin
			a_in = a;
			b_in = b;
			act_in = act;
			begin : sv2v_autoblock_1
				reg signed [31:0] k;
				for (k = 0; k < lc_ctrl_pkg_TxWidth; k = k + 1)
					if (act_in[k])
						out[k] = a_in[k] && b_in[k];
					else
						out[k] = a_in[k] || b_in[k];
			end
			lc_ctrl_pkg_lc_tx_and = out;
		end
	endfunction
	function automatic [3:0] lc_ctrl_pkg_lc_tx_and_hi;
		input reg [3:0] a;
		input reg [3:0] b;
		lc_ctrl_pkg_lc_tx_and_hi = lc_ctrl_pkg_lc_tx_and(a, b, sv2v_cast_A1913(4'b0101));
	endfunction
	assign fetch_enable = lc_ctrl_pkg_lc_tx_and_hi(local_fetch_enable_q, lc_ctrl_pkg_lc_tx_and_hi(lc_cpu_en[0+:lc_ctrl_pkg_TxWidth], pwrmgr_cpu_en[0+:lc_ctrl_pkg_TxWidth]));
	wire [159:0] crash_dump;
	function automatic [3:0] sv2v_cast_38B98;
		input reg [3:0] inp;
		sv2v_cast_38B98 = inp;
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_true_strict;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_true_strict = sv2v_cast_38B98(4'h6) == val;
	endfunction
	ibex_top #(
		.PMPEnable(PMPEnable),
		.PMPGranularity(PMPGranularity),
		.PMPNumRegions(PMPNumRegions),
		.MHPMCounterNum(MHPMCounterNum),
		.MHPMCounterWidth(MHPMCounterWidth),
		.RV32E(RV32E),
		.RV32M(RV32M),
		.RV32B(RV32B),
		.RegFile(RegFile),
		.BranchTargetALU(BranchTargetALU),
		.WritebackStage(WritebackStage),
		.ICache(ICache),
		.ICacheECC(ICacheECC),
		.ICacheScramble(ICacheScramble),
		.BranchPredictor(BranchPredictor),
		.DbgTriggerEn(DbgTriggerEn),
		.DbgHwBreakNum(DbgHwBreakNum),
		.SecureIbex(SecureIbex),
		.RndCnstLfsrSeed(RndCnstLfsrSeed),
		.RndCnstLfsrPerm(RndCnstLfsrPerm),
		.RndCnstIbexKey(RndCnstIbexKeyDefault),
		.RndCnstIbexNonce(RndCnstIbexNonceDefault),
		.DmHaltAddr(DmHaltAddr),
		.DmExceptionAddr(DmExceptionAddr)
	) u_core(
		.clk_i(ibex_top_clk_i),
		.rst_ni(rst_ni),
		.test_en_i(prim_mubi_pkg_mubi4_test_true_strict(scanmode_i)),
		.scan_rst_ni(scan_rst_ni),
		.ram_cfg_i(ram_cfg_i),
		.hart_id_i(hart_id_i),
		.boot_addr_i(boot_addr_i),
		.instr_req_o(instr_req),
		.instr_gnt_i(instr_gnt),
		.instr_rvalid_i(instr_rvalid),
		.instr_addr_o(instr_addr),
		.instr_rdata_i(instr_rdata),
		.instr_rdata_intg_i(instr_rdata_intg),
		.instr_err_i(instr_err),
		.data_req_o(data_req),
		.data_gnt_i(data_gnt),
		.data_rvalid_i(data_rvalid),
		.data_we_o(data_we),
		.data_be_o(data_be),
		.data_addr_o(data_addr),
		.data_wdata_o(data_wdata),
		.data_wdata_intg_o(data_wdata_intg),
		.data_rdata_i(data_rdata),
		.data_rdata_intg_i(data_rdata_intg),
		.data_err_i(data_err),
		.irq_software_i(irq_software),
		.irq_timer_i(irq_timer),
		.irq_external_i(irq_external),
		.irq_fast_i(1'sb0),
		.irq_nm_i(irq_nm),
		.debug_req_i(debug_req_i),
		.crash_dump_o(crash_dump),
		.scramble_key_valid_i(key_ack),
		.scramble_key_i(key),
		.scramble_nonce_i(nonce),
		.scramble_req_o(key_req),
		.double_fault_seen_o(double_fault),
		.fetch_enable_i(fetch_enable),
		.alert_minor_o(alert_minor),
		.alert_major_internal_o(alert_major_internal),
		.alert_major_bus_o(alert_major_bus),
		.core_sleep_o(core_sleep)
	);
	reg core_sleep_q;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			core_sleep_q <= 1'sb0;
		else
			core_sleep_q <= core_sleep;
	prim_buf #(.Width(1)) u_core_sleeping_buf(
		.in_i(core_sleep_q),
		.out_o(pwrmgr_o[0])
	);
	reg prev_valid;
	reg [31:0] prev_exception_pc;
	reg [31:0] prev_exception_addr;
	assign crash_dump_o[159-:160] = crash_dump;
	assign crash_dump_o[224] = prev_valid;
	assign crash_dump_o[223-:32] = prev_exception_pc;
	assign crash_dump_o[191-:32] = prev_exception_addr;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			prev_valid <= 1'sb0;
			prev_exception_pc <= 1'sb0;
			prev_exception_addr <= 1'sb0;
		end
		else if (double_fault) begin
			prev_valid <= 1'b1;
			prev_exception_pc <= crash_dump[63-:32];
			prev_exception_addr <= crash_dump[31-:32];
		end
	wire [31:0] instr_addr_trans;
	rv_core_addr_trans #(
		.AddrWidth(32),
		.NumRegions(rv_core_ibex_reg_pkg_NumRegions)
	) u_ibus_trans(
		.clk_i(clk_i),
		.rst_ni(addr_trans_rst_ni),
		.region_cfg_i(ibus_region_cfg),
		.addr_i(instr_addr),
		.addr_o(instr_addr_trans)
	);
	assign instr_err = 0;
	wire [6:0] instr_wdata_intg;
	wire [31:0] unused_data;
	function automatic [38:0] sv2v_cast_39;
		input reg [38:0] inp;
		sv2v_cast_39 = inp;
	endfunction
	function automatic [38:0] prim_secded_pkg_prim_secded_inv_39_32_enc;
		input reg [31:0] data_i;
		reg [38:0] data_o;
		begin
			data_o = sv2v_cast_39(data_i);
			data_o[32] = ^(data_o & 39'h002606bd25);
			data_o[33] = ^(data_o & 39'h00deba8050);
			data_o[34] = ^(data_o & 39'h00413d89aa);
			data_o[35] = ^(data_o & 39'h0031234ed1);
			data_o[36] = ^(data_o & 39'h00c2c1323b);
			data_o[37] = ^(data_o & 39'h002dcc624c);
			data_o[38] = ^(data_o & 39'h0098505586);
			data_o = data_o ^ 39'h2a00000000;
			prim_secded_pkg_prim_secded_inv_39_32_enc = data_o;
		end
	endfunction
	assign {instr_wdata_intg, unused_data} = prim_secded_pkg_prim_secded_inv_39_32_enc(instr_rdata);
	tlul_adapter_host #(
		.MAX_REQS(NumOutstandingReqs),
		.EnableDataIntgGen(~SecureIbex)
	) tl_adapter_host_i_ibex(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.req_i(instr_req),
		.instr_type_i(sv2v_cast_38B98(4'h6)),
		.gnt_o(instr_gnt),
		.addr_i(instr_addr_trans),
		.we_i(1'b0),
		.wdata_i(32'b00000000000000000000000000000000),
		.wdata_intg_i(instr_wdata_intg),
		.be_i(4'hf),
		.valid_o(instr_rvalid),
		.rdata_o(instr_rdata),
		.rdata_intg_o(instr_rdata_intg),
		.intg_err_o(ibus_intg_err),
		.tl_o(tl_i_ibex2fifo),
		.tl_i(tl_i_fifo2ibex)
	);
	tlul_fifo_sync #(
		.ReqPass(FifoPass),
		.RspPass(FifoPass),
		.ReqDepth(FifoDepth),
		.RspDepth(FifoDepth)
	) fifo_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_h_i(tl_i_ibex2fifo),
		.tl_h_o(tl_i_fifo2ibex),
		.tl_d_o(corei_tl_h_o),
		.tl_d_i(corei_tl_h_i),
		.spare_req_i(1'b0),
		.spare_rsp_i(1'b0)
	);
	wire [31:0] data_addr_trans;
	rv_core_addr_trans #(
		.AddrWidth(32),
		.NumRegions(rv_core_ibex_reg_pkg_NumRegions)
	) u_dbus_trans(
		.clk_i(clk_i),
		.rst_ni(addr_trans_rst_ni),
		.region_cfg_i(dbus_region_cfg),
		.addr_i(data_addr),
		.addr_o(data_addr_trans)
	);
	assign data_err = 0;
	tlul_adapter_host #(
		.MAX_REQS(2),
		.EnableDataIntgGen(~SecureIbex)
	) tl_adapter_host_d_ibex(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.req_i(data_req),
		.instr_type_i(sv2v_cast_38B98(4'h9)),
		.gnt_o(data_gnt),
		.addr_i(data_addr_trans),
		.we_i(data_we),
		.wdata_i(data_wdata),
		.wdata_intg_i(data_wdata_intg),
		.be_i(data_be),
		.valid_o(data_rvalid),
		.rdata_o(data_rdata),
		.rdata_intg_o(data_rdata_intg),
		.intg_err_o(dbus_intg_err),
		.tl_o(tl_d_ibex2fifo),
		.tl_i(tl_d_fifo2ibex)
	);
	tlul_fifo_sync #(
		.ReqPass(FifoPass),
		.RspPass(FifoPass),
		.ReqDepth(FifoDepth),
		.RspDepth(FifoDepth)
	) fifo_d(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_h_i(tl_d_ibex2fifo),
		.tl_h_o(tl_d_fifo2ibex),
		.tl_d_o(cored_tl_h_o),
		.tl_d_i(cored_tl_h_i),
		.spare_req_i(1'b0),
		.spare_rsp_i(1'b0)
	);
	wire intg_err;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_win_h2d;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_win_d2h;
	rv_core_ibex_cfg_reg_top u_reg_cfg(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(cfg_tl_d_i),
		.tl_o(cfg_tl_d_o),
		.reg2hw(reg2hw),
		.hw2reg(hw2reg),
		.intg_err_o(intg_err),
		.tl_win_o(tl_win_h2d),
		.tl_win_i(tl_win_d2h),
		.devmode_i(1'b1)
	);
	genvar i;
	generate
		for (i = 0; i < rv_core_ibex_reg_pkg_NumRegions; i = i + 1) begin : gen_ibus_region_cfgs
			assign ibus_region_cfg[(i * 65) + 64] = reg2hw[295 + i+:1];
			assign ibus_region_cfg[(i * 65) + 63-:32] = reg2hw[231 + (i * 32)+:32];
			assign ibus_region_cfg[(i * 65) + 31-:32] = reg2hw[167 + (i * 32)+:32];
		end
		for (i = 0; i < rv_core_ibex_reg_pkg_NumRegions; i = i + 1) begin : gen_dbus_region_cfgs
			assign dbus_region_cfg[(i * 65) + 64] = reg2hw[165 + i+:1];
			assign dbus_region_cfg[(i * 65) + 63-:32] = reg2hw[101 + (i * 32)+:32];
			assign dbus_region_cfg[(i * 65) + 31-:32] = reg2hw[37 + (i * 32)+:32];
		end
	endgenerate
	assign fatal_intg_err = fatal_intg_event;
	assign fatal_core_err = fatal_core_event;
	assign recov_core_err = recov_core_event;
	assign hw2reg[73] = 1'b1;
	assign hw2reg[72] = intg_err;
	assign hw2reg[71] = 1'b1;
	assign hw2reg[70] = fatal_intg_err;
	assign hw2reg[69] = 1'b1;
	assign hw2reg[68] = fatal_core_err;
	assign hw2reg[67] = 1'b1;
	assign hw2reg[66] = recov_core_err;
	wire [3:0] alert_test;
	assign alert_test[0] = reg2hw[312] & reg2hw[311];
	assign alert_test[1] = reg2hw[310] & reg2hw[309];
	assign alert_test[2] = reg2hw[308] & reg2hw[307];
	assign alert_test[3] = reg2hw[306] & reg2hw[305];
	localparam [3:0] AlertFatal = 4'b0101;
	wire [3:0] alert_events;
	wire [3:0] alert_acks;
	function automatic prim_mubi_pkg_mubi4_test_true_loose;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_true_loose = sv2v_cast_38B98(4'h9) != val;
	endfunction
	assign alert_events[0] = prim_mubi_pkg_mubi4_test_true_loose(sv2v_cast_38B98(reg2hw[300-:4]));
	assign alert_events[1] = prim_mubi_pkg_mubi4_test_true_loose(sv2v_cast_38B98(reg2hw[304-:4]));
	assign alert_events[2] = (intg_err | fatal_intg_err) | fatal_core_err;
	assign alert_events[3] = recov_core_err;
	wire unused_alert_acks;
	assign unused_alert_acks = |alert_acks;
	assign hw2reg[78] = alert_acks[1];
	assign hw2reg[82-:4] = sv2v_cast_38B98(4'h9);
	generate
		for (i = 0; i < rv_core_ibex_reg_pkg_NumAlerts; i = i + 1) begin : gen_alert_senders
			prim_alert_sender #(
				.AsyncOn(AlertAsyncOn[0]),
				.IsFatal(AlertFatal[i])
			) u_alert_sender(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.alert_test_i(alert_test[i]),
				.alert_req_i(alert_events[i]),
				.alert_ack_o(alert_acks[i]),
				.alert_rx_i(alert_rx_i[i * 4+:4]),
				.alert_tx_o(alert_tx_o[i * 2+:2])
			);
		end
	endgenerate
	reg [31:0] rnd_data_q;
	reg [31:0] rnd_data_d;
	reg rnd_valid_q;
	reg rnd_valid_d;
	reg rnd_fips_q;
	reg rnd_fips_d;
	wire edn_req;
	wire [31:0] edn_data;
	wire edn_ack;
	wire edn_fips;
	always @(*) begin
		rnd_valid_d = rnd_valid_q;
		rnd_data_d = rnd_data_q;
		rnd_fips_d = rnd_fips_q;
		if (reg2hw[0]) begin
			rnd_valid_d = 1'sb0;
			rnd_data_d = 1'sb0;
			rnd_fips_d = 1'sb0;
		end
		else if (edn_req && edn_ack) begin
			rnd_valid_d = 1'b1;
			rnd_data_d = edn_data;
			rnd_fips_d = edn_fips;
		end
	end
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			rnd_valid_q <= 1'sb0;
			rnd_data_q <= 1'sb0;
			rnd_fips_q <= 1'sb0;
		end
		else begin
			rnd_valid_q <= rnd_valid_d;
			rnd_data_q <= rnd_data_d;
			rnd_fips_q <= rnd_fips_d;
		end
	assign edn_req = ~rnd_valid_q;
	prim_edn_req #(.OutWidth(32)) u_edn_if(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.req_chk_i(1'b1),
		.req_i(edn_req),
		.ack_o(edn_ack),
		.data_o(edn_data),
		.fips_o(edn_fips),
		.clk_edn_i(clk_edn_i),
		.rst_edn_ni(rst_edn_ni),
		.edn_o(edn_o),
		.edn_i(edn_i)
	);
	assign hw2reg[65-:32] = rnd_data_q;
	assign hw2reg[33] = rnd_valid_q;
	assign hw2reg[32] = rnd_fips_q;
	wire unused_reg2hw;
	assign unused_reg2hw = |reg2hw[32-:32];
	assign hw2reg[31-:32] = fpga_info_i;
	localparam signed [31:0] TlH2DWidth = 1 * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24);
	localparam signed [31:0] TlD2HWidth = 1 * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2);
	wire [TlH2DWidth - 1:0] tl_win_h2d_int;
	wire [TlD2HWidth - 1:0] tl_win_d2h_int;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_win_d2h_err_rsp;
	prim_buf #(.Width(TlH2DWidth)) u_tlul_req_buf(
		.in_i(tl_win_h2d),
		.out_o(tl_win_h2d_int)
	);
	prim_buf #(.Width(TlD2HWidth)) u_tlul_rsp_buf(
		.in_i(tl_win_d2h_err_rsp),
		.out_o(tl_win_d2h_int)
	);
	function automatic [((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1)) - 1:0] sv2v_cast_51793;
		input reg [((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1)) - 1:0] inp;
		sv2v_cast_51793 = inp;
	endfunction
	assign tl_win_d2h = sv2v_cast_51793(tl_win_d2h_int);
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_win_h2d_int_tmp;
	function automatic [(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23)) - 1:0] sv2v_cast_E9713;
		input reg [(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23)) - 1:0] inp;
		sv2v_cast_E9713 = inp;
	endfunction
	assign tl_win_h2d_int_tmp = sv2v_cast_E9713(tl_win_h2d_int);
	tlul_err_resp u_sim_win_rsp(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_h_i(tl_win_h2d_int_tmp),
		.tl_h_o(tl_win_d2h_err_rsp)
	);
endmodule
module noerr_tlul_adapter_sram (
	clk_i,
	rst_ni,
	tl_i,
	tl_o,
	en_ifetch_i,
	req_o,
	req_type_o,
	gnt_i,
	we_o,
	addr_o,
	wdata_o,
	wmask_o,
	intg_error_o,
	rdata_i,
	rvalid_i,
	rerror_i
);
	parameter signed [31:0] SramAw = 12;
	parameter signed [31:0] SramDw = 32;
	parameter signed [31:0] Outstanding = 1;
	parameter [0:0] ByteAccess = 1;
	parameter [0:0] ErrOnWrite = 0;
	parameter [0:0] ErrOnRead = 0;
	parameter [0:0] CmdIntgCheck = 0;
	parameter [0:0] EnableRspIntgGen = 0;
	parameter [0:0] EnableDataIntgGen = 0;
	parameter [0:0] EnableDataIntgPt = 0;
	parameter [0:0] SecFifoPtr = 0;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] WidthMult = SramDw / top_pkg_TL_DW;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] IntgWidth = tlul_pkg_DataIntgWidth * WidthMult;
	localparam signed [31:0] DataOutW = (EnableDataIntgPt ? SramDw + IntgWidth : SramDw);
	input clk_i;
	input rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_i;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	input wire [3:0] en_ifetch_i;
	output wire req_o;
	output wire [3:0] req_type_o;
	input gnt_i;
	output wire we_o;
	output wire [SramAw - 1:0] addr_o;
	output wire [DataOutW - 1:0] wdata_o;
	output wire [DataOutW - 1:0] wmask_o;
	output wire intg_error_o;
	input [DataOutW - 1:0] rdata_i;
	input rvalid_i;
	input [1:0] rerror_i;
	localparam signed [31:0] SramByte = SramDw / 8;
	function automatic integer prim_util_pkg_vbits;
		input integer value;
		prim_util_pkg_vbits = (value == 1 ? 1 : $clog2(value));
	endfunction
	localparam signed [31:0] DataBitWidth = prim_util_pkg_vbits(SramByte);
	localparam signed [31:0] WoffsetWidth = (SramByte == top_pkg_TL_DBW ? 1 : DataBitWidth - prim_util_pkg_vbits(top_pkg_TL_DBW));
	wire error_det;
	wire error_internal;
	wire wr_attr_error;
	wire instr_error;
	wire wr_vld_error;
	wire rd_vld_error;
	wire rsp_fifo_error;
	wire intg_error;
	wire tlul_error;
	generate
		if (CmdIntgCheck) begin : gen_cmd_intg_check
			tlul_cmd_intg_chk u_cmd_intg_chk(
				.tl_i(tl_i),
				.err_o(intg_error)
			);
		end
		else begin : gen_no_cmd_intg_check
			assign intg_error = 1'sb0;
		end
	endgenerate
	reg intg_error_q;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			intg_error_q <= 1'sb0;
		else if (intg_error || rsp_fifo_error)
			intg_error_q <= 1'b1;
	assign intg_error_o = (intg_error | rsp_fifo_error) | intg_error_q;
	assign wr_attr_error = ((tl_i[6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) - (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))))) + 1 : ((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) - (6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))))) + 1)] == 3'h0) || (tl_i[6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) - (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))))) + 1 : ((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) - (6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))))) + 1)] == 3'h1) ? (ByteAccess == 0 ? (tl_i[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))] != {((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55)) * 1 {1'sb1}}) || (tl_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)] != 2'h2) : 1'b0) : 1'b0);
	function automatic [3:0] sv2v_cast_A2CB9;
		input reg [3:0] inp;
		sv2v_cast_A2CB9 = inp;
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_false_loose;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_false_loose = sv2v_cast_A2CB9(4'h6) != val;
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_invalid;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_invalid = ~(|{((sv2v_cast_A2CB9(4'h6) ^ (val ^ val)) === (val ^ (sv2v_cast_A2CB9(4'h6) ^ sv2v_cast_A2CB9(4'h6)))) & ((((val ^ val) ^ (sv2v_cast_A2CB9(4'h6) ^ sv2v_cast_A2CB9(4'h6))) === (sv2v_cast_A2CB9(4'h6) ^ sv2v_cast_A2CB9(4'h6))) | 1'bx), ((sv2v_cast_A2CB9(4'h9) ^ (val ^ val)) === (val ^ (sv2v_cast_A2CB9(4'h9) ^ sv2v_cast_A2CB9(4'h9)))) & ((((val ^ val) ^ (sv2v_cast_A2CB9(4'h9) ^ sv2v_cast_A2CB9(4'h9))) === (sv2v_cast_A2CB9(4'h9) ^ sv2v_cast_A2CB9(4'h9))) | 1'bx)});
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_true_strict;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_true_strict = sv2v_cast_A2CB9(4'h6) == val;
	endfunction
	assign instr_error = prim_mubi_pkg_mubi4_test_invalid(tl_i[18-:4]) | (prim_mubi_pkg_mubi4_test_true_strict(tl_i[18-:4]) & prim_mubi_pkg_mubi4_test_false_loose(en_ifetch_i));
	generate
		if (ErrOnWrite == 1) begin : gen_no_writes
			assign wr_vld_error = tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] != 3'h4;
		end
		else begin : gen_writes_allowed
			assign wr_vld_error = 1'b0;
		end
		if (ErrOnRead == 1) begin : gen_no_reads
			assign rd_vld_error = tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h4;
		end
		else begin : gen_reads_allowed
			assign rd_vld_error = 1'b0;
		end
	endgenerate
	tlul_err u_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_i),
		.err_o(tlul_error)
	);
	assign error_det = ((((wr_attr_error | wr_vld_error) | rd_vld_error) | instr_error) | tlul_error) | intg_error;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_i_int;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o_int;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_out;
	wire unused_tl_i_int;
	assign unused_tl_i_int = ^tl_i_int;
	tlul_rsp_intg_gen #(
		.EnableRspIntgGen(EnableRspIntgGen),
		.EnableDataIntgGen(EnableDataIntgGen)
	) u_rsp_gen(
		.tl_i(tl_out),
		.tl_o(tl_o)
	);
	assign error_internal = 0;
	tlul_sram_byte #(
		.EnableIntg((ByteAccess & EnableDataIntgPt) & !ErrOnWrite),
		.Outstanding(Outstanding)
	) u_sram_byte(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_i),
		.tl_o(tl_out),
		.tl_sram_o(tl_i_int),
		.tl_sram_i(tl_o_int),
		.error_i(error_det)
	);
	localparam signed [31:0] SramReqFifoWidth = top_pkg_TL_DBW + WoffsetWidth;
	localparam signed [31:0] ReqFifoWidth = (7 + top_pkg_TL_SZW) + top_pkg_TL_AIW;
	localparam signed [31:0] RspFifoWidth = (((top_pkg_TL_DW + tlul_pkg_DataIntgWidth) + 0) >= 0 ? (top_pkg_TL_DW + tlul_pkg_DataIntgWidth) + 1 : 1 - ((top_pkg_TL_DW + tlul_pkg_DataIntgWidth) + 0));
	wire reqfifo_wvalid;
	wire reqfifo_wready;
	wire reqfifo_rvalid;
	wire reqfifo_rready;
	wire [((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) - 1:0] reqfifo_wdata;
	wire [((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) - 1:0] reqfifo_rdata;
	wire sramreqfifo_wvalid;
	wire sramreqfifo_wready;
	wire sramreqfifo_rready;
	wire [(top_pkg_TL_DBW + WoffsetWidth) - 1:0] sramreqfifo_wdata;
	wire [(top_pkg_TL_DBW + WoffsetWidth) - 1:0] sramreqfifo_rdata;
	wire rspfifo_wvalid;
	wire rspfifo_wready;
	wire rspfifo_rvalid;
	wire rspfifo_rready;
	wire [(top_pkg_TL_DW + tlul_pkg_DataIntgWidth) + 0:0] rspfifo_wdata;
	wire [(top_pkg_TL_DW + tlul_pkg_DataIntgWidth) + 0:0] rspfifo_rdata;
	wire a_ack;
	wire d_ack;
	wire sram_ack;
	assign a_ack = tl_i_int[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & tl_o_int[0];
	assign d_ack = tl_o_int[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] & tl_i_int[0];
	assign sram_ack = req_o & gnt_i;
	reg d_valid;
	reg d_error;
	always @(*) begin
		d_valid = 1'b0;
		if (reqfifo_rvalid) begin
			if (reqfifo_rdata[1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))])
				d_valid = 1'b1;
			else if (reqfifo_rdata[3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))-:((7 + (top_pkg_TL_SZW + 7)) >= (5 + (top_pkg_TL_SZW + 8)) ? ((3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))) - (1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 8)))) + 1 : ((1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 8))) - (3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)))) + 1)] == 2'd1)
				d_valid = rspfifo_rvalid;
			else
				d_valid = 1'b1;
		end
		else
			d_valid = 1'b0;
	end
	always @(*) begin
		d_error = 1'b0;
		if (reqfifo_rvalid) begin
			if (reqfifo_rdata[3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))-:((7 + (top_pkg_TL_SZW + 7)) >= (5 + (top_pkg_TL_SZW + 8)) ? ((3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))) - (1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 8)))) + 1 : ((1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 8))) - (3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)))) + 1)] == 2'd1)
				d_error = rspfifo_rdata[0] | reqfifo_rdata[1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))];
			else
				d_error = reqfifo_rdata[1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))];
		end
		else
			d_error = 1'b0;
	end
	wire vld_rd_rsp;
	assign vld_rd_rsp = ((d_valid & reqfifo_rvalid) & rspfifo_rvalid) & (reqfifo_rdata[3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))-:((7 + (top_pkg_TL_SZW + 7)) >= (5 + (top_pkg_TL_SZW + 8)) ? ((3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))) - (1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 8)))) + 1 : ((1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 8))) - (3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)))) + 1)] == 2'd1);
	wire [31:0] error_blanking_data;
	localparam [31:0] tlul_pkg_DataWhenError = {top_pkg_TL_DW {1'b1}};
	localparam [31:0] tlul_pkg_DataWhenInstrError = 1'sb0;
	assign error_blanking_data = (prim_mubi_pkg_mubi4_test_true_strict(reqfifo_rdata[prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)-:((prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)) >= (top_pkg_TL_SZW + 8) ? ((prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)) - (top_pkg_TL_SZW + 8)) + 1 : ((top_pkg_TL_SZW + 8) - (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))) + 1)]) ? tlul_pkg_DataWhenInstrError : tlul_pkg_DataWhenError);
	wire [31:0] unused_instr;
	wire [31:0] unused_data;
	wire [6:0] error_instr_integ;
	wire [6:0] error_data_integ;
	localparam signed [31:0] tlul_pkg_DataMaxWidth = 32;
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	tlul_data_integ_enc u_tlul_data_integ_enc_instr(
		.data_i(sv2v_cast_32(tlul_pkg_DataWhenInstrError)),
		.data_intg_o({error_instr_integ, unused_instr})
	);
	tlul_data_integ_enc u_tlul_data_integ_enc_data(
		.data_i(sv2v_cast_32(tlul_pkg_DataWhenError)),
		.data_intg_o({error_data_integ, unused_data})
	);
	wire [6:0] error_blanking_integ;
	assign error_blanking_integ = (prim_mubi_pkg_mubi4_test_true_strict(reqfifo_rdata[prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)-:((prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)) >= (top_pkg_TL_SZW + 8) ? ((prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)) - (top_pkg_TL_SZW + 8)) + 1 : ((top_pkg_TL_SZW + 8) - (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))) + 1)]) ? error_instr_integ : error_data_integ);
	wire [31:0] d_data;
	assign d_data = (vld_rd_rsp & ~d_error ? rspfifo_rdata[39-:32] : error_blanking_data);
	wire [6:0] data_intg;
	localparam [6:0] prim_secded_pkg_SecdedInv3932ZeroEcc = 7'h2a;
	assign data_intg = (vld_rd_rsp && reqfifo_rdata[5 + (top_pkg_TL_SZW + 7)] ? error_blanking_integ : (vld_rd_rsp ? rspfifo_rdata[7-:7] : prim_secded_pkg_SecdedInv3932ZeroEcc));
	function automatic [6:0] sv2v_cast_5F39A;
		input reg [6:0] inp;
		sv2v_cast_5F39A = inp;
	endfunction
	function automatic [top_pkg_TL_SZW - 1:0] sv2v_cast_4660A;
		input reg [top_pkg_TL_SZW - 1:0] inp;
		sv2v_cast_4660A = inp;
	endfunction
	function automatic [7:0] sv2v_cast_964CB;
		input reg [7:0] inp;
		sv2v_cast_964CB = inp;
	endfunction
	function automatic [0:0] sv2v_cast_702AC;
		input reg [0:0] inp;
		sv2v_cast_702AC = inp;
	endfunction
	function automatic [31:0] sv2v_cast_35AE2;
		input reg [31:0] inp;
		sv2v_cast_35AE2 = inp;
	endfunction
	function automatic [(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 1:0] sv2v_cast_1D31F;
		input reg [(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 1:0] inp;
		sv2v_cast_1D31F = inp;
	endfunction
	assign tl_o_int = {d_valid, (d_valid && (reqfifo_rdata[7 + (top_pkg_TL_SZW + 7)-:((7 + (top_pkg_TL_SZW + 7)) >= (5 + (top_pkg_TL_SZW + 8)) ? ((7 + (top_pkg_TL_SZW + 7)) - (5 + (top_pkg_TL_SZW + 8))) + 1 : ((5 + (top_pkg_TL_SZW + 8)) - (7 + (top_pkg_TL_SZW + 7))) + 1)] != 2'd1) ? 3'h0 : 3'h1), 3'b000, sv2v_cast_4660A((d_valid ? reqfifo_rdata[top_pkg_TL_SZW + 7-:((top_pkg_TL_SZW + 7) >= 8 ? top_pkg_TL_SZW : 9 - (top_pkg_TL_SZW + 7))] : {((top_pkg_TL_SZW + 7) >= 8 ? top_pkg_TL_SZW : 9 - (top_pkg_TL_SZW + 7)) * 1 {1'sb0}})), sv2v_cast_964CB((d_valid ? reqfifo_rdata[7-:top_pkg_TL_AIW] : {8 {1'sb0}})), sv2v_cast_702AC(1'b0), sv2v_cast_35AE2(d_data), sv2v_cast_1D31F({sv2v_cast_5F39A(1'sb0), data_intg}), d_valid && d_error, ((gnt_i | error_internal) & reqfifo_wready) & sramreqfifo_wready};
	assign req_o = (tl_i_int[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & reqfifo_wready) & ~error_internal;
	assign req_type_o = tl_i_int[18-:4];
	assign we_o = tl_i_int[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & |{tl_i_int[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h0, tl_i_int[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h1};
	assign addr_o = (tl_i_int[7 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))] ? tl_i_int[(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (31 - DataBitWidth)+:SramAw] : {SramAw {1'sb0}});
	wire [WoffsetWidth - 1:0] woffset;
	generate
		if (top_pkg_TL_DW != SramDw) begin : gen_wordwidthadapt
			assign woffset = tl_i_int[(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (32 - DataBitWidth):(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (31 - prim_util_pkg_vbits(top_pkg_TL_DBW))];
		end
		else begin : gen_no_wordwidthadapt
			assign woffset = 1'sb0;
		end
	endgenerate
	localparam signed [31:0] DataWidth = (EnableDataIntgPt ? top_pkg_TL_DW + tlul_pkg_DataIntgWidth : top_pkg_TL_DW);
	wire [(WidthMult * DataWidth) - 1:0] wmask_combined;
	wire [(WidthMult * DataWidth) - 1:0] wdata_combined;
	reg [(WidthMult * top_pkg_TL_DW) - 1:0] wmask_int;
	reg [(WidthMult * top_pkg_TL_DW) - 1:0] wdata_int;
	reg [(WidthMult * tlul_pkg_DataIntgWidth) - 1:0] wmask_intg;
	reg [(WidthMult * tlul_pkg_DataIntgWidth) - 1:0] wdata_intg;
	always @(*) begin
		wmask_int = 1'sb0;
		wdata_int = 1'sb0;
		if (tl_i_int[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))]) begin : sv2v_autoblock_1
			reg signed [31:0] i;
			for (i = 0; i < 4; i = i + 1)
				begin
					wmask_int[(woffset * top_pkg_TL_DW) + (8 * i)+:8] = {8 {tl_i_int[(top_pkg_TL_DBW + 55) - ((top_pkg_TL_DBW - 1) - i)]}};
					wdata_int[(woffset * top_pkg_TL_DW) + (8 * i)+:8] = (tl_i_int[(top_pkg_TL_DBW + 55) - ((top_pkg_TL_DBW - 1) - i)] && we_o ? tl_i_int[24 + (8 * i)+:8] : {8 {1'sb0}});
				end
		end
	end
	always @(*) begin
		wmask_intg = 1'sb0;
		wdata_intg = 1'sb0;
		if (tl_i_int[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))]) begin
			wmask_intg[woffset * tlul_pkg_DataIntgWidth+:tlul_pkg_DataIntgWidth] = {tlul_pkg_DataIntgWidth {1'b1}};
			wdata_intg[woffset * tlul_pkg_DataIntgWidth+:tlul_pkg_DataIntgWidth] = tl_i_int[7-:tlul_pkg_DataIntgWidth];
		end
	end
	genvar i;
	generate
		for (i = 0; i < WidthMult; i = i + 1) begin : gen_write_output
			if (EnableDataIntgPt) begin : gen_combined_output
				assign wmask_combined[i * DataWidth+:DataWidth] = {wmask_intg[i * tlul_pkg_DataIntgWidth+:tlul_pkg_DataIntgWidth], wmask_int[i * top_pkg_TL_DW+:top_pkg_TL_DW]};
				assign wdata_combined[i * DataWidth+:DataWidth] = {wdata_intg[i * tlul_pkg_DataIntgWidth+:tlul_pkg_DataIntgWidth], wdata_int[i * top_pkg_TL_DW+:top_pkg_TL_DW]};
			end
			else begin : gen_ft_output
				wire unused_w;
				assign wmask_combined[i * DataWidth+:DataWidth] = wmask_int[i * top_pkg_TL_DW+:top_pkg_TL_DW];
				assign wdata_combined[i * DataWidth+:DataWidth] = wdata_int[i * top_pkg_TL_DW+:top_pkg_TL_DW];
				assign unused_w = |wmask_intg & |wdata_intg;
			end
		end
	endgenerate
	assign wmask_o = wmask_combined;
	assign wdata_o = wdata_combined;
	assign reqfifo_wvalid = a_ack;
	assign reqfifo_wdata = {(tl_i_int[6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) - (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))))) + 1 : ((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) - (6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))))) + 1)] != 3'h4 ? 2'd0 : 2'd1), error_internal, sv2v_cast_A2CB9(tl_i_int[18-:4]), tl_i_int[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)], tl_i_int[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) >= (32'sd32 + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 56)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1)]};
	assign reqfifo_rready = d_ack;
	assign sramreqfifo_wdata = {tl_i_int[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))], woffset};
	assign sramreqfifo_wvalid = sram_ack & ~we_o;
	assign sramreqfifo_rready = rspfifo_wvalid;
	assign rspfifo_wvalid = rvalid_i & reqfifo_rvalid;
	wire [(WidthMult * DataWidth) - 1:0] rdata_reshaped;
	reg [DataWidth - 1:0] rdata_tlword;
	assign rdata_reshaped = rdata_i;
	localparam [38:0] prim_secded_pkg_SecdedInv3932ZeroWord = 39'h2a00000000;
	generate
		if (EnableDataIntgPt) begin : gen_no_rmask
			always @(*) begin
				rdata_tlword = prim_secded_pkg_SecdedInv3932ZeroWord;
				if (|sramreqfifo_rdata[top_pkg_TL_DBW + (WoffsetWidth - 1)-:((top_pkg_TL_DBW + (WoffsetWidth - 1)) >= (WoffsetWidth + 0) ? ((top_pkg_TL_DBW + (WoffsetWidth - 1)) - (WoffsetWidth + 0)) + 1 : ((WoffsetWidth + 0) - (top_pkg_TL_DBW + (WoffsetWidth - 1))) + 1)])
					rdata_tlword = rdata_reshaped[sramreqfifo_rdata[WoffsetWidth - 1-:WoffsetWidth] * DataWidth+:DataWidth];
			end
		end
		else begin : gen_rmask
			reg [DataWidth - 1:0] rmask;
			always @(*) begin
				rmask = 1'sb0;
				begin : sv2v_autoblock_2
					reg signed [31:0] i;
					for (i = 0; i < 4; i = i + 1)
						rmask[8 * i+:8] = {8 {sramreqfifo_rdata[(top_pkg_TL_DBW + (WoffsetWidth - 1)) - ((top_pkg_TL_DBW - 1) - i)]}};
				end
			end
			wire [DataWidth:1] sv2v_tmp_037A0;
			assign sv2v_tmp_037A0 = rdata_reshaped[sramreqfifo_rdata[WoffsetWidth - 1-:WoffsetWidth] * DataWidth+:DataWidth] & rmask;
			always @(*) rdata_tlword = sv2v_tmp_037A0;
		end
	endgenerate
	function automatic [6:0] sv2v_cast_8DC45;
		input reg [6:0] inp;
		sv2v_cast_8DC45 = inp;
	endfunction
	assign rspfifo_wdata = {sv2v_cast_35AE2(rdata_tlword[31:0]), sv2v_cast_8DC45((EnableDataIntgPt ? rdata_tlword[DataWidth - 1-:tlul_pkg_DataIntgWidth] : {7 {1'sb0}})), rerror_i[1]};
	assign rspfifo_rready = ((reqfifo_rdata[7 + (top_pkg_TL_SZW + 7)-:((7 + (top_pkg_TL_SZW + 7)) >= (5 + (top_pkg_TL_SZW + 8)) ? ((7 + (top_pkg_TL_SZW + 7)) - (5 + (top_pkg_TL_SZW + 8))) + 1 : ((5 + (top_pkg_TL_SZW + 8)) - (7 + (top_pkg_TL_SZW + 7))) + 1)] == 2'd1) & ~reqfifo_rdata[5 + (top_pkg_TL_SZW + 7)] ? reqfifo_rready : 1'b0);
	wire unused_rerror;
	assign unused_rerror = rerror_i[0];
	prim_fifo_sync #(
		.Width(ReqFifoWidth),
		.Pass(1'b0),
		.Depth(Outstanding)
	) u_reqfifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(1'b0),
		.wvalid_i(reqfifo_wvalid),
		.wready_o(reqfifo_wready),
		.wdata_i(reqfifo_wdata),
		.rvalid_o(reqfifo_rvalid),
		.rready_i(reqfifo_rready),
		.rdata_o(reqfifo_rdata)
	);
	prim_fifo_sync #(
		.Width(SramReqFifoWidth),
		.Pass(1'b0),
		.Depth(Outstanding)
	) u_sramreqfifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(1'b0),
		.wvalid_i(sramreqfifo_wvalid),
		.wready_o(sramreqfifo_wready),
		.wdata_i(sramreqfifo_wdata),
		.rready_i(sramreqfifo_rready),
		.rdata_o(sramreqfifo_rdata)
	);
	prim_fifo_sync #(
		.Width(RspFifoWidth),
		.Pass(1'b1),
		.Depth(Outstanding),
		.Secure(SecFifoPtr)
	) u_rspfifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(1'b0),
		.wvalid_i(rspfifo_wvalid),
		.wready_o(rspfifo_wready),
		.wdata_i(rspfifo_wdata),
		.rvalid_o(rspfifo_rvalid),
		.rready_i(rspfifo_rready),
		.rdata_o(rspfifo_rdata),
		.err_o(rsp_fifo_error)
	);
endmodule
module prim_alert_receiver (
	clk_i,
	rst_ni,
	init_trig_i,
	ping_req_i,
	ping_ok_o,
	integ_fail_o,
	alert_o,
	alert_rx_o,
	alert_tx_i
);
	parameter [0:0] AsyncOn = 1'b0;
	input clk_i;
	input rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	input wire [3:0] init_trig_i;
	input ping_req_i;
	output reg ping_ok_o;
	output reg integ_fail_o;
	output reg alert_o;
	output wire [3:0] alert_rx_o;
	input wire [1:0] alert_tx_i;
	wire alert_level;
	wire alert_sigint;
	wire alert_p;
	wire alert_n;
	prim_sec_anchor_buf #(.Width(2)) u_prim_buf_in(
		.in_i({alert_tx_i[0], alert_tx_i[1]}),
		.out_o({alert_n, alert_p})
	);
	prim_diff_decode #(.AsyncOn(AsyncOn)) u_decode_alert(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.diff_pi(alert_p),
		.diff_ni(alert_n),
		.level_o(alert_level),
		.sigint_o(alert_sigint)
	);
	reg [2:0] state_d;
	reg [2:0] state_q;
	wire ping_rise;
	wire ping_tog_pd;
	wire ping_tog_pq;
	wire ping_tog_dn;
	wire ping_tog_nq;
	reg ack_pd;
	wire ack_pq;
	wire ack_dn;
	wire ack_nq;
	wire ping_req_d;
	reg ping_req_q;
	wire ping_pending_d;
	reg ping_pending_q;
	reg send_init;
	reg send_ping;
	assign ping_req_d = ping_req_i;
	assign ping_rise = ping_req_d && !ping_req_q;
	assign ping_tog_pd = (send_init ? 1'b0 : (send_ping ? ~ping_tog_pq : ping_tog_pq));
	assign ack_dn = (send_init ? ack_pd : ~ack_pd);
	assign ping_tog_dn = ~ping_tog_pd;
	prim_sec_anchor_flop #(
		.Width(2),
		.ResetValue(2'b10)
	) u_prim_generic_flop_ack(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i({ack_dn, ack_pd}),
		.q_o({ack_nq, ack_pq})
	);
	prim_sec_anchor_flop #(
		.Width(2),
		.ResetValue(2'b10)
	) u_prim_generic_flop_ping(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i({ping_tog_dn, ping_tog_pd}),
		.q_o({ping_tog_nq, ping_tog_pq})
	);
	assign ping_pending_d = ping_rise | ((~ping_ok_o & ping_req_i) & ping_pending_q);
	assign alert_rx_o[1] = ack_pq;
	assign alert_rx_o[0] = ack_nq;
	assign alert_rx_o[3] = ping_tog_pq;
	assign alert_rx_o[2] = ping_tog_nq;
	function automatic [3:0] sv2v_cast_25BC0;
		input reg [3:0] inp;
		sv2v_cast_25BC0 = inp;
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_true_strict;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_true_strict = sv2v_cast_25BC0(4'h6) == val;
	endfunction
	always @(*) begin : p_fsm
		state_d = state_q;
		ack_pd = 1'b0;
		ping_ok_o = 1'b0;
		integ_fail_o = 1'b0;
		alert_o = 1'b0;
		send_init = 1'b0;
		send_ping = ping_rise;
		case (state_q)
			3'd0:
				if (alert_level) begin
					state_d = 3'd1;
					ack_pd = 1'b1;
					if (ping_pending_q)
						ping_ok_o = 1'b1;
					else
						alert_o = 1'b1;
				end
			3'd1:
				if (!alert_level)
					state_d = 3'd2;
				else
					ack_pd = 1'b1;
			3'd2: state_d = 3'd3;
			3'd3: state_d = 3'd0;
			3'd4: begin
				send_init = 1'b1;
				send_ping = 1'b0;
				if (prim_mubi_pkg_mubi4_test_true_strict(init_trig_i))
					ping_ok_o = ping_pending_q;
				else if (alert_sigint)
					state_d = 3'd5;
			end
			3'd5: begin
				send_ping = 1'b0;
				if (!alert_sigint) begin
					state_d = 3'd2;
					send_ping = ping_rise || ping_pending_q;
				end
			end
			default: state_d = 3'd0;
		endcase
		if (!(|{state_q == 3'd4, state_q == 3'd5}))
			if (prim_mubi_pkg_mubi4_test_true_strict(init_trig_i)) begin
				state_d = 3'd4;
				ack_pd = 1'b0;
				ping_ok_o = 1'b0;
				integ_fail_o = 1'b0;
				alert_o = 1'b0;
				send_init = 1'b1;
			end
			else if (alert_sigint) begin
				state_d = 3'd0;
				ack_pd = 1'b0;
				ping_ok_o = 1'b0;
				integ_fail_o = 1'b1;
				alert_o = 1'b0;
			end
	end
	always @(posedge clk_i or negedge rst_ni) begin : p_reg
		if (!rst_ni) begin
			state_q <= 3'd4;
			ping_req_q <= 1'b0;
			ping_pending_q <= 1'b0;
		end
		else begin
			state_q <= state_d;
			ping_req_q <= ping_req_d;
			ping_pending_q <= ping_pending_d;
		end
	end
endmodule
module prim_alert_sender (
	clk_i,
	rst_ni,
	alert_test_i,
	alert_req_i,
	alert_ack_o,
	alert_state_o,
	alert_rx_i,
	alert_tx_o
);
	parameter [0:0] AsyncOn = 1'b1;
	parameter [0:0] IsFatal = 1'b0;
	input clk_i;
	input rst_ni;
	input alert_test_i;
	input alert_req_i;
	output wire alert_ack_o;
	output wire alert_state_o;
	input wire [3:0] alert_rx_i;
	output wire [1:0] alert_tx_o;
	wire ping_sigint;
	wire ping_event;
	wire ping_n;
	wire ping_p;
	prim_sec_anchor_buf #(.Width(2)) u_prim_buf_ping(
		.in_i({alert_rx_i[2], alert_rx_i[3]}),
		.out_o({ping_n, ping_p})
	);
	prim_diff_decode #(.AsyncOn(AsyncOn)) u_decode_ping(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.diff_pi(ping_p),
		.diff_ni(ping_n),
		.event_o(ping_event),
		.sigint_o(ping_sigint)
	);
	wire ack_sigint;
	wire ack_level;
	wire ack_n;
	wire ack_p;
	prim_sec_anchor_buf #(.Width(2)) u_prim_buf_ack(
		.in_i({alert_rx_i[0], alert_rx_i[1]}),
		.out_o({ack_n, ack_p})
	);
	prim_diff_decode #(.AsyncOn(AsyncOn)) u_decode_ack(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.diff_pi(ack_p),
		.diff_ni(ack_n),
		.level_o(ack_level),
		.sigint_o(ack_sigint)
	);
	reg [2:0] state_d;
	reg [2:0] state_q;
	wire alert_pq;
	wire alert_nq;
	reg alert_pd;
	reg alert_nd;
	wire sigint_detected;
	assign sigint_detected = ack_sigint | ping_sigint;
	assign alert_tx_o[1] = alert_pq;
	assign alert_tx_o[0] = alert_nq;
	wire alert_set_d;
	reg alert_set_q;
	reg alert_clr;
	wire alert_test_set_d;
	reg alert_test_set_q;
	wire ping_set_d;
	reg ping_set_q;
	reg ping_clr;
	wire alert_req_trigger;
	wire alert_test_trigger;
	wire ping_trigger;
	wire alert_req;
	prim_sec_anchor_buf #(.Width(1)) u_prim_buf_in_req(
		.in_i(alert_req_i),
		.out_o(alert_req)
	);
	assign alert_req_trigger = alert_req | alert_set_q;
	generate
		if (IsFatal) begin : gen_fatal
			assign alert_set_d = alert_req_trigger;
		end
		else begin : gen_recov
			assign alert_set_d = (alert_clr ? 1'b0 : alert_req_trigger);
		end
	endgenerate
	assign alert_test_trigger = alert_test_i | alert_test_set_q;
	assign alert_test_set_d = (alert_clr ? 1'b0 : alert_test_trigger);
	wire alert_trigger;
	assign alert_trigger = alert_req_trigger | alert_test_trigger;
	assign ping_trigger = ping_set_q | ping_event;
	assign ping_set_d = (ping_clr ? 1'b0 : ping_trigger);
	assign alert_ack_o = alert_clr & alert_set_q;
	assign alert_state_o = alert_set_q;
	always @(*) begin : p_fsm
		state_d = state_q;
		alert_pd = 1'b0;
		alert_nd = 1'b1;
		ping_clr = 1'b0;
		alert_clr = 1'b0;
		case (state_q)
			3'd0:
				if (alert_trigger || ping_trigger) begin
					state_d = (alert_trigger ? 3'd1 : 3'd3);
					alert_pd = 1'b1;
					alert_nd = 1'b0;
				end
			3'd1:
				if (ack_level)
					state_d = 3'd2;
				else begin
					alert_pd = 1'b1;
					alert_nd = 1'b0;
				end
			3'd2:
				if (!ack_level) begin
					state_d = 3'd5;
					alert_clr = 1'b1;
				end
			3'd3:
				if (ack_level)
					state_d = 3'd4;
				else begin
					alert_pd = 1'b1;
					alert_nd = 1'b0;
				end
			3'd4:
				if (!ack_level) begin
					ping_clr = 1'b1;
					state_d = 3'd5;
				end
			3'd5: state_d = 3'd6;
			3'd6: state_d = 3'd0;
			default: state_d = 3'd0;
		endcase
		if (sigint_detected) begin
			state_d = 3'd0;
			alert_pd = 1'b0;
			alert_nd = 1'b0;
			ping_clr = 1'b1;
			alert_clr = 1'b0;
		end
	end
	prim_sec_anchor_flop #(
		.Width(2),
		.ResetValue(2'b10)
	) u_prim_flop_alert(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i({alert_nd, alert_pd}),
		.q_o({alert_nq, alert_pq})
	);
	always @(posedge clk_i or negedge rst_ni) begin : p_reg
		if (!rst_ni) begin
			state_q <= 3'd0;
			alert_set_q <= 1'b0;
			alert_test_set_q <= 1'b0;
			ping_set_q <= 1'b0;
		end
		else begin
			state_q <= state_d;
			alert_set_q <= alert_set_d;
			alert_test_set_q <= alert_test_set_d;
			ping_set_q <= ping_set_d;
		end
	end
endmodule
module prim_and2 (
	in0_i,
	in1_i,
	out_o
);
	parameter signed [31:0] Width = 1;
	input [Width - 1:0] in0_i;
	input [Width - 1:0] in1_i;
	output wire [Width - 1:0] out_o;
	parameter integer Impl = 32'sd0;
	generate
		if (Impl == 32'sd2) begin : gen_xilinx
			prim_xilinx_and2 #(.Width(Width)) u_impl_xilinx(
				.in0_i(in0_i),
				.in1_i(in1_i),
				.out_o(out_o)
			);
		end
		else begin : gen_generic
			prim_generic_and2 #(.Width(Width)) u_impl_generic(
				.in0_i(in0_i),
				.in1_i(in1_i),
				.out_o(out_o)
			);
		end
	endgenerate
endmodule
module prim_arbiter_fixed (
	clk_i,
	rst_ni,
	req_i,
	data_i,
	gnt_o,
	idx_o,
	valid_o,
	data_o,
	ready_i
);
	parameter signed [31:0] N = 8;
	parameter signed [31:0] DW = 32;
	parameter [0:0] EnDataPort = 1;
	localparam signed [31:0] IdxW = $clog2(N);
	input clk_i;
	input rst_ni;
	input [N - 1:0] req_i;
	input [(N * DW) - 1:0] data_i;
	output wire [N - 1:0] gnt_o;
	output wire [IdxW - 1:0] idx_o;
	output wire valid_o;
	output wire [DW - 1:0] data_o;
	input ready_i;
	generate
		if (N == 1) begin : gen_degenerate_case
			assign valid_o = req_i[0];
			assign data_o = data_i[(N - 1) * DW+:DW];
			assign gnt_o[0] = valid_o & ready_i;
			assign idx_o = 1'sb0;
		end
		else begin : gen_normal_case
			reg [(2 ** (IdxW + 1)) - 2:0] req_tree;
			reg [(2 ** (IdxW + 1)) - 2:0] gnt_tree;
			reg [(((2 ** (IdxW + 1)) - 2) >= 0 ? (((2 ** (IdxW + 1)) - 1) * IdxW) - 1 : ((3 - (2 ** (IdxW + 1))) * IdxW) + ((((2 ** (IdxW + 1)) - 2) * IdxW) - 1)):(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : ((2 ** (IdxW + 1)) - 2) * IdxW)] idx_tree;
			reg [(((2 ** (IdxW + 1)) - 2) >= 0 ? (((2 ** (IdxW + 1)) - 1) * DW) - 1 : ((3 - (2 ** (IdxW + 1))) * DW) + ((((2 ** (IdxW + 1)) - 2) * DW) - 1)):(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : ((2 ** (IdxW + 1)) - 2) * DW)] data_tree;
			genvar level;
			for (level = 0; level < (IdxW + 1); level = level + 1) begin : gen_tree
				localparam signed [31:0] Base0 = (2 ** level) - 1;
				localparam signed [31:0] Base1 = (2 ** (level + 1)) - 1;
				genvar offset;
				for (offset = 0; offset < (2 ** level); offset = offset + 1) begin : gen_level
					localparam signed [31:0] Pa = Base0 + offset;
					localparam signed [31:0] C0 = Base1 + (2 * offset);
					localparam signed [31:0] C1 = (Base1 + (2 * offset)) + 1;
					if (level == IdxW) begin : gen_leafs
						if (offset < N) begin : gen_assign
							wire [1:1] sv2v_tmp_40210;
							assign sv2v_tmp_40210 = req_i[offset];
							always @(*) req_tree[Pa] = sv2v_tmp_40210;
							wire [IdxW * 1:1] sv2v_tmp_7E44F;
							assign sv2v_tmp_7E44F = offset;
							always @(*) idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * IdxW+:IdxW] = sv2v_tmp_7E44F;
							wire [DW * 1:1] sv2v_tmp_59E9C;
							assign sv2v_tmp_59E9C = data_i[((N - 1) - offset) * DW+:DW];
							always @(*) data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * DW+:DW] = sv2v_tmp_59E9C;
							assign gnt_o[offset] = gnt_tree[Pa];
						end
						else begin : gen_tie_off
							wire [1:1] sv2v_tmp_93CDE;
							assign sv2v_tmp_93CDE = 1'sb0;
							always @(*) req_tree[Pa] = sv2v_tmp_93CDE;
							wire [IdxW * 1:1] sv2v_tmp_0AB12;
							assign sv2v_tmp_0AB12 = 1'sb0;
							always @(*) idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * IdxW+:IdxW] = sv2v_tmp_0AB12;
							wire [DW * 1:1] sv2v_tmp_2EDCA;
							assign sv2v_tmp_2EDCA = 1'sb0;
							always @(*) data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * DW+:DW] = sv2v_tmp_2EDCA;
							wire unused_sigs;
							assign unused_sigs = gnt_tree[Pa];
						end
					end
					else begin : gen_nodes
						reg sel;
						always @(*) begin : p_node
							sel = ~req_tree[C0];
							req_tree[Pa] = req_tree[C0] | req_tree[C1];
							idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * IdxW+:IdxW] = (sel ? idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? C1 : ((2 ** (IdxW + 1)) - 2) - C1) * IdxW+:IdxW] : idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? C0 : ((2 ** (IdxW + 1)) - 2) - C0) * IdxW+:IdxW]);
							data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * DW+:DW] = (sel ? data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? C1 : ((2 ** (IdxW + 1)) - 2) - C1) * DW+:DW] : data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? C0 : ((2 ** (IdxW + 1)) - 2) - C0) * DW+:DW]);
							gnt_tree[C0] = gnt_tree[Pa] & ~sel;
							gnt_tree[C1] = gnt_tree[Pa] & sel;
						end
					end
				end
			end
			if (EnDataPort) begin : gen_data_port
				assign data_o = data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : (2 ** (IdxW + 1)) - 2) * DW+:DW];
			end
			else begin : gen_no_dataport
				wire [DW - 1:0] unused_data;
				assign unused_data = data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : (2 ** (IdxW + 1)) - 2) * DW+:DW];
				assign data_o = 1'sb1;
			end
			assign idx_o = idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : (2 ** (IdxW + 1)) - 2) * IdxW+:IdxW];
			assign valid_o = req_tree[0];
			wire [1:1] sv2v_tmp_C3EB5;
			assign sv2v_tmp_C3EB5 = valid_o & ready_i;
			always @(*) gnt_tree[0] = sv2v_tmp_C3EB5;
		end
	endgenerate
endmodule
module prim_arbiter_ppc (
	clk_i,
	rst_ni,
	req_chk_i,
	req_i,
	data_i,
	gnt_o,
	idx_o,
	valid_o,
	data_o,
	ready_i
);
	parameter [31:0] N = 8;
	parameter [31:0] DW = 32;
	parameter [0:0] EnDataPort = 1;
	localparam signed [31:0] IdxW = $clog2(N);
	input clk_i;
	input rst_ni;
	input req_chk_i;
	input [N - 1:0] req_i;
	input [(N * DW) - 1:0] data_i;
	output wire [N - 1:0] gnt_o;
	output reg [IdxW - 1:0] idx_o;
	output wire valid_o;
	output reg [DW - 1:0] data_o;
	input ready_i;
	wire unused_req_chk;
	assign unused_req_chk = req_chk_i;
	generate
		if (N == 1) begin : gen_degenerate_case
			assign valid_o = req_i[0];
			wire [DW:1] sv2v_tmp_B7B25;
			assign sv2v_tmp_B7B25 = data_i[(N - 1) * DW+:DW];
			always @(*) data_o = sv2v_tmp_B7B25;
			assign gnt_o[0] = valid_o & ready_i;
			wire [IdxW:1] sv2v_tmp_78DD8;
			assign sv2v_tmp_78DD8 = 1'sb0;
			always @(*) idx_o = sv2v_tmp_78DD8;
		end
		else begin : gen_normal_case
			wire [N - 1:0] masked_req;
			reg [N - 1:0] ppc_out;
			wire [N - 1:0] arb_req;
			reg [N - 1:0] mask;
			wire [N - 1:0] mask_next;
			wire [N - 1:0] winner;
			assign masked_req = mask & req_i;
			assign arb_req = (|masked_req ? masked_req : req_i);
			always @(*) begin
				ppc_out[0] = arb_req[0];
				begin : sv2v_autoblock_1
					reg signed [31:0] i;
					for (i = 1; i < N; i = i + 1)
						ppc_out[i] = ppc_out[i - 1] | arb_req[i];
				end
			end
			assign winner = ppc_out ^ {ppc_out[N - 2:0], 1'b0};
			assign gnt_o = (ready_i ? winner : {N {1'sb0}});
			assign valid_o = |req_i;
			assign mask_next = {ppc_out[N - 2:0], 1'b0};
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mask <= 1'sb0;
				else if (valid_o && ready_i)
					mask <= mask_next;
				else if (valid_o && !ready_i)
					mask <= ppc_out;
			if (EnDataPort == 1) begin : gen_datapath
				always @(*) begin
					data_o = 1'sb0;
					begin : sv2v_autoblock_2
						reg signed [31:0] i;
						for (i = 0; i < N; i = i + 1)
							if (winner[i])
								data_o = data_i[((N - 1) - i) * DW+:DW];
					end
				end
			end
			else begin : gen_nodatapath
				wire [DW:1] sv2v_tmp_3BABB;
				assign sv2v_tmp_3BABB = 1'sb1;
				always @(*) data_o = sv2v_tmp_3BABB;
				wire [(N * DW) - 1:0] unused_data;
				assign unused_data = data_i;
			end
			always @(*) begin
				idx_o = 1'sb0;
				begin : sv2v_autoblock_3
					reg [31:0] i;
					for (i = 0; i < N; i = i + 1)
						if (winner[i])
							idx_o = i[IdxW - 1:0];
				end
			end
		end
	endgenerate
endmodule
module prim_arbiter_tree (
	clk_i,
	rst_ni,
	req_chk_i,
	req_i,
	data_i,
	gnt_o,
	idx_o,
	valid_o,
	data_o,
	ready_i
);
	parameter signed [31:0] N = 8;
	parameter signed [31:0] DW = 32;
	parameter [0:0] EnDataPort = 1;
	localparam signed [31:0] IdxW = $clog2(N);
	input clk_i;
	input rst_ni;
	input req_chk_i;
	input [N - 1:0] req_i;
	input [(N * DW) - 1:0] data_i;
	output wire [N - 1:0] gnt_o;
	output wire [IdxW - 1:0] idx_o;
	output wire valid_o;
	output wire [DW - 1:0] data_o;
	input ready_i;
	wire unused_req_chk;
	assign unused_req_chk = req_chk_i;
	generate
		if (N == 1) begin : gen_degenerate_case
			assign valid_o = req_i[0];
			assign data_o = data_i[(N - 1) * DW+:DW];
			assign gnt_o[0] = valid_o & ready_i;
			assign idx_o = 1'sb0;
		end
		else begin : gen_normal_case
			wire [(2 ** (IdxW + 1)) - 2:0] req_tree;
			wire [(2 ** (IdxW + 1)) - 2:0] prio_tree;
			wire [(2 ** (IdxW + 1)) - 2:0] sel_tree;
			wire [(2 ** (IdxW + 1)) - 2:0] mask_tree;
			wire [(((2 ** (IdxW + 1)) - 2) >= 0 ? (((2 ** (IdxW + 1)) - 1) * IdxW) - 1 : ((3 - (2 ** (IdxW + 1))) * IdxW) + ((((2 ** (IdxW + 1)) - 2) * IdxW) - 1)):(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : ((2 ** (IdxW + 1)) - 2) * IdxW)] idx_tree;
			wire [(((2 ** (IdxW + 1)) - 2) >= 0 ? (((2 ** (IdxW + 1)) - 1) * DW) - 1 : ((3 - (2 ** (IdxW + 1))) * DW) + ((((2 ** (IdxW + 1)) - 2) * DW) - 1)):(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : ((2 ** (IdxW + 1)) - 2) * DW)] data_tree;
			wire [N - 1:0] prio_mask_d;
			reg [N - 1:0] prio_mask_q;
			genvar level;
			for (level = 0; level < (IdxW + 1); level = level + 1) begin : gen_tree
				localparam signed [31:0] Base0 = (2 ** level) - 1;
				localparam signed [31:0] Base1 = (2 ** (level + 1)) - 1;
				genvar offset;
				for (offset = 0; offset < (2 ** level); offset = offset + 1) begin : gen_level
					localparam signed [31:0] Pa = Base0 + offset;
					localparam signed [31:0] C0 = Base1 + (2 * offset);
					localparam signed [31:0] C1 = (Base1 + (2 * offset)) + 1;
					if (level == IdxW) begin : gen_leafs
						if (offset < N) begin : gen_assign
							assign req_tree[Pa] = req_i[offset];
							assign prio_tree[Pa] = req_i[offset] & prio_mask_q[offset];
							assign idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * IdxW+:IdxW] = offset;
							assign data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * DW+:DW] = data_i[((N - 1) - offset) * DW+:DW];
							assign gnt_o[offset] = (req_i[offset] & sel_tree[Pa]) & ready_i;
							assign prio_mask_d[offset] = (|req_i ? mask_tree[Pa] | (sel_tree[Pa] & ~ready_i) : prio_mask_q[offset]);
						end
						else begin : gen_tie_off
							assign req_tree[Pa] = 1'sb0;
							assign prio_tree[Pa] = 1'sb0;
							assign idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * IdxW+:IdxW] = 1'sb0;
							assign data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * DW+:DW] = 1'sb0;
							wire unused_sigs;
							assign unused_sigs = ^{mask_tree[Pa], sel_tree[Pa]};
						end
					end
					else begin : gen_nodes
						wire sel;
						assign sel = ~req_tree[C0] | (~prio_tree[C0] & prio_tree[C1]);
						assign req_tree[Pa] = req_tree[C0] | req_tree[C1];
						assign prio_tree[Pa] = prio_tree[C1] | prio_tree[C0];
						assign idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * IdxW+:IdxW] = (sel ? idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? C1 : ((2 ** (IdxW + 1)) - 2) - C1) * IdxW+:IdxW] : idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? C0 : ((2 ** (IdxW + 1)) - 2) - C0) * IdxW+:IdxW]);
						assign data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? Pa : ((2 ** (IdxW + 1)) - 2) - Pa) * DW+:DW] = (sel ? data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? C1 : ((2 ** (IdxW + 1)) - 2) - C1) * DW+:DW] : data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? C0 : ((2 ** (IdxW + 1)) - 2) - C0) * DW+:DW]);
						assign sel_tree[C0] = sel_tree[Pa] & ~sel;
						assign sel_tree[C1] = sel_tree[Pa] & sel;
						assign mask_tree[C0] = mask_tree[Pa];
						assign mask_tree[C1] = mask_tree[Pa] | sel_tree[C0];
					end
				end
			end
			if (EnDataPort) begin : gen_data_port
				assign data_o = data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : (2 ** (IdxW + 1)) - 2) * DW+:DW];
			end
			else begin : gen_no_dataport
				wire [DW - 1:0] unused_data;
				assign unused_data = data_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : (2 ** (IdxW + 1)) - 2) * DW+:DW];
				assign data_o = 1'sb1;
			end
			wire unused_prio_tree;
			assign unused_prio_tree = prio_tree[0];
			assign idx_o = idx_tree[(((2 ** (IdxW + 1)) - 2) >= 0 ? 0 : (2 ** (IdxW + 1)) - 2) * IdxW+:IdxW];
			assign valid_o = req_tree[0];
			assign sel_tree[0] = 1'b1;
			assign mask_tree[0] = 1'b0;
			always @(posedge clk_i or negedge rst_ni) begin : p_mask_reg
				if (!rst_ni)
					prio_mask_q <= 1'sb0;
				else
					prio_mask_q <= prio_mask_d;
			end
		end
	endgenerate
endmodule
module prim_arbiter_tree_dup (
	clk_i,
	rst_ni,
	req_chk_i,
	req_i,
	data_i,
	gnt_o,
	idx_o,
	valid_o,
	data_o,
	ready_i,
	err_o
);
	parameter signed [31:0] N = 8;
	parameter signed [31:0] DW = 32;
	parameter [0:0] EnDataPort = 1;
	parameter [0:0] FixedArb = 0;
	localparam signed [31:0] IdxW = $clog2(N);
	input clk_i;
	input rst_ni;
	input req_chk_i;
	input [N - 1:0] req_i;
	input [(N * DW) - 1:0] data_i;
	output wire [N - 1:0] gnt_o;
	output wire [IdxW - 1:0] idx_o;
	output wire valid_o;
	output wire [DW - 1:0] data_o;
	input ready_i;
	output wire err_o;
	localparam signed [31:0] ArbInstances = 2;
	wire [(ArbInstances * (((1 + N) + IdxW) + DW)) - 1:0] arb_output_buf;
	genvar i;
	generate
		for (i = 0; i < ArbInstances; i = i + 1) begin : gen_input_bufs
			wire [N - 1:0] req_buf;
			prim_buf #(.Width(N)) u_req_buf(
				.in_i(req_i),
				.out_o(req_buf)
			);
			wire [(N * DW) - 1:0] data_buf;
			genvar j;
			for (j = 0; j < N; j = j + 1) begin : gen_data_bufs
				prim_buf #(.Width(DW)) u_dat_buf(
					.in_i(data_i[((N - 1) - j) * DW+:DW]),
					.out_o(data_buf[((N - 1) - j) * DW+:DW])
				);
			end
			if (FixedArb) begin : gen_fixed_arbiter
				prim_arbiter_fixed #(
					.N(N),
					.DW(DW),
					.EnDataPort(EnDataPort)
				) u_arb(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.req_i(req_buf),
					.data_i(data_buf),
					.gnt_o(arb_output_buf[(i * (((1 + N) + IdxW) + DW)) + (N + (IdxW + (DW - 1)))-:((N + (IdxW + (DW - 1))) >= (IdxW + (DW + 0)) ? ((N + (IdxW + (DW - 1))) - (IdxW + (DW + 0))) + 1 : ((IdxW + (DW + 0)) - (N + (IdxW + (DW - 1)))) + 1)]),
					.idx_o(arb_output_buf[(i * (((1 + N) + IdxW) + DW)) + (IdxW + (DW - 1))-:((IdxW + (DW - 1)) >= (DW + 0) ? ((IdxW + (DW - 1)) - (DW + 0)) + 1 : ((DW + 0) - (IdxW + (DW - 1))) + 1)]),
					.valid_o(arb_output_buf[(i * (((1 + N) + IdxW) + DW)) + (1 + (N + (IdxW + (DW - 1))))]),
					.data_o(arb_output_buf[(i * (((1 + N) + IdxW) + DW)) + (DW - 1)-:DW]),
					.ready_i(ready_i)
				);
				wire unused_req_chk;
				assign unused_req_chk = req_chk_i;
			end
			else begin : gen_rr_arbiter
				prim_arbiter_tree #(
					.N(N),
					.DW(DW),
					.EnDataPort(EnDataPort)
				) u_arb(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.req_chk_i(req_chk_i),
					.req_i(req_buf),
					.data_i(data_buf),
					.gnt_o(arb_output_buf[(i * (((1 + N) + IdxW) + DW)) + (N + (IdxW + (DW - 1)))-:((N + (IdxW + (DW - 1))) >= (IdxW + (DW + 0)) ? ((N + (IdxW + (DW - 1))) - (IdxW + (DW + 0))) + 1 : ((IdxW + (DW + 0)) - (N + (IdxW + (DW - 1)))) + 1)]),
					.idx_o(arb_output_buf[(i * (((1 + N) + IdxW) + DW)) + (IdxW + (DW - 1))-:((IdxW + (DW - 1)) >= (DW + 0) ? ((IdxW + (DW - 1)) - (DW + 0)) + 1 : ((DW + 0) - (IdxW + (DW - 1))) + 1)]),
					.valid_o(arb_output_buf[(i * (((1 + N) + IdxW) + DW)) + (1 + (N + (IdxW + (DW - 1))))]),
					.data_o(arb_output_buf[(i * (((1 + N) + IdxW) + DW)) + (DW - 1)-:DW]),
					.ready_i(ready_i)
				);
			end
		end
	endgenerate
	assign gnt_o = arb_output_buf[(1 * (((1 + N) + IdxW) + DW)) + (N + (IdxW + (DW - 1)))-:((N + (IdxW + (DW - 1))) >= (IdxW + (DW + 0)) ? ((N + (IdxW + (DW - 1))) - (IdxW + (DW + 0))) + 1 : ((IdxW + (DW + 0)) - (N + (IdxW + (DW - 1)))) + 1)];
	assign idx_o = arb_output_buf[(1 * (((1 + N) + IdxW) + DW)) + (IdxW + (DW - 1))-:((IdxW + (DW - 1)) >= (DW + 0) ? ((IdxW + (DW - 1)) - (DW + 0)) + 1 : ((DW + 0) - (IdxW + (DW - 1))) + 1)];
	assign valid_o = arb_output_buf[(1 * (((1 + N) + IdxW) + DW)) + (1 + (N + (IdxW + (DW - 1))))];
	assign data_o = arb_output_buf[(1 * (((1 + N) + IdxW) + DW)) + (DW - 1)-:DW];
	wire [0:0] output_delta;
	generate
		for (i = 0; i < 1; i = i + 1) begin : gen_checks
			assign output_delta[i] = arb_output_buf[1 * (((1 + N) + IdxW) + DW)+:((1 + N) + IdxW) + DW] != arb_output_buf[i * (((1 + N) + IdxW) + DW)+:((1 + N) + IdxW) + DW];
		end
	endgenerate
	wire err_d;
	reg err_q;
	assign err_d = |output_delta;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			err_q <= 1'sb0;
		else
			err_q <= err_d | err_q;
	assign err_o = err_q;
endmodule
module prim_badbit_ram_1p (
	clk_i,
	req_i,
	write_i,
	addr_i,
	wdata_i,
	wmask_i,
	rdata_o
);
	parameter signed [31:0] Width = 32;
	parameter signed [31:0] Depth = 128;
	parameter signed [31:0] DataBitsPerMask = 1;
	parameter MemInitFile = "";
	localparam signed [31:0] Aw = $clog2(Depth);
	input wire clk_i;
	input wire req_i;
	input wire write_i;
	input wire [Aw - 1:0] addr_i;
	input wire [Width - 1:0] wdata_i;
	input wire [Width - 1:0] wmask_i;
	output wire [Width - 1:0] rdata_o;
	wire [Width - 1:0] sram_rdata;
	prim_generic_ram_1p #(
		.Width(Width),
		.Depth(Depth),
		.DataBitsPerMask(DataBitsPerMask),
		.MemInitFile(MemInitFile)
	) u_mem(
		.clk_i(clk_i),
		.cfg_i(1'sb0),
		.req_i(req_i),
		.write_i(write_i),
		.addr_i(addr_i),
		.wdata_i(wdata_i),
		.wmask_i(wmask_i),
		.rdata_o(sram_rdata)
	);
	wire [31:0] width;
	assign width = Width;
	wire [31:0] addr;
	wire [127:0] wdata;
	wire [127:0] wmask;
	wire [127:0] rdata;
	assign addr = {{32 - Aw {1'b0}}, addr_i};
	assign wdata = {{128 - Width {1'b0}}, wdata_i};
	assign wmask = {{128 - Width {1'b0}}, wmask_i};
	assign rdata = {{128 - Width {1'b0}}, sram_rdata};
	logic [127:0] bad_bit_mask;
	assign bad_bit_mask = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	assign rdata_o = sram_rdata ^ bad_bit_mask;
endmodule
module prim_blanker (
	in_i,
	en_i,
	out_o
);
	parameter signed [31:0] Width = 1;
	input wire [Width - 1:0] in_i;
	input wire en_i;
	output wire [Width - 1:0] out_o;
	prim_and2 #(.Width(Width)) u_blank_and(
		.in0_i(in_i),
		.in1_i({Width {en_i}}),
		.out_o(out_o)
	);
endmodule
module prim_buf (
	in_i,
	out_o
);
	parameter signed [31:0] Width = 1;
	input [Width - 1:0] in_i;
	output wire [Width - 1:0] out_o;
	parameter integer Impl = 32'sd0;
	generate
		if (Impl == 32'sd2) begin : gen_xilinx
			prim_xilinx_buf #(.Width(Width)) u_impl_xilinx(
				.in_i(in_i),
				.out_o(out_o)
			);
		end
		else begin : gen_generic
			prim_generic_buf #(.Width(Width)) u_impl_generic(
				.in_i(in_i),
				.out_o(out_o)
			);
		end
	endgenerate
endmodule
module prim_cdc_rand_delay (
	clk_i,
	rst_ni,
	prev_data_i,
	src_data_i,
	dst_data_o
);
	parameter signed [31:0] DataWidth = 1;
	parameter [0:0] Enable = 1;
	input wire clk_i;
	input wire rst_ni;
	input wire [DataWidth - 1:0] prev_data_i;
	input wire [DataWidth - 1:0] src_data_i;
	output wire [DataWidth - 1:0] dst_data_o;
	assign dst_data_o = src_data_i;
endmodule
module prim_clock_gating (
	clk_i,
	en_i,
	test_en_i,
	clk_o
);
	parameter [0:0] NoFpgaGate = 1'b0;
	parameter [0:0] FpgaBufGlobal = 1'b1;
	input clk_i;
	input en_i;
	input test_en_i;
	output wire clk_o;
	parameter integer Impl = 32'sd0;
	generate
		if (Impl == 32'sd2) begin : gen_xilinx
			prim_xilinx_clock_gating #(
				.FpgaBufGlobal(FpgaBufGlobal),
				.NoFpgaGate(NoFpgaGate)
			) u_impl_xilinx(
				.clk_i(clk_i),
				.en_i(en_i),
				.test_en_i(test_en_i),
				.clk_o(clk_o)
			);
		end
		else begin : gen_generic
			prim_generic_clock_gating #(
				.FpgaBufGlobal(FpgaBufGlobal),
				.NoFpgaGate(NoFpgaGate)
			) u_impl_generic(
				.clk_i(clk_i),
				.en_i(en_i),
				.test_en_i(test_en_i),
				.clk_o(clk_o)
			);
		end
	endgenerate
endmodule
module prim_clock_gating_sync (
	clk_i,
	rst_ni,
	test_en_i,
	async_en_i,
	en_o,
	clk_o
);
	input clk_i;
	input rst_ni;
	input test_en_i;
	input async_en_i;
	output wire en_o;
	output wire clk_o;
	prim_flop_2sync #(.Width(1)) i_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(async_en_i),
		.q_o(en_o)
	);
	prim_clock_gating i_cg(
		.clk_i(clk_i),
		.en_i(en_o),
		.test_en_i(test_en_i),
		.clk_o(clk_o)
	);
endmodule
module prim_clock_mux2 (
	clk0_i,
	clk1_i,
	sel_i,
	clk_o
);
	parameter [0:0] NoFpgaBufG = 1'b0;
	input clk0_i;
	input clk1_i;
	input sel_i;
	output wire clk_o;
	parameter integer Impl = 32'sd0;
	generate
		if (Impl == 32'sd2) begin : gen_xilinx
			prim_xilinx_clock_mux2 #(.NoFpgaBufG(NoFpgaBufG)) u_impl_xilinx(
				.clk0_i(clk0_i),
				.clk1_i(clk1_i),
				.sel_i(sel_i),
				.clk_o(clk_o)
			);
		end
		else begin : gen_generic
			prim_generic_clock_mux2 #(.NoFpgaBufG(NoFpgaBufG)) u_impl_generic(
				.clk0_i(clk0_i),
				.clk1_i(clk1_i),
				.sel_i(sel_i),
				.clk_o(clk_o)
			);
		end
	endgenerate
endmodule
module prim_count (
	clk_i,
	rst_ni,
	clr_i,
	set_i,
	set_cnt_i,
	incr_en_i,
	decr_en_i,
	step_i,
	cnt_o,
	cnt_next_o,
	err_o
);
	parameter signed [31:0] Width = 2;
	parameter [Width - 1:0] ResetValue = 1'sb0;
	parameter [0:0] EnableAlertTriggerSVA = 1;
	input clk_i;
	input rst_ni;
	input clr_i;
	input set_i;
	input [Width - 1:0] set_cnt_i;
	input incr_en_i;
	input decr_en_i;
	input [Width - 1:0] step_i;
	output wire [Width - 1:0] cnt_o;
	output wire [Width - 1:0] cnt_next_o;
	output wire err_o;
	localparam signed [31:0] NumCnt = 2;
	localparam [(NumCnt * Width) - 1:0] ResetValues = {{Width {1'b1}} - ResetValue, ResetValue};
	wire [(NumCnt * Width) - 1:0] cnt_d;
	wire [(NumCnt * Width) - 1:0] cnt_q;
	wire [(NumCnt * Width) - 1:0] fpv_force;
	assign fpv_force = 1'sb0;
	genvar k;
	generate
		for (k = 0; k < NumCnt; k = k + 1) begin : gen_cnts
			wire incr_en;
			wire decr_en;
			wire [Width - 1:0] set_val;
			if (k == 0) begin : gen_up_cnt
				assign incr_en = incr_en_i;
				assign decr_en = decr_en_i;
				assign set_val = set_cnt_i;
			end
			else begin : gen_dn_cnt
				assign incr_en = decr_en_i;
				assign decr_en = incr_en_i;
				assign set_val = {Width {1'b1}} - set_cnt_i;
			end
			wire [Width:0] ext_cnt;
			assign ext_cnt = (decr_en ? {1'b0, cnt_q[k * Width+:Width]} - {1'b0, step_i} : (incr_en ? {1'b0, cnt_q[k * Width+:Width]} + {1'b0, step_i} : {1'b0, cnt_q[k * Width+:Width]}));
			wire uflow;
			wire oflow;
			assign oflow = incr_en && ext_cnt[Width];
			assign uflow = decr_en && ext_cnt[Width];
			wire [Width - 1:0] cnt_sat;
			assign cnt_sat = (uflow ? {Width {1'sb0}} : (oflow ? {Width {1'b1}} : ext_cnt[Width - 1:0]));
			wire cnt_en;
			assign cnt_en = (incr_en ^ decr_en) && ((incr_en && !(&cnt_q[k * Width+:Width])) || (decr_en && (cnt_q[k * Width+:Width] != {Width * 1 {1'sb0}})));
			assign cnt_d[k * Width+:Width] = (clr_i ? ResetValues[k * Width+:Width] : (set_i ? set_val : (cnt_en ? cnt_sat : cnt_q[k * Width+:Width])));
			wire [Width - 1:0] cnt_unforced_q;
			prim_flop #(
				.Width(Width),
				.ResetValue(ResetValues[k * Width+:Width])
			) u_cnt_flop(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(cnt_d[k * Width+:Width]),
				.q_o(cnt_unforced_q)
			);
			assign cnt_q[k * Width+:Width] = fpv_force[k * Width+:Width] + cnt_unforced_q;
		end
	endgenerate
	wire [Width:0] sum;
	assign sum = cnt_q[0+:Width] + cnt_q[Width+:Width];
	assign err_o = sum != {1'b0, {Width {1'b1}}};
	assign cnt_o = cnt_q[0+:Width];
	assign cnt_next_o = cnt_d[0+:Width];
endmodule
module prim_diff_decode (
	clk_i,
	rst_ni,
	diff_pi,
	diff_ni,
	level_o,
	rise_o,
	fall_o,
	event_o,
	sigint_o
);
	parameter [0:0] AsyncOn = 1'b0;
	input clk_i;
	input rst_ni;
	input diff_pi;
	input diff_ni;
	output wire level_o;
	output reg rise_o;
	output reg fall_o;
	output wire event_o;
	output reg sigint_o;
	reg level_d;
	reg level_q;
	generate
		if (AsyncOn) begin : gen_async
			reg [1:0] state_d;
			reg [1:0] state_q;
			wire diff_p_edge;
			wire diff_n_edge;
			wire diff_check_ok;
			wire level;
			reg diff_pq;
			reg diff_nq;
			wire diff_pd;
			wire diff_nd;
			prim_flop_2sync #(
				.Width(1),
				.ResetValue(1'sb0)
			) i_sync_p(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(diff_pi),
				.q_o(diff_pd)
			);
			prim_flop_2sync #(
				.Width(1),
				.ResetValue(1'b1)
			) i_sync_n(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(diff_ni),
				.q_o(diff_nd)
			);
			assign diff_p_edge = diff_pq ^ diff_pd;
			assign diff_n_edge = diff_nq ^ diff_nd;
			assign diff_check_ok = diff_pd ^ diff_nd;
			assign level = diff_pd;
			assign level_o = level_d;
			assign event_o = rise_o | fall_o;
			always @(*) begin : p_diff_fsm
				state_d = state_q;
				level_d = level_q;
				rise_o = 1'b0;
				fall_o = 1'b0;
				sigint_o = 1'b0;
				case (state_q)
					2'd0:
						if (diff_check_ok) begin
							level_d = level;
							if (diff_p_edge && diff_n_edge)
								if (level)
									rise_o = 1'b1;
								else
									fall_o = 1'b1;
						end
						else if (diff_p_edge || diff_n_edge)
							state_d = 2'd1;
						else begin
							state_d = 2'd2;
							sigint_o = 1'b1;
						end
					2'd1:
						if (diff_check_ok) begin
							state_d = 2'd0;
							level_d = level;
							if (level)
								rise_o = 1'b1;
							else
								fall_o = 1'b1;
						end
						else begin
							state_d = 2'd2;
							sigint_o = 1'b1;
						end
					2'd2: begin
						sigint_o = 1'b1;
						if (diff_check_ok) begin
							state_d = 2'd0;
							sigint_o = 1'b0;
						end
					end
					default:
						;
				endcase
			end
			always @(posedge clk_i or negedge rst_ni) begin : p_sync_reg
				if (!rst_ni) begin
					state_q <= 2'd0;
					diff_pq <= 1'b0;
					diff_nq <= 1'b1;
					level_q <= 1'b0;
				end
				else begin
					state_q <= state_d;
					diff_pq <= diff_pd;
					diff_nq <= diff_nd;
					level_q <= level_d;
				end
			end
		end
		else begin : gen_no_async
			reg diff_pq;
			wire diff_pd;
			assign diff_pd = diff_pi;
			wire [1:1] sv2v_tmp_E2CC7;
			assign sv2v_tmp_E2CC7 = ~(diff_pi ^ diff_ni);
			always @(*) sigint_o = sv2v_tmp_E2CC7;
			assign level_o = (sigint_o ? level_q : diff_pi);
			wire [1:1] sv2v_tmp_75F4D;
			assign sv2v_tmp_75F4D = level_o;
			always @(*) level_d = sv2v_tmp_75F4D;
			wire [1:1] sv2v_tmp_97BB0;
			assign sv2v_tmp_97BB0 = (~diff_pq & diff_pi) & ~sigint_o;
			always @(*) rise_o = sv2v_tmp_97BB0;
			wire [1:1] sv2v_tmp_B4F46;
			assign sv2v_tmp_B4F46 = (diff_pq & ~diff_pi) & ~sigint_o;
			always @(*) fall_o = sv2v_tmp_B4F46;
			assign event_o = rise_o | fall_o;
			always @(posedge clk_i or negedge rst_ni) begin : p_edge_reg
				if (!rst_ni) begin
					diff_pq <= 1'b0;
					level_q <= 1'b0;
				end
				else begin
					diff_pq <= diff_pd;
					level_q <= level_d;
				end
			end
		end
	endgenerate
endmodule
module prim_edn_req (
	clk_i,
	rst_ni,
	req_chk_i,
	req_i,
	ack_o,
	data_o,
	fips_o,
	err_o,
	clk_edn_i,
	rst_edn_ni,
	edn_o,
	edn_i
);
	parameter signed [31:0] OutWidth = 32;
	parameter [0:0] RepCheck = 0;
	parameter [0:0] EnRstChks = 0;
	parameter [31:0] MaxLatency = 0;
	input clk_i;
	input rst_ni;
	input req_chk_i;
	input req_i;
	output wire ack_o;
	output wire [OutWidth - 1:0] data_o;
	output wire fips_o;
	output wire err_o;
	input clk_edn_i;
	input rst_edn_ni;
	output wire [0:0] edn_o;
	localparam [31:0] edn_pkg_ENDPOINT_BUS_WIDTH = 32;
	input wire [33:0] edn_i;
	wire word_req;
	wire word_ack;
	assign word_req = req_i & ~ack_o;
	wire [31:0] word_data;
	wire word_fips;
	localparam signed [31:0] SyncWidth = 33;
	prim_sync_reqack_data #(
		.Width(SyncWidth),
		.EnRstChks(EnRstChks),
		.DataSrc2Dst(1'b0),
		.DataReg(1'b0)
	) u_prim_sync_reqack_data(
		.clk_src_i(clk_i),
		.rst_src_ni(rst_ni),
		.clk_dst_i(clk_edn_i),
		.rst_dst_ni(rst_edn_ni),
		.req_chk_i(req_chk_i),
		.src_req_i(word_req),
		.src_ack_o(word_ack),
		.dst_req_o(edn_o[0]),
		.dst_ack_i(edn_i[33]),
		.data_i({edn_i[32], edn_i[31-:edn_pkg_ENDPOINT_BUS_WIDTH]}),
		.data_o({word_fips, word_data})
	);
	generate
		if (RepCheck) begin : gen_rep_chk
			reg [31:0] word_data_q;
			always @(posedge clk_i)
				if (word_ack)
					word_data_q <= word_data;
			reg chk_rep;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					chk_rep <= 1'sb0;
				else if (word_ack)
					chk_rep <= 1'b1;
			wire err_d;
			reg err_q;
			assign err_d = (req_i && ack_o ? 1'b0 : ((chk_rep && word_ack) && (word_data == word_data_q) ? 1'b1 : err_q));
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					err_q <= 1'b0;
				else
					err_q <= err_d;
			assign err_o = err_q;
		end
		else begin : gen_no_rep_chk
			assign err_o = 1'sb0;
		end
	endgenerate
	prim_packer_fifo #(
		.InW(edn_pkg_ENDPOINT_BUS_WIDTH),
		.OutW(OutWidth),
		.ClearOnRead(1'b0)
	) u_prim_packer_fifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(1'b0),
		.wvalid_i(word_ack),
		.wdata_i(word_data),
		.rvalid_o(ack_o),
		.rdata_o(data_o),
		.rready_i(1'b1)
	);
	wire fips_d;
	reg fips_q;
	assign fips_d = (req_i && ack_o ? 1'b1 : (word_ack ? fips_q & word_fips : fips_q));
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			fips_q <= 1'b1;
		else
			fips_q <= fips_d;
	assign fips_o = fips_q;
	wire unused_param_maxlatency;
	assign unused_param_maxlatency = ^MaxLatency;
endmodule
module prim_esc_receiver (
	clk_i,
	rst_ni,
	esc_req_o,
	esc_rx_o,
	esc_tx_i
);
	parameter signed [31:0] N_ESC_SEV = 4;
	parameter signed [31:0] PING_CNT_DW = 16;
	localparam signed [31:0] MarginFactor = 4;
	localparam signed [31:0] NumWaitCounts = 2;
	localparam signed [31:0] NumTimeoutCounts = 2;
	parameter signed [31:0] TimeoutCntDw = ((2 + $clog2(N_ESC_SEV)) + 2) + PING_CNT_DW;
	input clk_i;
	input rst_ni;
	output wire esc_req_o;
	output wire [1:0] esc_rx_o;
	input wire [1:0] esc_tx_i;
	wire esc_level;
	wire esc_p;
	wire esc_n;
	wire sigint_detected;
	prim_buf #(.Width(2)) u_prim_buf_esc(
		.in_i({esc_tx_i[0], esc_tx_i[1]}),
		.out_o({esc_n, esc_p})
	);
	prim_diff_decode #(.AsyncOn(1'b0)) u_decode_esc(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.diff_pi(esc_p),
		.diff_ni(esc_n),
		.level_o(esc_level),
		.sigint_o(sigint_detected)
	);
	reg ping_en;
	wire timeout_cnt_error;
	wire timeout_cnt_set;
	wire timeout_cnt_en;
	wire [TimeoutCntDw - 1:0] timeout_cnt;
	assign timeout_cnt_set = ping_en && !(&timeout_cnt);
	assign timeout_cnt_en = (timeout_cnt > {TimeoutCntDw {1'sb0}}) && !(&timeout_cnt);
	function automatic signed [TimeoutCntDw - 1:0] sv2v_cast_1053F_signed;
		input reg signed [TimeoutCntDw - 1:0] inp;
		sv2v_cast_1053F_signed = inp;
	endfunction
	prim_count #(
		.Width(TimeoutCntDw),
		.EnableAlertTriggerSVA(0)
	) u_prim_count(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(1'b0),
		.set_i(timeout_cnt_set),
		.set_cnt_i(sv2v_cast_1053F_signed(1)),
		.incr_en_i(timeout_cnt_en),
		.decr_en_i(1'b0),
		.step_i(sv2v_cast_1053F_signed(1)),
		.cnt_o(timeout_cnt),
		.err_o(timeout_cnt_error)
	);
	reg esc_req;
	prim_sec_anchor_buf #(.Width(1)) u_prim_buf_esc_req(
		.in_i((esc_req || &timeout_cnt) || timeout_cnt_error),
		.out_o(esc_req_o)
	);
	reg [2:0] state_d;
	reg [2:0] state_q;
	reg resp_pd;
	wire resp_pq;
	reg resp_nd;
	wire resp_nq;
	prim_sec_anchor_flop #(
		.Width(2),
		.ResetValue(2'b10)
	) u_prim_flop_esc(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i({resp_nd, resp_pd}),
		.q_o({resp_nq, resp_pq})
	);
	assign esc_rx_o[1] = resp_pq;
	assign esc_rx_o[0] = resp_nq;
	always @(*) begin : p_fsm
		state_d = state_q;
		resp_pd = 1'b0;
		resp_nd = 1'b1;
		esc_req = 1'b0;
		ping_en = 1'b0;
		case (state_q)
			3'd0:
				if (esc_level) begin
					state_d = 3'd1;
					resp_pd = ~resp_pq;
					resp_nd = resp_pq;
				end
			3'd1: begin
				state_d = 3'd2;
				resp_pd = ~resp_pq;
				resp_nd = resp_pq;
				if (esc_level) begin
					state_d = 3'd3;
					esc_req = 1'b1;
				end
			end
			3'd2: begin
				state_d = 3'd0;
				resp_pd = ~resp_pq;
				resp_nd = resp_pq;
				ping_en = 1'b1;
				if (esc_level) begin
					state_d = 3'd3;
					esc_req = 1'b1;
				end
			end
			3'd3: begin
				state_d = 3'd0;
				if (esc_level) begin
					state_d = 3'd3;
					resp_pd = ~resp_pq;
					resp_nd = resp_pq;
					esc_req = 1'b1;
				end
			end
			3'd4: begin
				state_d = 3'd0;
				esc_req = 1'b1;
				if (sigint_detected) begin
					state_d = 3'd4;
					resp_pd = ~resp_pq;
					resp_nd = ~resp_pq;
				end
			end
			default: state_d = 3'd0;
		endcase
		if (sigint_detected && (state_q != 3'd4)) begin
			state_d = 3'd4;
			resp_pd = 1'b0;
			resp_nd = 1'b0;
		end
	end
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		if (!rst_ni)
			state_q <= 3'd0;
		else
			state_q <= state_d;
	end
endmodule
module prim_esc_sender (
	clk_i,
	rst_ni,
	ping_req_i,
	ping_ok_o,
	integ_fail_o,
	esc_req_i,
	esc_rx_i,
	esc_tx_o
);
	input clk_i;
	input rst_ni;
	input ping_req_i;
	output reg ping_ok_o;
	output reg integ_fail_o;
	input esc_req_i;
	input wire [1:0] esc_rx_i;
	output wire [1:0] esc_tx_o;
	wire resp;
	wire resp_n;
	wire resp_p;
	wire sigint_detected;
	prim_sec_anchor_buf #(.Width(2)) u_prim_buf_resp(
		.in_i({esc_rx_i[0], esc_rx_i[1]}),
		.out_o({resp_n, resp_p})
	);
	prim_diff_decode #(.AsyncOn(1'b0)) u_decode_resp(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.diff_pi(resp_p),
		.diff_ni(resp_n),
		.level_o(resp),
		.sigint_o(sigint_detected)
	);
	wire ping_req_d;
	reg ping_req_q;
	wire esc_req_d;
	reg esc_req_q;
	reg esc_req_q1;
	assign ping_req_d = ping_req_i;
	assign esc_req_d = esc_req_i;
	wire esc_p;
	assign esc_p = (esc_req_i | esc_req_q) | (ping_req_d & ~ping_req_q);
	prim_sec_anchor_buf #(.Width(2)) u_prim_buf_esc(
		.in_i({~esc_p, esc_p}),
		.out_o({esc_tx_o[0], esc_tx_o[1]})
	);
	reg [2:0] state_d;
	reg [2:0] state_q;
	always @(*) begin : p_fsm
		state_d = state_q;
		ping_ok_o = 1'b0;
		integ_fail_o = sigint_detected;
		case (state_q)
			3'd0: begin
				if (esc_req_i)
					state_d = 3'd2;
				else if (ping_req_d & ~ping_req_q)
					state_d = 3'd3;
				if (resp)
					integ_fail_o = 1'b1;
			end
			3'd1: begin
				state_d = 3'd2;
				if (!esc_tx_o[1] || resp) begin
					state_d = 3'd0;
					integ_fail_o = sigint_detected | resp;
				end
			end
			3'd2: begin
				state_d = 3'd1;
				if (!esc_tx_o[1] || !resp) begin
					state_d = 3'd0;
					integ_fail_o = sigint_detected | ~resp;
				end
			end
			3'd3: begin
				state_d = 3'd4;
				if (esc_req_i)
					state_d = 3'd1;
				else if (!resp) begin
					state_d = 3'd0;
					integ_fail_o = 1'b1;
				end
			end
			3'd4: begin
				state_d = 3'd5;
				if (esc_req_i)
					state_d = 3'd2;
				else if (resp) begin
					state_d = 3'd0;
					integ_fail_o = 1'b1;
				end
			end
			3'd5: begin
				state_d = 3'd6;
				if (esc_req_i)
					state_d = 3'd1;
				else if (!resp) begin
					state_d = 3'd0;
					integ_fail_o = 1'b1;
				end
			end
			3'd6: begin
				state_d = 3'd0;
				if (esc_req_i)
					state_d = 3'd2;
				else if (resp)
					integ_fail_o = 1'b1;
				else
					ping_ok_o = ping_req_i;
			end
			default: state_d = 3'd0;
		endcase
		if (sigint_detected) begin
			ping_ok_o = 1'b0;
			state_d = 3'd0;
		end
		if (((esc_req_i || esc_req_q) || esc_req_q1) && ping_req_i)
			ping_ok_o = 1'b1;
	end
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		if (!rst_ni) begin
			state_q <= 3'd0;
			esc_req_q <= 1'b0;
			esc_req_q1 <= 1'b0;
			ping_req_q <= 1'b0;
		end
		else begin
			state_q <= state_d;
			esc_req_q <= esc_req_d;
			esc_req_q1 <= esc_req_q;
			ping_req_q <= ping_req_d;
		end
	end
endmodule
module prim_fifo_async (
	clk_wr_i,
	rst_wr_ni,
	wvalid_i,
	wready_o,
	wdata_i,
	wdepth_o,
	clk_rd_i,
	rst_rd_ni,
	rvalid_o,
	rready_i,
	rdata_o,
	rdepth_o
);
	parameter [31:0] Width = 16;
	parameter [31:0] Depth = 4;
	parameter [0:0] OutputZeroIfEmpty = 1'b0;
	parameter [0:0] OutputZeroIfInvalid = 1'b0;
	localparam [31:0] DepthW = $clog2(Depth + 1);
	input wire clk_wr_i;
	input wire rst_wr_ni;
	input wire wvalid_i;
	output wire wready_o;
	input wire [Width - 1:0] wdata_i;
	output wire [DepthW - 1:0] wdepth_o;
	input wire clk_rd_i;
	input wire rst_rd_ni;
	output wire rvalid_o;
	input wire rready_i;
	output wire [Width - 1:0] rdata_o;
	output wire [DepthW - 1:0] rdepth_o;
	localparam [31:0] PTRV_W = (Depth == 1 ? 1 : $clog2(Depth));
	localparam [31:0] PTR_WIDTH = (Depth == 1 ? 1 : PTRV_W + 1);
	reg [PTR_WIDTH - 1:0] fifo_wptr_q;
	wire [PTR_WIDTH - 1:0] fifo_wptr_d;
	reg [PTR_WIDTH - 1:0] fifo_rptr_q;
	wire [PTR_WIDTH - 1:0] fifo_rptr_d;
	wire [PTR_WIDTH - 1:0] fifo_wptr_sync_combi;
	wire [PTR_WIDTH - 1:0] fifo_rptr_sync_combi;
	wire [PTR_WIDTH - 1:0] fifo_wptr_gray_sync;
	wire [PTR_WIDTH - 1:0] fifo_rptr_gray_sync;
	reg [PTR_WIDTH - 1:0] fifo_rptr_sync_q;
	reg [PTR_WIDTH - 1:0] fifo_wptr_gray_q;
	wire [PTR_WIDTH - 1:0] fifo_wptr_gray_d;
	reg [PTR_WIDTH - 1:0] fifo_rptr_gray_q;
	wire [PTR_WIDTH - 1:0] fifo_rptr_gray_d;
	wire fifo_incr_wptr;
	wire fifo_incr_rptr;
	wire full_wclk;
	wire full_rclk;
	wire empty_rclk;
	reg [Width - 1:0] storage [0:Depth - 1];
	assign fifo_incr_wptr = wvalid_i & wready_o;
	function automatic [PTR_WIDTH - 1:0] sv2v_cast_06624;
		input reg [PTR_WIDTH - 1:0] inp;
		sv2v_cast_06624 = inp;
	endfunction
	assign fifo_wptr_d = fifo_wptr_q + sv2v_cast_06624(1'b1);
	always @(posedge clk_wr_i or negedge rst_wr_ni)
		if (!rst_wr_ni)
			fifo_wptr_q <= 1'sb0;
		else if (fifo_incr_wptr)
			fifo_wptr_q <= fifo_wptr_d;
	always @(posedge clk_wr_i or negedge rst_wr_ni)
		if (!rst_wr_ni)
			fifo_wptr_gray_q <= 1'sb0;
		else if (fifo_incr_wptr)
			fifo_wptr_gray_q <= fifo_wptr_gray_d;
	prim_flop_2sync #(.Width(PTR_WIDTH)) sync_wptr(
		.clk_i(clk_rd_i),
		.rst_ni(rst_rd_ni),
		.d_i(fifo_wptr_gray_q),
		.q_o(fifo_wptr_gray_sync)
	);
	assign fifo_incr_rptr = rvalid_o & rready_i;
	assign fifo_rptr_d = fifo_rptr_q + sv2v_cast_06624(1'b1);
	always @(posedge clk_rd_i or negedge rst_rd_ni)
		if (!rst_rd_ni)
			fifo_rptr_q <= 1'sb0;
		else if (fifo_incr_rptr)
			fifo_rptr_q <= fifo_rptr_d;
	always @(posedge clk_rd_i or negedge rst_rd_ni)
		if (!rst_rd_ni)
			fifo_rptr_gray_q <= 1'sb0;
		else if (fifo_incr_rptr)
			fifo_rptr_gray_q <= fifo_rptr_gray_d;
	prim_flop_2sync #(.Width(PTR_WIDTH)) sync_rptr(
		.clk_i(clk_wr_i),
		.rst_ni(rst_wr_ni),
		.d_i(fifo_rptr_gray_q),
		.q_o(fifo_rptr_gray_sync)
	);
	always @(posedge clk_wr_i or negedge rst_wr_ni)
		if (!rst_wr_ni)
			fifo_rptr_sync_q <= 1'sb0;
		else
			fifo_rptr_sync_q <= fifo_rptr_sync_combi;
	wire [PTR_WIDTH - 1:0] xor_mask;
	assign xor_mask = sv2v_cast_06624(1'b1) << (PTR_WIDTH - 1);
	assign full_wclk = fifo_wptr_q == (fifo_rptr_sync_q ^ xor_mask);
	assign full_rclk = fifo_wptr_sync_combi == (fifo_rptr_q ^ xor_mask);
	assign empty_rclk = fifo_wptr_sync_combi == fifo_rptr_q;
	function automatic [DepthW - 1:0] sv2v_cast_00304;
		input reg [DepthW - 1:0] inp;
		sv2v_cast_00304 = inp;
	endfunction
	generate
		if (Depth > 1) begin : g_depth_calc
			wire wptr_msb;
			wire rptr_sync_msb;
			wire [PTRV_W - 1:0] wptr_value;
			wire [PTRV_W - 1:0] rptr_sync_value;
			assign wptr_msb = fifo_wptr_q[PTR_WIDTH - 1];
			assign rptr_sync_msb = fifo_rptr_sync_q[PTR_WIDTH - 1];
			assign wptr_value = fifo_wptr_q[0+:PTRV_W];
			assign rptr_sync_value = fifo_rptr_sync_q[0+:PTRV_W];
			assign wdepth_o = (full_wclk ? sv2v_cast_00304(Depth) : (wptr_msb == rptr_sync_msb ? sv2v_cast_00304(wptr_value) - sv2v_cast_00304(rptr_sync_value) : (sv2v_cast_00304(Depth) - sv2v_cast_00304(rptr_sync_value)) + sv2v_cast_00304(wptr_value)));
			wire rptr_msb;
			wire wptr_sync_msb;
			wire [PTRV_W - 1:0] rptr_value;
			wire [PTRV_W - 1:0] wptr_sync_value;
			assign wptr_sync_msb = fifo_wptr_sync_combi[PTR_WIDTH - 1];
			assign rptr_msb = fifo_rptr_q[PTR_WIDTH - 1];
			assign wptr_sync_value = fifo_wptr_sync_combi[0+:PTRV_W];
			assign rptr_value = fifo_rptr_q[0+:PTRV_W];
			assign rdepth_o = (full_rclk ? sv2v_cast_00304(Depth) : (wptr_sync_msb == rptr_msb ? sv2v_cast_00304(wptr_sync_value) - sv2v_cast_00304(rptr_value) : (sv2v_cast_00304(Depth) - sv2v_cast_00304(rptr_value)) + sv2v_cast_00304(wptr_sync_value)));
		end
		else begin : g_no_depth_calc
			assign rdepth_o = full_rclk;
			assign wdepth_o = full_wclk;
		end
	endgenerate
	assign wready_o = ~full_wclk;
	assign rvalid_o = ~empty_rclk;
	wire [Width - 1:0] rdata_int;
	generate
		if (Depth > 1) begin : g_storage_mux
			always @(posedge clk_wr_i)
				if (fifo_incr_wptr)
					storage[fifo_wptr_q[PTRV_W - 1:0]] <= wdata_i;
			assign rdata_int = storage[fifo_rptr_q[PTRV_W - 1:0]];
		end
		else begin : g_storage_simple
			always @(posedge clk_wr_i)
				if (fifo_incr_wptr)
					storage[0] <= wdata_i;
			assign rdata_int = storage[0];
		end
		if (OutputZeroIfEmpty == 1'b1) begin : gen_output_zero
			if (OutputZeroIfInvalid == 1'b1) begin : gen_invalid_zero
				assign rdata_o = (empty_rclk ? {Width {1'sb0}} : (rvalid_o ? rdata_int : {Width {1'sb0}}));
			end
			else begin : gen_invalid_non_zero
				assign rdata_o = (empty_rclk ? {Width {1'sb0}} : rdata_int);
			end
		end
		else begin : gen_no_output_zero
			if (OutputZeroIfInvalid == 1'b1) begin : gen_invalid_zero
				assign rdata_o = (rvalid_o ? rdata_int : {Width {1'sb0}});
			end
			else begin : gen_invalid_non_zero
				assign rdata_o = rdata_int;
			end
		end
		if (Depth > 2) begin : g_full_gray_conversion
			function automatic [PTR_WIDTH - 1:0] dec2gray;
				input reg [PTR_WIDTH - 1:0] decval;
				reg [PTR_WIDTH - 1:0] decval_sub;
				reg [PTR_WIDTH - 1:0] decval_in;
				reg unused_decval_msb;
				begin
					decval_sub = (sv2v_cast_06624(Depth) - {1'b0, decval[PTR_WIDTH - 2:0]}) - 1'b1;
					decval_in = (decval[PTR_WIDTH - 1] ? decval_sub : decval);
					unused_decval_msb = decval_in[PTR_WIDTH - 1];
					decval_in[PTR_WIDTH - 1] = 1'b0;
					dec2gray = decval_in;
					dec2gray = dec2gray ^ (decval_in >> 1);
					dec2gray[PTR_WIDTH - 1] = decval[PTR_WIDTH - 1];
				end
			endfunction
			function automatic [PTR_WIDTH - 1:0] gray2dec;
				input reg [PTR_WIDTH - 1:0] grayval;
				reg [PTR_WIDTH - 1:0] dec_tmp;
				reg [PTR_WIDTH - 1:0] dec_tmp_sub;
				reg unused_decsub_msb;
				begin
					dec_tmp = 1'sb0;
					begin : sv2v_autoblock_1
						reg signed [31:0] i;
						for (i = PTR_WIDTH - 2; i >= 0; i = i - 1)
							dec_tmp[i] = dec_tmp[i + 1] ^ grayval[i];
					end
					dec_tmp_sub = (sv2v_cast_06624(Depth) - dec_tmp) - 1'b1;
					if (grayval[PTR_WIDTH - 1]) begin
						gray2dec = dec_tmp_sub;
						gray2dec[PTR_WIDTH - 1] = 1'b1;
						unused_decsub_msb = dec_tmp_sub[PTR_WIDTH - 1];
					end
					else
						gray2dec = dec_tmp;
				end
			endfunction
			assign fifo_rptr_sync_combi = gray2dec(fifo_rptr_gray_sync);
			assign fifo_wptr_sync_combi = gray2dec(fifo_wptr_gray_sync);
			assign fifo_rptr_gray_d = dec2gray(fifo_rptr_d);
			assign fifo_wptr_gray_d = dec2gray(fifo_wptr_d);
		end
		else if (Depth == 2) begin : g_simple_gray_conversion
			assign fifo_rptr_sync_combi = {fifo_rptr_gray_sync[PTR_WIDTH - 1], ^fifo_rptr_gray_sync};
			assign fifo_wptr_sync_combi = {fifo_wptr_gray_sync[PTR_WIDTH - 1], ^fifo_wptr_gray_sync};
			assign fifo_rptr_gray_d = {fifo_rptr_d[PTR_WIDTH - 1], ^fifo_rptr_d};
			assign fifo_wptr_gray_d = {fifo_wptr_d[PTR_WIDTH - 1], ^fifo_wptr_d};
		end
		else begin : g_no_gray_conversion
			assign fifo_rptr_sync_combi = fifo_rptr_gray_sync;
			assign fifo_wptr_sync_combi = fifo_wptr_gray_sync;
			assign fifo_rptr_gray_d = fifo_rptr_d;
			assign fifo_wptr_gray_d = fifo_wptr_d;
		end
	endgenerate
endmodule
module prim_fifo_async_simple (
	clk_wr_i,
	rst_wr_ni,
	wvalid_i,
	wready_o,
	wdata_i,
	clk_rd_i,
	rst_rd_ni,
	rvalid_o,
	rready_i,
	rdata_o
);
	parameter [31:0] Width = 16;
	parameter [0:0] EnRstChks = 1'b0;
	parameter [0:0] EnRzHs = 1'b0;
	input wire clk_wr_i;
	input wire rst_wr_ni;
	input wire wvalid_i;
	output wire wready_o;
	input wire [Width - 1:0] wdata_i;
	input wire clk_rd_i;
	input wire rst_rd_ni;
	output wire rvalid_o;
	input wire rready_i;
	output wire [Width - 1:0] rdata_o;
	wire wr_en;
	wire src_req;
	wire src_ack;
	wire pending_d;
	reg pending_q;
	reg not_in_reset_q;
	assign wready_o = !pending_q && not_in_reset_q;
	assign wr_en = wvalid_i && wready_o;
	assign src_req = pending_q || wvalid_i;
	assign pending_d = (src_ack ? 1'b0 : (wr_en ? 1'b1 : pending_q));
	wire dst_req;
	wire dst_ack;
	assign rvalid_o = dst_req;
	assign dst_ack = dst_req && rready_i;
	always @(posedge clk_wr_i or negedge rst_wr_ni)
		if (!rst_wr_ni) begin
			pending_q <= 1'b0;
			not_in_reset_q <= 1'b0;
		end
		else begin
			pending_q <= pending_d;
			not_in_reset_q <= 1'b1;
		end
	prim_sync_reqack #(
		.EnRstChks(EnRstChks),
		.EnRzHs(EnRzHs)
	) u_prim_sync_reqack(
		.clk_src_i(clk_wr_i),
		.rst_src_ni(rst_wr_ni),
		.clk_dst_i(clk_rd_i),
		.rst_dst_ni(rst_rd_ni),
		.req_chk_i(1'b0),
		.src_req_i(src_req),
		.src_ack_o(src_ack),
		.dst_req_o(dst_req),
		.dst_ack_i(dst_ack)
	);
	reg [Width - 1:0] data_q;
	always @(posedge clk_wr_i)
		if (wr_en)
			data_q <= wdata_i;
	assign rdata_o = data_q;
endmodule
module prim_fifo_async_sram_adapter (
	clk_wr_i,
	rst_wr_ni,
	wvalid_i,
	wready_o,
	wdata_i,
	wdepth_o,
	clk_rd_i,
	rst_rd_ni,
	rvalid_o,
	rready_i,
	rdata_o,
	rdepth_o,
	r_full_o,
	r_notempty_o,
	w_full_o,
	w_sram_req_o,
	w_sram_gnt_i,
	w_sram_write_o,
	w_sram_addr_o,
	w_sram_wdata_o,
	w_sram_wmask_o,
	w_sram_rvalid_i,
	w_sram_rdata_i,
	w_sram_rerror_i,
	r_sram_req_o,
	r_sram_gnt_i,
	r_sram_write_o,
	r_sram_addr_o,
	r_sram_wdata_o,
	r_sram_wmask_o,
	r_sram_rvalid_i,
	r_sram_rdata_i,
	r_sram_rerror_i
);
	parameter [31:0] Width = 32;
	parameter [31:0] Depth = 16;
	parameter [31:0] SramAw = 16;
	parameter [31:0] SramDw = 32;
	parameter [SramAw - 1:0] SramBaseAddr = 'h0;
	localparam [31:0] DepthW = $clog2(Depth + 1);
	input clk_wr_i;
	input rst_wr_ni;
	input wvalid_i;
	output wire wready_o;
	input [Width - 1:0] wdata_i;
	output wire [DepthW - 1:0] wdepth_o;
	input clk_rd_i;
	input rst_rd_ni;
	output wire rvalid_o;
	input rready_i;
	output wire [Width - 1:0] rdata_o;
	output wire [DepthW - 1:0] rdepth_o;
	output wire r_full_o;
	output wire r_notempty_o;
	output wire w_full_o;
	output wire w_sram_req_o;
	input w_sram_gnt_i;
	output wire w_sram_write_o;
	output wire [SramAw - 1:0] w_sram_addr_o;
	output wire [SramDw - 1:0] w_sram_wdata_o;
	output wire [SramDw - 1:0] w_sram_wmask_o;
	input w_sram_rvalid_i;
	input [SramDw - 1:0] w_sram_rdata_i;
	input [1:0] w_sram_rerror_i;
	output reg r_sram_req_o;
	input r_sram_gnt_i;
	output wire r_sram_write_o;
	output wire [SramAw - 1:0] r_sram_addr_o;
	output wire [SramDw - 1:0] r_sram_wdata_o;
	output wire [SramDw - 1:0] r_sram_wmask_o;
	input r_sram_rvalid_i;
	input [SramDw - 1:0] r_sram_rdata_i;
	input [1:0] r_sram_rerror_i;
	localparam [31:0] PtrVW = $clog2(Depth);
	localparam [31:0] PtrW = PtrVW + 1;
	reg [PtrW - 1:0] w_wptr_q;
	wire [PtrW - 1:0] w_wptr_d;
	wire [PtrW - 1:0] w_wptr_gray_d;
	reg [PtrW - 1:0] w_wptr_gray_q;
	wire [PtrW - 1:0] r_wptr_gray;
	wire [PtrW - 1:0] r_wptr;
	wire [PtrVW - 1:0] w_wptr_v;
	wire [PtrVW - 1:0] r_wptr_v;
	wire w_wptr_p;
	wire r_wptr_p;
	reg [PtrW - 1:0] r_rptr_q;
	wire [PtrW - 1:0] r_rptr_d;
	wire [PtrW - 1:0] r_rptr_gray_d;
	reg [PtrW - 1:0] r_rptr_gray_q;
	wire [PtrW - 1:0] w_rptr_gray;
	wire [PtrW - 1:0] w_rptr;
	wire [PtrVW - 1:0] r_rptr_v;
	wire [PtrVW - 1:0] w_rptr_v;
	wire r_rptr_p;
	wire w_rptr_p;
	wire w_wptr_inc;
	wire r_rptr_inc;
	wire w_full;
	wire r_full;
	wire r_empty;
	reg stored;
	reg [Width - 1:0] rdata_q;
	wire [Width - 1:0] rdata_d;
	wire r_sram_rptr_inc;
	reg [PtrW - 1:0] r_sram_rptr;
	wire r_sramrptr_empty;
	wire rfifo_ack;
	wire rsram_ack;
	assign w_wptr_inc = wvalid_i & wready_o;
	function automatic signed [PtrW - 1:0] sv2v_cast_7A7B7_signed;
		input reg signed [PtrW - 1:0] inp;
		sv2v_cast_7A7B7_signed = inp;
	endfunction
	assign w_wptr_d = w_wptr_q + sv2v_cast_7A7B7_signed(1);
	always @(posedge clk_wr_i or negedge rst_wr_ni)
		if (!rst_wr_ni) begin
			w_wptr_q <= sv2v_cast_7A7B7_signed(0);
			w_wptr_gray_q <= sv2v_cast_7A7B7_signed(0);
		end
		else if (w_wptr_inc) begin
			w_wptr_q <= w_wptr_d;
			w_wptr_gray_q <= w_wptr_gray_d;
		end
	assign w_wptr_v = w_wptr_q[0+:PtrVW];
	assign w_wptr_p = w_wptr_q[PtrW - 1];
	function automatic [PtrW - 1:0] sv2v_cast_7A7B7;
		input reg [PtrW - 1:0] inp;
		sv2v_cast_7A7B7 = inp;
	endfunction
	function automatic [PtrW - 1:0] dec2gray;
		input reg [PtrW - 1:0] decval;
		reg [PtrW - 1:0] decval_sub;
		reg [PtrW - 1:0] decval_in;
		reg unused_decval_msb;
		begin
			decval_sub = (sv2v_cast_7A7B7(Depth) - {1'b0, decval[PtrW - 2:0]}) - 1'b1;
			decval_in = (decval[PtrW - 1] ? decval_sub : decval);
			unused_decval_msb = decval_in[PtrW - 1];
			decval_in[PtrW - 1] = 1'b0;
			dec2gray = decval_in;
			dec2gray = dec2gray ^ (decval_in >> 1);
			dec2gray[PtrW - 1] = decval[PtrW - 1];
		end
	endfunction
	assign w_wptr_gray_d = dec2gray(w_wptr_d);
	prim_flop_2sync #(.Width(PtrW)) u_sync_wptr_gray(
		.clk_i(clk_rd_i),
		.rst_ni(rst_rd_ni),
		.d_i(w_wptr_gray_q),
		.q_o(r_wptr_gray)
	);
	function automatic [PtrW - 1:0] gray2dec;
		input reg [PtrW - 1:0] grayval;
		reg [PtrW - 1:0] dec_tmp;
		reg [PtrW - 1:0] dec_tmp_sub;
		reg unused_decsub_msb;
		begin
			dec_tmp = 1'sb0;
			begin : sv2v_autoblock_1
				reg signed [31:0] i;
				for (i = PtrW - 2; i >= 0; i = i - 1)
					dec_tmp[i] = dec_tmp[i + 1] ^ grayval[i];
			end
			dec_tmp_sub = (sv2v_cast_7A7B7(Depth) - dec_tmp) - 1'b1;
			if (grayval[PtrW - 1]) begin
				gray2dec = dec_tmp_sub;
				gray2dec[PtrW - 1] = 1'b1;
				unused_decsub_msb = dec_tmp_sub[PtrW - 1];
			end
			else
				gray2dec = dec_tmp;
		end
	endfunction
	assign r_wptr = gray2dec(r_wptr_gray);
	assign r_wptr_p = r_wptr[PtrW - 1];
	assign r_wptr_v = r_wptr[0+:PtrVW];
	function automatic [DepthW - 1:0] sv2v_cast_00304;
		input reg [DepthW - 1:0] inp;
		sv2v_cast_00304 = inp;
	endfunction
	assign wdepth_o = (w_wptr_p == w_rptr_p ? sv2v_cast_00304(w_wptr_v - w_rptr_v) : sv2v_cast_00304({1'b1, w_wptr_v} - {1'b0, w_rptr_v}));
	assign r_rptr_inc = rfifo_ack;
	assign r_rptr_d = r_rptr_q + sv2v_cast_7A7B7_signed(1);
	always @(posedge clk_rd_i or negedge rst_rd_ni)
		if (!rst_rd_ni) begin
			r_rptr_q <= sv2v_cast_7A7B7_signed(0);
			r_rptr_gray_q <= sv2v_cast_7A7B7_signed(0);
		end
		else if (r_rptr_inc) begin
			r_rptr_q <= r_rptr_d;
			r_rptr_gray_q <= r_rptr_gray_d;
		end
	assign r_rptr_v = r_rptr_q[0+:PtrVW];
	assign r_rptr_p = r_rptr_q[PtrW - 1];
	assign r_rptr_gray_d = dec2gray(r_rptr_d);
	prim_flop_2sync #(.Width(PtrW)) u_sync_rptr_gray(
		.clk_i(clk_wr_i),
		.rst_ni(rst_wr_ni),
		.d_i(r_rptr_gray_q),
		.q_o(w_rptr_gray)
	);
	assign w_rptr = gray2dec(w_rptr_gray);
	assign w_rptr_p = w_rptr[PtrW - 1];
	assign w_rptr_v = w_rptr[0+:PtrVW];
	assign rdepth_o = (r_wptr_p == r_rptr_p ? sv2v_cast_00304(r_wptr_v - r_rptr_v) : sv2v_cast_00304({1'b1, r_wptr_v} - {1'b0, r_rptr_v}));
	assign r_sram_rptr_inc = rsram_ack;
	always @(posedge clk_rd_i or negedge rst_rd_ni)
		if (!rst_rd_ni)
			r_sram_rptr <= sv2v_cast_7A7B7_signed(0);
		else if (r_sram_rptr_inc)
			r_sram_rptr <= r_sram_rptr + sv2v_cast_7A7B7_signed(1);
	assign r_sramrptr_empty = r_wptr == r_sram_rptr;
	localparam [PtrW - 1:0] XorMask = {1'b1, {PtrW - 1 {1'b0}}};
	assign w_full = w_wptr_q == (w_rptr ^ XorMask);
	assign r_full = r_wptr == (r_rptr_q ^ XorMask);
	assign r_empty = r_wptr == r_rptr_q;
	wire unused_r_empty;
	assign unused_r_empty = r_empty;
	assign r_full_o = r_full;
	assign w_full_o = w_full;
	assign r_notempty_o = rvalid_o;
	assign rsram_ack = r_sram_req_o && r_sram_gnt_i;
	assign rfifo_ack = rvalid_o && rready_i;
	assign w_sram_req_o = wvalid_i && !w_full;
	assign wready_o = !w_full && w_sram_gnt_i;
	assign w_sram_write_o = 1'b1;
	function automatic [SramAw - 1:0] sv2v_cast_576AD;
		input reg [SramAw - 1:0] inp;
		sv2v_cast_576AD = inp;
	endfunction
	assign w_sram_addr_o = SramBaseAddr + sv2v_cast_576AD(w_wptr_v);
	function automatic [SramDw - 1:0] sv2v_cast_24298;
		input reg [SramDw - 1:0] inp;
		sv2v_cast_24298 = inp;
	endfunction
	assign w_sram_wdata_o = sv2v_cast_24298(wdata_i);
	assign w_sram_wmask_o = sv2v_cast_24298({Width {1'b1}});
	wire unused_w_sram;
	assign unused_w_sram = ^{w_sram_rvalid_i, w_sram_rdata_i, w_sram_rerror_i};
	always @(*) begin : r_sram_req
		r_sram_req_o = 1'b0;
		if (stored)
			r_sram_req_o = !r_sramrptr_empty && rfifo_ack;
		else
			r_sram_req_o = !r_sramrptr_empty && !(r_sram_rvalid_i ^ rfifo_ack);
	end
	assign rvalid_o = stored || r_sram_rvalid_i;
	assign r_sram_write_o = 1'b0;
	assign r_sram_wdata_o = 1'sb0;
	assign r_sram_wmask_o = 1'sb0;
	assign r_sram_addr_o = SramBaseAddr + sv2v_cast_576AD(r_sram_rptr[0+:PtrVW]);
	function automatic signed [Width - 1:0] sv2v_cast_92C3D_signed;
		input reg signed [Width - 1:0] inp;
		sv2v_cast_92C3D_signed = inp;
	endfunction
	assign rdata_d = (r_sram_rvalid_i ? r_sram_rdata_i[0+:Width] : sv2v_cast_92C3D_signed(0));
	assign rdata_o = (stored ? rdata_q : rdata_d);
	wire unused_rsram;
	assign unused_rsram = ^{r_sram_rerror_i};
	generate
		if (Width < SramDw) begin : g_unused_rdata
			wire unused_rdata;
			assign unused_rdata = ^r_sram_rdata_i[SramDw - 1:Width];
		end
	endgenerate
	wire store_en;
	assign store_en = r_sram_rvalid_i && !(stored ^ rfifo_ack);
	always @(posedge clk_rd_i or negedge rst_rd_ni)
		if (!rst_rd_ni) begin
			stored <= 1'b0;
			rdata_q <= sv2v_cast_92C3D_signed(0);
		end
		else if (store_en) begin
			stored <= 1'b1;
			rdata_q <= rdata_d;
		end
		else if (!r_sram_rvalid_i && rfifo_ack) begin
			stored <= 1'b0;
			rdata_q <= sv2v_cast_92C3D_signed(0);
		end
endmodule
module prim_fifo_sync (
	clk_i,
	rst_ni,
	clr_i,
	wvalid_i,
	wready_o,
	wdata_i,
	rvalid_o,
	rready_i,
	rdata_o,
	full_o,
	depth_o,
	err_o
);
	parameter [31:0] Width = 16;
	parameter [0:0] Pass = 1'b1;
	parameter [31:0] Depth = 4;
	parameter [0:0] OutputZeroIfEmpty = 1'b1;
	parameter [0:0] Secure = 1'b0;
	function automatic integer prim_util_pkg_vbits;
		input integer value;
		prim_util_pkg_vbits = (value == 1 ? 1 : $clog2(value));
	endfunction
	localparam signed [31:0] DepthW = prim_util_pkg_vbits(Depth + 1);
	input clk_i;
	input rst_ni;
	input clr_i;
	input wvalid_i;
	output wire wready_o;
	input [Width - 1:0] wdata_i;
	output wire rvalid_o;
	input rready_i;
	output wire [Width - 1:0] rdata_o;
	output wire full_o;
	output wire [DepthW - 1:0] depth_o;
	output wire err_o;
	function automatic [DepthW - 1:0] sv2v_cast_00304;
		input reg [DepthW - 1:0] inp;
		sv2v_cast_00304 = inp;
	endfunction
	generate
		if (Depth == 0) begin : gen_passthru_fifo
			assign depth_o = 1'b0;
			assign rvalid_o = wvalid_i;
			assign rdata_o = wdata_i;
			assign wready_o = rready_i;
			assign full_o = rready_i;
			wire unused_clr;
			assign unused_clr = clr_i;
			assign err_o = 1'b0;
		end
		else begin : gen_normal_fifo
			localparam [31:0] PTRV_W = prim_util_pkg_vbits(Depth);
			localparam [31:0] PTR_WIDTH = PTRV_W + 1;
			wire [PTR_WIDTH - 1:0] fifo_wptr;
			wire [PTR_WIDTH - 1:0] fifo_rptr;
			wire fifo_incr_wptr;
			wire fifo_incr_rptr;
			wire fifo_empty;
			reg under_rst;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					under_rst <= 1'b1;
				else if (under_rst)
					under_rst <= ~under_rst;
			wire full;
			wire empty;
			wire wptr_msb;
			wire rptr_msb;
			wire [PTRV_W - 1:0] wptr_value;
			wire [PTRV_W - 1:0] rptr_value;
			assign wptr_msb = fifo_wptr[PTR_WIDTH - 1];
			assign rptr_msb = fifo_rptr[PTR_WIDTH - 1];
			assign wptr_value = fifo_wptr[0+:PTRV_W];
			assign rptr_value = fifo_rptr[0+:PTRV_W];
			assign depth_o = (full ? sv2v_cast_00304(Depth) : (wptr_msb == rptr_msb ? sv2v_cast_00304(wptr_value) - sv2v_cast_00304(rptr_value) : (sv2v_cast_00304(Depth) - sv2v_cast_00304(rptr_value)) + sv2v_cast_00304(wptr_value)));
			assign fifo_incr_wptr = (wvalid_i & wready_o) & ~under_rst;
			assign fifo_incr_rptr = (rvalid_o & rready_i) & ~under_rst;
			assign wready_o = ~full & ~under_rst;
			assign full_o = full;
			assign rvalid_o = ~empty & ~under_rst;
			prim_fifo_sync_cnt #(
				.Width(PTR_WIDTH),
				.Depth(Depth),
				.Secure(Secure)
			) u_fifo_cnt(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.clr_i(clr_i),
				.incr_wptr_i(fifo_incr_wptr),
				.incr_rptr_i(fifo_incr_rptr),
				.wptr_o(fifo_wptr),
				.rptr_o(fifo_rptr),
				.err_o(err_o)
			);
			assign full = fifo_wptr == (fifo_rptr ^ {1'b1, {PTR_WIDTH - 1 {1'b0}}});
			assign fifo_empty = fifo_wptr == fifo_rptr;
			reg [(Depth * Width) - 1:0] storage;
			wire [Width - 1:0] storage_rdata;
			if (Depth == 1) begin : gen_depth_eq1
				assign storage_rdata = storage[0+:Width];
				always @(posedge clk_i)
					if (fifo_incr_wptr)
						storage[0+:Width] <= wdata_i;
			end
			else begin : gen_depth_gt1
				assign storage_rdata = storage[fifo_rptr[PTR_WIDTH - 2:0] * Width+:Width];
				always @(posedge clk_i)
					if (fifo_incr_wptr)
						storage[fifo_wptr[PTR_WIDTH - 2:0] * Width+:Width] <= wdata_i;
			end
			wire [Width - 1:0] rdata_int;
			if (Pass == 1'b1) begin : gen_pass
				assign rdata_int = (fifo_empty && wvalid_i ? wdata_i : storage_rdata);
				assign empty = fifo_empty & ~wvalid_i;
			end
			else begin : gen_nopass
				assign rdata_int = storage_rdata;
				assign empty = fifo_empty;
			end
			if (OutputZeroIfEmpty == 1'b1) begin : gen_output_zero
				assign rdata_o = (empty ? 'b0 : rdata_int);
			end
			else begin : gen_no_output_zero
				assign rdata_o = rdata_int;
			end
		end
	endgenerate
endmodule
module prim_fifo_sync_cnt (
	clk_i,
	rst_ni,
	clr_i,
	incr_wptr_i,
	incr_rptr_i,
	wptr_o,
	rptr_o,
	err_o
);
	parameter signed [31:0] Depth = 4;
	parameter signed [31:0] Width = 16;
	parameter [0:0] Secure = 1'b0;
	input clk_i;
	input rst_ni;
	input clr_i;
	input incr_wptr_i;
	input incr_rptr_i;
	output reg [Width - 1:0] wptr_o;
	output reg [Width - 1:0] rptr_o;
	output wire err_o;
	wire wptr_wrap;
	wire [Width - 1:0] wptr_wrap_cnt;
	wire rptr_wrap;
	wire [Width - 1:0] rptr_wrap_cnt;
	function automatic signed [((Width - 2) >= 0 ? Width - 1 : 3 - Width) - 1:0] sv2v_cast_582D5_signed;
		input reg signed [((Width - 2) >= 0 ? Width - 1 : 3 - Width) - 1:0] inp;
		sv2v_cast_582D5_signed = inp;
	endfunction
	assign wptr_wrap = incr_wptr_i & (wptr_o[Width - 2:0] == $unsigned(sv2v_cast_582D5_signed(Depth - 1)));
	assign rptr_wrap = incr_rptr_i & (rptr_o[Width - 2:0] == $unsigned(sv2v_cast_582D5_signed(Depth - 1)));
	assign wptr_wrap_cnt = {~wptr_o[Width - 1], {Width - 1 {1'b0}}};
	assign rptr_wrap_cnt = {~rptr_o[Width - 1], {Width - 1 {1'b0}}};
	function automatic [Width - 1:0] sv2v_cast_92C3D;
		input reg [Width - 1:0] inp;
		sv2v_cast_92C3D = inp;
	endfunction
	generate
		if (Secure) begin : gen_secure_ptrs
			wire wptr_err;
			wire [Width:1] sv2v_tmp_u_wptr_cnt_o;
			always @(*) wptr_o = sv2v_tmp_u_wptr_cnt_o;
			prim_count #(.Width(Width)) u_wptr(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.clr_i(clr_i),
				.set_i(wptr_wrap),
				.set_cnt_i(wptr_wrap_cnt),
				.incr_en_i(incr_wptr_i),
				.decr_en_i(1'b0),
				.step_i(sv2v_cast_92C3D(1'b1)),
				.cnt_o(sv2v_tmp_u_wptr_cnt_o),
				.err_o(wptr_err)
			);
			wire rptr_err;
			wire [Width:1] sv2v_tmp_u_rptr_cnt_o;
			always @(*) rptr_o = sv2v_tmp_u_rptr_cnt_o;
			prim_count #(.Width(Width)) u_rptr(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.clr_i(clr_i),
				.set_i(rptr_wrap),
				.set_cnt_i(rptr_wrap_cnt),
				.incr_en_i(incr_rptr_i),
				.decr_en_i(1'b0),
				.step_i(sv2v_cast_92C3D(1'b1)),
				.cnt_o(sv2v_tmp_u_rptr_cnt_o),
				.err_o(rptr_err)
			);
			assign err_o = wptr_err | rptr_err;
		end
		else begin : gen_normal_ptrs
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					wptr_o <= {Width {1'b0}};
				else if (clr_i)
					wptr_o <= {Width {1'b0}};
				else if (wptr_wrap)
					wptr_o <= wptr_wrap_cnt;
				else if (incr_wptr_i)
					wptr_o <= wptr_o + {{Width - 1 {1'b0}}, 1'b1};
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					rptr_o <= {Width {1'b0}};
				else if (clr_i)
					rptr_o <= {Width {1'b0}};
				else if (rptr_wrap)
					rptr_o <= rptr_wrap_cnt;
				else if (incr_rptr_i)
					rptr_o <= rptr_o + {{Width - 1 {1'b0}}, 1'b1};
			assign err_o = 1'sb0;
		end
	endgenerate
endmodule
module prim_filter (
	clk_i,
	rst_ni,
	enable_i,
	filter_i,
	filter_o
);
	parameter [0:0] AsyncOn = 0;
	parameter [31:0] Cycles = 4;
	input clk_i;
	input rst_ni;
	input enable_i;
	input filter_i;
	output wire filter_o;
	reg [Cycles - 1:0] stored_vector_q;
	wire [Cycles - 1:0] stored_vector_d;
	reg stored_value_q;
	wire update_stored_value;
	wire unused_stored_vector_q_msb;
	wire filter_synced;
	generate
		if (AsyncOn) begin : gen_async
			prim_flop_2sync #(.Width(1)) prim_flop_2sync(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(filter_i),
				.q_o(filter_synced)
			);
		end
		else begin : gen_sync
			assign filter_synced = filter_i;
		end
	endgenerate
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			stored_value_q <= 1'b0;
		else if (update_stored_value)
			stored_value_q <= filter_synced;
	assign stored_vector_d = {stored_vector_q[Cycles - 2:0], filter_synced};
	assign unused_stored_vector_q_msb = stored_vector_q[Cycles - 1];
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			stored_vector_q <= 1'sb0;
		else
			stored_vector_q <= stored_vector_d;
	assign update_stored_value = (stored_vector_d == {Cycles {1'b0}}) | (stored_vector_d == {Cycles {1'b1}});
	assign filter_o = (enable_i ? stored_value_q : filter_synced);
endmodule
module prim_filter_ctr (
	clk_i,
	rst_ni,
	enable_i,
	filter_i,
	thresh_i,
	filter_o
);
	parameter [0:0] AsyncOn = 0;
	parameter [31:0] CntWidth = 2;
	input clk_i;
	input rst_ni;
	input enable_i;
	input filter_i;
	input [CntWidth - 1:0] thresh_i;
	output wire filter_o;
	reg [CntWidth - 1:0] diff_ctr_q;
	wire [CntWidth - 1:0] diff_ctr_d;
	reg filter_q;
	reg stored_value_q;
	wire update_stored_value;
	wire filter_synced;
	generate
		if (AsyncOn) begin : gen_async
			prim_flop_2sync #(.Width(1)) prim_flop_2sync(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(filter_i),
				.q_o(filter_synced)
			);
		end
		else begin : gen_sync
			assign filter_synced = filter_i;
		end
	endgenerate
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			filter_q <= 1'b0;
		else
			filter_q <= filter_synced;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			stored_value_q <= 1'b0;
		else if (update_stored_value)
			stored_value_q <= filter_synced;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			diff_ctr_q <= 1'sb0;
		else
			diff_ctr_q <= diff_ctr_d;
	assign update_stored_value = diff_ctr_d == thresh_i;
	assign diff_ctr_d = (filter_synced != filter_q ? {CntWidth {1'sb0}} : (diff_ctr_q >= thresh_i ? thresh_i : diff_ctr_q + 1'b1));
	assign filter_o = (enable_i ? stored_value_q : filter_synced);
endmodule
module prim_flop (
	clk_i,
	rst_ni,
	d_i,
	q_o
);
	parameter signed [31:0] Width = 1;
	parameter [Width - 1:0] ResetValue = 0;
	input clk_i;
	input rst_ni;
	input [Width - 1:0] d_i;
	output wire [Width - 1:0] q_o;
	parameter integer Impl = 32'sd0;
	generate
		if (Impl == 32'sd2) begin : gen_xilinx
			prim_xilinx_flop #(
				.ResetValue(ResetValue),
				.Width(Width)
			) u_impl_xilinx(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(d_i),
				.q_o(q_o)
			);
		end
		else begin : gen_generic
			prim_generic_flop #(
				.ResetValue(ResetValue),
				.Width(Width)
			) u_impl_generic(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(d_i),
				.q_o(q_o)
			);
		end
	endgenerate
endmodule
module prim_flop_2sync (
	clk_i,
	rst_ni,
	d_i,
	q_o
);
	parameter signed [31:0] Width = 16;
	parameter [Width - 1:0] ResetValue = 1'sb0;
	parameter [0:0] EnablePrimCdcRand = 1;
	input clk_i;
	input rst_ni;
	input [Width - 1:0] d_i;
	output wire [Width - 1:0] q_o;
	reg [Width - 1:0] d_o;
	wire [Width - 1:0] intq;
	wire unused_sig;
	assign unused_sig = EnablePrimCdcRand;
	always @(*) d_o = d_i;
	prim_flop #(
		.Width(Width),
		.ResetValue(ResetValue)
	) u_sync_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(d_o),
		.q_o(intq)
	);
	prim_flop #(
		.Width(Width),
		.ResetValue(ResetValue)
	) u_sync_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(intq),
		.q_o(q_o)
	);
endmodule
module prim_flop_en (
	clk_i,
	rst_ni,
	en_i,
	d_i,
	q_o
);
	parameter signed [31:0] Width = 1;
	parameter [0:0] EnSecBuf = 0;
	parameter [Width - 1:0] ResetValue = 0;
	input clk_i;
	input rst_ni;
	input en_i;
	input [Width - 1:0] d_i;
	output wire [Width - 1:0] q_o;
	parameter integer Impl = 32'sd0;
	generate
		if (Impl == 32'sd2) begin : gen_xilinx
			prim_xilinx_flop_en #(
				.EnSecBuf(EnSecBuf),
				.ResetValue(ResetValue),
				.Width(Width)
			) u_impl_xilinx(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.en_i(en_i),
				.d_i(d_i),
				.q_o(q_o)
			);
		end
		else begin : gen_generic
			prim_generic_flop_en #(
				.EnSecBuf(EnSecBuf),
				.ResetValue(ResetValue),
				.Width(Width)
			) u_impl_generic(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.en_i(en_i),
				.d_i(d_i),
				.q_o(q_o)
			);
		end
	endgenerate
endmodule
module prim_gate_gen (
	clk_i,
	rst_ni,
	valid_i,
	data_i,
	data_o,
	valid_o
);
	parameter signed [31:0] DataWidth = 32;
	parameter signed [31:0] NumGates = 1000;
	input clk_i;
	input rst_ni;
	input valid_i;
	input [DataWidth - 1:0] data_i;
	output wire [DataWidth - 1:0] data_o;
	output wire valid_o;
	localparam signed [31:0] NumInnerRounds = 2;
	localparam signed [31:0] GatesPerRound = DataWidth * 14;
	localparam signed [31:0] NumOuterRounds = (NumGates + (GatesPerRound / 2)) / GatesPerRound;
	wire [(NumOuterRounds * DataWidth) - 1:0] regs_d;
	reg [(NumOuterRounds * DataWidth) - 1:0] regs_q;
	wire [NumOuterRounds - 1:0] valid_d;
	reg [NumOuterRounds - 1:0] valid_q;
	genvar k;
	localparam [63:0] prim_cipher_pkg_PRINCE_SBOX4 = 64'h4d5e087619ca23fb;
	function automatic [7:0] prim_cipher_pkg_sbox4_8bit;
		input reg [7:0] state_in;
		input reg [63:0] sbox4;
		reg [7:0] state_out;
		begin
			begin : sv2v_autoblock_1
				reg signed [31:0] k;
				for (k = 0; k < 2; k = k + 1)
					state_out[k * 4+:4] = sbox4[state_in[k * 4+:4] * 4+:4];
			end
			prim_cipher_pkg_sbox4_8bit = state_out;
		end
	endfunction
	function automatic [31:0] prim_cipher_pkg_sbox4_32bit;
		input reg [31:0] state_in;
		input reg [63:0] sbox4;
		reg [31:0] state_out;
		begin
			begin : sv2v_autoblock_2
				reg signed [31:0] k;
				for (k = 0; k < 4; k = k + 1)
					state_out[k * 8+:8] = prim_cipher_pkg_sbox4_8bit(state_in[k * 8+:8], sbox4);
			end
			prim_cipher_pkg_sbox4_32bit = state_out;
		end
	endfunction
	generate
		for (k = 0; k < NumOuterRounds; k = k + 1) begin : gen_outer_round
			wire [(3 * DataWidth) - 1:0] inner_data;
			if (k == 0) begin : gen_first
				assign inner_data[0+:DataWidth] = data_i;
				assign valid_d[0] = valid_i;
			end
			else begin : gen_others
				assign inner_data[0+:DataWidth] = regs_q[(k - 1) * DataWidth+:DataWidth];
				assign valid_d[k] = valid_q[k - 1];
			end
			genvar l;
			for (l = 0; l < NumInnerRounds; l = l + 1) begin : gen_inner
				assign inner_data[(l + 1) * DataWidth+:DataWidth] = prim_cipher_pkg_sbox4_32bit({inner_data[(l * DataWidth) + 1-:2], inner_data[(l * DataWidth) + ((DataWidth - 1) >= 2 ? DataWidth - 1 : ((DataWidth - 1) + ((DataWidth - 1) >= 2 ? DataWidth - 2 : 4 - DataWidth)) - 1)-:((DataWidth - 1) >= 2 ? DataWidth - 2 : 4 - DataWidth)]}, prim_cipher_pkg_PRINCE_SBOX4);
			end
			assign regs_d[k * DataWidth+:DataWidth] = inner_data[NumInnerRounds * DataWidth+:DataWidth];
		end
	endgenerate
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		if (!rst_ni) begin
			regs_q <= 1'sb0;
			valid_q <= 1'sb0;
		end
		else begin
			valid_q <= valid_d;
			begin : sv2v_autoblock_3
				reg signed [31:0] k;
				for (k = 0; k < NumOuterRounds; k = k + 1)
					if (valid_d[k])
						regs_q[k * DataWidth+:DataWidth] <= regs_d[k * DataWidth+:DataWidth];
			end
		end
	end
	assign data_o = regs_q[(NumOuterRounds - 1) * DataWidth+:DataWidth];
	assign valid_o = valid_q[NumOuterRounds - 1];
endmodule
module prim_generic_and2 (
	in0_i,
	in1_i,
	out_o
);
	parameter signed [31:0] Width = 1;
	input [Width - 1:0] in0_i;
	input [Width - 1:0] in1_i;
	output wire [Width - 1:0] out_o;
	assign out_o = in0_i & in1_i;
endmodule
module prim_generic_buf (
	in_i,
	out_o
);
	parameter signed [31:0] Width = 1;
	input [Width - 1:0] in_i;
	output wire [Width - 1:0] out_o;
	wire [Width - 1:0] inv;
	assign inv = ~in_i;
	assign out_o = ~inv;
endmodule
module prim_generic_clock_gating (
	clk_i,
	en_i,
	test_en_i,
	clk_o
);
	parameter [0:0] NoFpgaGate = 1'b0;
	parameter [0:0] FpgaBufGlobal = 1'b1;
	input clk_i;
	input en_i;
	input test_en_i;
	output wire clk_o;
	reg en_latch;
	always @(*)
		if (!clk_i)
			en_latch = en_i | test_en_i;
	assign clk_o = en_latch & clk_i;
endmodule
module prim_generic_clock_mux2 (
	clk0_i,
	clk1_i,
	sel_i,
	clk_o
);
	parameter [0:0] NoFpgaBufG = 1'b0;
	input clk0_i;
	input clk1_i;
	input sel_i;
	output wire clk_o;
	assign clk_o = (sel_i & clk1_i) | (~sel_i & clk0_i);
endmodule
module prim_generic_flop (
	clk_i,
	rst_ni,
	d_i,
	q_o
);
	parameter signed [31:0] Width = 1;
	parameter [Width - 1:0] ResetValue = 0;
	input clk_i;
	input rst_ni;
	input [Width - 1:0] d_i;
	output reg [Width - 1:0] q_o;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			q_o <= ResetValue;
		else
			q_o <= d_i;
endmodule
module prim_generic_flop_en (
	clk_i,
	rst_ni,
	en_i,
	d_i,
	q_o
);
	parameter signed [31:0] Width = 1;
	parameter [0:0] EnSecBuf = 0;
	parameter [Width - 1:0] ResetValue = 0;
	input clk_i;
	input rst_ni;
	input en_i;
	input [Width - 1:0] d_i;
	output reg [Width - 1:0] q_o;
	wire en;
	generate
		if (EnSecBuf) begin : gen_en_sec_buf
			prim_sec_anchor_buf #(.Width(1)) u_en_buf(
				.in_i(en_i),
				.out_o(en)
			);
		end
		else begin : gen_en_no_sec_buf
			assign en = en_i;
		end
	endgenerate
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			q_o <= ResetValue;
		else if (en)
			q_o <= d_i;
endmodule
module prim_generic_ram_1p (
	clk_i,
	req_i,
	write_i,
	addr_i,
	wdata_i,
	wmask_i,
	rdata_o,
	cfg_i
);
	parameter signed [31:0] Width = 32;
	parameter signed [31:0] Depth = 128;
	parameter signed [31:0] DataBitsPerMask = 1;
	parameter MemInitFile = "";
	localparam signed [31:0] Aw = $clog2(Depth);
	input wire clk_i;
	input wire req_i;
	input wire write_i;
	input wire [Aw - 1:0] addr_i;
	input wire [Width - 1:0] wdata_i;
	input wire [Width - 1:0] wmask_i;
	output reg [Width - 1:0] rdata_o;
	input wire [9:0] cfg_i;
	wire unused_cfg;
	assign unused_cfg = ^cfg_i;
	localparam signed [31:0] MaskWidth = Width / DataBitsPerMask;
	reg [Width - 1:0] mem [0:Depth - 1];
	wire [MaskWidth - 1:0] wmask;
	genvar k;
	generate
		for (k = 0; k < MaskWidth; k = k + 1) begin : gen_wmask
			assign wmask[k] = &wmask_i[k * DataBitsPerMask+:DataBitsPerMask];
		end
	endgenerate
	always @(posedge clk_i)
		if (req_i)
			if (write_i) begin : sv2v_autoblock_1
				reg signed [31:0] i;
				for (i = 0; i < MaskWidth; i = i + 1)
					if (wmask[i])
						mem[addr_i][i * DataBitsPerMask+:DataBitsPerMask] <= wdata_i[i * DataBitsPerMask+:DataBitsPerMask];
			end
			else
				rdata_o <= mem[addr_i];
	initial begin : sv2v_autoblock_2
		reg show_mem_paths;
		if (MemInitFile != "") begin : gen_meminit
			$display("Initializing memory %m from file '%s'.", MemInitFile);
			$readmemh(MemInitFile, mem);
		end
	end
endmodule
module prim_generic_xnor2 (
	in0_i,
	in1_i,
	out_o
);
	parameter signed [31:0] Width = 1;
	input [Width - 1:0] in0_i;
	input [Width - 1:0] in1_i;
	output wire [Width - 1:0] out_o;
	assign out_o = !(in0_i ^ in1_i);
endmodule
module prim_generic_xor2 (
	in0_i,
	in1_i,
	out_o
);
	parameter signed [31:0] Width = 1;
	input [Width - 1:0] in0_i;
	input [Width - 1:0] in1_i;
	output wire [Width - 1:0] out_o;
	assign out_o = in0_i ^ in1_i;
endmodule
module prim_intr_hw (
	clk_i,
	rst_ni,
	event_intr_i,
	reg2hw_intr_enable_q_i,
	reg2hw_intr_test_q_i,
	reg2hw_intr_test_qe_i,
	reg2hw_intr_state_q_i,
	hw2reg_intr_state_de_o,
	hw2reg_intr_state_d_o,
	intr_o
);
	parameter [31:0] Width = 1;
	parameter [0:0] FlopOutput = 1;
	parameter IntrT = "Event";
	input clk_i;
	input rst_ni;
	input [Width - 1:0] event_intr_i;
	input [Width - 1:0] reg2hw_intr_enable_q_i;
	input [Width - 1:0] reg2hw_intr_test_q_i;
	input reg2hw_intr_test_qe_i;
	input [Width - 1:0] reg2hw_intr_state_q_i;
	output wire hw2reg_intr_state_de_o;
	output wire [Width - 1:0] hw2reg_intr_state_d_o;
	output reg [Width - 1:0] intr_o;
	wire [Width - 1:0] status;
	generate
		if (IntrT == "Event") begin : g_intr_event
			wire [Width - 1:0] new_event;
			assign new_event = ({Width {reg2hw_intr_test_qe_i}} & reg2hw_intr_test_q_i) | event_intr_i;
			assign hw2reg_intr_state_de_o = |new_event;
			assign hw2reg_intr_state_d_o = new_event | reg2hw_intr_state_q_i;
			assign status = reg2hw_intr_state_q_i;
		end
		else if (IntrT == "Status") begin : g_intr_status
			reg [Width - 1:0] test_q;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					test_q <= 1'sb0;
				else if (reg2hw_intr_test_qe_i)
					test_q <= reg2hw_intr_test_q_i;
			assign hw2reg_intr_state_de_o = 1'b1;
			assign hw2reg_intr_state_d_o = event_intr_i | test_q;
			assign status = event_intr_i | test_q;
			wire unused_reg2hw;
			assign unused_reg2hw = ^reg2hw_intr_state_q_i;
		end
		if (FlopOutput == 1) begin : gen_flop_intr_output
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					intr_o <= 1'sb0;
				else
					intr_o <= status & reg2hw_intr_enable_q_i;
		end
		else begin : gen_intr_passthrough_output
			wire unused_clk;
			wire unused_rst_n;
			assign unused_clk = clk_i;
			assign unused_rst_n = rst_ni;
			wire [Width:1] sv2v_tmp_EDC5D;
			assign sv2v_tmp_EDC5D = reg2hw_intr_state_q_i & reg2hw_intr_enable_q_i;
			always @(*) intr_o = sv2v_tmp_EDC5D;
		end
	endgenerate
endmodule
module prim_keccak (
	rnd_i,
	s_i,
	s_o
);
	parameter signed [31:0] Width = 1600;
	localparam signed [31:0] W = Width / 25;
	localparam signed [31:0] L = $clog2(W);
	localparam signed [31:0] MaxRound = 12 + (2 * L);
	localparam signed [31:0] RndW = $clog2(MaxRound + 1);
	input [RndW - 1:0] rnd_i;
	input [Width - 1:0] s_i;
	output wire [Width - 1:0] s_o;
	wire [(25 * W) - 1:0] state_in;
	wire [(25 * W) - 1:0] keccak_f;
	wire [(25 * W) - 1:0] theta_data;
	wire [(25 * W) - 1:0] rho_data;
	wire [(25 * W) - 1:0] pi_data;
	wire [(25 * W) - 1:0] chi_data;
	wire [(25 * W) - 1:0] iota_data;
	function automatic [(25 * W) - 1:0] bitarray_to_box;
		input reg [Width - 1:0] s_in;
		reg [(25 * W) - 1:0] box;
		begin
			begin : sv2v_autoblock_1
				reg signed [31:0] y;
				for (y = 0; y < 5; y = y + 1)
					begin : sv2v_autoblock_2
						reg signed [31:0] x;
						for (x = 0; x < 5; x = x + 1)
							begin : sv2v_autoblock_3
								reg signed [31:0] z;
								for (z = 0; z < W; z = z + 1)
									box[(((x * 5) + y) * W) + z] = s_in[(W * ((5 * y) + x)) + z];
							end
					end
			end
			bitarray_to_box = box;
		end
	endfunction
	assign state_in = bitarray_to_box(s_i);
	function automatic [(25 * W) - 1:0] theta;
		input reg [(25 * W) - 1:0] state;
		reg [(5 * W) - 1:0] c;
		reg [(5 * W) - 1:0] d;
		reg [(25 * W) - 1:0] result;
		begin
			begin : sv2v_autoblock_4
				reg signed [31:0] x;
				for (x = 0; x < 5; x = x + 1)
					begin : sv2v_autoblock_5
						reg signed [31:0] z;
						for (z = 0; z < W; z = z + 1)
							c[(x * W) + z] = (((state[((x * 5) * W) + z] ^ state[(((x * 5) + 1) * W) + z]) ^ state[(((x * 5) + 2) * W) + z]) ^ state[(((x * 5) + 3) * W) + z]) ^ state[(((x * 5) + 4) * W) + z];
					end
			end
			begin : sv2v_autoblock_6
				reg signed [31:0] x;
				for (x = 0; x < 5; x = x + 1)
					begin : sv2v_autoblock_7
						reg signed [31:0] index_x1;
						reg signed [31:0] index_x2;
						index_x1 = (x == 0 ? 4 : x - 1);
						index_x2 = (x == 4 ? 0 : x + 1);
						begin : sv2v_autoblock_8
							reg signed [31:0] z;
							for (z = 0; z < W; z = z + 1)
								begin : sv2v_autoblock_9
									reg signed [31:0] index_z;
									index_z = (z == 0 ? W - 1 : z - 1);
									d[(x * W) + z] = c[(index_x1 * W) + z] ^ c[(index_x2 * W) + index_z];
								end
						end
					end
			end
			begin : sv2v_autoblock_10
				reg signed [31:0] x;
				for (x = 0; x < 5; x = x + 1)
					begin : sv2v_autoblock_11
						reg signed [31:0] y;
						for (y = 0; y < 5; y = y + 1)
							begin : sv2v_autoblock_12
								reg signed [31:0] z;
								for (z = 0; z < W; z = z + 1)
									result[(((x * 5) + y) * W) + z] = state[(((x * 5) + y) * W) + z] ^ d[(x * W) + z];
							end
					end
			end
			theta = result;
		end
	endfunction
	assign theta_data = theta(state_in);
	localparam signed [799:0] PiRotate = 800'h30000000100000004000000020000000100000004000000020000000000000003000000020000000000000003000000010000000400000003000000010000000400000002000000000000000400000002000000000000000300000001;
	function automatic [(25 * W) - 1:0] pi;
		input reg [(25 * W) - 1:0] state;
		reg [(25 * W) - 1:0] result;
		begin
			begin : sv2v_autoblock_13
				reg signed [31:0] x;
				for (x = 0; x < 5; x = x + 1)
					begin : sv2v_autoblock_14
						reg signed [31:0] y;
						for (y = 0; y < 5; y = y + 1)
							begin : sv2v_autoblock_15
								reg signed [31:0] index_x;
								result[(((x * 5) + y) * W) + (W - 1)-:W] = state[(((PiRotate[(((4 - x) * 5) + (4 - y)) * 32+:32] * 5) + x) * W) + (W - 1)-:W];
							end
					end
			end
			pi = result;
		end
	endfunction
	assign pi_data = pi(rho_data);
	function automatic [(25 * W) - 1:0] chi;
		input reg [(25 * W) - 1:0] state;
		reg [(25 * W) - 1:0] result;
		begin
			begin : sv2v_autoblock_16
				reg signed [31:0] x;
				for (x = 0; x < 5; x = x + 1)
					begin : sv2v_autoblock_17
						reg signed [31:0] index_x1;
						reg signed [31:0] index_x2;
						index_x1 = (x == 4 ? 0 : x + 1);
						index_x2 = (x >= 3 ? x - 3 : x + 2);
						begin : sv2v_autoblock_18
							reg signed [31:0] y;
							for (y = 0; y < 5; y = y + 1)
								begin : sv2v_autoblock_19
									reg signed [31:0] z;
									for (z = 0; z < W; z = z + 1)
										result[(((x * 5) + y) * W) + z] = state[(((x * 5) + y) * W) + z] ^ (~state[(((index_x1 * 5) + y) * W) + z] & state[(((index_x2 * 5) + y) * W) + z]);
								end
						end
					end
			end
			chi = result;
		end
	endfunction
	assign chi_data = chi(pi_data);
	localparam [1535:0] RC = 1536'h10000000000008082800000000000808a8000000080008000000000000000808b000000008000000180000000800080818000000000008009000000000000008a00000000000000880000000080008009000000008000000a000000008000808b800000000000008b8000000000008089800000000000800380000000000080028000000000000080000000000000800a800000008000000a8000000080008081800000000000808000000000800000018000000080008008;
	function automatic [(25 * W) - 1:0] iota;
		input reg [(25 * W) - 1:0] state;
		input reg [RndW - 1:0] rnd;
		reg [(25 * W) - 1:0] result;
		begin
			result = state;
			result[W - 1-:W] = state[W - 1-:W] ^ RC[((23 - rnd) * 64) + (W - 1)-:W];
			iota = result;
		end
	endfunction
	assign iota_data = iota(chi_data, rnd_i);
	assign keccak_f = iota_data;
	function automatic [Width - 1:0] box_to_bitarray;
		input reg [(25 * W) - 1:0] state;
		reg [Width - 1:0] bitarray;
		begin
			begin : sv2v_autoblock_20
				reg signed [31:0] y;
				for (y = 0; y < 5; y = y + 1)
					begin : sv2v_autoblock_21
						reg signed [31:0] x;
						for (x = 0; x < 5; x = x + 1)
							begin : sv2v_autoblock_22
								reg signed [31:0] z;
								for (z = 0; z < W; z = z + 1)
									bitarray[(W * ((5 * y) + x)) + z] = state[(((x * 5) + y) * W) + z];
							end
					end
			end
			box_to_bitarray = bitarray;
		end
	endfunction
	assign s_o = box_to_bitarray(keccak_f);
	localparam signed [799:0] RhoOffset = 800'h240000000300000069000000d2000000010000012c0000000a0000002d00000042000000be00000006000000ab0000000f000000fd0000001c000000370000009900000015000000780000005b00000114000000e7000000880000004e;
	genvar x;
	generate
		for (x = 0; x < 5; x = x + 1) begin : gen_rho_x
			genvar y;
			for (y = 0; y < 5; y = y + 1) begin : gen_rho_y
				localparam signed [31:0] Offset = RhoOffset[(((4 - x) * 5) + (4 - y)) * 32+:32] % W;
				localparam signed [31:0] ShiftAmt = W - Offset;
				if (Offset == 0) begin : gen_offset0
					assign rho_data[(((x * 5) + y) * W) + (W - 1)-:W] = theta_data[(((x * 5) + y) * W) + (W - 1)-:W];
				end
				else begin : gen_others
					assign rho_data[(((x * 5) + y) * W) + (W - 1)-:W] = {theta_data[((x * 5) + y) * W+:ShiftAmt], theta_data[(((x * 5) + y) * W) + ShiftAmt+:Offset]};
				end
			end
		end
	endgenerate
endmodule
module prim_lc_sender (
	clk_i,
	rst_ni,
	lc_en_i,
	lc_en_o
);
	parameter [0:0] AsyncOn = 1;
	parameter [0:0] ResetValueIsOn = 0;
	input clk_i;
	input rst_ni;
	localparam signed [31:0] lc_ctrl_pkg_TxWidth = 4;
	input wire [3:0] lc_en_i;
	output wire [3:0] lc_en_o;
	function automatic [3:0] sv2v_cast_01D55;
		input reg [3:0] inp;
		sv2v_cast_01D55 = inp;
	endfunction
	localparam [3:0] ResetValue = (ResetValueIsOn ? sv2v_cast_01D55(4'b0101) : sv2v_cast_01D55(4'b1010));
	wire [3:0] lc_en;
	wire [3:0] lc_en_out;
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	assign lc_en = sv2v_cast_4(lc_en_i);
	generate
		if (AsyncOn) begin : gen_flops
			prim_sec_anchor_flop #(
				.Width(lc_ctrl_pkg_TxWidth),
				.ResetValue(sv2v_cast_4(ResetValue))
			) u_prim_flop(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(lc_en),
				.q_o(lc_en_out)
			);
		end
		else begin : gen_no_flops
			genvar k;
			for (k = 0; k < lc_ctrl_pkg_TxWidth; k = k + 1) begin : gen_bits
				prim_sec_anchor_buf u_prim_buf(
					.in_i(lc_en[k]),
					.out_o(lc_en_out[k])
				);
			end
			reg [3:0] unused_logic;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					unused_logic <= sv2v_cast_01D55(4'b1010);
				else
					unused_logic <= lc_en_i;
		end
	endgenerate
	assign lc_en_o = lc_en_out;
endmodule
module prim_lc_sync (
	clk_i,
	rst_ni,
	lc_en_i,
	lc_en_o
);
	parameter signed [31:0] NumCopies = 1;
	parameter [0:0] AsyncOn = 1;
	parameter [0:0] ResetValueIsOn = 0;
	input clk_i;
	input rst_ni;
	localparam signed [31:0] lc_ctrl_pkg_TxWidth = 4;
	input wire [3:0] lc_en_i;
	output wire [(NumCopies * lc_ctrl_pkg_TxWidth) - 1:0] lc_en_o;
	function automatic [3:0] sv2v_cast_EFDF5;
		input reg [3:0] inp;
		sv2v_cast_EFDF5 = inp;
	endfunction
	localparam [3:0] LcResetValue = (ResetValueIsOn ? sv2v_cast_EFDF5(4'b0101) : sv2v_cast_EFDF5(4'b1010));
	wire [3:0] lc_en;
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	generate
		if (AsyncOn) begin : gen_flops
			prim_flop_2sync #(
				.Width(lc_ctrl_pkg_TxWidth),
				.ResetValue(sv2v_cast_4(LcResetValue))
			) u_prim_flop_2sync(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(lc_en_i),
				.q_o(lc_en)
			);
		end
		else begin : gen_no_flops
			reg [3:0] unused_logic;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					unused_logic <= sv2v_cast_EFDF5(4'b1010);
				else
					unused_logic <= lc_en_i;
			assign lc_en = lc_en_i;
		end
	endgenerate
	genvar j;
	generate
		for (j = 0; j < NumCopies; j = j + 1) begin : gen_buffs
			wire [3:0] lc_en_out;
			genvar k;
			for (k = 0; k < lc_ctrl_pkg_TxWidth; k = k + 1) begin : gen_bits
				prim_sec_anchor_buf u_prim_buf(
					.in_i(lc_en[k]),
					.out_o(lc_en_out[k])
				);
			end
			assign lc_en_o[j * lc_ctrl_pkg_TxWidth+:lc_ctrl_pkg_TxWidth] = lc_en_out;
		end
	endgenerate
endmodule
module prim_lfsr (
	clk_i,
	rst_ni,
	seed_en_i,
	seed_i,
	lfsr_en_i,
	entropy_i,
	state_o
);
	parameter LfsrType = "GAL_XOR";
	parameter [31:0] LfsrDw = 32;
	localparam [31:0] LfsrIdxDw = $clog2(LfsrDw);
	parameter [31:0] EntropyDw = 8;
	parameter [31:0] StateOutDw = 8;
	function automatic signed [LfsrDw - 1:0] sv2v_cast_B0C40_signed;
		input reg signed [LfsrDw - 1:0] inp;
		sv2v_cast_B0C40_signed = inp;
	endfunction
	parameter [LfsrDw - 1:0] DefaultSeed = sv2v_cast_B0C40_signed(1);
	parameter [LfsrDw - 1:0] CustomCoeffs = 1'sb0;
	parameter [0:0] StatePermEn = 1'b0;
	parameter [(LfsrDw * LfsrIdxDw) - 1:0] StatePerm = 1'sb0;
	parameter [0:0] MaxLenSVA = 1'b1;
	parameter [0:0] LockupSVA = 1'b1;
	parameter [0:0] ExtSeedSVA = 1'b1;
	parameter [0:0] NonLinearOut = 1'b0;
	input clk_i;
	input rst_ni;
	input seed_en_i;
	input [LfsrDw - 1:0] seed_i;
	input lfsr_en_i;
	input [EntropyDw - 1:0] entropy_i;
	output wire [StateOutDw - 1:0] state_o;
	localparam [31:0] GAL_XOR_LUT_OFF = 4;
	localparam [3903:0] GAL_XOR_COEFFS = 3904'h9000000000000001200000000000000210000000000000041000000000000008e0000000000000108000000000000020400000000000004020000000000000829000000000000100d0000000000002015000000000000400100000000000080160000000000010004000000000002001300000000000400130000000000080004000000000010000200000000002000010000000000400010000000000080000d00000000010000040000000002000023000000000400001300000000080000040000000010000002000000002000002900000000400000040000000080000057000000010000002900000002000000730000000400000002000000080000003b000000100000001f00000020000000310000004000000008000000800000001c0000010000000004000002000000001f000004000000002c0000080000000032000010000000000d00002000000000970000400000000010000080000000005b0001000000000038000200000000000e000400000000002500080000000000040010000000000023002000000000003e0040000000000023008000000000004a01000000000000160200000000000031040000000000003d0800000000000001100000000000001320000000000000344000000000000001800000000000000d;
	localparam [31:0] FIB_XNOR_LUT_OFF = 3;
	localparam [27887:0] FIB_XNOR_COEFFS = 27888'h600000000000000000000000000000000000000000c0000000000000000000000000000000000000000140000000000000000000000000000000000000000300000000000000000000000000000000000000000600000000000000000000000000000000000000000b800000000000000000000000000000000000000011000000000000000000000000000000000000000024000000000000000000000000000000000000000050000000000000000000000000000000000000000082900000000000000000000000000000000000000100d00000000000000000000000000000000000000201500000000000000000000000000000000000000600000000000000000000000000000000000000000d008000000000000000000000000000000000000012000000000000000000000000000000000000000020400000000000000000000000000000000000000040023000000000000000000000000000000000000090000000000000000000000000000000000000000140000000000000000000000000000000000000000300000000000000000000000000000000000000000420000000000000000000000000000000000000000e1000000000000000000000000000000000000000120000000000000000000000000000000000000000200002300000000000000000000000000000000000400001300000000000000000000000000000000000900000000000000000000000000000000000000001400000000000000000000000000000000000000002000002900000000000000000000000000000000004800000000000000000000000000000000000000008020000300000000000000000000000000000000010008000000000000000000000000000000000000020400000300000000000000000000000000000000050000000000000000000000000000000000000000080100000000000000000000000000000000000000100000001f00000000000000000000000000000000200000003100000000000000000000000000000000440000000000000000000000000000000000000000a0001400000000000000000000000000000000000120000000000000000000000000000000000000000300000c00000000000000000000000000000000000630000000000000000000000000000000000000000c00000300000000000000000000000000000000001b0000000000000000000000000000000000000000300003000000000000000000000000000000000000420000000000000000000000000000000000000000c00000180000000000000000000000000000000001008000000000000000000000000000000000000003000000c00000000000000000000000000000000006000c000000000000000000000000000000000000090000000000000000000000000000000000000000180030000000000000000000000000000000000000300000000300000000000000000000000000000000400000400000000000000000000000000000000000c0000600000000000000000000000000000000000102000000000000000000000000000000000000000200004000000000000000000000000000000000000600003000000000000000000000000000000000000c0000000000000000000000000000000000000000180030000000000000000000000000000000000000300000000000003000000000000000000000000000600000000000000000000000000000000000000000d80000000000000000000000000000000000000001000040000000000000000000000000000000000003018000000000000000000000000000000000000006030000000000000000000000000000000000000008040000000000000000000000000000000000000014000002800000000000000000000000000000000030006000000000000000000000000000000000000041000000000000000000000000000000000000000082000000000104000000000000000000000000000100000080000000000000000000000000000000000300060000000000000000000000000000000000000601800000000000000000000000000000000000000c0000000180000000000000000000000000000000180000006000000000000000000000000000000000300006000000000000000000000000000000000000402000000000000000000000000000000000000000c000000006000000000000000000000000000000011000000000000000000000000000000000000000024000000048000000000000000000000000000000060000000000300000000000000000000000000000080040000000000000000000000000000000000000180000030000000000000000000000000000000000300300000000000000000000000000000000000000400200000000000000000000000000000000000000c000000000000000018000000000000000000000010000000004000000000000000000000000000000030000c000000000000000000000000000000000000600000000000000000000c00000000000000000000c00c0000000000000000000000000000000000000140000000000000000000000000000000000000000200001000000000000000000000000000000000000400800000000000000000000000000000000000000a00000000001400000000000000000000000000001040000000000000000000000000000000000000002004000000000000000000000000000000000000005000000000028000000000000000000000000000008000000004000000000000000000000000000000018600000000000000000000000000000000000000030000000000000000c000000000000000000000000402000000000000000000000000000000000000000c03000000000000000000000000000000000000001000100000000000000000000000000000000000002000400000000000000000000000000000000000005000000000000000a000000000000000000000000080000001000000000000000000000000000000000186000000000000000000000000000000000000000300300000000000000000000000000000000000000401000000000000000000000000000000000000000a0000000001400000000000000000000000000000100800000000000000000000000000000000000000300000000000000000001800000000000000000000600180000000000000000000000000000000000000c00000000000000003000000000000000000000001400050000000000000000000000000000000000002000000010000000000000000000000000000000004040000000000000000000000000000000000000008100000000000000000000000001020000000000010000400000000000000000000000000000000000030000000000000060000000000000000000000000050000000000000000000000000000000000000000080000000040000000000000000000000000000000180000000000000000000000000300000000000000300000000300000000000000000000000000000000600000000000000000000000000000000000000000a0000014000000000000000000000000000000000108000000000000000000000000000000000000000240000000000000000000000000000000000000000600000000000c0000000000000000000000000000080000004000000000000000000000000000000000180000000000030000000000000000000000000000200000000000001000000000000000000000000000400800000000000000000000000000000000000000c00000000000000000000000000000060000000001000008000000000000000000000000000000000003060000000000000000000000000000000000000004a400000000000000000000000000000000000000080000004000000000000000000000000000000000180000003000000000000000000000000000000000200001000000000000000000000000000000000000600006000000000000000000000000000000000000c0000000000000000600000000000000000000000100000000000010000000000000000000000000000300000000000000600000000000000000000000000600000000300000000000000000000000000000000800000100000000000000000000000000000000001800000000000000000000000000c0000000000000200000000000010000000000000000000000000000480000000000000000000000000000000000000000c000000000000000600000000000000000000000018000000000000000000000000000000000000000028000000000000000000000000000000500000000060000000c000000000000000000000000000000000c00000000000000000000000000018000000000001800000600000000000000000000000000000000003000000c0000000000000000000000000000000000400000008000000000000000000000000000000000c0003000000000000000000000000000000000000100004000000000000000000000000000000000000300000000000000000000060000000000000000000600000000000000c00000000000000000000000000c00600000000000000000000000000000000000001800000060000000000000000000000000000000003000000000c0000000000000000000000000000000410000000000000000000000000000000000000000a00140000000000000000000000000000000000000;
	wire lockup;
	wire [LfsrDw - 1:0] lfsr_d;
	reg [LfsrDw - 1:0] lfsr_q;
	wire [LfsrDw - 1:0] next_lfsr_state;
	wire [LfsrDw - 1:0] coeffs;
	localparam [LfsrDw - 1:0] DefaultSeedLocal = DefaultSeed;
	function automatic [LfsrDw - 1:0] sv2v_cast_B0C40;
		input reg [LfsrDw - 1:0] inp;
		sv2v_cast_B0C40 = inp;
	endfunction
	function automatic [63:0] sv2v_cast_64;
		input reg [63:0] inp;
		sv2v_cast_64 = inp;
	endfunction
	generate
		if (sv2v_cast_64(LfsrType) == sv2v_cast_64("GAL_XOR")) begin : gen_gal_xor
			if (CustomCoeffs > 0) begin : gen_custom
				assign coeffs = CustomCoeffs[LfsrDw - 1:0];
			end
			else begin : gen_lut
				assign coeffs = GAL_XOR_COEFFS[((60 - (LfsrDw - GAL_XOR_LUT_OFF)) * 64) + (LfsrDw - 1)-:LfsrDw];
			end
			assign next_lfsr_state = (sv2v_cast_B0C40(entropy_i) ^ ({LfsrDw {lfsr_q[0]}} & coeffs)) ^ (lfsr_q >> 1);
			assign lockup = ~(|lfsr_q);
		end
		else if (sv2v_cast_64(LfsrType) == "FIB_XNOR") begin : gen_fib_xnor
			if (CustomCoeffs > 0) begin : gen_custom
				assign coeffs = CustomCoeffs[LfsrDw - 1:0];
			end
			else begin : gen_lut
				assign coeffs = FIB_XNOR_COEFFS[((165 - (LfsrDw - FIB_XNOR_LUT_OFF)) * 168) + (LfsrDw - 1)-:LfsrDw];
			end
			assign next_lfsr_state = sv2v_cast_B0C40(entropy_i) ^ {lfsr_q[LfsrDw - 2:0], ~(^(lfsr_q & coeffs))};
			assign lockup = &lfsr_q;
		end
		else begin : gen_unknown_type
			assign coeffs = 1'sb0;
			assign next_lfsr_state = 1'sb0;
			assign lockup = 1'b0;
		end
	endgenerate
	assign lfsr_d = (seed_en_i ? seed_i : (lfsr_en_i && lockup ? DefaultSeedLocal : (lfsr_en_i ? next_lfsr_state : lfsr_q)));
	wire [LfsrDw - 1:0] sbox_out;
	localparam [63:0] prim_cipher_pkg_PRINCE_SBOX4 = 64'h4d5e087619ca23fb;
	generate
		if (NonLinearOut) begin : gen_out_non_linear
			localparam signed [31:0] NumSboxes = LfsrDw / 4;
			wire [((4 * NumSboxes) * LfsrIdxDw) - 1:0] matrix_indices;
			genvar j;
			for (j = 0; j < LfsrDw; j = j + 1) begin : gen_input_idx_map
				assign matrix_indices[(((j / NumSboxes) * NumSboxes) + (j % NumSboxes)) * LfsrIdxDw+:LfsrIdxDw] = j;
			end
			reg [((4 * NumSboxes) * LfsrIdxDw) - 1:0] matrix_rotrev_indices;
			function automatic [(NumSboxes * LfsrIdxDw) - 1:0] lrotcol;
				input reg [(NumSboxes * LfsrIdxDw) - 1:0] col;
				input integer shift;
				reg [(NumSboxes * LfsrIdxDw) - 1:0] out;
				begin
					begin : sv2v_autoblock_1
						reg signed [31:0] k;
						for (k = 0; k < NumSboxes; k = k + 1)
							out[((k + shift) % NumSboxes) * LfsrIdxDw+:LfsrIdxDw] = col[k * LfsrIdxDw+:LfsrIdxDw];
					end
					lrotcol = out;
				end
			endfunction
			function automatic [(NumSboxes * LfsrIdxDw) - 1:0] revcol;
				input reg [(NumSboxes * LfsrIdxDw) - 1:0] col;
				begin : sv2v_autoblock_2
					reg [(0 + (NumSboxes * LfsrIdxDw)) - 1:0] _sv2v_strm_C393D_inp;
					reg [(0 + (NumSboxes * LfsrIdxDw)) - 1:0] _sv2v_strm_C393D_out;
					integer _sv2v_strm_C393D_idx;
					_sv2v_strm_C393D_inp = {col};
					for (_sv2v_strm_C393D_idx = 0; _sv2v_strm_C393D_idx <= ((0 + (NumSboxes * LfsrIdxDw)) - LfsrIdxDw); _sv2v_strm_C393D_idx = _sv2v_strm_C393D_idx + LfsrIdxDw)
						_sv2v_strm_C393D_out[((0 + (NumSboxes * LfsrIdxDw)) - 1) - _sv2v_strm_C393D_idx-:LfsrIdxDw] = _sv2v_strm_C393D_inp[_sv2v_strm_C393D_idx+:LfsrIdxDw];
					if (((0 + (NumSboxes * LfsrIdxDw)) % LfsrIdxDw) > 0)
						_sv2v_strm_C393D_out[0+:(0 + (NumSboxes * LfsrIdxDw)) % LfsrIdxDw] = _sv2v_strm_C393D_inp[_sv2v_strm_C393D_idx+:(0 + (NumSboxes * LfsrIdxDw)) % LfsrIdxDw];
					revcol = ((0 + (NumSboxes * LfsrIdxDw)) <= (NumSboxes * LfsrIdxDw) ? _sv2v_strm_C393D_out << ((NumSboxes * LfsrIdxDw) - (0 + (NumSboxes * LfsrIdxDw))) : _sv2v_strm_C393D_out >> ((0 + (NumSboxes * LfsrIdxDw)) - (NumSboxes * LfsrIdxDw)));
				end
			endfunction
			always @(*) begin : p_rotrev
				matrix_rotrev_indices[0+:LfsrIdxDw * NumSboxes] = matrix_indices[0+:LfsrIdxDw * NumSboxes];
				matrix_rotrev_indices[LfsrIdxDw * NumSboxes+:LfsrIdxDw * NumSboxes] = lrotcol(matrix_indices[LfsrIdxDw * NumSboxes+:LfsrIdxDw * NumSboxes], NumSboxes / 2);
				matrix_rotrev_indices[LfsrIdxDw * (2 * NumSboxes)+:LfsrIdxDw * NumSboxes] = revcol(matrix_indices[LfsrIdxDw * (2 * NumSboxes)+:LfsrIdxDw * NumSboxes]);
				matrix_rotrev_indices[LfsrIdxDw * (3 * NumSboxes)+:LfsrIdxDw * NumSboxes] = revcol(lrotcol(matrix_indices[LfsrIdxDw * (3 * NumSboxes)+:LfsrIdxDw * NumSboxes], 1));
			end
			wire [(LfsrDw * LfsrIdxDw) - 1:0] sbox_in_indices;
			genvar k;
			for (k = 0; k < LfsrDw; k = k + 1) begin : gen_reverse_upper
				assign sbox_in_indices[k * LfsrIdxDw+:LfsrIdxDw] = matrix_rotrev_indices[(((k % 4) * NumSboxes) + (k / 4)) * LfsrIdxDw+:LfsrIdxDw];
			end
			for (k = 0; k < NumSboxes; k = k + 1) begin : gen_sboxes
				wire [3:0] sbox_in;
				assign sbox_in = {lfsr_q[sbox_in_indices[((k * 4) + 3) * LfsrIdxDw+:LfsrIdxDw]], lfsr_q[sbox_in_indices[((k * 4) + 2) * LfsrIdxDw+:LfsrIdxDw]], lfsr_q[sbox_in_indices[((k * 4) + 1) * LfsrIdxDw+:LfsrIdxDw]], lfsr_q[sbox_in_indices[((k * 4) + 0) * LfsrIdxDw+:LfsrIdxDw]]};
				assign sbox_out[k * 4+:4] = prim_cipher_pkg_PRINCE_SBOX4[sbox_in * 4+:4];
			end
		end
		else begin : gen_out_passthru
			assign sbox_out = lfsr_q;
		end
	endgenerate
	function automatic [StateOutDw - 1:0] sv2v_cast_23274;
		input reg [StateOutDw - 1:0] inp;
		sv2v_cast_23274 = inp;
	endfunction
	generate
		if (StatePermEn) begin : gen_state_perm
			genvar k;
			for (k = 0; k < StateOutDw; k = k + 1) begin : gen_perm_loop
				assign state_o[k] = sbox_out[StatePerm[k * LfsrIdxDw+:LfsrIdxDw]];
			end
			if (LfsrDw > StateOutDw) begin : gen_tieoff_unused
				wire unused_sbox_out;
				assign unused_sbox_out = ^sbox_out;
			end
		end
		else begin : gen_no_state_perm
			assign state_o = sv2v_cast_23274(sbox_out);
		end
	endgenerate
	always @(posedge clk_i or negedge rst_ni) begin : p_reg
		if (!rst_ni)
			lfsr_q <= DefaultSeedLocal;
		else
			lfsr_q <= lfsr_d;
	end
endmodule
module prim_mubi12_dec (
	mubi_i,
	mubi_dec_o
);
	parameter [0:0] TestTrue = 1;
	parameter [0:0] TestStrict = 1;
	localparam signed [31:0] prim_mubi_pkg_MuBi12Width = 12;
	input wire [11:0] mubi_i;
	output wire mubi_dec_o;
	wire [11:0] mubi;
	wire [11:0] mubi_out;
	function automatic [11:0] sv2v_cast_12;
		input reg [11:0] inp;
		sv2v_cast_12 = inp;
	endfunction
	assign mubi = sv2v_cast_12(mubi_i);
	genvar k;
	generate
		for (k = 0; k < prim_mubi_pkg_MuBi12Width; k = k + 1) begin : gen_bits
			prim_buf u_prim_buf(
				.in_i(mubi[k]),
				.out_o(mubi_out[k])
			);
		end
	endgenerate
	function automatic [11:0] sv2v_cast_514AD;
		input reg [11:0] inp;
		sv2v_cast_514AD = inp;
	endfunction
	function automatic prim_mubi_pkg_mubi12_test_false_loose;
		input reg [11:0] val;
		prim_mubi_pkg_mubi12_test_false_loose = sv2v_cast_514AD(12'h696) != val;
	endfunction
	function automatic prim_mubi_pkg_mubi12_test_false_strict;
		input reg [11:0] val;
		prim_mubi_pkg_mubi12_test_false_strict = sv2v_cast_514AD(12'h969) == val;
	endfunction
	function automatic prim_mubi_pkg_mubi12_test_true_loose;
		input reg [11:0] val;
		prim_mubi_pkg_mubi12_test_true_loose = sv2v_cast_514AD(12'h969) != val;
	endfunction
	function automatic prim_mubi_pkg_mubi12_test_true_strict;
		input reg [11:0] val;
		prim_mubi_pkg_mubi12_test_true_strict = sv2v_cast_514AD(12'h696) == val;
	endfunction
	generate
		if (TestTrue && TestStrict) begin : gen_test_true_strict
			assign mubi_dec_o = prim_mubi_pkg_mubi12_test_true_strict(mubi_out);
		end
		else if (TestTrue && !TestStrict) begin : gen_test_true_loose
			assign mubi_dec_o = prim_mubi_pkg_mubi12_test_true_loose(mubi_out);
		end
		else if (!TestTrue && TestStrict) begin : gen_test_false_strict
			assign mubi_dec_o = prim_mubi_pkg_mubi12_test_false_strict(mubi_out);
		end
		else if (!TestTrue && !TestStrict) begin : gen_test_false_loose
			assign mubi_dec_o = prim_mubi_pkg_mubi12_test_false_loose(mubi_out);
		end
	endgenerate
endmodule
module prim_mubi12_sender (
	clk_i,
	rst_ni,
	mubi_i,
	mubi_o
);
	parameter [0:0] AsyncOn = 1;
	parameter [0:0] EnSecBuf = 0;
	localparam signed [31:0] prim_mubi_pkg_MuBi12Width = 12;
	function automatic [11:0] sv2v_cast_29745;
		input reg [11:0] inp;
		sv2v_cast_29745 = inp;
	endfunction
	parameter [11:0] ResetValue = sv2v_cast_29745(12'h969);
	input clk_i;
	input rst_ni;
	input wire [11:0] mubi_i;
	output wire [11:0] mubi_o;
	wire [11:0] mubi;
	wire [11:0] mubi_int;
	wire [11:0] mubi_out;
	function automatic [11:0] sv2v_cast_12;
		input reg [11:0] inp;
		sv2v_cast_12 = inp;
	endfunction
	assign mubi = sv2v_cast_12(mubi_i);
	generate
		if (AsyncOn) begin : gen_flops
			prim_flop #(
				.Width(prim_mubi_pkg_MuBi12Width),
				.ResetValue(sv2v_cast_12(ResetValue))
			) u_prim_flop(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(mubi),
				.q_o(mubi_int)
			);
		end
		else begin : gen_no_flops
			assign mubi_int = mubi;
			reg [11:0] unused_logic;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					unused_logic <= sv2v_cast_29745(12'h969);
				else
					unused_logic <= mubi_i;
		end
		if (EnSecBuf) begin : gen_sec_buf
			prim_sec_anchor_buf #(.Width(12)) u_prim_sec_buf(
				.in_i(mubi_int),
				.out_o(mubi_out)
			);
		end
		else if (!AsyncOn) begin : gen_prim_buf
			prim_buf #(.Width(12)) u_prim_buf(
				.in_i(mubi_int),
				.out_o(mubi_out)
			);
		end
		else begin : gen_feedthru
			assign mubi_out = mubi_int;
		end
	endgenerate
	assign mubi_o = mubi_out;
endmodule
module prim_mubi12_sync (
	clk_i,
	rst_ni,
	mubi_i,
	mubi_o
);
	parameter signed [31:0] NumCopies = 1;
	parameter [0:0] AsyncOn = 1;
	parameter [0:0] StabilityCheck = 0;
	localparam signed [31:0] prim_mubi_pkg_MuBi12Width = 12;
	function automatic [11:0] sv2v_cast_43D25;
		input reg [11:0] inp;
		sv2v_cast_43D25 = inp;
	endfunction
	parameter [11:0] ResetValue = sv2v_cast_43D25(12'h969);
	input clk_i;
	input rst_ni;
	input wire [11:0] mubi_i;
	output wire [(NumCopies * prim_mubi_pkg_MuBi12Width) - 1:0] mubi_o;
	wire [11:0] mubi;
	function automatic [11:0] sv2v_cast_12;
		input reg [11:0] inp;
		sv2v_cast_12 = inp;
	endfunction
	generate
		if (AsyncOn) begin : gen_flops
			wire [11:0] mubi_sync;
			prim_flop_2sync #(
				.Width(prim_mubi_pkg_MuBi12Width),
				.ResetValue(sv2v_cast_12(ResetValue))
			) u_prim_flop_2sync(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(sv2v_cast_12(mubi_i)),
				.q_o(mubi_sync)
			);
			if (StabilityCheck) begin : gen_stable_chks
				wire [11:0] mubi_q;
				prim_flop #(
					.Width(prim_mubi_pkg_MuBi12Width),
					.ResetValue(sv2v_cast_12(ResetValue))
				) u_prim_flop_3rd_stage(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.d_i(mubi_sync),
					.q_o(mubi_q)
				);
				wire [11:0] sig_unstable;
				prim_xor2 #(.Width(prim_mubi_pkg_MuBi12Width)) u_mubi_xor(
					.in0_i(mubi_sync),
					.in1_i(mubi_q),
					.out_o(sig_unstable)
				);
				wire [11:0] reset_value;
				assign reset_value = ResetValue;
				genvar k;
				for (k = 0; k < prim_mubi_pkg_MuBi12Width; k = k + 1) begin : gen_bufs_muxes
					wire [11:0] sig_unstable_buf;
					prim_sec_anchor_buf #(.Width(prim_mubi_pkg_MuBi12Width)) u_sig_unstable_buf(
						.in_i(sig_unstable),
						.out_o(sig_unstable_buf)
					);
					assign mubi[k] = (|sig_unstable_buf ? reset_value[k] : mubi_q[k]);
				end
			end
			else begin : gen_no_stable_chks
				assign mubi = mubi_sync;
			end
		end
		else begin : gen_no_flops
			reg [11:0] unused_logic;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					unused_logic <= sv2v_cast_43D25(12'h969);
				else
					unused_logic <= mubi_i;
			assign mubi = sv2v_cast_12(mubi_i);
		end
	endgenerate
	genvar j;
	generate
		for (j = 0; j < NumCopies; j = j + 1) begin : gen_buffs
			wire [11:0] mubi_out;
			genvar k;
			for (k = 0; k < prim_mubi_pkg_MuBi12Width; k = k + 1) begin : gen_bits
				prim_buf u_prim_buf(
					.in_i(mubi[k]),
					.out_o(mubi_out[k])
				);
			end
			assign mubi_o[j * prim_mubi_pkg_MuBi12Width+:prim_mubi_pkg_MuBi12Width] = mubi_out;
		end
	endgenerate
endmodule
module prim_mubi16_dec (
	mubi_i,
	mubi_dec_o
);
	parameter [0:0] TestTrue = 1;
	parameter [0:0] TestStrict = 1;
	localparam signed [31:0] prim_mubi_pkg_MuBi16Width = 16;
	input wire [15:0] mubi_i;
	output wire mubi_dec_o;
	wire [15:0] mubi;
	wire [15:0] mubi_out;
	function automatic [15:0] sv2v_cast_16;
		input reg [15:0] inp;
		sv2v_cast_16 = inp;
	endfunction
	assign mubi = sv2v_cast_16(mubi_i);
	genvar k;
	generate
		for (k = 0; k < prim_mubi_pkg_MuBi16Width; k = k + 1) begin : gen_bits
			prim_buf u_prim_buf(
				.in_i(mubi[k]),
				.out_o(mubi_out[k])
			);
		end
	endgenerate
	function automatic [15:0] sv2v_cast_6CE35;
		input reg [15:0] inp;
		sv2v_cast_6CE35 = inp;
	endfunction
	function automatic prim_mubi_pkg_mubi16_test_false_loose;
		input reg [15:0] val;
		prim_mubi_pkg_mubi16_test_false_loose = sv2v_cast_6CE35(16'h9696) != val;
	endfunction
	function automatic prim_mubi_pkg_mubi16_test_false_strict;
		input reg [15:0] val;
		prim_mubi_pkg_mubi16_test_false_strict = sv2v_cast_6CE35(16'h6969) == val;
	endfunction
	function automatic prim_mubi_pkg_mubi16_test_true_loose;
		input reg [15:0] val;
		prim_mubi_pkg_mubi16_test_true_loose = sv2v_cast_6CE35(16'h6969) != val;
	endfunction
	function automatic prim_mubi_pkg_mubi16_test_true_strict;
		input reg [15:0] val;
		prim_mubi_pkg_mubi16_test_true_strict = sv2v_cast_6CE35(16'h9696) == val;
	endfunction
	generate
		if (TestTrue && TestStrict) begin : gen_test_true_strict
			assign mubi_dec_o = prim_mubi_pkg_mubi16_test_true_strict(mubi_out);
		end
		else if (TestTrue && !TestStrict) begin : gen_test_true_loose
			assign mubi_dec_o = prim_mubi_pkg_mubi16_test_true_loose(mubi_out);
		end
		else if (!TestTrue && TestStrict) begin : gen_test_false_strict
			assign mubi_dec_o = prim_mubi_pkg_mubi16_test_false_strict(mubi_out);
		end
		else if (!TestTrue && !TestStrict) begin : gen_test_false_loose
			assign mubi_dec_o = prim_mubi_pkg_mubi16_test_false_loose(mubi_out);
		end
	endgenerate
endmodule
module prim_mubi16_sender (
	clk_i,
	rst_ni,
	mubi_i,
	mubi_o
);
	parameter [0:0] AsyncOn = 1;
	parameter [0:0] EnSecBuf = 0;
	localparam signed [31:0] prim_mubi_pkg_MuBi16Width = 16;
	function automatic [15:0] sv2v_cast_75CDD;
		input reg [15:0] inp;
		sv2v_cast_75CDD = inp;
	endfunction
	parameter [15:0] ResetValue = sv2v_cast_75CDD(16'h6969);
	input clk_i;
	input rst_ni;
	input wire [15:0] mubi_i;
	output wire [15:0] mubi_o;
	wire [15:0] mubi;
	wire [15:0] mubi_int;
	wire [15:0] mubi_out;
	function automatic [15:0] sv2v_cast_16;
		input reg [15:0] inp;
		sv2v_cast_16 = inp;
	endfunction
	assign mubi = sv2v_cast_16(mubi_i);
	generate
		if (AsyncOn) begin : gen_flops
			prim_flop #(
				.Width(prim_mubi_pkg_MuBi16Width),
				.ResetValue(sv2v_cast_16(ResetValue))
			) u_prim_flop(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(mubi),
				.q_o(mubi_int)
			);
		end
		else begin : gen_no_flops
			assign mubi_int = mubi;
			reg [15:0] unused_logic;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					unused_logic <= sv2v_cast_75CDD(16'h6969);
				else
					unused_logic <= mubi_i;
		end
		if (EnSecBuf) begin : gen_sec_buf
			prim_sec_anchor_buf #(.Width(16)) u_prim_sec_buf(
				.in_i(mubi_int),
				.out_o(mubi_out)
			);
		end
		else if (!AsyncOn) begin : gen_prim_buf
			prim_buf #(.Width(16)) u_prim_buf(
				.in_i(mubi_int),
				.out_o(mubi_out)
			);
		end
		else begin : gen_feedthru
			assign mubi_out = mubi_int;
		end
	endgenerate
	assign mubi_o = mubi_out;
endmodule
module prim_mubi16_sync (
	clk_i,
	rst_ni,
	mubi_i,
	mubi_o
);
	parameter signed [31:0] NumCopies = 1;
	parameter [0:0] AsyncOn = 1;
	parameter [0:0] StabilityCheck = 0;
	localparam signed [31:0] prim_mubi_pkg_MuBi16Width = 16;
	function automatic [15:0] sv2v_cast_0F4D5;
		input reg [15:0] inp;
		sv2v_cast_0F4D5 = inp;
	endfunction
	parameter [15:0] ResetValue = sv2v_cast_0F4D5(16'h6969);
	input clk_i;
	input rst_ni;
	input wire [15:0] mubi_i;
	output wire [(NumCopies * prim_mubi_pkg_MuBi16Width) - 1:0] mubi_o;
	wire [15:0] mubi;
	function automatic [15:0] sv2v_cast_16;
		input reg [15:0] inp;
		sv2v_cast_16 = inp;
	endfunction
	generate
		if (AsyncOn) begin : gen_flops
			wire [15:0] mubi_sync;
			prim_flop_2sync #(
				.Width(prim_mubi_pkg_MuBi16Width),
				.ResetValue(sv2v_cast_16(ResetValue))
			) u_prim_flop_2sync(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(sv2v_cast_16(mubi_i)),
				.q_o(mubi_sync)
			);
			if (StabilityCheck) begin : gen_stable_chks
				wire [15:0] mubi_q;
				prim_flop #(
					.Width(prim_mubi_pkg_MuBi16Width),
					.ResetValue(sv2v_cast_16(ResetValue))
				) u_prim_flop_3rd_stage(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.d_i(mubi_sync),
					.q_o(mubi_q)
				);
				wire [15:0] sig_unstable;
				prim_xor2 #(.Width(prim_mubi_pkg_MuBi16Width)) u_mubi_xor(
					.in0_i(mubi_sync),
					.in1_i(mubi_q),
					.out_o(sig_unstable)
				);
				wire [15:0] reset_value;
				assign reset_value = ResetValue;
				genvar k;
				for (k = 0; k < prim_mubi_pkg_MuBi16Width; k = k + 1) begin : gen_bufs_muxes
					wire [15:0] sig_unstable_buf;
					prim_sec_anchor_buf #(.Width(prim_mubi_pkg_MuBi16Width)) u_sig_unstable_buf(
						.in_i(sig_unstable),
						.out_o(sig_unstable_buf)
					);
					assign mubi[k] = (|sig_unstable_buf ? reset_value[k] : mubi_q[k]);
				end
			end
			else begin : gen_no_stable_chks
				assign mubi = mubi_sync;
			end
		end
		else begin : gen_no_flops
			reg [15:0] unused_logic;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					unused_logic <= sv2v_cast_0F4D5(16'h6969);
				else
					unused_logic <= mubi_i;
			assign mubi = sv2v_cast_16(mubi_i);
		end
	endgenerate
	genvar j;
	generate
		for (j = 0; j < NumCopies; j = j + 1) begin : gen_buffs
			wire [15:0] mubi_out;
			genvar k;
			for (k = 0; k < prim_mubi_pkg_MuBi16Width; k = k + 1) begin : gen_bits
				prim_buf u_prim_buf(
					.in_i(mubi[k]),
					.out_o(mubi_out[k])
				);
			end
			assign mubi_o[j * prim_mubi_pkg_MuBi16Width+:prim_mubi_pkg_MuBi16Width] = mubi_out;
		end
	endgenerate
endmodule
module prim_mubi4_dec (
	mubi_i,
	mubi_dec_o
);
	parameter [0:0] TestTrue = 1;
	parameter [0:0] TestStrict = 1;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	input wire [3:0] mubi_i;
	output wire mubi_dec_o;
	wire [3:0] mubi;
	wire [3:0] mubi_out;
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	assign mubi = sv2v_cast_4(mubi_i);
	genvar k;
	generate
		for (k = 0; k < prim_mubi_pkg_MuBi4Width; k = k + 1) begin : gen_bits
			prim_buf u_prim_buf(
				.in_i(mubi[k]),
				.out_o(mubi_out[k])
			);
		end
	endgenerate
	function automatic [3:0] sv2v_cast_555F9;
		input reg [3:0] inp;
		sv2v_cast_555F9 = inp;
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_false_loose;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_false_loose = sv2v_cast_555F9(4'h6) != val;
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_false_strict;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_false_strict = sv2v_cast_555F9(4'h9) == val;
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_true_loose;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_true_loose = sv2v_cast_555F9(4'h9) != val;
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_true_strict;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_true_strict = sv2v_cast_555F9(4'h6) == val;
	endfunction
	generate
		if (TestTrue && TestStrict) begin : gen_test_true_strict
			assign mubi_dec_o = prim_mubi_pkg_mubi4_test_true_strict(mubi_out);
		end
		else if (TestTrue && !TestStrict) begin : gen_test_true_loose
			assign mubi_dec_o = prim_mubi_pkg_mubi4_test_true_loose(mubi_out);
		end
		else if (!TestTrue && TestStrict) begin : gen_test_false_strict
			assign mubi_dec_o = prim_mubi_pkg_mubi4_test_false_strict(mubi_out);
		end
		else if (!TestTrue && !TestStrict) begin : gen_test_false_loose
			assign mubi_dec_o = prim_mubi_pkg_mubi4_test_false_loose(mubi_out);
		end
	endgenerate
endmodule
module prim_mubi4_sender (
	clk_i,
	rst_ni,
	mubi_i,
	mubi_o
);
	parameter [0:0] AsyncOn = 1;
	parameter [0:0] EnSecBuf = 0;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	function automatic [3:0] sv2v_cast_024A9;
		input reg [3:0] inp;
		sv2v_cast_024A9 = inp;
	endfunction
	parameter [3:0] ResetValue = sv2v_cast_024A9(4'h9);
	input clk_i;
	input rst_ni;
	input wire [3:0] mubi_i;
	output wire [3:0] mubi_o;
	wire [3:0] mubi;
	wire [3:0] mubi_int;
	wire [3:0] mubi_out;
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	assign mubi = sv2v_cast_4(mubi_i);
	generate
		if (AsyncOn) begin : gen_flops
			prim_flop #(
				.Width(prim_mubi_pkg_MuBi4Width),
				.ResetValue(sv2v_cast_4(ResetValue))
			) u_prim_flop(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(mubi),
				.q_o(mubi_int)
			);
		end
		else begin : gen_no_flops
			assign mubi_int = mubi;
			reg [3:0] unused_logic;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					unused_logic <= sv2v_cast_024A9(4'h9);
				else
					unused_logic <= mubi_i;
		end
		if (EnSecBuf) begin : gen_sec_buf
			prim_sec_anchor_buf #(.Width(4)) u_prim_sec_buf(
				.in_i(mubi_int),
				.out_o(mubi_out)
			);
		end
		else if (!AsyncOn) begin : gen_prim_buf
			prim_buf #(.Width(4)) u_prim_buf(
				.in_i(mubi_int),
				.out_o(mubi_out)
			);
		end
		else begin : gen_feedthru
			assign mubi_out = mubi_int;
		end
	endgenerate
	assign mubi_o = mubi_out;
endmodule
module prim_mubi4_sync (
	clk_i,
	rst_ni,
	mubi_i,
	mubi_o
);
	parameter signed [31:0] NumCopies = 1;
	parameter [0:0] AsyncOn = 1;
	parameter [0:0] StabilityCheck = 0;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	function automatic [3:0] sv2v_cast_2C9C5;
		input reg [3:0] inp;
		sv2v_cast_2C9C5 = inp;
	endfunction
	parameter [3:0] ResetValue = sv2v_cast_2C9C5(4'h9);
	input clk_i;
	input rst_ni;
	input wire [3:0] mubi_i;
	output wire [(NumCopies * prim_mubi_pkg_MuBi4Width) - 1:0] mubi_o;
	wire [3:0] mubi;
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	generate
		if (AsyncOn) begin : gen_flops
			wire [3:0] mubi_sync;
			prim_flop_2sync #(
				.Width(prim_mubi_pkg_MuBi4Width),
				.ResetValue(sv2v_cast_4(ResetValue))
			) u_prim_flop_2sync(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(sv2v_cast_4(mubi_i)),
				.q_o(mubi_sync)
			);
			if (StabilityCheck) begin : gen_stable_chks
				wire [3:0] mubi_q;
				prim_flop #(
					.Width(prim_mubi_pkg_MuBi4Width),
					.ResetValue(sv2v_cast_4(ResetValue))
				) u_prim_flop_3rd_stage(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.d_i(mubi_sync),
					.q_o(mubi_q)
				);
				wire [3:0] sig_unstable;
				prim_xor2 #(.Width(prim_mubi_pkg_MuBi4Width)) u_mubi_xor(
					.in0_i(mubi_sync),
					.in1_i(mubi_q),
					.out_o(sig_unstable)
				);
				wire [3:0] reset_value;
				assign reset_value = ResetValue;
				genvar k;
				for (k = 0; k < prim_mubi_pkg_MuBi4Width; k = k + 1) begin : gen_bufs_muxes
					wire [3:0] sig_unstable_buf;
					prim_sec_anchor_buf #(.Width(prim_mubi_pkg_MuBi4Width)) u_sig_unstable_buf(
						.in_i(sig_unstable),
						.out_o(sig_unstable_buf)
					);
					assign mubi[k] = (|sig_unstable_buf ? reset_value[k] : mubi_q[k]);
				end
			end
			else begin : gen_no_stable_chks
				assign mubi = mubi_sync;
			end
		end
		else begin : gen_no_flops
			reg [3:0] unused_logic;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					unused_logic <= sv2v_cast_2C9C5(4'h9);
				else
					unused_logic <= mubi_i;
			assign mubi = sv2v_cast_4(mubi_i);
		end
	endgenerate
	genvar j;
	generate
		for (j = 0; j < NumCopies; j = j + 1) begin : gen_buffs
			wire [3:0] mubi_out;
			genvar k;
			for (k = 0; k < prim_mubi_pkg_MuBi4Width; k = k + 1) begin : gen_bits
				prim_buf u_prim_buf(
					.in_i(mubi[k]),
					.out_o(mubi_out[k])
				);
			end
			assign mubi_o[j * prim_mubi_pkg_MuBi4Width+:prim_mubi_pkg_MuBi4Width] = mubi_out;
		end
	endgenerate
endmodule
module prim_mubi8_dec (
	mubi_i,
	mubi_dec_o
);
	parameter [0:0] TestTrue = 1;
	parameter [0:0] TestStrict = 1;
	localparam signed [31:0] prim_mubi_pkg_MuBi8Width = 8;
	input wire [7:0] mubi_i;
	output wire mubi_dec_o;
	wire [7:0] mubi;
	wire [7:0] mubi_out;
	function automatic [7:0] sv2v_cast_8;
		input reg [7:0] inp;
		sv2v_cast_8 = inp;
	endfunction
	assign mubi = sv2v_cast_8(mubi_i);
	genvar k;
	generate
		for (k = 0; k < prim_mubi_pkg_MuBi8Width; k = k + 1) begin : gen_bits
			prim_buf u_prim_buf(
				.in_i(mubi[k]),
				.out_o(mubi_out[k])
			);
		end
	endgenerate
	function automatic [7:0] sv2v_cast_42311;
		input reg [7:0] inp;
		sv2v_cast_42311 = inp;
	endfunction
	function automatic prim_mubi_pkg_mubi8_test_false_loose;
		input reg [7:0] val;
		prim_mubi_pkg_mubi8_test_false_loose = sv2v_cast_42311(8'h96) != val;
	endfunction
	function automatic prim_mubi_pkg_mubi8_test_false_strict;
		input reg [7:0] val;
		prim_mubi_pkg_mubi8_test_false_strict = sv2v_cast_42311(8'h69) == val;
	endfunction
	function automatic prim_mubi_pkg_mubi8_test_true_loose;
		input reg [7:0] val;
		prim_mubi_pkg_mubi8_test_true_loose = sv2v_cast_42311(8'h69) != val;
	endfunction
	function automatic prim_mubi_pkg_mubi8_test_true_strict;
		input reg [7:0] val;
		prim_mubi_pkg_mubi8_test_true_strict = sv2v_cast_42311(8'h96) == val;
	endfunction
	generate
		if (TestTrue && TestStrict) begin : gen_test_true_strict
			assign mubi_dec_o = prim_mubi_pkg_mubi8_test_true_strict(mubi_out);
		end
		else if (TestTrue && !TestStrict) begin : gen_test_true_loose
			assign mubi_dec_o = prim_mubi_pkg_mubi8_test_true_loose(mubi_out);
		end
		else if (!TestTrue && TestStrict) begin : gen_test_false_strict
			assign mubi_dec_o = prim_mubi_pkg_mubi8_test_false_strict(mubi_out);
		end
		else if (!TestTrue && !TestStrict) begin : gen_test_false_loose
			assign mubi_dec_o = prim_mubi_pkg_mubi8_test_false_loose(mubi_out);
		end
	endgenerate
endmodule
module prim_mubi8_sender (
	clk_i,
	rst_ni,
	mubi_i,
	mubi_o
);
	parameter [0:0] AsyncOn = 1;
	parameter [0:0] EnSecBuf = 0;
	localparam signed [31:0] prim_mubi_pkg_MuBi8Width = 8;
	function automatic [7:0] sv2v_cast_E7611;
		input reg [7:0] inp;
		sv2v_cast_E7611 = inp;
	endfunction
	parameter [7:0] ResetValue = sv2v_cast_E7611(8'h69);
	input clk_i;
	input rst_ni;
	input wire [7:0] mubi_i;
	output wire [7:0] mubi_o;
	wire [7:0] mubi;
	wire [7:0] mubi_int;
	wire [7:0] mubi_out;
	function automatic [7:0] sv2v_cast_8;
		input reg [7:0] inp;
		sv2v_cast_8 = inp;
	endfunction
	assign mubi = sv2v_cast_8(mubi_i);
	generate
		if (AsyncOn) begin : gen_flops
			prim_flop #(
				.Width(prim_mubi_pkg_MuBi8Width),
				.ResetValue(sv2v_cast_8(ResetValue))
			) u_prim_flop(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(mubi),
				.q_o(mubi_int)
			);
		end
		else begin : gen_no_flops
			assign mubi_int = mubi;
			reg [7:0] unused_logic;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					unused_logic <= sv2v_cast_E7611(8'h69);
				else
					unused_logic <= mubi_i;
		end
		if (EnSecBuf) begin : gen_sec_buf
			prim_sec_anchor_buf #(.Width(8)) u_prim_sec_buf(
				.in_i(mubi_int),
				.out_o(mubi_out)
			);
		end
		else if (!AsyncOn) begin : gen_prim_buf
			prim_buf #(.Width(8)) u_prim_buf(
				.in_i(mubi_int),
				.out_o(mubi_out)
			);
		end
		else begin : gen_feedthru
			assign mubi_out = mubi_int;
		end
	endgenerate
	assign mubi_o = mubi_out;
endmodule
module prim_mubi8_sync (
	clk_i,
	rst_ni,
	mubi_i,
	mubi_o
);
	parameter signed [31:0] NumCopies = 1;
	parameter [0:0] AsyncOn = 1;
	parameter [0:0] StabilityCheck = 0;
	localparam signed [31:0] prim_mubi_pkg_MuBi8Width = 8;
	function automatic [7:0] sv2v_cast_E2F65;
		input reg [7:0] inp;
		sv2v_cast_E2F65 = inp;
	endfunction
	parameter [7:0] ResetValue = sv2v_cast_E2F65(8'h69);
	input clk_i;
	input rst_ni;
	input wire [7:0] mubi_i;
	output wire [(NumCopies * prim_mubi_pkg_MuBi8Width) - 1:0] mubi_o;
	wire [7:0] mubi;
	function automatic [7:0] sv2v_cast_8;
		input reg [7:0] inp;
		sv2v_cast_8 = inp;
	endfunction
	generate
		if (AsyncOn) begin : gen_flops
			wire [7:0] mubi_sync;
			prim_flop_2sync #(
				.Width(prim_mubi_pkg_MuBi8Width),
				.ResetValue(sv2v_cast_8(ResetValue))
			) u_prim_flop_2sync(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.d_i(sv2v_cast_8(mubi_i)),
				.q_o(mubi_sync)
			);
			if (StabilityCheck) begin : gen_stable_chks
				wire [7:0] mubi_q;
				prim_flop #(
					.Width(prim_mubi_pkg_MuBi8Width),
					.ResetValue(sv2v_cast_8(ResetValue))
				) u_prim_flop_3rd_stage(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.d_i(mubi_sync),
					.q_o(mubi_q)
				);
				wire [7:0] sig_unstable;
				prim_xor2 #(.Width(prim_mubi_pkg_MuBi8Width)) u_mubi_xor(
					.in0_i(mubi_sync),
					.in1_i(mubi_q),
					.out_o(sig_unstable)
				);
				wire [7:0] reset_value;
				assign reset_value = ResetValue;
				genvar k;
				for (k = 0; k < prim_mubi_pkg_MuBi8Width; k = k + 1) begin : gen_bufs_muxes
					wire [7:0] sig_unstable_buf;
					prim_sec_anchor_buf #(.Width(prim_mubi_pkg_MuBi8Width)) u_sig_unstable_buf(
						.in_i(sig_unstable),
						.out_o(sig_unstable_buf)
					);
					assign mubi[k] = (|sig_unstable_buf ? reset_value[k] : mubi_q[k]);
				end
			end
			else begin : gen_no_stable_chks
				assign mubi = mubi_sync;
			end
		end
		else begin : gen_no_flops
			reg [7:0] unused_logic;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					unused_logic <= sv2v_cast_E2F65(8'h69);
				else
					unused_logic <= mubi_i;
			assign mubi = sv2v_cast_8(mubi_i);
		end
	endgenerate
	genvar j;
	generate
		for (j = 0; j < NumCopies; j = j + 1) begin : gen_buffs
			wire [7:0] mubi_out;
			genvar k;
			for (k = 0; k < prim_mubi_pkg_MuBi8Width; k = k + 1) begin : gen_bits
				prim_buf u_prim_buf(
					.in_i(mubi[k]),
					.out_o(mubi_out[k])
				);
			end
			assign mubi_o[j * prim_mubi_pkg_MuBi8Width+:prim_mubi_pkg_MuBi8Width] = mubi_out;
		end
	endgenerate
endmodule
module prim_onehot_check (
	clk_i,
	rst_ni,
	oh_i,
	addr_i,
	en_i,
	err_o
);
	parameter [31:0] AddrWidth = 5;
	parameter [31:0] OneHotWidth = 2 ** AddrWidth;
	parameter [0:0] AddrCheck = 1;
	parameter [0:0] EnableCheck = 1;
	parameter [0:0] StrictCheck = 1;
	parameter [0:0] EnableAlertTriggerSVA = 1;
	input clk_i;
	input rst_ni;
	input wire [OneHotWidth - 1:0] oh_i;
	input wire [AddrWidth - 1:0] addr_i;
	input wire en_i;
	output wire err_o;
	localparam signed [31:0] NumLevels = AddrWidth;
	wire [(2 ** (NumLevels + 1)) - 2:0] or_tree;
	wire [(2 ** (NumLevels + 1)) - 2:0] and_tree;
	wire [(2 ** (NumLevels + 1)) - 2:0] err_tree;
	genvar level;
	generate
		for (level = 0; level < (NumLevels + 1); level = level + 1) begin : gen_tree
			localparam signed [31:0] Base0 = (2 ** level) - 1;
			localparam signed [31:0] Base1 = (2 ** (level + 1)) - 1;
			genvar offset;
			for (offset = 0; offset < (2 ** level); offset = offset + 1) begin : gen_level
				localparam signed [31:0] Pa = Base0 + offset;
				localparam signed [31:0] C0 = Base1 + (2 * offset);
				localparam signed [31:0] C1 = (Base1 + (2 * offset)) + 1;
				if (level == NumLevels) begin : gen_leafs
					if (offset < OneHotWidth) begin : gen_assign
						assign or_tree[Pa] = oh_i[offset];
						assign and_tree[Pa] = oh_i[offset];
					end
					else begin : gen_tie_off
						assign or_tree[Pa] = 1'b0;
						assign and_tree[Pa] = 1'b0;
					end
					assign err_tree[Pa] = 1'b0;
				end
				else begin : gen_nodes
					assign or_tree[Pa] = or_tree[C0] || or_tree[C1];
					assign and_tree[Pa] = (!addr_i[(AddrWidth - 1) - level] && and_tree[C0]) || (addr_i[(AddrWidth - 1) - level] && and_tree[C1]);
					assign err_tree[Pa] = ((or_tree[C0] && or_tree[C1]) || err_tree[C0]) || err_tree[C1];
				end
			end
		end
	endgenerate
	wire enable_err;
	wire addr_err;
	wire oh0_err;
	assign err_o = (oh0_err || enable_err) || addr_err;
	assign oh0_err = err_tree[0];
	generate
		if (EnableCheck) begin : gen_enable_check
			if (StrictCheck) begin : gen_strict
				assign enable_err = or_tree[0] ^ en_i;
			end
			else begin : gen_not_strict
				assign enable_err = !en_i && or_tree[0];
			end
		end
		else begin : gen_no_enable_check
			wire unused_or_tree;
			assign unused_or_tree = ^or_tree;
			assign enable_err = 1'b0;
		end
		if (AddrCheck) begin : gen_addr_check_strict
			assign addr_err = or_tree[0] ^ and_tree[0];
		end
		else begin : gen_no_addr_check_strict
			wire unused_and_tree;
			assign unused_and_tree = ^and_tree;
			assign addr_err = 1'b0;
		end
	endgenerate
endmodule
module prim_packer (
	clk_i,
	rst_ni,
	valid_i,
	data_i,
	mask_i,
	ready_o,
	valid_o,
	data_o,
	mask_o,
	ready_i,
	flush_i,
	flush_done_o,
	err_o
);
	parameter [31:0] InW = 32;
	parameter [31:0] OutW = 32;
	parameter signed [31:0] HintByteData = 0;
	parameter [0:0] EnProtection = 1'b0;
	input clk_i;
	input rst_ni;
	input valid_i;
	input [InW - 1:0] data_i;
	input [InW - 1:0] mask_i;
	output wire ready_o;
	output wire valid_o;
	output wire [OutW - 1:0] data_o;
	output wire [OutW - 1:0] mask_o;
	input ready_i;
	input flush_i;
	output wire flush_done_o;
	output wire err_o;
	localparam [31:0] Width = InW + OutW;
	localparam [31:0] ConcatW = Width + InW;
	localparam [31:0] PtrW = $clog2(ConcatW + 1);
	function automatic integer prim_util_pkg_vbits;
		input integer value;
		prim_util_pkg_vbits = (value == 1 ? 1 : $clog2(value));
	endfunction
	localparam [31:0] IdxW = prim_util_pkg_vbits(InW);
	localparam [31:0] OnesCntW = $clog2(InW + 1);
	wire valid_next;
	wire ready_next;
	reg [Width - 1:0] stored_data;
	reg [Width - 1:0] stored_mask;
	wire [ConcatW - 1:0] concat_data;
	wire [ConcatW - 1:0] concat_mask;
	wire [ConcatW - 1:0] shiftl_data;
	wire [ConcatW - 1:0] shiftl_mask;
	wire [InW - 1:0] shiftr_data;
	wire [InW - 1:0] shiftr_mask;
	reg [PtrW - 1:0] pos_q;
	reg [IdxW - 1:0] lod_idx;
	reg [OnesCntW - 1:0] inmask_ones;
	wire ack_in;
	wire ack_out;
	reg flush_valid;
	reg flush_done;
	function automatic [OnesCntW - 1:0] sv2v_cast_A9CD9;
		input reg [OnesCntW - 1:0] inp;
		sv2v_cast_A9CD9 = inp;
	endfunction
	always @(*) begin
		inmask_ones = 1'sb0;
		begin : sv2v_autoblock_1
			reg signed [31:0] i;
			for (i = 0; i < InW; i = i + 1)
				inmask_ones = inmask_ones + sv2v_cast_A9CD9(mask_i[i]);
		end
	end
	wire [PtrW - 1:0] pos_with_input;
	function automatic [PtrW - 1:0] sv2v_cast_7A7B7;
		input reg [PtrW - 1:0] inp;
		sv2v_cast_7A7B7 = inp;
	endfunction
	assign pos_with_input = pos_q + sv2v_cast_7A7B7(inmask_ones);
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		if (EnProtection == 1'b0) begin : g_pos_nodup
			reg [PtrW - 1:0] pos_d;
			always @(*) begin
				pos_d = pos_q;
				case ({ack_in, ack_out})
					2'b00: pos_d = pos_q;
					2'b01: pos_d = (sv2v_cast_32_signed(pos_q) <= OutW ? {PtrW {1'sb0}} : pos_q - sv2v_cast_7A7B7(OutW));
					2'b10: pos_d = pos_with_input;
					2'b11: pos_d = (sv2v_cast_32_signed(pos_with_input) <= OutW ? {PtrW {1'sb0}} : pos_with_input - sv2v_cast_7A7B7(OutW));
					default: pos_d = pos_q;
				endcase
			end
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					pos_q <= 1'sb0;
				else if (flush_done)
					pos_q <= 1'sb0;
				else
					pos_q <= pos_d;
			assign err_o = 1'b0;
		end
		else begin : g_pos_dupcnt
			wire cnt_incr_en;
			wire cnt_decr_en;
			wire cnt_set_en;
			wire [PtrW - 1:0] cnt_step;
			reg [PtrW - 1:0] cnt_set;
			assign cnt_incr_en = ack_in && !ack_out;
			assign cnt_decr_en = !ack_in && ack_out;
			assign cnt_set_en = ack_in && ack_out;
			assign cnt_step = (cnt_incr_en ? sv2v_cast_7A7B7(inmask_ones) : sv2v_cast_7A7B7(OutW));
			always @(*) begin : cnt_set_logic
				cnt_set = 1'sb0;
				if (pos_with_input > sv2v_cast_7A7B7(OutW))
					cnt_set = pos_with_input - sv2v_cast_7A7B7(OutW);
			end
			wire [PtrW:1] sv2v_tmp_u_pos_cnt_o;
			always @(*) pos_q = sv2v_tmp_u_pos_cnt_o;
			prim_count #(
				.Width(PtrW),
				.ResetValue(1'sb0)
			) u_pos(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.clr_i(flush_done),
				.set_i(cnt_set_en),
				.set_cnt_i(cnt_set),
				.incr_en_i(cnt_incr_en),
				.decr_en_i(cnt_decr_en),
				.step_i(cnt_step),
				.cnt_o(sv2v_tmp_u_pos_cnt_o),
				.err_o(err_o)
			);
		end
	endgenerate
	function automatic [IdxW - 1:0] sv2v_cast_ADF40;
		input reg [IdxW - 1:0] inp;
		sv2v_cast_ADF40 = inp;
	endfunction
	always @(*) begin
		lod_idx = 0;
		begin : sv2v_autoblock_2
			reg signed [31:0] i;
			for (i = InW - 1; i >= 0; i = i - 1)
				if (mask_i[i] == 1'b1)
					lod_idx = sv2v_cast_ADF40($unsigned(i));
		end
	end
	assign ack_in = valid_i & ready_o;
	assign ack_out = valid_o & ready_i;
	assign shiftr_data = (valid_i ? data_i >> lod_idx : {InW {1'sb0}});
	assign shiftr_mask = (valid_i ? mask_i >> lod_idx : {InW {1'sb0}});
	function automatic [ConcatW - 1:0] sv2v_cast_2EE66;
		input reg [ConcatW - 1:0] inp;
		sv2v_cast_2EE66 = inp;
	endfunction
	assign shiftl_data = sv2v_cast_2EE66(shiftr_data) << pos_q;
	assign shiftl_mask = sv2v_cast_2EE66(shiftr_mask) << pos_q;
	assign concat_data = {{InW {1'b0}}, stored_data & stored_mask} | (shiftl_data & shiftl_mask);
	assign concat_mask = {{InW {1'b0}}, stored_mask} | shiftl_mask;
	reg [Width - 1:0] stored_data_next;
	reg [Width - 1:0] stored_mask_next;
	always @(*)
		case ({ack_in, ack_out})
			2'b00: begin
				stored_data_next = stored_data;
				stored_mask_next = stored_mask;
			end
			2'b01: begin
				stored_data_next = {{OutW {1'b0}}, stored_data[Width - 1:OutW]};
				stored_mask_next = {{OutW {1'b0}}, stored_mask[Width - 1:OutW]};
			end
			2'b10: begin
				stored_data_next = concat_data[0+:Width];
				stored_mask_next = concat_mask[0+:Width];
			end
			2'b11: begin
				stored_data_next = concat_data[ConcatW - 1:OutW];
				stored_mask_next = concat_mask[ConcatW - 1:OutW];
			end
			default: begin
				stored_data_next = stored_data;
				stored_mask_next = stored_mask;
			end
		endcase
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			stored_data <= 1'sb0;
			stored_mask <= 1'sb0;
		end
		else if (flush_done) begin
			stored_data <= 1'sb0;
			stored_mask <= 1'sb0;
		end
		else begin
			stored_data <= stored_data_next;
			stored_mask <= stored_mask_next;
		end
	reg flush_st;
	reg flush_st_next;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			flush_st <= 1'd0;
		else
			flush_st <= flush_st_next;
	always @(*) begin
		flush_st_next = 1'd0;
		flush_valid = 1'b0;
		flush_done = 1'b0;
		case (flush_st)
			1'd0:
				if (flush_i)
					flush_st_next = 1'd1;
				else
					flush_st_next = 1'd0;
			1'd1:
				if (pos_q == {PtrW {1'sb0}}) begin
					flush_st_next = 1'd0;
					flush_valid = 1'b0;
					flush_done = 1'b1;
				end
				else begin
					flush_st_next = 1'd1;
					flush_valid = 1'b1;
					flush_done = 1'b0;
				end
			default: begin
				flush_st_next = 1'd0;
				flush_valid = 1'b0;
				flush_done = 1'b0;
			end
		endcase
	end
	assign flush_done_o = flush_done;
	assign valid_next = (sv2v_cast_32_signed(pos_q) >= OutW ? 1'b1 : flush_valid);
	assign ready_next = sv2v_cast_32_signed(pos_q) <= OutW;
	assign valid_o = valid_next;
	assign data_o = stored_data[OutW - 1:0];
	assign mask_o = stored_mask[OutW - 1:0];
	assign ready_o = ready_next;
	generate
		if (HintByteData != 0) begin : g_byte_assert
			genvar i;
		end
	endgenerate
endmodule
module prim_packer_fifo (
	clk_i,
	rst_ni,
	clr_i,
	wvalid_i,
	wdata_i,
	wready_o,
	rvalid_o,
	rdata_o,
	rready_i,
	depth_o
);
	parameter signed [31:0] InW = 32;
	parameter signed [31:0] OutW = 8;
	parameter [0:0] ClearOnRead = 1'b1;
	localparam signed [31:0] MaxW = (InW > OutW ? InW : OutW);
	localparam signed [31:0] MinW = (InW < OutW ? InW : OutW);
	localparam signed [31:0] DepthW = $clog2(MaxW / MinW);
	input wire clk_i;
	input wire rst_ni;
	input wire clr_i;
	input wire wvalid_i;
	input wire [InW - 1:0] wdata_i;
	output wire wready_o;
	output wire rvalid_o;
	output wire [OutW - 1:0] rdata_o;
	input wire rready_i;
	output wire [DepthW:0] depth_o;
	localparam [31:0] WidthRatio = MaxW / MinW;
	localparam [DepthW:0] FullDepth = WidthRatio[DepthW:0];
	wire load_data;
	wire clear_data;
	wire clear_status;
	reg [DepthW:0] depth_q;
	wire [DepthW:0] depth_d;
	reg [MaxW - 1:0] data_q;
	wire [MaxW - 1:0] data_d;
	reg clr_q;
	wire clr_d;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			depth_q <= 1'sb0;
			data_q <= 1'sb0;
			clr_q <= 1'b1;
		end
		else begin
			depth_q <= depth_d;
			data_q <= data_d;
			clr_q <= clr_d;
		end
	assign clr_d = clr_i;
	assign depth_o = depth_q;
	generate
		if (InW < OutW) begin : gen_pack_mode
			wire [MaxW - 1:0] wdata_shifted;
			assign wdata_shifted = {{OutW - InW {1'b0}}, wdata_i} << (depth_q * InW);
			assign clear_status = (rready_i && rvalid_o) || clr_q;
			assign clear_data = (ClearOnRead && clear_status) || clr_q;
			assign load_data = wvalid_i && wready_o;
			assign depth_d = (clear_status ? {(DepthW >= 0 ? DepthW + 1 : 1 - DepthW) {1'sb0}} : (load_data ? depth_q + 1 : depth_q));
			assign data_d = (clear_data ? {MaxW {1'sb0}} : (load_data ? wdata_shifted | (depth_q == 0 ? {MaxW {1'sb0}} : data_q) : data_q));
			assign wready_o = (depth_q != FullDepth) && !clr_q;
			assign rdata_o = data_q;
			assign rvalid_o = (depth_q == FullDepth) && !clr_q;
		end
		else begin : gen_unpack_mode
			wire [MaxW - 1:0] rdata_shifted;
			wire pull_data;
			reg [DepthW:0] ptr_q;
			wire [DepthW:0] ptr_d;
			wire [DepthW:0] lsb_is_one;
			wire [DepthW:0] max_value;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					ptr_q <= 1'sb0;
				else
					ptr_q <= ptr_d;
			assign lsb_is_one = {{DepthW {1'b0}}, 1'b1};
			assign max_value = FullDepth;
			assign rdata_shifted = data_q >> (ptr_q * OutW);
			assign clear_status = (rready_i && (depth_q == lsb_is_one)) || clr_q;
			assign clear_data = (ClearOnRead && clear_status) || clr_q;
			assign load_data = wvalid_i && wready_o;
			assign pull_data = rvalid_o && rready_i;
			assign depth_d = (clear_status ? {(DepthW >= 0 ? DepthW + 1 : 1 - DepthW) {1'sb0}} : (load_data ? max_value : (pull_data ? depth_q - 1 : depth_q)));
			assign ptr_d = (clear_status ? {(DepthW >= 0 ? DepthW + 1 : 1 - DepthW) {1'sb0}} : (pull_data ? ptr_q + 1 : ptr_q));
			assign data_d = (clear_data ? {MaxW {1'sb0}} : (load_data ? wdata_i : data_q));
			assign wready_o = (depth_q == {(DepthW >= 0 ? DepthW + 1 : 1 - DepthW) {1'sb0}}) && !clr_q;
			assign rdata_o = rdata_shifted[OutW - 1:0];
			assign rvalid_o = (depth_q != {(DepthW >= 0 ? DepthW + 1 : 1 - DepthW) {1'sb0}}) && !clr_q;
			if (InW > OutW) begin : gen_unused
				wire [(MaxW - MinW) - 1:0] unused_rdata_shifted;
				assign unused_rdata_shifted = rdata_shifted[MaxW - 1:MinW];
			end
		end
	endgenerate
endmodule
module prim_present (
	data_i,
	key_i,
	idx_i,
	data_o,
	key_o,
	idx_o
);
	parameter signed [31:0] DataWidth = 64;
	parameter signed [31:0] KeyWidth = 128;
	parameter signed [31:0] NumRounds = 31;
	parameter signed [31:0] NumPhysRounds = NumRounds;
	parameter [0:0] Decrypt = 0;
	input [DataWidth - 1:0] data_i;
	input [KeyWidth - 1:0] key_i;
	input [4:0] idx_i;
	output wire [DataWidth - 1:0] data_o;
	output wire [KeyWidth - 1:0] key_o;
	output wire [4:0] idx_o;
	wire [(NumPhysRounds >= 0 ? ((NumPhysRounds + 1) * DataWidth) - 1 : ((1 - NumPhysRounds) * DataWidth) + ((NumPhysRounds * DataWidth) - 1)):(NumPhysRounds >= 0 ? 0 : NumPhysRounds * DataWidth)] data_state;
	wire [(NumPhysRounds >= 0 ? ((NumPhysRounds + 1) * KeyWidth) - 1 : ((1 - NumPhysRounds) * KeyWidth) + ((NumPhysRounds * KeyWidth) - 1)):(NumPhysRounds >= 0 ? 0 : NumPhysRounds * KeyWidth)] round_key;
	wire [(NumPhysRounds >= 0 ? ((NumPhysRounds + 1) * 5) - 1 : ((1 - NumPhysRounds) * 5) + ((NumPhysRounds * 5) - 1)):(NumPhysRounds >= 0 ? 0 : NumPhysRounds * 5)] round_idx;
	assign data_state[(NumPhysRounds >= 0 ? 0 : NumPhysRounds) * DataWidth+:DataWidth] = data_i;
	assign round_key[(NumPhysRounds >= 0 ? 0 : NumPhysRounds) * KeyWidth+:KeyWidth] = key_i;
	assign round_idx[(NumPhysRounds >= 0 ? 0 : NumPhysRounds) * 5+:5] = idx_i;
	genvar k;
	localparam [159:0] prim_cipher_pkg_PRESENT_PERM32 = 160'hfdde7f59c6ed5a5e5184dcd63d4942cc521c4100;
	localparam [159:0] prim_cipher_pkg_PRESENT_PERM32_INV = 160'hfeef37ace3f6ad2728c2ee6b16a4a1e629062080;
	localparam [383:0] prim_cipher_pkg_PRESENT_PERM64 = 384'hfef7cffae78ef6d74df2c70ceeb6cbeaa68ae69649e28608de75c7da6586d65545d24504ce34c3ca2482c61441c20400;
	localparam [383:0] prim_cipher_pkg_PRESENT_PERM64_INV = 384'hffbdf3beb9e37db5d33cb1c3fbadb2baa9a279a59238a182f79d71b69961759551349141f38d30b28920718510308100;
	localparam [63:0] prim_cipher_pkg_PRESENT_SBOX4 = 64'h21748fe3da09b65c;
	localparam [63:0] prim_cipher_pkg_PRESENT_SBOX4_INV = 64'ha970364bd21c8fe5;
	function automatic [31:0] prim_cipher_pkg_perm_32bit;
		input reg [31:0] state_in;
		input reg [159:0] perm;
		reg [31:0] state_out;
		begin
			begin : sv2v_autoblock_1
				reg signed [31:0] k;
				for (k = 0; k < 32; k = k + 1)
					state_out[perm[k * 5+:5]] = state_in[k];
			end
			prim_cipher_pkg_perm_32bit = state_out;
		end
	endfunction
	function automatic [63:0] prim_cipher_pkg_perm_64bit;
		input reg [63:0] state_in;
		input reg [383:0] perm;
		reg [63:0] state_out;
		begin
			begin : sv2v_autoblock_2
				reg signed [31:0] k;
				for (k = 0; k < 64; k = k + 1)
					state_out[perm[k * 6+:6]] = state_in[k];
			end
			prim_cipher_pkg_perm_64bit = state_out;
		end
	endfunction
	function automatic [127:0] prim_cipher_pkg_present_inv_update_key128;
		input reg [127:0] key_in;
		input reg [4:0] round_idx;
		reg [127:0] key_out;
		begin
			key_out = key_in;
			key_out[66:62] = key_out[66:62] ^ round_idx;
			key_out[123-:4] = prim_cipher_pkg_PRESENT_SBOX4_INV[key_out[123-:4] * 4+:4];
			key_out[127-:4] = prim_cipher_pkg_PRESENT_SBOX4_INV[key_out[127-:4] * 4+:4];
			key_out = {key_out[60:0], key_out[127:61]};
			prim_cipher_pkg_present_inv_update_key128 = key_out;
		end
	endfunction
	function automatic [63:0] prim_cipher_pkg_present_inv_update_key64;
		input reg [63:0] key_in;
		input reg [4:0] round_idx;
		reg [63:0] key_out;
		begin
			key_out = key_in;
			key_out[19:15] = key_out[19:15] ^ round_idx;
			key_out[63-:4] = prim_cipher_pkg_PRESENT_SBOX4_INV[key_out[63-:4] * 4+:4];
			key_out = {key_out[60:0], key_out[63:61]};
			prim_cipher_pkg_present_inv_update_key64 = key_out;
		end
	endfunction
	function automatic [79:0] prim_cipher_pkg_present_inv_update_key80;
		input reg [79:0] key_in;
		input reg [4:0] round_idx;
		reg [79:0] key_out;
		begin
			key_out = key_in;
			key_out[19:15] = key_out[19:15] ^ round_idx;
			key_out[79-:4] = prim_cipher_pkg_PRESENT_SBOX4_INV[key_out[79-:4] * 4+:4];
			key_out = {key_out[60:0], key_out[79:61]};
			prim_cipher_pkg_present_inv_update_key80 = key_out;
		end
	endfunction
	function automatic [127:0] prim_cipher_pkg_present_update_key128;
		input reg [127:0] key_in;
		input reg [4:0] round_idx;
		reg [127:0] key_out;
		begin
			key_out = {key_in[66:0], key_in[127:67]};
			key_out[127-:4] = prim_cipher_pkg_PRESENT_SBOX4[key_out[127-:4] * 4+:4];
			key_out[123-:4] = prim_cipher_pkg_PRESENT_SBOX4[key_out[123-:4] * 4+:4];
			key_out[66:62] = key_out[66:62] ^ round_idx;
			prim_cipher_pkg_present_update_key128 = key_out;
		end
	endfunction
	function automatic [63:0] prim_cipher_pkg_present_update_key64;
		input reg [63:0] key_in;
		input reg [4:0] round_idx;
		reg [63:0] key_out;
		begin
			key_out = {key_in[2:0], key_in[63:3]};
			key_out[63-:4] = prim_cipher_pkg_PRESENT_SBOX4[key_out[63-:4] * 4+:4];
			key_out[19:15] = key_out[19:15] ^ round_idx;
			prim_cipher_pkg_present_update_key64 = key_out;
		end
	endfunction
	function automatic [79:0] prim_cipher_pkg_present_update_key80;
		input reg [79:0] key_in;
		input reg [4:0] round_idx;
		reg [79:0] key_out;
		begin
			key_out = {key_in[18:0], key_in[79:19]};
			key_out[79-:4] = prim_cipher_pkg_PRESENT_SBOX4[key_out[79-:4] * 4+:4];
			key_out[19:15] = key_out[19:15] ^ round_idx;
			prim_cipher_pkg_present_update_key80 = key_out;
		end
	endfunction
	function automatic [7:0] prim_cipher_pkg_sbox4_8bit;
		input reg [7:0] state_in;
		input reg [63:0] sbox4;
		reg [7:0] state_out;
		begin
			begin : sv2v_autoblock_3
				reg signed [31:0] k;
				for (k = 0; k < 2; k = k + 1)
					state_out[k * 4+:4] = sbox4[state_in[k * 4+:4] * 4+:4];
			end
			prim_cipher_pkg_sbox4_8bit = state_out;
		end
	endfunction
	function automatic [31:0] prim_cipher_pkg_sbox4_32bit;
		input reg [31:0] state_in;
		input reg [63:0] sbox4;
		reg [31:0] state_out;
		begin
			begin : sv2v_autoblock_4
				reg signed [31:0] k;
				for (k = 0; k < 4; k = k + 1)
					state_out[k * 8+:8] = prim_cipher_pkg_sbox4_8bit(state_in[k * 8+:8], sbox4);
			end
			prim_cipher_pkg_sbox4_32bit = state_out;
		end
	endfunction
	function automatic [63:0] prim_cipher_pkg_sbox4_64bit;
		input reg [63:0] state_in;
		input reg [63:0] sbox4;
		reg [63:0] state_out;
		begin
			begin : sv2v_autoblock_5
				reg signed [31:0] k;
				for (k = 0; k < 8; k = k + 1)
					state_out[k * 8+:8] = prim_cipher_pkg_sbox4_8bit(state_in[k * 8+:8], sbox4);
			end
			prim_cipher_pkg_sbox4_64bit = state_out;
		end
	endfunction
	generate
		for (k = 0; k < NumPhysRounds; k = k + 1) begin : gen_round
			wire [DataWidth - 1:0] data_state_xor;
			wire [DataWidth - 1:0] data_state_sbox;
			assign data_state_xor = data_state[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * DataWidth+:DataWidth] ^ round_key[((NumPhysRounds >= 0 ? k : NumPhysRounds - k) * KeyWidth) + ((KeyWidth - 1) >= (KeyWidth - DataWidth) ? KeyWidth - 1 : ((KeyWidth - 1) + ((KeyWidth - 1) >= (KeyWidth - DataWidth) ? ((KeyWidth - 1) - (KeyWidth - DataWidth)) + 1 : ((KeyWidth - DataWidth) - (KeyWidth - 1)) + 1)) - 1)-:((KeyWidth - 1) >= (KeyWidth - DataWidth) ? ((KeyWidth - 1) - (KeyWidth - DataWidth)) + 1 : ((KeyWidth - DataWidth) - (KeyWidth - 1)) + 1)];
			if (Decrypt) begin : gen_dec
				assign round_idx[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * 5+:5] = round_idx[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * 5+:5] - 1'b1;
				if (DataWidth == 64) begin : gen_d64
					assign data_state_sbox = prim_cipher_pkg_perm_64bit(data_state_xor, prim_cipher_pkg_PRESENT_PERM64_INV);
					assign data_state[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * DataWidth+:DataWidth] = prim_cipher_pkg_sbox4_64bit(data_state_sbox, prim_cipher_pkg_PRESENT_SBOX4_INV);
				end
				else begin : gen_d32
					assign data_state_sbox = prim_cipher_pkg_perm_32bit(data_state_xor, prim_cipher_pkg_PRESENT_PERM32_INV);
					assign data_state[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * DataWidth+:DataWidth] = prim_cipher_pkg_sbox4_32bit(data_state_sbox, prim_cipher_pkg_PRESENT_SBOX4_INV);
				end
				if (KeyWidth == 128) begin : gen_k128
					assign round_key[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * KeyWidth+:KeyWidth] = prim_cipher_pkg_present_inv_update_key128(round_key[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * KeyWidth+:KeyWidth], round_idx[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * 5+:5]);
				end
				else if (KeyWidth == 80) begin : gen_k80
					assign round_key[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * KeyWidth+:KeyWidth] = prim_cipher_pkg_present_inv_update_key80(round_key[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * KeyWidth+:KeyWidth], round_idx[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * 5+:5]);
				end
				else begin : gen_k64
					assign round_key[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * KeyWidth+:KeyWidth] = prim_cipher_pkg_present_inv_update_key64(round_key[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * KeyWidth+:KeyWidth], round_idx[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * 5+:5]);
				end
			end
			else begin : gen_enc
				assign round_idx[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * 5+:5] = round_idx[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * 5+:5] + 1'b1;
				if (DataWidth == 64) begin : gen_d64
					assign data_state_sbox = prim_cipher_pkg_sbox4_64bit(data_state_xor, prim_cipher_pkg_PRESENT_SBOX4);
					assign data_state[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * DataWidth+:DataWidth] = prim_cipher_pkg_perm_64bit(data_state_sbox, prim_cipher_pkg_PRESENT_PERM64);
				end
				else begin : gen_d32
					assign data_state_sbox = prim_cipher_pkg_sbox4_32bit(data_state_xor, prim_cipher_pkg_PRESENT_SBOX4);
					assign data_state[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * DataWidth+:DataWidth] = prim_cipher_pkg_perm_32bit(data_state_sbox, prim_cipher_pkg_PRESENT_PERM32);
				end
				if (KeyWidth == 128) begin : gen_k128
					assign round_key[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * KeyWidth+:KeyWidth] = prim_cipher_pkg_present_update_key128(round_key[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * KeyWidth+:KeyWidth], round_idx[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * 5+:5]);
				end
				else if (KeyWidth == 80) begin : gen_k80
					assign round_key[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * KeyWidth+:KeyWidth] = prim_cipher_pkg_present_update_key80(round_key[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * KeyWidth+:KeyWidth], round_idx[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * 5+:5]);
				end
				else begin : gen_k64
					assign round_key[(NumPhysRounds >= 0 ? k + 1 : NumPhysRounds - (k + 1)) * KeyWidth+:KeyWidth] = prim_cipher_pkg_present_update_key64(round_key[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * KeyWidth+:KeyWidth], round_idx[(NumPhysRounds >= 0 ? k : NumPhysRounds - k) * 5+:5]);
				end
			end
		end
	endgenerate
	localparam signed [31:0] LastRoundIdx = ((Decrypt != 0) || (NumRounds == 31) ? 0 : NumRounds + 1);
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	assign data_o = (sv2v_cast_32_signed(idx_o) == LastRoundIdx ? data_state[(NumPhysRounds >= 0 ? NumPhysRounds : NumPhysRounds - NumPhysRounds) * DataWidth+:DataWidth] ^ round_key[((NumPhysRounds >= 0 ? NumPhysRounds : NumPhysRounds - NumPhysRounds) * KeyWidth) + ((KeyWidth - 1) >= (KeyWidth - DataWidth) ? KeyWidth - 1 : ((KeyWidth - 1) + ((KeyWidth - 1) >= (KeyWidth - DataWidth) ? ((KeyWidth - 1) - (KeyWidth - DataWidth)) + 1 : ((KeyWidth - DataWidth) - (KeyWidth - 1)) + 1)) - 1)-:((KeyWidth - 1) >= (KeyWidth - DataWidth) ? ((KeyWidth - 1) - (KeyWidth - DataWidth)) + 1 : ((KeyWidth - DataWidth) - (KeyWidth - 1)) + 1)] : data_state[(NumPhysRounds >= 0 ? NumPhysRounds : NumPhysRounds - NumPhysRounds) * DataWidth+:DataWidth]);
	assign key_o = round_key[(NumPhysRounds >= 0 ? NumPhysRounds : NumPhysRounds - NumPhysRounds) * KeyWidth+:KeyWidth];
	assign idx_o = round_idx[(NumPhysRounds >= 0 ? NumPhysRounds : NumPhysRounds - NumPhysRounds) * 5+:5];
endmodule
module prim_prince (
	clk_i,
	rst_ni,
	valid_i,
	data_i,
	key_i,
	dec_i,
	valid_o,
	data_o
);
	parameter signed [31:0] DataWidth = 64;
	parameter signed [31:0] KeyWidth = 128;
	parameter signed [31:0] NumRoundsHalf = 5;
	parameter [0:0] UseOldKeySched = 1'b0;
	parameter [0:0] HalfwayDataReg = 1'b0;
	parameter [0:0] HalfwayKeyReg = 1'b0;
	input clk_i;
	input rst_ni;
	input valid_i;
	input [DataWidth - 1:0] data_i;
	input [KeyWidth - 1:0] key_i;
	input dec_i;
	output wire valid_o;
	output reg [DataWidth - 1:0] data_o;
	reg [DataWidth - 1:0] k0;
	reg [DataWidth - 1:0] k0_prime_d;
	reg [DataWidth - 1:0] k1_d;
	reg [DataWidth - 1:0] k0_new_d;
	reg [DataWidth - 1:0] k0_prime_q;
	reg [DataWidth - 1:0] k1_q;
	reg [DataWidth - 1:0] k0_new_q;
	localparam [63:0] prim_cipher_pkg_PRINCE_ALPHA_CONST = 64'hc0ac29b7c97c50dd;
	always @(*) begin : p_key_expansion
		k0 = key_i[(2 * DataWidth) - 1:DataWidth];
		k0_prime_d = {k0[0], k0[DataWidth - 1:2], k0[DataWidth - 1] ^ k0[1]};
		k1_d = key_i[DataWidth - 1:0];
		if (dec_i) begin
			k0 = k0_prime_d;
			k0_prime_d = key_i[(2 * DataWidth) - 1:DataWidth];
			k1_d = k1_d ^ prim_cipher_pkg_PRINCE_ALPHA_CONST[DataWidth - 1:0];
		end
	end
	generate
		if (UseOldKeySched) begin : gen_legacy_keyschedule
			wire [DataWidth:1] sv2v_tmp_A4614;
			assign sv2v_tmp_A4614 = k1_d;
			always @(*) k0_new_d = sv2v_tmp_A4614;
		end
		else begin : gen_new_keyschedule
			always @(*) begin : p_new_keyschedule_k0_alpha
				k0_new_d = key_i[(2 * DataWidth) - 1:DataWidth];
				if (dec_i)
					k0_new_d = k0_new_d ^ prim_cipher_pkg_PRINCE_ALPHA_CONST[DataWidth - 1:0];
			end
		end
		if (HalfwayKeyReg) begin : gen_key_reg
			always @(posedge clk_i or negedge rst_ni) begin : p_key_reg
				if (!rst_ni) begin
					k1_q <= 1'sb0;
					k0_prime_q <= 1'sb0;
					k0_new_q <= 1'sb0;
				end
				else if (valid_i) begin
					k1_q <= k1_d;
					k0_prime_q <= k0_prime_d;
					k0_new_q <= k0_new_d;
				end
			end
		end
		else begin : gen_no_key_reg
			wire [DataWidth:1] sv2v_tmp_BDE31;
			assign sv2v_tmp_BDE31 = k1_d;
			always @(*) k1_q = sv2v_tmp_BDE31;
			wire [DataWidth:1] sv2v_tmp_ECEAB;
			assign sv2v_tmp_ECEAB = k0_prime_d;
			always @(*) k0_prime_q = sv2v_tmp_ECEAB;
			wire [DataWidth:1] sv2v_tmp_CB365;
			assign sv2v_tmp_CB365 = k0_new_d;
			always @(*) k0_new_q = sv2v_tmp_CB365;
		end
	endgenerate
	reg [(((NumRoundsHalf * 2) + 1) >= 0 ? (((NumRoundsHalf * 2) + 2) * DataWidth) - 1 : ((1 - ((NumRoundsHalf * 2) + 1)) * DataWidth) + ((((NumRoundsHalf * 2) + 1) * DataWidth) - 1)):(((NumRoundsHalf * 2) + 1) >= 0 ? 0 : ((NumRoundsHalf * 2) + 1) * DataWidth)] data_state;
	localparam [767:0] prim_cipher_pkg_PRINCE_ROUND_CONST = 768'hc0ac29b7c97c50ddd3b5a399ca0c239964a51195e0e3610dc882d32f25323c5485840851f1ac43aa7ef84f78fd955cb1be5466cf34e90c6c452821e638d01377082efa98ec4e6c89a4093822299f31d013198a2e037073440000000000000000;
	always @(*) begin : p_pre_round_xor
		data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? 0 : (NumRoundsHalf * 2) + 1) * DataWidth+:DataWidth] = data_i ^ k0;
		data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? 0 : (NumRoundsHalf * 2) + 1) * DataWidth+:DataWidth] = data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? 0 : (NumRoundsHalf * 2) + 1) * DataWidth+:DataWidth] ^ k1_d;
		data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? 0 : (NumRoundsHalf * 2) + 1) * DataWidth+:DataWidth] = data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? 0 : (NumRoundsHalf * 2) + 1) * DataWidth+:DataWidth] ^ prim_cipher_pkg_PRINCE_ROUND_CONST[DataWidth - 1-:DataWidth];
	end
	genvar k;
	localparam [63:0] prim_cipher_pkg_PRINCE_SBOX4 = 64'h4d5e087619ca23fb;
	localparam [63:0] prim_cipher_pkg_PRINCE_SHIFT_ROWS64 = 64'hfa50b61c72d83e94;
	localparam [15:0] prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST0 = 16'h7bde;
	localparam [15:0] prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST1 = 16'hbde7;
	localparam [15:0] prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST2 = 16'hde7b;
	localparam [15:0] prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST3 = 16'he7bd;
	function automatic [3:0] prim_cipher_pkg_prince_nibble_red16;
		input reg [15:0] vect;
		prim_cipher_pkg_prince_nibble_red16 = ((vect[0+:4] ^ vect[4+:4]) ^ vect[8+:4]) ^ vect[12+:4];
	endfunction
	function automatic [31:0] prim_cipher_pkg_prince_mult_prime_32bit;
		input reg [31:0] state_in;
		reg [31:0] state_out;
		begin
			state_out[0+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[0+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST3);
			state_out[4+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[0+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST2);
			state_out[8+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[0+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST1);
			state_out[12+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[0+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST0);
			state_out[16+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[16+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST0);
			state_out[20+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[16+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST3);
			state_out[24+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[16+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST2);
			state_out[28+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[16+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST1);
			prim_cipher_pkg_prince_mult_prime_32bit = state_out;
		end
	endfunction
	function automatic [63:0] prim_cipher_pkg_prince_mult_prime_64bit;
		input reg [63:0] state_in;
		reg [63:0] state_out;
		begin
			state_out[0+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[0+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST3);
			state_out[4+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[0+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST2);
			state_out[8+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[0+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST1);
			state_out[12+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[0+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST0);
			state_out[16+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[16+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST0);
			state_out[20+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[16+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST3);
			state_out[24+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[16+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST2);
			state_out[28+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[16+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST1);
			state_out[32+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[32+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST0);
			state_out[36+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[32+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST3);
			state_out[40+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[32+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST2);
			state_out[44+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[32+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST1);
			state_out[48+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[48+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST3);
			state_out[52+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[48+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST2);
			state_out[56+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[48+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST1);
			state_out[60+:4] = prim_cipher_pkg_prince_nibble_red16(state_in[48+:16] & prim_cipher_pkg_PRINCE_SHIFT_ROWS_CONST0);
			prim_cipher_pkg_prince_mult_prime_64bit = state_out;
		end
	endfunction
	function automatic [31:0] prim_cipher_pkg_prince_shiftrows_32bit;
		input reg [31:0] state_in;
		input reg [63:0] shifts;
		reg [31:0] state_out;
		begin
			begin : sv2v_autoblock_1
				reg signed [31:0] k;
				for (k = 0; k < 16; k = k + 1)
					state_out[k * 2+:2] = state_in[shifts[k * 4+:4] * 2+:2];
			end
			prim_cipher_pkg_prince_shiftrows_32bit = state_out;
		end
	endfunction
	function automatic [63:0] prim_cipher_pkg_prince_shiftrows_64bit;
		input reg [63:0] state_in;
		input reg [63:0] shifts;
		reg [63:0] state_out;
		begin
			begin : sv2v_autoblock_2
				reg signed [31:0] k;
				for (k = 0; k < 16; k = k + 1)
					state_out[k * 4+:4] = state_in[shifts[k * 4+:4] * 4+:4];
			end
			prim_cipher_pkg_prince_shiftrows_64bit = state_out;
		end
	endfunction
	function automatic [7:0] prim_cipher_pkg_sbox4_8bit;
		input reg [7:0] state_in;
		input reg [63:0] sbox4;
		reg [7:0] state_out;
		begin
			begin : sv2v_autoblock_3
				reg signed [31:0] k;
				for (k = 0; k < 2; k = k + 1)
					state_out[k * 4+:4] = sbox4[state_in[k * 4+:4] * 4+:4];
			end
			prim_cipher_pkg_sbox4_8bit = state_out;
		end
	endfunction
	function automatic [31:0] prim_cipher_pkg_sbox4_32bit;
		input reg [31:0] state_in;
		input reg [63:0] sbox4;
		reg [31:0] state_out;
		begin
			begin : sv2v_autoblock_4
				reg signed [31:0] k;
				for (k = 0; k < 4; k = k + 1)
					state_out[k * 8+:8] = prim_cipher_pkg_sbox4_8bit(state_in[k * 8+:8], sbox4);
			end
			prim_cipher_pkg_sbox4_32bit = state_out;
		end
	endfunction
	function automatic [63:0] prim_cipher_pkg_sbox4_64bit;
		input reg [63:0] state_in;
		input reg [63:0] sbox4;
		reg [63:0] state_out;
		begin
			begin : sv2v_autoblock_5
				reg signed [31:0] k;
				for (k = 0; k < 8; k = k + 1)
					state_out[k * 8+:8] = prim_cipher_pkg_sbox4_8bit(state_in[k * 8+:8], sbox4);
			end
			prim_cipher_pkg_sbox4_64bit = state_out;
		end
	endfunction
	generate
		for (k = 1; k <= NumRoundsHalf; k = k + 1) begin : gen_fwd_pass
			reg [DataWidth - 1:0] data_state_round;
			if (DataWidth == 64) begin : gen_fwd_d64
				always @(*) begin : p_fwd_d64
					data_state_round = prim_cipher_pkg_sbox4_64bit(data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? k - 1 : ((NumRoundsHalf * 2) + 1) - (k - 1)) * DataWidth+:DataWidth], prim_cipher_pkg_PRINCE_SBOX4);
					data_state_round = prim_cipher_pkg_prince_mult_prime_64bit(data_state_round);
					data_state_round = prim_cipher_pkg_prince_shiftrows_64bit(data_state_round, prim_cipher_pkg_PRINCE_SHIFT_ROWS64);
				end
			end
			else begin : gen_fwd_d32
				always @(*) begin : p_fwd_d32
					data_state_round = prim_cipher_pkg_sbox4_32bit(data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? k - 1 : ((NumRoundsHalf * 2) + 1) - (k - 1)) * DataWidth+:DataWidth], prim_cipher_pkg_PRINCE_SBOX4);
					data_state_round = prim_cipher_pkg_prince_mult_prime_32bit(data_state_round);
					data_state_round = prim_cipher_pkg_prince_shiftrows_32bit(data_state_round, prim_cipher_pkg_PRINCE_SHIFT_ROWS64);
				end
			end
			wire [DataWidth - 1:0] data_state_xor;
			assign data_state_xor = data_state_round ^ prim_cipher_pkg_PRINCE_ROUND_CONST[(k * 64) + (DataWidth - 1)-:DataWidth];
			if ((k % 2) == 1) begin : gen_fwd_key_odd
				wire [DataWidth * 1:1] sv2v_tmp_6C890;
				assign sv2v_tmp_6C890 = data_state_xor ^ k0_new_d;
				always @(*) data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? k : ((NumRoundsHalf * 2) + 1) - k) * DataWidth+:DataWidth] = sv2v_tmp_6C890;
			end
			else begin : gen_fwd_key_even
				wire [DataWidth * 1:1] sv2v_tmp_9028E;
				assign sv2v_tmp_9028E = data_state_xor ^ k1_d;
				always @(*) data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? k : ((NumRoundsHalf * 2) + 1) - k) * DataWidth+:DataWidth] = sv2v_tmp_9028E;
			end
		end
	endgenerate
	reg [DataWidth - 1:0] data_state_middle_d;
	reg [DataWidth - 1:0] data_state_middle_q;
	reg [DataWidth - 1:0] data_state_middle;
	localparam [63:0] prim_cipher_pkg_PRINCE_SBOX4_INV = 64'h1ce5046a98df237b;
	generate
		if (DataWidth == 64) begin : gen_middle_d64
			always @(*) begin : p_middle_d64
				data_state_middle_d = prim_cipher_pkg_sbox4_64bit(data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? NumRoundsHalf : ((NumRoundsHalf * 2) + 1) - NumRoundsHalf) * DataWidth+:DataWidth], prim_cipher_pkg_PRINCE_SBOX4);
				data_state_middle = prim_cipher_pkg_prince_mult_prime_64bit(data_state_middle_q);
				data_state_middle = prim_cipher_pkg_sbox4_64bit(data_state_middle, prim_cipher_pkg_PRINCE_SBOX4_INV);
			end
		end
		else begin : gen_middle_d32
			always @(*) begin : p_middle_d32
				data_state_middle_d = prim_cipher_pkg_sbox4_32bit(data_state_middle[NumRoundsHalf], prim_cipher_pkg_PRINCE_SBOX4);
				data_state_middle = prim_cipher_pkg_prince_mult_prime_32bit(data_state_middle_q);
				data_state_middle = prim_cipher_pkg_sbox4_32bit(data_state_middle, prim_cipher_pkg_PRINCE_SBOX4_INV);
			end
		end
		if (HalfwayDataReg) begin : gen_data_reg
			reg valid_q;
			always @(posedge clk_i or negedge rst_ni) begin : p_data_reg
				if (!rst_ni) begin
					valid_q <= 1'b0;
					data_state_middle_q <= 1'sb0;
				end
				else begin
					valid_q <= valid_i;
					if (valid_i)
						data_state_middle_q <= data_state_middle_d;
				end
			end
			assign valid_o = valid_q;
		end
		else begin : gen_no_data_reg
			wire [DataWidth:1] sv2v_tmp_F6B27;
			assign sv2v_tmp_F6B27 = data_state_middle_d;
			always @(*) data_state_middle_q = sv2v_tmp_F6B27;
			assign valid_o = valid_i;
		end
	endgenerate
	wire [DataWidth * 1:1] sv2v_tmp_54D8E;
	assign sv2v_tmp_54D8E = data_state_middle;
	always @(*) data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? NumRoundsHalf + 1 : ((NumRoundsHalf * 2) + 1) - (NumRoundsHalf + 1)) * DataWidth+:DataWidth] = sv2v_tmp_54D8E;
	localparam [63:0] prim_cipher_pkg_PRINCE_SHIFT_ROWS64_INV = 64'hf258be147ad0369c;
	generate
		for (k = 1; k <= NumRoundsHalf; k = k + 1) begin : gen_bwd_pass
			wire [DataWidth - 1:0] data_state_xor0;
			wire [DataWidth - 1:0] data_state_xor1;
			if ((((NumRoundsHalf + k) + 1) % 2) == 1) begin : gen_bkwd_key_odd
				assign data_state_xor0 = data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? NumRoundsHalf + k : ((NumRoundsHalf * 2) + 1) - (NumRoundsHalf + k)) * DataWidth+:DataWidth] ^ k0_new_q;
			end
			else begin : gen_bkwd_key_even
				assign data_state_xor0 = data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? NumRoundsHalf + k : ((NumRoundsHalf * 2) + 1) - (NumRoundsHalf + k)) * DataWidth+:DataWidth] ^ k1_q;
			end
			assign data_state_xor1 = data_state_xor0 ^ prim_cipher_pkg_PRINCE_ROUND_CONST[(((10 - NumRoundsHalf) + k) * 64) + (DataWidth - 1)-:DataWidth];
			reg [DataWidth - 1:0] data_state_bwd;
			if (DataWidth == 64) begin : gen_bwd_d64
				always @(*) begin : p_bwd_d64
					data_state_bwd = prim_cipher_pkg_prince_shiftrows_64bit(data_state_xor1, prim_cipher_pkg_PRINCE_SHIFT_ROWS64_INV);
					data_state_bwd = prim_cipher_pkg_prince_mult_prime_64bit(data_state_bwd);
					data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? (NumRoundsHalf + k) + 1 : ((NumRoundsHalf * 2) + 1) - ((NumRoundsHalf + k) + 1)) * DataWidth+:DataWidth] = prim_cipher_pkg_sbox4_64bit(data_state_bwd, prim_cipher_pkg_PRINCE_SBOX4_INV);
				end
			end
			else begin : gen_bwd_d32
				always @(*) begin : p_bwd_d32
					data_state_bwd = prim_cipher_pkg_prince_shiftrows_32bit(data_state_xor1, prim_cipher_pkg_PRINCE_SHIFT_ROWS64_INV);
					data_state_bwd = prim_cipher_pkg_prince_mult_prime_32bit(data_state_bwd);
					data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? (NumRoundsHalf + k) + 1 : ((NumRoundsHalf * 2) + 1) - ((NumRoundsHalf + k) + 1)) * DataWidth+:DataWidth] = prim_cipher_pkg_sbox4_32bit(data_state_bwd, prim_cipher_pkg_PRINCE_SBOX4_INV);
				end
			end
		end
	endgenerate
	always @(*) begin : p_post_round_xor
		data_o = data_state[(((NumRoundsHalf * 2) + 1) >= 0 ? (2 * NumRoundsHalf) + 1 : ((NumRoundsHalf * 2) + 1) - ((2 * NumRoundsHalf) + 1)) * DataWidth+:DataWidth] ^ prim_cipher_pkg_PRINCE_ROUND_CONST[DataWidth + 703-:DataWidth];
		data_o = data_o ^ k1_q;
		data_o = data_o ^ k0_prime_q;
	end
endmodule
module prim_pulse_sync (
	clk_src_i,
	rst_src_ni,
	src_pulse_i,
	clk_dst_i,
	rst_dst_ni,
	dst_pulse_o
);
	input wire clk_src_i;
	input wire rst_src_ni;
	input wire src_pulse_i;
	input wire clk_dst_i;
	input wire rst_dst_ni;
	output wire dst_pulse_o;
	reg src_level;
	always @(posedge clk_src_i or negedge rst_src_ni)
		if (!rst_src_ni)
			src_level <= 1'b0;
		else
			src_level <= src_level ^ src_pulse_i;
	wire dst_level;
	prim_flop_2sync #(.Width(1)) prim_flop_2sync(
		.d_i(src_level),
		.clk_i(clk_dst_i),
		.rst_ni(rst_dst_ni),
		.q_o(dst_level)
	);
	reg dst_level_q;
	always @(posedge clk_dst_i or negedge rst_dst_ni)
		if (!rst_dst_ni)
			dst_level_q <= 1'b0;
		else
			dst_level_q <= dst_level;
	assign dst_pulse_o = dst_level_q ^ dst_level;
endmodule
module prim_ram_1p (
	clk_i,
	req_i,
	write_i,
	addr_i,
	wdata_i,
	wmask_i,
	rdata_o,
	cfg_i
);
	parameter signed [31:0] Width = 32;
	parameter signed [31:0] Depth = 128;
	parameter signed [31:0] DataBitsPerMask = 1;
	parameter MemInitFile = "";
	localparam signed [31:0] Aw = $clog2(Depth);
	input wire clk_i;
	input wire req_i;
	input wire write_i;
	input wire [Aw - 1:0] addr_i;
	input wire [Width - 1:0] wdata_i;
	input wire [Width - 1:0] wmask_i;
	output wire [Width - 1:0] rdata_o;
	input wire [9:0] cfg_i;
	parameter integer Impl = 32'sd0;
	generate
		if (Impl == 32'sd1) begin : gen_badbit
			prim_badbit_ram_1p #(
				.DataBitsPerMask(DataBitsPerMask),
				.Depth(Depth),
				.MemInitFile(MemInitFile),
				.Width(Width)
			) u_impl_badbit(
				.clk_i(clk_i),
				.req_i(req_i),
				.write_i(write_i),
				.addr_i(addr_i),
				.wdata_i(wdata_i),
				.wmask_i(wmask_i),
				.rdata_o(rdata_o)
			);
		end
		else begin : gen_generic
			prim_generic_ram_1p #(
				.DataBitsPerMask(DataBitsPerMask),
				.Depth(Depth),
				.MemInitFile(MemInitFile),
				.Width(Width)
			) u_impl_generic(
				.clk_i(clk_i),
				.req_i(req_i),
				.write_i(write_i),
				.addr_i(addr_i),
				.wdata_i(wdata_i),
				.wmask_i(wmask_i),
				.rdata_o(rdata_o),
				.cfg_i(cfg_i)
			);
		end
	endgenerate
endmodule
module prim_ram_1p_adv (
	clk_i,
	rst_ni,
	req_i,
	write_i,
	addr_i,
	wdata_i,
	wmask_i,
	rdata_o,
	rvalid_o,
	rerror_o,
	cfg_i
);
	parameter signed [31:0] Depth = 512;
	parameter signed [31:0] Width = 32;
	parameter signed [31:0] DataBitsPerMask = 1;
	parameter MemInitFile = "";
	parameter [0:0] EnableECC = 0;
	parameter [0:0] EnableParity = 0;
	parameter [0:0] EnableInputPipeline = 0;
	parameter [0:0] EnableOutputPipeline = 0;
	parameter [0:0] HammingECC = 0;
	function automatic integer prim_util_pkg_vbits;
		input integer value;
		prim_util_pkg_vbits = (value == 1 ? 1 : $clog2(value));
	endfunction
	localparam signed [31:0] Aw = prim_util_pkg_vbits(Depth);
	input clk_i;
	input rst_ni;
	input req_i;
	input write_i;
	input [Aw - 1:0] addr_i;
	input [Width - 1:0] wdata_i;
	input [Width - 1:0] wmask_i;
	output wire [Width - 1:0] rdata_o;
	output wire rvalid_o;
	output wire [1:0] rerror_o;
	input wire [9:0] cfg_i;
	localparam signed [31:0] ParWidth = (EnableParity ? Width / 8 : (!EnableECC ? 0 : (Width <= 4 ? 4 : (Width <= 11 ? 5 : (Width <= 26 ? 6 : (Width <= 57 ? 7 : (Width <= 120 ? 8 : 8)))))));
	localparam signed [31:0] TotalWidth = Width + ParWidth;
	localparam signed [31:0] LocalDataBitsPerMask = (EnableParity ? 9 : (EnableECC ? TotalWidth : DataBitsPerMask));
	reg req_q;
	wire req_d;
	reg write_q;
	wire write_d;
	reg [Aw - 1:0] addr_q;
	wire [Aw - 1:0] addr_d;
	reg [TotalWidth - 1:0] wdata_q;
	reg [TotalWidth - 1:0] wdata_d;
	reg [TotalWidth - 1:0] wmask_q;
	reg [TotalWidth - 1:0] wmask_d;
	reg rvalid_q;
	wire rvalid_d;
	reg rvalid_sram_q;
	reg [Width - 1:0] rdata_q;
	reg [Width - 1:0] rdata_d;
	wire [TotalWidth - 1:0] rdata_sram;
	reg [1:0] rerror_q;
	reg [1:0] rerror_d;
	prim_ram_1p #(
		.MemInitFile(MemInitFile),
		.Width(TotalWidth),
		.Depth(Depth),
		.DataBitsPerMask(LocalDataBitsPerMask)
	) u_mem(
		.clk_i(clk_i),
		.req_i(req_q),
		.write_i(write_q),
		.addr_i(addr_q),
		.wdata_i(wdata_q),
		.wmask_i(wmask_q),
		.rdata_o(rdata_sram),
		.cfg_i(cfg_i)
	);
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			rvalid_sram_q <= 1'b0;
		else
			rvalid_sram_q <= req_q & ~write_q;
	assign req_d = req_i;
	assign write_d = write_i;
	assign addr_d = addr_i;
	assign rvalid_o = rvalid_q;
	assign rdata_o = rdata_q;
	assign rerror_o = rerror_q;
	generate
		if ((EnableParity == 0) && EnableECC) begin : gen_secded
			wire unused_wmask;
			assign unused_wmask = ^wmask_i;
			wire [TotalWidth:1] sv2v_tmp_48FEB;
			assign sv2v_tmp_48FEB = {TotalWidth {1'b1}};
			always @(*) wmask_d = sv2v_tmp_48FEB;
			if (Width == 16) begin : gen_secded_22_16
				if (HammingECC) begin : gen_hamming
					wire [TotalWidth:1] sv2v_tmp_u_enc_data_o;
					always @(*) wdata_d = sv2v_tmp_u_enc_data_o;
					prim_secded_inv_hamming_22_16_enc u_enc(
						.data_i(wdata_i),
						.data_o(sv2v_tmp_u_enc_data_o)
					);
					wire [Width * 1:1] sv2v_tmp_u_dec_data_o;
					always @(*) rdata_d[0+:Width] = sv2v_tmp_u_dec_data_o;
					wire [2:1] sv2v_tmp_u_dec_err_o;
					always @(*) rerror_d = sv2v_tmp_u_dec_err_o;
					prim_secded_inv_hamming_22_16_dec u_dec(
						.data_i(rdata_sram),
						.data_o(sv2v_tmp_u_dec_data_o),
						.err_o(sv2v_tmp_u_dec_err_o)
					);
				end
				else begin : gen_hsiao
					wire [TotalWidth:1] sv2v_tmp_u_enc_data_o;
					always @(*) wdata_d = sv2v_tmp_u_enc_data_o;
					prim_secded_inv_22_16_enc u_enc(
						.data_i(wdata_i),
						.data_o(sv2v_tmp_u_enc_data_o)
					);
					wire [Width * 1:1] sv2v_tmp_u_dec_data_o;
					always @(*) rdata_d[0+:Width] = sv2v_tmp_u_dec_data_o;
					wire [2:1] sv2v_tmp_u_dec_err_o;
					always @(*) rerror_d = sv2v_tmp_u_dec_err_o;
					prim_secded_inv_22_16_dec u_dec(
						.data_i(rdata_sram),
						.data_o(sv2v_tmp_u_dec_data_o),
						.err_o(sv2v_tmp_u_dec_err_o)
					);
				end
			end
			else if (Width == 32) begin : gen_secded_39_32
				if (HammingECC) begin : gen_hamming
					wire [TotalWidth:1] sv2v_tmp_u_enc_data_o;
					always @(*) wdata_d = sv2v_tmp_u_enc_data_o;
					prim_secded_inv_hamming_39_32_enc u_enc(
						.data_i(wdata_i),
						.data_o(sv2v_tmp_u_enc_data_o)
					);
					wire [Width * 1:1] sv2v_tmp_u_dec_data_o;
					always @(*) rdata_d[0+:Width] = sv2v_tmp_u_dec_data_o;
					wire [2:1] sv2v_tmp_u_dec_err_o;
					always @(*) rerror_d = sv2v_tmp_u_dec_err_o;
					prim_secded_inv_hamming_39_32_dec u_dec(
						.data_i(rdata_sram),
						.data_o(sv2v_tmp_u_dec_data_o),
						.err_o(sv2v_tmp_u_dec_err_o)
					);
				end
				else begin : gen_hsiao
					wire [TotalWidth:1] sv2v_tmp_u_enc_data_o;
					always @(*) wdata_d = sv2v_tmp_u_enc_data_o;
					prim_secded_inv_39_32_enc u_enc(
						.data_i(wdata_i),
						.data_o(sv2v_tmp_u_enc_data_o)
					);
					wire [Width * 1:1] sv2v_tmp_u_dec_data_o;
					always @(*) rdata_d[0+:Width] = sv2v_tmp_u_dec_data_o;
					wire [2:1] sv2v_tmp_u_dec_err_o;
					always @(*) rerror_d = sv2v_tmp_u_dec_err_o;
					prim_secded_inv_39_32_dec u_dec(
						.data_i(rdata_sram),
						.data_o(sv2v_tmp_u_dec_data_o),
						.err_o(sv2v_tmp_u_dec_err_o)
					);
				end
			end
		end
		else if (EnableParity) begin : gen_byte_parity
			always @(*) begin : p_parity
				rerror_d = 1'sb0;
				begin : sv2v_autoblock_1
					reg signed [31:0] i;
					for (i = 0; i < (Width / 8); i = i + 1)
						begin
							wmask_d[i * 9+:8] = wmask_i[i * 8+:8];
							wdata_d[i * 9+:8] = wdata_i[i * 8+:8];
							rdata_d[i * 8+:8] = rdata_sram[i * 9+:8];
							wdata_d[(i * 9) + 8] = ~(^wdata_i[i * 8+:8]);
							wmask_d[(i * 9) + 8] = &wmask_i[i * 8+:8];
							rerror_d[1] = rerror_d[1] | ~(^{rdata_sram[i * 9+:8], rdata_sram[(i * 9) + 8]});
						end
				end
			end
		end
		else begin : gen_nosecded_noparity
			wire [TotalWidth:1] sv2v_tmp_36DB7;
			assign sv2v_tmp_36DB7 = wmask_i;
			always @(*) wmask_d = sv2v_tmp_36DB7;
			wire [TotalWidth:1] sv2v_tmp_957FF;
			assign sv2v_tmp_957FF = wdata_i;
			always @(*) wdata_d = sv2v_tmp_957FF;
			wire [Width:1] sv2v_tmp_49613;
			assign sv2v_tmp_49613 = rdata_sram[0+:Width];
			always @(*) rdata_d = sv2v_tmp_49613;
			wire [2:1] sv2v_tmp_3E32B;
			assign sv2v_tmp_3E32B = 1'sb0;
			always @(*) rerror_d = sv2v_tmp_3E32B;
		end
	endgenerate
	assign rvalid_d = rvalid_sram_q;
	generate
		if (EnableInputPipeline) begin : gen_regslice_input
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni) begin
					req_q <= 1'sb0;
					write_q <= 1'sb0;
					addr_q <= 1'sb0;
					wdata_q <= 1'sb0;
					wmask_q <= 1'sb0;
				end
				else begin
					req_q <= req_d;
					write_q <= write_d;
					addr_q <= addr_d;
					wdata_q <= wdata_d;
					wmask_q <= wmask_d;
				end
		end
		else begin : gen_dirconnect_input
			wire [1:1] sv2v_tmp_48E47;
			assign sv2v_tmp_48E47 = req_d;
			always @(*) req_q = sv2v_tmp_48E47;
			wire [1:1] sv2v_tmp_988DF;
			assign sv2v_tmp_988DF = write_d;
			always @(*) write_q = sv2v_tmp_988DF;
			wire [Aw:1] sv2v_tmp_81E67;
			assign sv2v_tmp_81E67 = addr_d;
			always @(*) addr_q = sv2v_tmp_81E67;
			wire [TotalWidth:1] sv2v_tmp_D5C8F;
			assign sv2v_tmp_D5C8F = wdata_d;
			always @(*) wdata_q = sv2v_tmp_D5C8F;
			wire [TotalWidth:1] sv2v_tmp_7BD63;
			assign sv2v_tmp_7BD63 = wmask_d;
			always @(*) wmask_q = sv2v_tmp_7BD63;
		end
		if (EnableOutputPipeline) begin : gen_regslice_output
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni) begin
					rvalid_q <= 1'sb0;
					rdata_q <= 1'sb0;
					rerror_q <= 1'sb0;
				end
				else begin
					rvalid_q <= rvalid_d;
					rdata_q <= rdata_d;
					rerror_q <= rerror_d & {2 {rvalid_d}};
				end
		end
		else begin : gen_dirconnect_output
			wire [1:1] sv2v_tmp_2C5C9;
			assign sv2v_tmp_2C5C9 = rvalid_d;
			always @(*) rvalid_q = sv2v_tmp_2C5C9;
			wire [Width:1] sv2v_tmp_5A93F;
			assign sv2v_tmp_5A93F = rdata_d;
			always @(*) rdata_q = sv2v_tmp_5A93F;
			wire [2:1] sv2v_tmp_7B225;
			assign sv2v_tmp_7B225 = rerror_d & {2 {rvalid_d}};
			always @(*) rerror_q = sv2v_tmp_7B225;
		end
	endgenerate
endmodule
module prim_ram_1p_scr (
	clk_i,
	rst_ni,
	key_valid_i,
	key_i,
	nonce_i,
	req_i,
	gnt_o,
	write_i,
	addr_i,
	wdata_i,
	wmask_i,
	intg_error_i,
	rdata_o,
	rvalid_o,
	rerror_o,
	raddr_o,
	cfg_i
);
	parameter signed [31:0] Depth = 16384;
	parameter signed [31:0] Width = 32;
	parameter signed [31:0] DataBitsPerMask = 8;
	parameter [0:0] EnableParity = 1;
	parameter signed [31:0] NumPrinceRoundsHalf = 2;
	parameter signed [31:0] NumDiffRounds = 2;
	parameter signed [31:0] DiffWidth = DataBitsPerMask;
	parameter signed [31:0] NumAddrScrRounds = 2;
	parameter [0:0] ReplicateKeyStream = 1'b0;
	function automatic integer prim_util_pkg_vbits;
		input integer value;
		prim_util_pkg_vbits = (value == 1 ? 1 : $clog2(value));
	endfunction
	localparam signed [31:0] AddrWidth = prim_util_pkg_vbits(Depth);
	localparam signed [31:0] NumParScr = (ReplicateKeyStream ? 1 : (Width + 63) / 64);
	localparam signed [31:0] NumParKeystr = (ReplicateKeyStream ? (Width + 63) / 64 : 1);
	localparam signed [31:0] DataKeyWidth = 128;
	localparam signed [31:0] NonceWidth = 64 * NumParScr;
	input clk_i;
	input rst_ni;
	input key_valid_i;
	input [127:0] key_i;
	input [NonceWidth - 1:0] nonce_i;
	input req_i;
	output wire gnt_o;
	input write_i;
	input [AddrWidth - 1:0] addr_i;
	input [Width - 1:0] wdata_i;
	input [Width - 1:0] wmask_i;
	input intg_error_i;
	output reg [Width - 1:0] rdata_o;
	output reg rvalid_o;
	output wire [1:0] rerror_o;
	output wire [31:0] raddr_o;
	input wire [9:0] cfg_i;
	wire read_en;
	wire write_en_d;
	reg write_en_q;
	assign gnt_o = req_i & key_valid_i;
	assign read_en = gnt_o & ~write_i;
	assign write_en_d = gnt_o & write_i;
	reg write_pending_q;
	wire addr_collision_d;
	reg addr_collision_q;
	wire [AddrWidth - 1:0] addr_scr;
	reg [AddrWidth - 1:0] waddr_scr_q;
	assign addr_collision_d = (read_en & (write_en_q | write_pending_q)) & (addr_scr == waddr_scr_q);
	wire intg_error_buf;
	reg intg_error_w_q;
	prim_buf u_intg_error(
		.in_i(intg_error_i),
		.out_o(intg_error_buf)
	);
	wire macro_req;
	assign macro_req = (~intg_error_w_q & ~intg_error_buf) & ((read_en | write_en_q) | write_pending_q);
	wire macro_write;
	assign macro_write = ((write_en_q | write_pending_q) & ~read_en) & ~intg_error_w_q;
	wire rw_collision;
	assign rw_collision = write_en_q & read_en;
	wire [AddrWidth - 1:0] addr_mux;
	assign addr_mux = (read_en ? addr_scr : waddr_scr_q);
	generate
		if (NumAddrScrRounds > 0) begin : gen_addr_scr
			wire [AddrWidth - 1:0] addr_scr_nonce;
			assign addr_scr_nonce = nonce_i[NonceWidth - AddrWidth+:AddrWidth];
			prim_subst_perm #(
				.DataWidth(AddrWidth),
				.NumRounds(NumAddrScrRounds),
				.Decrypt(0)
			) u_prim_subst_perm(
				.data_i(addr_i),
				.key_i(addr_scr_nonce),
				.data_o(addr_scr)
			);
		end
		else begin : gen_no_addr_scr
			assign addr_scr = addr_i;
		end
	endgenerate
	reg [AddrWidth - 1:0] raddr_q;
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	assign raddr_o = sv2v_cast_32(raddr_q);
	localparam signed [31:0] DataNonceWidth = 64 - AddrWidth;
	wire [(NumParScr * 64) - 1:0] keystream;
	wire [(NumParScr * DataNonceWidth) - 1:0] data_scr_nonce;
	genvar k;
	generate
		for (k = 0; k < NumParScr; k = k + 1) begin : gen_par_scr
			assign data_scr_nonce[k * DataNonceWidth+:DataNonceWidth] = nonce_i[k * DataNonceWidth+:DataNonceWidth];
			prim_prince #(
				.DataWidth(64),
				.KeyWidth(128),
				.NumRoundsHalf(NumPrinceRoundsHalf),
				.UseOldKeySched(1'b0),
				.HalfwayDataReg(1'b1),
				.HalfwayKeyReg(1'b0)
			) u_prim_prince(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.valid_i(gnt_o),
				.data_i({data_scr_nonce[k * DataNonceWidth+:DataNonceWidth], addr_i}),
				.key_i(key_i),
				.dec_i(1'b0),
				.data_o(keystream[k * 64+:64])
			);
			if ((k == (NumParKeystr - 1)) && ((Width % 64) > 0)) begin : gen_unread_last
				localparam signed [31:0] UnusedWidth = 64 - (Width % 64);
				wire [UnusedWidth - 1:0] unused_keystream;
				assign unused_keystream = keystream[((k + 1) * 64) - 1-:UnusedWidth];
			end
		end
	endgenerate
	wire [Width - 1:0] keystream_repl;
	function automatic [Width - 1:0] sv2v_cast_92C3D;
		input reg [Width - 1:0] inp;
		sv2v_cast_92C3D = inp;
	endfunction
	assign keystream_repl = sv2v_cast_92C3D({NumParKeystr {keystream}});
	wire [Width - 1:0] rdata_scr;
	wire [Width - 1:0] rdata;
	wire [Width - 1:0] wdata_scr_d;
	reg [Width - 1:0] wdata_scr_q;
	reg [Width - 1:0] wdata_q;
	generate
		for (k = 0; k < (((Width + DiffWidth) - 1) / DiffWidth); k = k + 1) begin : gen_diffuse_data
			localparam signed [31:0] LocalWidth = ((Width - (k * DiffWidth)) >= DiffWidth ? DiffWidth : Width - (k * DiffWidth));
			wire [LocalWidth - 1:0] wdata_xor;
			assign wdata_xor = wdata_q[k * DiffWidth+:LocalWidth] ^ keystream_repl[k * DiffWidth+:LocalWidth];
			prim_subst_perm #(
				.DataWidth(LocalWidth),
				.NumRounds(NumDiffRounds),
				.Decrypt(0)
			) u_prim_subst_perm_enc(
				.data_i(wdata_xor),
				.key_i(1'sb0),
				.data_o(wdata_scr_d[k * DiffWidth+:LocalWidth])
			);
			wire [LocalWidth - 1:0] rdata_xor;
			prim_subst_perm #(
				.DataWidth(LocalWidth),
				.NumRounds(NumDiffRounds),
				.Decrypt(1)
			) u_prim_subst_perm_dec(
				.data_i(rdata_scr[k * DiffWidth+:LocalWidth]),
				.key_i(1'sb0),
				.data_o(rdata_xor)
			);
			assign rdata[k * DiffWidth+:LocalWidth] = rdata_xor ^ keystream_repl[k * DiffWidth+:LocalWidth];
		end
	endgenerate
	wire write_scr_pending_d;
	assign write_scr_pending_d = (macro_write ? 1'b0 : (rw_collision ? 1'b1 : write_pending_q));
	wire [Width - 1:0] wdata_scr;
	assign wdata_scr = (write_pending_q ? wdata_scr_q : wdata_scr_d);
	reg rvalid_q;
	reg intg_error_r_q;
	reg [Width - 1:0] wmask_q;
	always @(*) begin : p_forward_mux
		rdata_o = 1'sb0;
		rvalid_o = 1'b0;
		if (!intg_error_r_q && rvalid_q) begin
			rvalid_o = 1'b1;
			if (addr_collision_q) begin : sv2v_autoblock_1
				reg signed [31:0] k;
				for (k = 0; k < Width; k = k + 1)
					if (wmask_q[k])
						rdata_o[k] = wdata_q[k];
					else
						rdata_o[k] = rdata[k];
			end
			else
				rdata_o = rdata;
		end
	end
	always @(posedge clk_i or negedge rst_ni) begin : p_wdata_buf
		if (!rst_ni) begin
			write_pending_q <= 1'b0;
			addr_collision_q <= 1'b0;
			rvalid_q <= 1'b0;
			write_en_q <= 1'b0;
			intg_error_r_q <= 1'b0;
			intg_error_w_q <= 1'b0;
			raddr_q <= 1'sb0;
			waddr_scr_q <= 1'sb0;
			wmask_q <= 1'sb0;
			wdata_q <= 1'sb0;
			wdata_scr_q <= 1'sb0;
		end
		else begin
			write_pending_q <= write_scr_pending_d;
			addr_collision_q <= addr_collision_d;
			rvalid_q <= read_en;
			write_en_q <= write_en_d;
			intg_error_r_q <= intg_error_buf;
			if (read_en)
				raddr_q <= addr_i;
			if (write_en_d) begin
				waddr_scr_q <= addr_scr;
				wmask_q <= wmask_i;
				wdata_q <= wdata_i;
				intg_error_w_q <= intg_error_buf;
			end
			if (rw_collision)
				wdata_scr_q <= wdata_scr_d;
		end
	end
	prim_ram_1p_adv #(
		.Depth(Depth),
		.Width(Width),
		.DataBitsPerMask(DataBitsPerMask),
		.EnableECC(1'b0),
		.EnableParity(EnableParity),
		.EnableInputPipeline(1'b0),
		.EnableOutputPipeline(1'b0)
	) u_prim_ram_1p_adv(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.req_i(macro_req),
		.write_i(macro_write),
		.addr_i(addr_mux),
		.wdata_i(wdata_scr),
		.wmask_i(wmask_q),
		.rdata_o(rdata_scr),
		.rerror_o(rerror_o),
		.cfg_i(cfg_i)
	);
endmodule
module prim_reg_cdc (
	clk_src_i,
	rst_src_ni,
	clk_dst_i,
	rst_dst_ni,
	src_regwen_i,
	src_we_i,
	src_re_i,
	src_wd_i,
	src_busy_o,
	src_qs_o,
	dst_ds_i,
	dst_qs_i,
	dst_update_i,
	dst_we_o,
	dst_re_o,
	dst_regwen_o,
	dst_wd_o
);
	parameter signed [31:0] DataWidth = 32;
	parameter [DataWidth - 1:0] ResetVal = 32'h00000000;
	parameter [DataWidth - 1:0] BitMask = 32'hffffffff;
	parameter [0:0] DstWrReq = 0;
	input clk_src_i;
	input rst_src_ni;
	input clk_dst_i;
	input rst_dst_ni;
	input src_regwen_i;
	input src_we_i;
	input src_re_i;
	input [DataWidth - 1:0] src_wd_i;
	output wire src_busy_o;
	output wire [DataWidth - 1:0] src_qs_o;
	input [DataWidth - 1:0] dst_ds_i;
	input [DataWidth - 1:0] dst_qs_i;
	input dst_update_i;
	output wire dst_we_o;
	output wire dst_re_o;
	output wire dst_regwen_o;
	output wire [DataWidth - 1:0] dst_wd_o;
	localparam signed [31:0] TxnWidth = 3;
	wire src_ack;
	reg src_busy_q;
	reg [DataWidth - 1:0] src_q;
	reg [2:0] txn_bits_q;
	wire src_req;
	assign src_req = src_we_i | src_re_i;
	always @(posedge clk_src_i or negedge rst_src_ni)
		if (!rst_src_ni)
			src_busy_q <= 1'sb0;
		else if (src_req)
			src_busy_q <= 1'b1;
		else if (src_ack)
			src_busy_q <= 1'b0;
	assign src_busy_o = src_busy_q;
	wire busy;
	assign busy = src_busy_q & !src_ack;
	wire [DataWidth - 1:0] dst_qs;
	wire src_update;
	always @(posedge clk_src_i or negedge rst_src_ni)
		if (!rst_src_ni) begin
			src_q <= ResetVal;
			txn_bits_q <= 1'sb0;
		end
		else if (src_req) begin
			src_q <= src_wd_i & BitMask;
			txn_bits_q <= {src_we_i, src_re_i, src_regwen_i};
		end
		else if ((src_busy_q && src_ack) || (src_update && !busy)) begin
			src_q <= dst_qs;
			txn_bits_q <= 1'sb0;
		end
	wire unused_wd;
	assign unused_wd = ^src_wd_i;
	assign src_qs_o = src_q;
	assign dst_wd_o = src_q;
	wire dst_req_from_src;
	wire dst_req;
	prim_pulse_sync u_src_to_dst_req(
		.clk_src_i(clk_src_i),
		.rst_src_ni(rst_src_ni),
		.clk_dst_i(clk_dst_i),
		.rst_dst_ni(rst_dst_ni),
		.src_pulse_i(src_req),
		.dst_pulse_o(dst_req_from_src)
	);
	prim_reg_cdc_arb #(
		.DataWidth(DataWidth),
		.ResetVal(ResetVal),
		.DstWrReq(DstWrReq)
	) u_arb(
		.clk_src_i(clk_src_i),
		.rst_src_ni(rst_src_ni),
		.clk_dst_i(clk_dst_i),
		.rst_dst_ni(rst_dst_ni),
		.src_ack_o(src_ack),
		.src_update_o(src_update),
		.dst_req_i(dst_req_from_src),
		.dst_req_o(dst_req),
		.dst_update_i(dst_update_i),
		.dst_ds_i(dst_ds_i),
		.dst_qs_i(dst_qs_i),
		.dst_qs_o(dst_qs)
	);
	assign {dst_we_o, dst_re_o, dst_regwen_o} = txn_bits_q & {TxnWidth {dst_req}};
endmodule
module prim_reg_cdc_arb (
	clk_src_i,
	rst_src_ni,
	clk_dst_i,
	rst_dst_ni,
	src_ack_o,
	src_update_o,
	dst_req_i,
	dst_req_o,
	dst_update_i,
	dst_ds_i,
	dst_qs_i,
	dst_qs_o
);
	parameter signed [31:0] DataWidth = 32;
	parameter [DataWidth - 1:0] ResetVal = 32'h00000000;
	parameter [0:0] DstWrReq = 0;
	input clk_src_i;
	input rst_src_ni;
	input clk_dst_i;
	input rst_dst_ni;
	output wire src_ack_o;
	output wire src_update_o;
	input dst_req_i;
	output wire dst_req_o;
	input dst_update_i;
	input [DataWidth - 1:0] dst_ds_i;
	input [DataWidth - 1:0] dst_qs_i;
	output reg [DataWidth - 1:0] dst_qs_o;
	wire dst_update;
	assign dst_update = dst_update_i & (dst_qs_o != dst_ds_i);
	generate
		if (DstWrReq) begin : gen_wr_req
			reg dst_lat_q;
			reg dst_lat_d;
			wire dst_update_req;
			wire dst_update_ack;
			reg id_q;
			reg [1:0] state_q;
			reg [1:0] state_d;
			always @(posedge clk_dst_i or negedge rst_dst_ni)
				if (!rst_dst_ni)
					state_q <= 2'd0;
				else
					state_q <= state_d;
			reg busy;
			reg dst_req_q;
			wire dst_req;
			always @(posedge clk_dst_i or negedge rst_dst_ni)
				if (!rst_dst_ni)
					dst_req_q <= 1'sb0;
				else if (dst_req_q && dst_lat_d)
					dst_req_q <= 1'sb0;
				else if ((dst_req_i && !dst_req_q) && busy)
					dst_req_q <= 1'b1;
			assign dst_req = dst_req_q | dst_req_i;
			always @(posedge clk_dst_i or negedge rst_dst_ni)
				if (!rst_dst_ni)
					dst_qs_o <= ResetVal;
				else if (dst_lat_d)
					dst_qs_o <= dst_ds_i;
				else if (dst_lat_q)
					dst_qs_o <= dst_qs_i;
			always @(posedge clk_dst_i or negedge rst_dst_ni)
				if (!rst_dst_ni)
					id_q <= 1'd0;
				else if (dst_update_req && dst_update_ack)
					id_q <= 1'd0;
				else if (dst_req && dst_lat_d)
					id_q <= 1'd0;
				else if (!dst_req && dst_lat_d)
					id_q <= 1'd1;
				else if (dst_lat_q)
					id_q <= 1'd1;
			assign dst_req_o = ~busy & dst_req;
			reg dst_hold_req;
			always @(*) begin
				state_d = state_q;
				dst_hold_req = 1'sb0;
				dst_lat_q = 1'sb0;
				dst_lat_d = 1'sb0;
				busy = 1'b1;
				case (state_q)
					2'd0: begin
						busy = 1'sb0;
						if (dst_req) begin
							state_d = 2'd1;
							dst_lat_d = 1'b1;
						end
						else if (dst_update) begin
							state_d = 2'd1;
							dst_lat_d = 1'b1;
						end
						else if (dst_qs_o != dst_qs_i) begin
							state_d = 2'd1;
							dst_lat_q = 1'b1;
						end
					end
					2'd1: begin
						dst_hold_req = 1'b1;
						if (dst_update_ack)
							state_d = 2'd0;
					end
					default: state_d = 2'd0;
				endcase
			end
			assign dst_update_req = (dst_hold_req | dst_lat_d) | dst_lat_q;
			wire src_req;
			prim_sync_reqack u_dst_update_sync(
				.clk_src_i(clk_dst_i),
				.rst_src_ni(rst_dst_ni),
				.clk_dst_i(clk_src_i),
				.rst_dst_ni(rst_src_ni),
				.req_chk_i(1'b1),
				.src_req_i(dst_update_req),
				.src_ack_o(dst_update_ack),
				.dst_req_o(src_req),
				.dst_ack_i(src_req)
			);
			assign src_ack_o = src_req & (id_q == 1'd0);
			assign src_update_o = src_req & (id_q == 1'd1);
		end
		else begin : gen_passthru
			wire [DataWidth:1] sv2v_tmp_0FEB6;
			assign sv2v_tmp_0FEB6 = dst_qs_i;
			always @(*) dst_qs_o = sv2v_tmp_0FEB6;
			assign dst_req_o = dst_req_i;
			assign src_update_o = 1'sb0;
			prim_pulse_sync u_dst_to_src_ack(
				.clk_src_i(clk_dst_i),
				.rst_src_ni(rst_dst_ni),
				.clk_dst_i(clk_src_i),
				.rst_dst_ni(rst_src_ni),
				.src_pulse_i(dst_req_i),
				.dst_pulse_o(src_ack_o)
			);
			wire unused_sigs;
			assign unused_sigs = |{dst_ds_i, dst_update};
		end
	endgenerate
endmodule
module prim_reg_we_check (
	clk_i,
	rst_ni,
	oh_i,
	en_i,
	err_o
);
	parameter [31:0] OneHotWidth = 32;
	input clk_i;
	input rst_ni;
	input wire [OneHotWidth - 1:0] oh_i;
	input wire en_i;
	output wire err_o;
	wire [OneHotWidth - 1:0] oh_buf;
	prim_buf #(.Width(OneHotWidth)) u_prim_buf(
		.in_i(oh_i),
		.out_o(oh_buf)
	);
	function automatic integer prim_util_pkg_vbits;
		input integer value;
		prim_util_pkg_vbits = (value == 1 ? 1 : $clog2(value));
	endfunction
	prim_onehot_check #(
		.OneHotWidth(OneHotWidth),
		.AddrWidth(prim_util_pkg_vbits(OneHotWidth)),
		.EnableCheck(1),
		.AddrCheck(0),
		.StrictCheck(0)
	) u_prim_onehot_check(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.oh_i(oh_buf),
		.addr_i(1'sb0),
		.en_i(en_i),
		.err_o(err_o)
	);
endmodule
module prim_rst_sync (
	clk_i,
	d_i,
	q_o,
	scan_rst_ni,
	scanmode_i
);
	parameter [0:0] ActiveHigh = 1'b0;
	parameter [0:0] SkipScan = 1'b0;
	input clk_i;
	input d_i;
	output wire q_o;
	input scan_rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	input wire [3:0] scanmode_i;
	wire async_rst_n;
	wire scan_rst;
	wire rst_sync;
	generate
		if (ActiveHigh == 1'b1) begin : g_rst_inv
			assign async_rst_n = ~d_i;
			assign scan_rst = ~scan_rst_ni;
		end
		else begin : g_rst_direct
			assign async_rst_n = d_i;
			assign scan_rst = scan_rst_ni;
		end
	endgenerate
	prim_flop_2sync #(
		.Width(1),
		.ResetValue(ActiveHigh)
	) u_sync(
		.clk_i(clk_i),
		.rst_ni(async_rst_n),
		.d_i(!ActiveHigh),
		.q_o(rst_sync)
	);
	function automatic [3:0] sv2v_cast_E830B;
		input reg [3:0] inp;
		sv2v_cast_E830B = inp;
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_true_strict;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_true_strict = sv2v_cast_E830B(4'h6) == val;
	endfunction
	generate
		if (SkipScan) begin : g_skip_scan
			wire unused_scan;
			assign unused_scan = ^{scan_rst, scanmode_i};
			assign q_o = rst_sync;
		end
		else begin : g_scan_mux
			prim_clock_mux2 #(.NoFpgaBufG(1'b1)) u_scan_mux(
				.clk0_i(rst_sync),
				.clk1_i(scan_rst),
				.sel_i(prim_mubi_pkg_mubi4_test_true_strict(scanmode_i)),
				.clk_o(q_o)
			);
		end
	endgenerate
endmodule
module prim_sec_anchor_buf (
	in_i,
	out_o
);
	parameter signed [31:0] Width = 1;
	input [Width - 1:0] in_i;
	output wire [Width - 1:0] out_o;
	prim_buf #(.Width(Width)) u_secure_anchor_buf(
		.in_i(in_i),
		.out_o(out_o)
	);
endmodule
module prim_sec_anchor_flop (
	clk_i,
	rst_ni,
	d_i,
	q_o
);
	parameter signed [31:0] Width = 1;
	parameter [Width - 1:0] ResetValue = 0;
	input clk_i;
	input rst_ni;
	input [Width - 1:0] d_i;
	output wire [Width - 1:0] q_o;
	prim_flop #(
		.Width(Width),
		.ResetValue(ResetValue)
	) u_secure_anchor_flop(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(d_i),
		.q_o(q_o)
	);
endmodule
module prim_secded_22_16_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [21:0] data_i;
	output reg [15:0] data_o;
	output reg [5:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^(data_i & 22'h01496e);
		syndrome_o[1] = ^(data_i & 22'h02f20b);
		syndrome_o[2] = ^(data_i & 22'h048ed8);
		syndrome_o[3] = ^(data_i & 22'h087714);
		syndrome_o[4] = ^(data_i & 22'h10aca5);
		syndrome_o[5] = ^(data_i & 22'h2011f3);
		data_o[0] = (syndrome_o == 6'h32) ^ data_i[0];
		data_o[1] = (syndrome_o == 6'h23) ^ data_i[1];
		data_o[2] = (syndrome_o == 6'h19) ^ data_i[2];
		data_o[3] = (syndrome_o == 6'h07) ^ data_i[3];
		data_o[4] = (syndrome_o == 6'h2c) ^ data_i[4];
		data_o[5] = (syndrome_o == 6'h31) ^ data_i[5];
		data_o[6] = (syndrome_o == 6'h25) ^ data_i[6];
		data_o[7] = (syndrome_o == 6'h34) ^ data_i[7];
		data_o[8] = (syndrome_o == 6'h29) ^ data_i[8];
		data_o[9] = (syndrome_o == 6'h0e) ^ data_i[9];
		data_o[10] = (syndrome_o == 6'h1c) ^ data_i[10];
		data_o[11] = (syndrome_o == 6'h15) ^ data_i[11];
		data_o[12] = (syndrome_o == 6'h2a) ^ data_i[12];
		data_o[13] = (syndrome_o == 6'h1a) ^ data_i[13];
		data_o[14] = (syndrome_o == 6'h0b) ^ data_i[14];
		data_o[15] = (syndrome_o == 6'h16) ^ data_i[15];
		err_o[0] = ^syndrome_o;
		err_o[1] = ~err_o[0] & |syndrome_o;
	end
endmodule
module prim_secded_22_16_enc (
	data_i,
	data_o
);
	input [15:0] data_i;
	output reg [21:0] data_o;
	function automatic [21:0] sv2v_cast_22;
		input reg [21:0] inp;
		sv2v_cast_22 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_22(data_i);
		data_o[16] = ^(data_o & 22'h00496e);
		data_o[17] = ^(data_o & 22'h00f20b);
		data_o[18] = ^(data_o & 22'h008ed8);
		data_o[19] = ^(data_o & 22'h007714);
		data_o[20] = ^(data_o & 22'h00aca5);
		data_o[21] = ^(data_o & 22'h0011f3);
	end
endmodule
module prim_secded_28_22_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [27:0] data_i;
	output reg [21:0] data_o;
	output reg [5:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^(data_i & 28'h07003ff);
		syndrome_o[1] = ^(data_i & 28'h090fc0f);
		syndrome_o[2] = ^(data_i & 28'h1271c71);
		syndrome_o[3] = ^(data_i & 28'h23b6592);
		syndrome_o[4] = ^(data_i & 28'h43daaa4);
		syndrome_o[5] = ^(data_i & 28'h83ed348);
		data_o[0] = (syndrome_o == 6'h07) ^ data_i[0];
		data_o[1] = (syndrome_o == 6'h0b) ^ data_i[1];
		data_o[2] = (syndrome_o == 6'h13) ^ data_i[2];
		data_o[3] = (syndrome_o == 6'h23) ^ data_i[3];
		data_o[4] = (syndrome_o == 6'h0d) ^ data_i[4];
		data_o[5] = (syndrome_o == 6'h15) ^ data_i[5];
		data_o[6] = (syndrome_o == 6'h25) ^ data_i[6];
		data_o[7] = (syndrome_o == 6'h19) ^ data_i[7];
		data_o[8] = (syndrome_o == 6'h29) ^ data_i[8];
		data_o[9] = (syndrome_o == 6'h31) ^ data_i[9];
		data_o[10] = (syndrome_o == 6'h0e) ^ data_i[10];
		data_o[11] = (syndrome_o == 6'h16) ^ data_i[11];
		data_o[12] = (syndrome_o == 6'h26) ^ data_i[12];
		data_o[13] = (syndrome_o == 6'h1a) ^ data_i[13];
		data_o[14] = (syndrome_o == 6'h2a) ^ data_i[14];
		data_o[15] = (syndrome_o == 6'h32) ^ data_i[15];
		data_o[16] = (syndrome_o == 6'h1c) ^ data_i[16];
		data_o[17] = (syndrome_o == 6'h2c) ^ data_i[17];
		data_o[18] = (syndrome_o == 6'h34) ^ data_i[18];
		data_o[19] = (syndrome_o == 6'h38) ^ data_i[19];
		data_o[20] = (syndrome_o == 6'h3b) ^ data_i[20];
		data_o[21] = (syndrome_o == 6'h3d) ^ data_i[21];
		err_o[0] = ^syndrome_o;
		err_o[1] = ~err_o[0] & |syndrome_o;
	end
endmodule
module prim_secded_28_22_enc (
	data_i,
	data_o
);
	input [21:0] data_i;
	output reg [27:0] data_o;
	function automatic [27:0] sv2v_cast_28;
		input reg [27:0] inp;
		sv2v_cast_28 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_28(data_i);
		data_o[22] = ^(data_o & 28'h03003ff);
		data_o[23] = ^(data_o & 28'h010fc0f);
		data_o[24] = ^(data_o & 28'h0271c71);
		data_o[25] = ^(data_o & 28'h03b6592);
		data_o[26] = ^(data_o & 28'h03daaa4);
		data_o[27] = ^(data_o & 28'h03ed348);
	end
endmodule
module prim_secded_39_32_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [38:0] data_i;
	output reg [31:0] data_o;
	output reg [6:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^(data_i & 39'h012606bd25);
		syndrome_o[1] = ^(data_i & 39'h02deba8050);
		syndrome_o[2] = ^(data_i & 39'h04413d89aa);
		syndrome_o[3] = ^(data_i & 39'h0831234ed1);
		syndrome_o[4] = ^(data_i & 39'h10c2c1323b);
		syndrome_o[5] = ^(data_i & 39'h202dcc624c);
		syndrome_o[6] = ^(data_i & 39'h4098505586);
		data_o[0] = (syndrome_o == 7'h19) ^ data_i[0];
		data_o[1] = (syndrome_o == 7'h54) ^ data_i[1];
		data_o[2] = (syndrome_o == 7'h61) ^ data_i[2];
		data_o[3] = (syndrome_o == 7'h34) ^ data_i[3];
		data_o[4] = (syndrome_o == 7'h1a) ^ data_i[4];
		data_o[5] = (syndrome_o == 7'h15) ^ data_i[5];
		data_o[6] = (syndrome_o == 7'h2a) ^ data_i[6];
		data_o[7] = (syndrome_o == 7'h4c) ^ data_i[7];
		data_o[8] = (syndrome_o == 7'h45) ^ data_i[8];
		data_o[9] = (syndrome_o == 7'h38) ^ data_i[9];
		data_o[10] = (syndrome_o == 7'h49) ^ data_i[10];
		data_o[11] = (syndrome_o == 7'h0d) ^ data_i[11];
		data_o[12] = (syndrome_o == 7'h51) ^ data_i[12];
		data_o[13] = (syndrome_o == 7'h31) ^ data_i[13];
		data_o[14] = (syndrome_o == 7'h68) ^ data_i[14];
		data_o[15] = (syndrome_o == 7'h07) ^ data_i[15];
		data_o[16] = (syndrome_o == 7'h1c) ^ data_i[16];
		data_o[17] = (syndrome_o == 7'h0b) ^ data_i[17];
		data_o[18] = (syndrome_o == 7'h25) ^ data_i[18];
		data_o[19] = (syndrome_o == 7'h26) ^ data_i[19];
		data_o[20] = (syndrome_o == 7'h46) ^ data_i[20];
		data_o[21] = (syndrome_o == 7'h0e) ^ data_i[21];
		data_o[22] = (syndrome_o == 7'h70) ^ data_i[22];
		data_o[23] = (syndrome_o == 7'h32) ^ data_i[23];
		data_o[24] = (syndrome_o == 7'h2c) ^ data_i[24];
		data_o[25] = (syndrome_o == 7'h13) ^ data_i[25];
		data_o[26] = (syndrome_o == 7'h23) ^ data_i[26];
		data_o[27] = (syndrome_o == 7'h62) ^ data_i[27];
		data_o[28] = (syndrome_o == 7'h4a) ^ data_i[28];
		data_o[29] = (syndrome_o == 7'h29) ^ data_i[29];
		data_o[30] = (syndrome_o == 7'h16) ^ data_i[30];
		data_o[31] = (syndrome_o == 7'h52) ^ data_i[31];
		err_o[0] = ^syndrome_o;
		err_o[1] = ~err_o[0] & |syndrome_o;
	end
endmodule
module prim_secded_39_32_enc (
	data_i,
	data_o
);
	input [31:0] data_i;
	output reg [38:0] data_o;
	function automatic [38:0] sv2v_cast_39;
		input reg [38:0] inp;
		sv2v_cast_39 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_39(data_i);
		data_o[32] = ^(data_o & 39'h002606bd25);
		data_o[33] = ^(data_o & 39'h00deba8050);
		data_o[34] = ^(data_o & 39'h00413d89aa);
		data_o[35] = ^(data_o & 39'h0031234ed1);
		data_o[36] = ^(data_o & 39'h00c2c1323b);
		data_o[37] = ^(data_o & 39'h002dcc624c);
		data_o[38] = ^(data_o & 39'h0098505586);
	end
endmodule
module prim_secded_64_57_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [63:0] data_i;
	output reg [56:0] data_o;
	output reg [6:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^(data_i & 64'h0303fff800007fff);
		syndrome_o[1] = ^(data_i & 64'h057c1ff801ff801f);
		syndrome_o[2] = ^(data_i & 64'h09bde1f87e0781e1);
		syndrome_o[3] = ^(data_i & 64'h11deee3b8e388e22);
		syndrome_o[4] = ^(data_i & 64'h21ef76cdb2c93244);
		syndrome_o[5] = ^(data_i & 64'h41f7bb56d5525488);
		syndrome_o[6] = ^(data_i & 64'h81fbdda769a46910);
		data_o[0] = (syndrome_o == 7'h07) ^ data_i[0];
		data_o[1] = (syndrome_o == 7'h0b) ^ data_i[1];
		data_o[2] = (syndrome_o == 7'h13) ^ data_i[2];
		data_o[3] = (syndrome_o == 7'h23) ^ data_i[3];
		data_o[4] = (syndrome_o == 7'h43) ^ data_i[4];
		data_o[5] = (syndrome_o == 7'h0d) ^ data_i[5];
		data_o[6] = (syndrome_o == 7'h15) ^ data_i[6];
		data_o[7] = (syndrome_o == 7'h25) ^ data_i[7];
		data_o[8] = (syndrome_o == 7'h45) ^ data_i[8];
		data_o[9] = (syndrome_o == 7'h19) ^ data_i[9];
		data_o[10] = (syndrome_o == 7'h29) ^ data_i[10];
		data_o[11] = (syndrome_o == 7'h49) ^ data_i[11];
		data_o[12] = (syndrome_o == 7'h31) ^ data_i[12];
		data_o[13] = (syndrome_o == 7'h51) ^ data_i[13];
		data_o[14] = (syndrome_o == 7'h61) ^ data_i[14];
		data_o[15] = (syndrome_o == 7'h0e) ^ data_i[15];
		data_o[16] = (syndrome_o == 7'h16) ^ data_i[16];
		data_o[17] = (syndrome_o == 7'h26) ^ data_i[17];
		data_o[18] = (syndrome_o == 7'h46) ^ data_i[18];
		data_o[19] = (syndrome_o == 7'h1a) ^ data_i[19];
		data_o[20] = (syndrome_o == 7'h2a) ^ data_i[20];
		data_o[21] = (syndrome_o == 7'h4a) ^ data_i[21];
		data_o[22] = (syndrome_o == 7'h32) ^ data_i[22];
		data_o[23] = (syndrome_o == 7'h52) ^ data_i[23];
		data_o[24] = (syndrome_o == 7'h62) ^ data_i[24];
		data_o[25] = (syndrome_o == 7'h1c) ^ data_i[25];
		data_o[26] = (syndrome_o == 7'h2c) ^ data_i[26];
		data_o[27] = (syndrome_o == 7'h4c) ^ data_i[27];
		data_o[28] = (syndrome_o == 7'h34) ^ data_i[28];
		data_o[29] = (syndrome_o == 7'h54) ^ data_i[29];
		data_o[30] = (syndrome_o == 7'h64) ^ data_i[30];
		data_o[31] = (syndrome_o == 7'h38) ^ data_i[31];
		data_o[32] = (syndrome_o == 7'h58) ^ data_i[32];
		data_o[33] = (syndrome_o == 7'h68) ^ data_i[33];
		data_o[34] = (syndrome_o == 7'h70) ^ data_i[34];
		data_o[35] = (syndrome_o == 7'h1f) ^ data_i[35];
		data_o[36] = (syndrome_o == 7'h2f) ^ data_i[36];
		data_o[37] = (syndrome_o == 7'h4f) ^ data_i[37];
		data_o[38] = (syndrome_o == 7'h37) ^ data_i[38];
		data_o[39] = (syndrome_o == 7'h57) ^ data_i[39];
		data_o[40] = (syndrome_o == 7'h67) ^ data_i[40];
		data_o[41] = (syndrome_o == 7'h3b) ^ data_i[41];
		data_o[42] = (syndrome_o == 7'h5b) ^ data_i[42];
		data_o[43] = (syndrome_o == 7'h6b) ^ data_i[43];
		data_o[44] = (syndrome_o == 7'h73) ^ data_i[44];
		data_o[45] = (syndrome_o == 7'h3d) ^ data_i[45];
		data_o[46] = (syndrome_o == 7'h5d) ^ data_i[46];
		data_o[47] = (syndrome_o == 7'h6d) ^ data_i[47];
		data_o[48] = (syndrome_o == 7'h75) ^ data_i[48];
		data_o[49] = (syndrome_o == 7'h79) ^ data_i[49];
		data_o[50] = (syndrome_o == 7'h3e) ^ data_i[50];
		data_o[51] = (syndrome_o == 7'h5e) ^ data_i[51];
		data_o[52] = (syndrome_o == 7'h6e) ^ data_i[52];
		data_o[53] = (syndrome_o == 7'h76) ^ data_i[53];
		data_o[54] = (syndrome_o == 7'h7a) ^ data_i[54];
		data_o[55] = (syndrome_o == 7'h7c) ^ data_i[55];
		data_o[56] = (syndrome_o == 7'h7f) ^ data_i[56];
		err_o[0] = ^syndrome_o;
		err_o[1] = ~err_o[0] & |syndrome_o;
	end
endmodule
module prim_secded_64_57_enc (
	data_i,
	data_o
);
	input [56:0] data_i;
	output reg [63:0] data_o;
	function automatic [63:0] sv2v_cast_64;
		input reg [63:0] inp;
		sv2v_cast_64 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_64(data_i);
		data_o[57] = ^(data_o & 64'h0103fff800007fff);
		data_o[58] = ^(data_o & 64'h017c1ff801ff801f);
		data_o[59] = ^(data_o & 64'h01bde1f87e0781e1);
		data_o[60] = ^(data_o & 64'h01deee3b8e388e22);
		data_o[61] = ^(data_o & 64'h01ef76cdb2c93244);
		data_o[62] = ^(data_o & 64'h01f7bb56d5525488);
		data_o[63] = ^(data_o & 64'h01fbdda769a46910);
	end
endmodule
module prim_secded_72_64_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [71:0] data_i;
	output reg [63:0] data_o;
	output reg [7:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^(data_i & 72'h01b9000000001fffff);
		syndrome_o[1] = ^(data_i & 72'h025e00000fffe0003f);
		syndrome_o[2] = ^(data_i & 72'h0467003ff003e007c1);
		syndrome_o[3] = ^(data_i & 72'h08cd0fc0f03c207842);
		syndrome_o[4] = ^(data_i & 72'h10b671c711c4438884);
		syndrome_o[5] = ^(data_i & 72'h20b5b65926488c9108);
		syndrome_o[6] = ^(data_i & 72'h40cbdaaa4a91152210);
		syndrome_o[7] = ^(data_i & 72'h807aed348d221a4420);
		data_o[0] = (syndrome_o == 8'h07) ^ data_i[0];
		data_o[1] = (syndrome_o == 8'h0b) ^ data_i[1];
		data_o[2] = (syndrome_o == 8'h13) ^ data_i[2];
		data_o[3] = (syndrome_o == 8'h23) ^ data_i[3];
		data_o[4] = (syndrome_o == 8'h43) ^ data_i[4];
		data_o[5] = (syndrome_o == 8'h83) ^ data_i[5];
		data_o[6] = (syndrome_o == 8'h0d) ^ data_i[6];
		data_o[7] = (syndrome_o == 8'h15) ^ data_i[7];
		data_o[8] = (syndrome_o == 8'h25) ^ data_i[8];
		data_o[9] = (syndrome_o == 8'h45) ^ data_i[9];
		data_o[10] = (syndrome_o == 8'h85) ^ data_i[10];
		data_o[11] = (syndrome_o == 8'h19) ^ data_i[11];
		data_o[12] = (syndrome_o == 8'h29) ^ data_i[12];
		data_o[13] = (syndrome_o == 8'h49) ^ data_i[13];
		data_o[14] = (syndrome_o == 8'h89) ^ data_i[14];
		data_o[15] = (syndrome_o == 8'h31) ^ data_i[15];
		data_o[16] = (syndrome_o == 8'h51) ^ data_i[16];
		data_o[17] = (syndrome_o == 8'h91) ^ data_i[17];
		data_o[18] = (syndrome_o == 8'h61) ^ data_i[18];
		data_o[19] = (syndrome_o == 8'ha1) ^ data_i[19];
		data_o[20] = (syndrome_o == 8'hc1) ^ data_i[20];
		data_o[21] = (syndrome_o == 8'h0e) ^ data_i[21];
		data_o[22] = (syndrome_o == 8'h16) ^ data_i[22];
		data_o[23] = (syndrome_o == 8'h26) ^ data_i[23];
		data_o[24] = (syndrome_o == 8'h46) ^ data_i[24];
		data_o[25] = (syndrome_o == 8'h86) ^ data_i[25];
		data_o[26] = (syndrome_o == 8'h1a) ^ data_i[26];
		data_o[27] = (syndrome_o == 8'h2a) ^ data_i[27];
		data_o[28] = (syndrome_o == 8'h4a) ^ data_i[28];
		data_o[29] = (syndrome_o == 8'h8a) ^ data_i[29];
		data_o[30] = (syndrome_o == 8'h32) ^ data_i[30];
		data_o[31] = (syndrome_o == 8'h52) ^ data_i[31];
		data_o[32] = (syndrome_o == 8'h92) ^ data_i[32];
		data_o[33] = (syndrome_o == 8'h62) ^ data_i[33];
		data_o[34] = (syndrome_o == 8'ha2) ^ data_i[34];
		data_o[35] = (syndrome_o == 8'hc2) ^ data_i[35];
		data_o[36] = (syndrome_o == 8'h1c) ^ data_i[36];
		data_o[37] = (syndrome_o == 8'h2c) ^ data_i[37];
		data_o[38] = (syndrome_o == 8'h4c) ^ data_i[38];
		data_o[39] = (syndrome_o == 8'h8c) ^ data_i[39];
		data_o[40] = (syndrome_o == 8'h34) ^ data_i[40];
		data_o[41] = (syndrome_o == 8'h54) ^ data_i[41];
		data_o[42] = (syndrome_o == 8'h94) ^ data_i[42];
		data_o[43] = (syndrome_o == 8'h64) ^ data_i[43];
		data_o[44] = (syndrome_o == 8'ha4) ^ data_i[44];
		data_o[45] = (syndrome_o == 8'hc4) ^ data_i[45];
		data_o[46] = (syndrome_o == 8'h38) ^ data_i[46];
		data_o[47] = (syndrome_o == 8'h58) ^ data_i[47];
		data_o[48] = (syndrome_o == 8'h98) ^ data_i[48];
		data_o[49] = (syndrome_o == 8'h68) ^ data_i[49];
		data_o[50] = (syndrome_o == 8'ha8) ^ data_i[50];
		data_o[51] = (syndrome_o == 8'hc8) ^ data_i[51];
		data_o[52] = (syndrome_o == 8'h70) ^ data_i[52];
		data_o[53] = (syndrome_o == 8'hb0) ^ data_i[53];
		data_o[54] = (syndrome_o == 8'hd0) ^ data_i[54];
		data_o[55] = (syndrome_o == 8'he0) ^ data_i[55];
		data_o[56] = (syndrome_o == 8'h6d) ^ data_i[56];
		data_o[57] = (syndrome_o == 8'hd6) ^ data_i[57];
		data_o[58] = (syndrome_o == 8'h3e) ^ data_i[58];
		data_o[59] = (syndrome_o == 8'hcb) ^ data_i[59];
		data_o[60] = (syndrome_o == 8'hb3) ^ data_i[60];
		data_o[61] = (syndrome_o == 8'hb5) ^ data_i[61];
		data_o[62] = (syndrome_o == 8'hce) ^ data_i[62];
		data_o[63] = (syndrome_o == 8'h79) ^ data_i[63];
		err_o[0] = ^syndrome_o;
		err_o[1] = ~err_o[0] & |syndrome_o;
	end
endmodule
module prim_secded_72_64_enc (
	data_i,
	data_o
);
	input [63:0] data_i;
	output reg [71:0] data_o;
	function automatic [71:0] sv2v_cast_72;
		input reg [71:0] inp;
		sv2v_cast_72 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_72(data_i);
		data_o[64] = ^(data_o & 72'h00b9000000001fffff);
		data_o[65] = ^(data_o & 72'h005e00000fffe0003f);
		data_o[66] = ^(data_o & 72'h0067003ff003e007c1);
		data_o[67] = ^(data_o & 72'h00cd0fc0f03c207842);
		data_o[68] = ^(data_o & 72'h00b671c711c4438884);
		data_o[69] = ^(data_o & 72'h00b5b65926488c9108);
		data_o[70] = ^(data_o & 72'h00cbdaaa4a91152210);
		data_o[71] = ^(data_o & 72'h007aed348d221a4420);
	end
endmodule
module prim_secded_hamming_22_16_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [21:0] data_i;
	output reg [15:0] data_o;
	output reg [5:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^(data_i & 22'h01ad5b);
		syndrome_o[1] = ^(data_i & 22'h02366d);
		syndrome_o[2] = ^(data_i & 22'h04c78e);
		syndrome_o[3] = ^(data_i & 22'h0807f0);
		syndrome_o[4] = ^(data_i & 22'h10f800);
		syndrome_o[5] = ^(data_i & 22'h3fffff);
		data_o[0] = (syndrome_o == 6'h23) ^ data_i[0];
		data_o[1] = (syndrome_o == 6'h25) ^ data_i[1];
		data_o[2] = (syndrome_o == 6'h26) ^ data_i[2];
		data_o[3] = (syndrome_o == 6'h27) ^ data_i[3];
		data_o[4] = (syndrome_o == 6'h29) ^ data_i[4];
		data_o[5] = (syndrome_o == 6'h2a) ^ data_i[5];
		data_o[6] = (syndrome_o == 6'h2b) ^ data_i[6];
		data_o[7] = (syndrome_o == 6'h2c) ^ data_i[7];
		data_o[8] = (syndrome_o == 6'h2d) ^ data_i[8];
		data_o[9] = (syndrome_o == 6'h2e) ^ data_i[9];
		data_o[10] = (syndrome_o == 6'h2f) ^ data_i[10];
		data_o[11] = (syndrome_o == 6'h31) ^ data_i[11];
		data_o[12] = (syndrome_o == 6'h32) ^ data_i[12];
		data_o[13] = (syndrome_o == 6'h33) ^ data_i[13];
		data_o[14] = (syndrome_o == 6'h34) ^ data_i[14];
		data_o[15] = (syndrome_o == 6'h35) ^ data_i[15];
		err_o[0] = syndrome_o[5];
		err_o[1] = |syndrome_o[4:0] & ~syndrome_o[5];
	end
endmodule
module prim_secded_hamming_22_16_enc (
	data_i,
	data_o
);
	input [15:0] data_i;
	output reg [21:0] data_o;
	function automatic [21:0] sv2v_cast_22;
		input reg [21:0] inp;
		sv2v_cast_22 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_22(data_i);
		data_o[16] = ^(data_o & 22'h00ad5b);
		data_o[17] = ^(data_o & 22'h00366d);
		data_o[18] = ^(data_o & 22'h00c78e);
		data_o[19] = ^(data_o & 22'h0007f0);
		data_o[20] = ^(data_o & 22'h00f800);
		data_o[21] = ^(data_o & 22'h1fffff);
	end
endmodule
module prim_secded_hamming_39_32_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [38:0] data_i;
	output reg [31:0] data_o;
	output reg [6:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^(data_i & 39'h0156aaad5b);
		syndrome_o[1] = ^(data_i & 39'h029b33366d);
		syndrome_o[2] = ^(data_i & 39'h04e3c3c78e);
		syndrome_o[3] = ^(data_i & 39'h0803fc07f0);
		syndrome_o[4] = ^(data_i & 39'h1003fff800);
		syndrome_o[5] = ^(data_i & 39'h20fc000000);
		syndrome_o[6] = ^(data_i & 39'h7fffffffff);
		data_o[0] = (syndrome_o == 7'h43) ^ data_i[0];
		data_o[1] = (syndrome_o == 7'h45) ^ data_i[1];
		data_o[2] = (syndrome_o == 7'h46) ^ data_i[2];
		data_o[3] = (syndrome_o == 7'h47) ^ data_i[3];
		data_o[4] = (syndrome_o == 7'h49) ^ data_i[4];
		data_o[5] = (syndrome_o == 7'h4a) ^ data_i[5];
		data_o[6] = (syndrome_o == 7'h4b) ^ data_i[6];
		data_o[7] = (syndrome_o == 7'h4c) ^ data_i[7];
		data_o[8] = (syndrome_o == 7'h4d) ^ data_i[8];
		data_o[9] = (syndrome_o == 7'h4e) ^ data_i[9];
		data_o[10] = (syndrome_o == 7'h4f) ^ data_i[10];
		data_o[11] = (syndrome_o == 7'h51) ^ data_i[11];
		data_o[12] = (syndrome_o == 7'h52) ^ data_i[12];
		data_o[13] = (syndrome_o == 7'h53) ^ data_i[13];
		data_o[14] = (syndrome_o == 7'h54) ^ data_i[14];
		data_o[15] = (syndrome_o == 7'h55) ^ data_i[15];
		data_o[16] = (syndrome_o == 7'h56) ^ data_i[16];
		data_o[17] = (syndrome_o == 7'h57) ^ data_i[17];
		data_o[18] = (syndrome_o == 7'h58) ^ data_i[18];
		data_o[19] = (syndrome_o == 7'h59) ^ data_i[19];
		data_o[20] = (syndrome_o == 7'h5a) ^ data_i[20];
		data_o[21] = (syndrome_o == 7'h5b) ^ data_i[21];
		data_o[22] = (syndrome_o == 7'h5c) ^ data_i[22];
		data_o[23] = (syndrome_o == 7'h5d) ^ data_i[23];
		data_o[24] = (syndrome_o == 7'h5e) ^ data_i[24];
		data_o[25] = (syndrome_o == 7'h5f) ^ data_i[25];
		data_o[26] = (syndrome_o == 7'h61) ^ data_i[26];
		data_o[27] = (syndrome_o == 7'h62) ^ data_i[27];
		data_o[28] = (syndrome_o == 7'h63) ^ data_i[28];
		data_o[29] = (syndrome_o == 7'h64) ^ data_i[29];
		data_o[30] = (syndrome_o == 7'h65) ^ data_i[30];
		data_o[31] = (syndrome_o == 7'h66) ^ data_i[31];
		err_o[0] = syndrome_o[6];
		err_o[1] = |syndrome_o[5:0] & ~syndrome_o[6];
	end
endmodule
module prim_secded_hamming_39_32_enc (
	data_i,
	data_o
);
	input [31:0] data_i;
	output reg [38:0] data_o;
	function automatic [38:0] sv2v_cast_39;
		input reg [38:0] inp;
		sv2v_cast_39 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_39(data_i);
		data_o[32] = ^(data_o & 39'h0056aaad5b);
		data_o[33] = ^(data_o & 39'h009b33366d);
		data_o[34] = ^(data_o & 39'h00e3c3c78e);
		data_o[35] = ^(data_o & 39'h0003fc07f0);
		data_o[36] = ^(data_o & 39'h0003fff800);
		data_o[37] = ^(data_o & 39'h00fc000000);
		data_o[38] = ^(data_o & 39'h3fffffffff);
	end
endmodule
module prim_secded_hamming_72_64_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [71:0] data_i;
	output reg [63:0] data_o;
	output reg [7:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^(data_i & 72'h01ab55555556aaad5b);
		syndrome_o[1] = ^(data_i & 72'h02cd9999999b33366d);
		syndrome_o[2] = ^(data_i & 72'h04f1e1e1e1e3c3c78e);
		syndrome_o[3] = ^(data_i & 72'h0801fe01fe03fc07f0);
		syndrome_o[4] = ^(data_i & 72'h1001fffe0003fff800);
		syndrome_o[5] = ^(data_i & 72'h2001fffffffc000000);
		syndrome_o[6] = ^(data_i & 72'h40fe00000000000000);
		syndrome_o[7] = ^(data_i & 72'hffffffffffffffffff);
		data_o[0] = (syndrome_o == 8'h83) ^ data_i[0];
		data_o[1] = (syndrome_o == 8'h85) ^ data_i[1];
		data_o[2] = (syndrome_o == 8'h86) ^ data_i[2];
		data_o[3] = (syndrome_o == 8'h87) ^ data_i[3];
		data_o[4] = (syndrome_o == 8'h89) ^ data_i[4];
		data_o[5] = (syndrome_o == 8'h8a) ^ data_i[5];
		data_o[6] = (syndrome_o == 8'h8b) ^ data_i[6];
		data_o[7] = (syndrome_o == 8'h8c) ^ data_i[7];
		data_o[8] = (syndrome_o == 8'h8d) ^ data_i[8];
		data_o[9] = (syndrome_o == 8'h8e) ^ data_i[9];
		data_o[10] = (syndrome_o == 8'h8f) ^ data_i[10];
		data_o[11] = (syndrome_o == 8'h91) ^ data_i[11];
		data_o[12] = (syndrome_o == 8'h92) ^ data_i[12];
		data_o[13] = (syndrome_o == 8'h93) ^ data_i[13];
		data_o[14] = (syndrome_o == 8'h94) ^ data_i[14];
		data_o[15] = (syndrome_o == 8'h95) ^ data_i[15];
		data_o[16] = (syndrome_o == 8'h96) ^ data_i[16];
		data_o[17] = (syndrome_o == 8'h97) ^ data_i[17];
		data_o[18] = (syndrome_o == 8'h98) ^ data_i[18];
		data_o[19] = (syndrome_o == 8'h99) ^ data_i[19];
		data_o[20] = (syndrome_o == 8'h9a) ^ data_i[20];
		data_o[21] = (syndrome_o == 8'h9b) ^ data_i[21];
		data_o[22] = (syndrome_o == 8'h9c) ^ data_i[22];
		data_o[23] = (syndrome_o == 8'h9d) ^ data_i[23];
		data_o[24] = (syndrome_o == 8'h9e) ^ data_i[24];
		data_o[25] = (syndrome_o == 8'h9f) ^ data_i[25];
		data_o[26] = (syndrome_o == 8'ha1) ^ data_i[26];
		data_o[27] = (syndrome_o == 8'ha2) ^ data_i[27];
		data_o[28] = (syndrome_o == 8'ha3) ^ data_i[28];
		data_o[29] = (syndrome_o == 8'ha4) ^ data_i[29];
		data_o[30] = (syndrome_o == 8'ha5) ^ data_i[30];
		data_o[31] = (syndrome_o == 8'ha6) ^ data_i[31];
		data_o[32] = (syndrome_o == 8'ha7) ^ data_i[32];
		data_o[33] = (syndrome_o == 8'ha8) ^ data_i[33];
		data_o[34] = (syndrome_o == 8'ha9) ^ data_i[34];
		data_o[35] = (syndrome_o == 8'haa) ^ data_i[35];
		data_o[36] = (syndrome_o == 8'hab) ^ data_i[36];
		data_o[37] = (syndrome_o == 8'hac) ^ data_i[37];
		data_o[38] = (syndrome_o == 8'had) ^ data_i[38];
		data_o[39] = (syndrome_o == 8'hae) ^ data_i[39];
		data_o[40] = (syndrome_o == 8'haf) ^ data_i[40];
		data_o[41] = (syndrome_o == 8'hb0) ^ data_i[41];
		data_o[42] = (syndrome_o == 8'hb1) ^ data_i[42];
		data_o[43] = (syndrome_o == 8'hb2) ^ data_i[43];
		data_o[44] = (syndrome_o == 8'hb3) ^ data_i[44];
		data_o[45] = (syndrome_o == 8'hb4) ^ data_i[45];
		data_o[46] = (syndrome_o == 8'hb5) ^ data_i[46];
		data_o[47] = (syndrome_o == 8'hb6) ^ data_i[47];
		data_o[48] = (syndrome_o == 8'hb7) ^ data_i[48];
		data_o[49] = (syndrome_o == 8'hb8) ^ data_i[49];
		data_o[50] = (syndrome_o == 8'hb9) ^ data_i[50];
		data_o[51] = (syndrome_o == 8'hba) ^ data_i[51];
		data_o[52] = (syndrome_o == 8'hbb) ^ data_i[52];
		data_o[53] = (syndrome_o == 8'hbc) ^ data_i[53];
		data_o[54] = (syndrome_o == 8'hbd) ^ data_i[54];
		data_o[55] = (syndrome_o == 8'hbe) ^ data_i[55];
		data_o[56] = (syndrome_o == 8'hbf) ^ data_i[56];
		data_o[57] = (syndrome_o == 8'hc1) ^ data_i[57];
		data_o[58] = (syndrome_o == 8'hc2) ^ data_i[58];
		data_o[59] = (syndrome_o == 8'hc3) ^ data_i[59];
		data_o[60] = (syndrome_o == 8'hc4) ^ data_i[60];
		data_o[61] = (syndrome_o == 8'hc5) ^ data_i[61];
		data_o[62] = (syndrome_o == 8'hc6) ^ data_i[62];
		data_o[63] = (syndrome_o == 8'hc7) ^ data_i[63];
		err_o[0] = syndrome_o[7];
		err_o[1] = |syndrome_o[6:0] & ~syndrome_o[7];
	end
endmodule
module prim_secded_hamming_72_64_enc (
	data_i,
	data_o
);
	input [63:0] data_i;
	output reg [71:0] data_o;
	function automatic [71:0] sv2v_cast_72;
		input reg [71:0] inp;
		sv2v_cast_72 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_72(data_i);
		data_o[64] = ^(data_o & 72'h00ab55555556aaad5b);
		data_o[65] = ^(data_o & 72'h00cd9999999b33366d);
		data_o[66] = ^(data_o & 72'h00f1e1e1e1e3c3c78e);
		data_o[67] = ^(data_o & 72'h0001fe01fe03fc07f0);
		data_o[68] = ^(data_o & 72'h0001fffe0003fff800);
		data_o[69] = ^(data_o & 72'h0001fffffffc000000);
		data_o[70] = ^(data_o & 72'h00fe00000000000000);
		data_o[71] = ^(data_o & 72'h7fffffffffffffffff);
	end
endmodule
module prim_secded_hamming_76_68_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [75:0] data_i;
	output reg [67:0] data_o;
	output reg [7:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^(data_i & 76'h01aab55555556aaad5b);
		syndrome_o[1] = ^(data_i & 76'h02ccd9999999b33366d);
		syndrome_o[2] = ^(data_i & 76'h040f1e1e1e1e3c3c78e);
		syndrome_o[3] = ^(data_i & 76'h08f01fe01fe03fc07f0);
		syndrome_o[4] = ^(data_i & 76'h10001fffe0003fff800);
		syndrome_o[5] = ^(data_i & 76'h20001fffffffc000000);
		syndrome_o[6] = ^(data_i & 76'h40ffe00000000000000);
		syndrome_o[7] = ^(data_i & 76'hfffffffffffffffffff);
		data_o[0] = (syndrome_o == 8'h83) ^ data_i[0];
		data_o[1] = (syndrome_o == 8'h85) ^ data_i[1];
		data_o[2] = (syndrome_o == 8'h86) ^ data_i[2];
		data_o[3] = (syndrome_o == 8'h87) ^ data_i[3];
		data_o[4] = (syndrome_o == 8'h89) ^ data_i[4];
		data_o[5] = (syndrome_o == 8'h8a) ^ data_i[5];
		data_o[6] = (syndrome_o == 8'h8b) ^ data_i[6];
		data_o[7] = (syndrome_o == 8'h8c) ^ data_i[7];
		data_o[8] = (syndrome_o == 8'h8d) ^ data_i[8];
		data_o[9] = (syndrome_o == 8'h8e) ^ data_i[9];
		data_o[10] = (syndrome_o == 8'h8f) ^ data_i[10];
		data_o[11] = (syndrome_o == 8'h91) ^ data_i[11];
		data_o[12] = (syndrome_o == 8'h92) ^ data_i[12];
		data_o[13] = (syndrome_o == 8'h93) ^ data_i[13];
		data_o[14] = (syndrome_o == 8'h94) ^ data_i[14];
		data_o[15] = (syndrome_o == 8'h95) ^ data_i[15];
		data_o[16] = (syndrome_o == 8'h96) ^ data_i[16];
		data_o[17] = (syndrome_o == 8'h97) ^ data_i[17];
		data_o[18] = (syndrome_o == 8'h98) ^ data_i[18];
		data_o[19] = (syndrome_o == 8'h99) ^ data_i[19];
		data_o[20] = (syndrome_o == 8'h9a) ^ data_i[20];
		data_o[21] = (syndrome_o == 8'h9b) ^ data_i[21];
		data_o[22] = (syndrome_o == 8'h9c) ^ data_i[22];
		data_o[23] = (syndrome_o == 8'h9d) ^ data_i[23];
		data_o[24] = (syndrome_o == 8'h9e) ^ data_i[24];
		data_o[25] = (syndrome_o == 8'h9f) ^ data_i[25];
		data_o[26] = (syndrome_o == 8'ha1) ^ data_i[26];
		data_o[27] = (syndrome_o == 8'ha2) ^ data_i[27];
		data_o[28] = (syndrome_o == 8'ha3) ^ data_i[28];
		data_o[29] = (syndrome_o == 8'ha4) ^ data_i[29];
		data_o[30] = (syndrome_o == 8'ha5) ^ data_i[30];
		data_o[31] = (syndrome_o == 8'ha6) ^ data_i[31];
		data_o[32] = (syndrome_o == 8'ha7) ^ data_i[32];
		data_o[33] = (syndrome_o == 8'ha8) ^ data_i[33];
		data_o[34] = (syndrome_o == 8'ha9) ^ data_i[34];
		data_o[35] = (syndrome_o == 8'haa) ^ data_i[35];
		data_o[36] = (syndrome_o == 8'hab) ^ data_i[36];
		data_o[37] = (syndrome_o == 8'hac) ^ data_i[37];
		data_o[38] = (syndrome_o == 8'had) ^ data_i[38];
		data_o[39] = (syndrome_o == 8'hae) ^ data_i[39];
		data_o[40] = (syndrome_o == 8'haf) ^ data_i[40];
		data_o[41] = (syndrome_o == 8'hb0) ^ data_i[41];
		data_o[42] = (syndrome_o == 8'hb1) ^ data_i[42];
		data_o[43] = (syndrome_o == 8'hb2) ^ data_i[43];
		data_o[44] = (syndrome_o == 8'hb3) ^ data_i[44];
		data_o[45] = (syndrome_o == 8'hb4) ^ data_i[45];
		data_o[46] = (syndrome_o == 8'hb5) ^ data_i[46];
		data_o[47] = (syndrome_o == 8'hb6) ^ data_i[47];
		data_o[48] = (syndrome_o == 8'hb7) ^ data_i[48];
		data_o[49] = (syndrome_o == 8'hb8) ^ data_i[49];
		data_o[50] = (syndrome_o == 8'hb9) ^ data_i[50];
		data_o[51] = (syndrome_o == 8'hba) ^ data_i[51];
		data_o[52] = (syndrome_o == 8'hbb) ^ data_i[52];
		data_o[53] = (syndrome_o == 8'hbc) ^ data_i[53];
		data_o[54] = (syndrome_o == 8'hbd) ^ data_i[54];
		data_o[55] = (syndrome_o == 8'hbe) ^ data_i[55];
		data_o[56] = (syndrome_o == 8'hbf) ^ data_i[56];
		data_o[57] = (syndrome_o == 8'hc1) ^ data_i[57];
		data_o[58] = (syndrome_o == 8'hc2) ^ data_i[58];
		data_o[59] = (syndrome_o == 8'hc3) ^ data_i[59];
		data_o[60] = (syndrome_o == 8'hc4) ^ data_i[60];
		data_o[61] = (syndrome_o == 8'hc5) ^ data_i[61];
		data_o[62] = (syndrome_o == 8'hc6) ^ data_i[62];
		data_o[63] = (syndrome_o == 8'hc7) ^ data_i[63];
		data_o[64] = (syndrome_o == 8'hc8) ^ data_i[64];
		data_o[65] = (syndrome_o == 8'hc9) ^ data_i[65];
		data_o[66] = (syndrome_o == 8'hca) ^ data_i[66];
		data_o[67] = (syndrome_o == 8'hcb) ^ data_i[67];
		err_o[0] = syndrome_o[7];
		err_o[1] = |syndrome_o[6:0] & ~syndrome_o[7];
	end
endmodule
module prim_secded_hamming_76_68_enc (
	data_i,
	data_o
);
	input [67:0] data_i;
	output reg [75:0] data_o;
	function automatic [75:0] sv2v_cast_76;
		input reg [75:0] inp;
		sv2v_cast_76 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_76(data_i);
		data_o[68] = ^(data_o & 76'h00aab55555556aaad5b);
		data_o[69] = ^(data_o & 76'h00ccd9999999b33366d);
		data_o[70] = ^(data_o & 76'h000f1e1e1e1e3c3c78e);
		data_o[71] = ^(data_o & 76'h00f01fe01fe03fc07f0);
		data_o[72] = ^(data_o & 76'h00001fffe0003fff800);
		data_o[73] = ^(data_o & 76'h00001fffffffc000000);
		data_o[74] = ^(data_o & 76'h00ffe00000000000000);
		data_o[75] = ^(data_o & 76'h7ffffffffffffffffff);
	end
endmodule
module prim_secded_inv_22_16_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [21:0] data_i;
	output reg [15:0] data_o;
	output reg [5:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^((data_i ^ 22'h2a0000) & 22'h01496e);
		syndrome_o[1] = ^((data_i ^ 22'h2a0000) & 22'h02f20b);
		syndrome_o[2] = ^((data_i ^ 22'h2a0000) & 22'h048ed8);
		syndrome_o[3] = ^((data_i ^ 22'h2a0000) & 22'h087714);
		syndrome_o[4] = ^((data_i ^ 22'h2a0000) & 22'h10aca5);
		syndrome_o[5] = ^((data_i ^ 22'h2a0000) & 22'h2011f3);
		data_o[0] = (syndrome_o == 6'h32) ^ data_i[0];
		data_o[1] = (syndrome_o == 6'h23) ^ data_i[1];
		data_o[2] = (syndrome_o == 6'h19) ^ data_i[2];
		data_o[3] = (syndrome_o == 6'h07) ^ data_i[3];
		data_o[4] = (syndrome_o == 6'h2c) ^ data_i[4];
		data_o[5] = (syndrome_o == 6'h31) ^ data_i[5];
		data_o[6] = (syndrome_o == 6'h25) ^ data_i[6];
		data_o[7] = (syndrome_o == 6'h34) ^ data_i[7];
		data_o[8] = (syndrome_o == 6'h29) ^ data_i[8];
		data_o[9] = (syndrome_o == 6'h0e) ^ data_i[9];
		data_o[10] = (syndrome_o == 6'h1c) ^ data_i[10];
		data_o[11] = (syndrome_o == 6'h15) ^ data_i[11];
		data_o[12] = (syndrome_o == 6'h2a) ^ data_i[12];
		data_o[13] = (syndrome_o == 6'h1a) ^ data_i[13];
		data_o[14] = (syndrome_o == 6'h0b) ^ data_i[14];
		data_o[15] = (syndrome_o == 6'h16) ^ data_i[15];
		err_o[0] = ^syndrome_o;
		err_o[1] = ~err_o[0] & |syndrome_o;
	end
endmodule
module prim_secded_inv_22_16_enc (
	data_i,
	data_o
);
	input [15:0] data_i;
	output reg [21:0] data_o;
	function automatic [21:0] sv2v_cast_22;
		input reg [21:0] inp;
		sv2v_cast_22 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_22(data_i);
		data_o[16] = ^(data_o & 22'h00496e);
		data_o[17] = ^(data_o & 22'h00f20b);
		data_o[18] = ^(data_o & 22'h008ed8);
		data_o[19] = ^(data_o & 22'h007714);
		data_o[20] = ^(data_o & 22'h00aca5);
		data_o[21] = ^(data_o & 22'h0011f3);
		data_o = data_o ^ 22'h2a0000;
	end
endmodule
module prim_secded_inv_28_22_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [27:0] data_i;
	output reg [21:0] data_o;
	output reg [5:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^((data_i ^ 28'ha800000) & 28'h07003ff);
		syndrome_o[1] = ^((data_i ^ 28'ha800000) & 28'h090fc0f);
		syndrome_o[2] = ^((data_i ^ 28'ha800000) & 28'h1271c71);
		syndrome_o[3] = ^((data_i ^ 28'ha800000) & 28'h23b6592);
		syndrome_o[4] = ^((data_i ^ 28'ha800000) & 28'h43daaa4);
		syndrome_o[5] = ^((data_i ^ 28'ha800000) & 28'h83ed348);
		data_o[0] = (syndrome_o == 6'h07) ^ data_i[0];
		data_o[1] = (syndrome_o == 6'h0b) ^ data_i[1];
		data_o[2] = (syndrome_o == 6'h13) ^ data_i[2];
		data_o[3] = (syndrome_o == 6'h23) ^ data_i[3];
		data_o[4] = (syndrome_o == 6'h0d) ^ data_i[4];
		data_o[5] = (syndrome_o == 6'h15) ^ data_i[5];
		data_o[6] = (syndrome_o == 6'h25) ^ data_i[6];
		data_o[7] = (syndrome_o == 6'h19) ^ data_i[7];
		data_o[8] = (syndrome_o == 6'h29) ^ data_i[8];
		data_o[9] = (syndrome_o == 6'h31) ^ data_i[9];
		data_o[10] = (syndrome_o == 6'h0e) ^ data_i[10];
		data_o[11] = (syndrome_o == 6'h16) ^ data_i[11];
		data_o[12] = (syndrome_o == 6'h26) ^ data_i[12];
		data_o[13] = (syndrome_o == 6'h1a) ^ data_i[13];
		data_o[14] = (syndrome_o == 6'h2a) ^ data_i[14];
		data_o[15] = (syndrome_o == 6'h32) ^ data_i[15];
		data_o[16] = (syndrome_o == 6'h1c) ^ data_i[16];
		data_o[17] = (syndrome_o == 6'h2c) ^ data_i[17];
		data_o[18] = (syndrome_o == 6'h34) ^ data_i[18];
		data_o[19] = (syndrome_o == 6'h38) ^ data_i[19];
		data_o[20] = (syndrome_o == 6'h3b) ^ data_i[20];
		data_o[21] = (syndrome_o == 6'h3d) ^ data_i[21];
		err_o[0] = ^syndrome_o;
		err_o[1] = ~err_o[0] & |syndrome_o;
	end
endmodule
module prim_secded_inv_28_22_enc (
	data_i,
	data_o
);
	input [21:0] data_i;
	output reg [27:0] data_o;
	function automatic [27:0] sv2v_cast_28;
		input reg [27:0] inp;
		sv2v_cast_28 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_28(data_i);
		data_o[22] = ^(data_o & 28'h03003ff);
		data_o[23] = ^(data_o & 28'h010fc0f);
		data_o[24] = ^(data_o & 28'h0271c71);
		data_o[25] = ^(data_o & 28'h03b6592);
		data_o[26] = ^(data_o & 28'h03daaa4);
		data_o[27] = ^(data_o & 28'h03ed348);
		data_o = data_o ^ 28'ha800000;
	end
endmodule
module prim_secded_inv_39_32_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [38:0] data_i;
	output reg [31:0] data_o;
	output reg [6:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^((data_i ^ 39'h2a00000000) & 39'h012606bd25);
		syndrome_o[1] = ^((data_i ^ 39'h2a00000000) & 39'h02deba8050);
		syndrome_o[2] = ^((data_i ^ 39'h2a00000000) & 39'h04413d89aa);
		syndrome_o[3] = ^((data_i ^ 39'h2a00000000) & 39'h0831234ed1);
		syndrome_o[4] = ^((data_i ^ 39'h2a00000000) & 39'h10c2c1323b);
		syndrome_o[5] = ^((data_i ^ 39'h2a00000000) & 39'h202dcc624c);
		syndrome_o[6] = ^((data_i ^ 39'h2a00000000) & 39'h4098505586);
		data_o[0] = (syndrome_o == 7'h19) ^ data_i[0];
		data_o[1] = (syndrome_o == 7'h54) ^ data_i[1];
		data_o[2] = (syndrome_o == 7'h61) ^ data_i[2];
		data_o[3] = (syndrome_o == 7'h34) ^ data_i[3];
		data_o[4] = (syndrome_o == 7'h1a) ^ data_i[4];
		data_o[5] = (syndrome_o == 7'h15) ^ data_i[5];
		data_o[6] = (syndrome_o == 7'h2a) ^ data_i[6];
		data_o[7] = (syndrome_o == 7'h4c) ^ data_i[7];
		data_o[8] = (syndrome_o == 7'h45) ^ data_i[8];
		data_o[9] = (syndrome_o == 7'h38) ^ data_i[9];
		data_o[10] = (syndrome_o == 7'h49) ^ data_i[10];
		data_o[11] = (syndrome_o == 7'h0d) ^ data_i[11];
		data_o[12] = (syndrome_o == 7'h51) ^ data_i[12];
		data_o[13] = (syndrome_o == 7'h31) ^ data_i[13];
		data_o[14] = (syndrome_o == 7'h68) ^ data_i[14];
		data_o[15] = (syndrome_o == 7'h07) ^ data_i[15];
		data_o[16] = (syndrome_o == 7'h1c) ^ data_i[16];
		data_o[17] = (syndrome_o == 7'h0b) ^ data_i[17];
		data_o[18] = (syndrome_o == 7'h25) ^ data_i[18];
		data_o[19] = (syndrome_o == 7'h26) ^ data_i[19];
		data_o[20] = (syndrome_o == 7'h46) ^ data_i[20];
		data_o[21] = (syndrome_o == 7'h0e) ^ data_i[21];
		data_o[22] = (syndrome_o == 7'h70) ^ data_i[22];
		data_o[23] = (syndrome_o == 7'h32) ^ data_i[23];
		data_o[24] = (syndrome_o == 7'h2c) ^ data_i[24];
		data_o[25] = (syndrome_o == 7'h13) ^ data_i[25];
		data_o[26] = (syndrome_o == 7'h23) ^ data_i[26];
		data_o[27] = (syndrome_o == 7'h62) ^ data_i[27];
		data_o[28] = (syndrome_o == 7'h4a) ^ data_i[28];
		data_o[29] = (syndrome_o == 7'h29) ^ data_i[29];
		data_o[30] = (syndrome_o == 7'h16) ^ data_i[30];
		data_o[31] = (syndrome_o == 7'h52) ^ data_i[31];
		err_o[0] = ^syndrome_o;
		err_o[1] = ~err_o[0] & |syndrome_o;
	end
endmodule
module prim_secded_inv_39_32_enc (
	data_i,
	data_o
);
	input [31:0] data_i;
	output reg [38:0] data_o;
	function automatic [38:0] sv2v_cast_39;
		input reg [38:0] inp;
		sv2v_cast_39 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_39(data_i);
		data_o[32] = ^(data_o & 39'h002606bd25);
		data_o[33] = ^(data_o & 39'h00deba8050);
		data_o[34] = ^(data_o & 39'h00413d89aa);
		data_o[35] = ^(data_o & 39'h0031234ed1);
		data_o[36] = ^(data_o & 39'h00c2c1323b);
		data_o[37] = ^(data_o & 39'h002dcc624c);
		data_o[38] = ^(data_o & 39'h0098505586);
		data_o = data_o ^ 39'h2a00000000;
	end
endmodule
module prim_secded_inv_64_57_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [63:0] data_i;
	output reg [56:0] data_o;
	output reg [6:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^((data_i ^ 64'h5400000000000000) & 64'h0303fff800007fff);
		syndrome_o[1] = ^((data_i ^ 64'h5400000000000000) & 64'h057c1ff801ff801f);
		syndrome_o[2] = ^((data_i ^ 64'h5400000000000000) & 64'h09bde1f87e0781e1);
		syndrome_o[3] = ^((data_i ^ 64'h5400000000000000) & 64'h11deee3b8e388e22);
		syndrome_o[4] = ^((data_i ^ 64'h5400000000000000) & 64'h21ef76cdb2c93244);
		syndrome_o[5] = ^((data_i ^ 64'h5400000000000000) & 64'h41f7bb56d5525488);
		syndrome_o[6] = ^((data_i ^ 64'h5400000000000000) & 64'h81fbdda769a46910);
		data_o[0] = (syndrome_o == 7'h07) ^ data_i[0];
		data_o[1] = (syndrome_o == 7'h0b) ^ data_i[1];
		data_o[2] = (syndrome_o == 7'h13) ^ data_i[2];
		data_o[3] = (syndrome_o == 7'h23) ^ data_i[3];
		data_o[4] = (syndrome_o == 7'h43) ^ data_i[4];
		data_o[5] = (syndrome_o == 7'h0d) ^ data_i[5];
		data_o[6] = (syndrome_o == 7'h15) ^ data_i[6];
		data_o[7] = (syndrome_o == 7'h25) ^ data_i[7];
		data_o[8] = (syndrome_o == 7'h45) ^ data_i[8];
		data_o[9] = (syndrome_o == 7'h19) ^ data_i[9];
		data_o[10] = (syndrome_o == 7'h29) ^ data_i[10];
		data_o[11] = (syndrome_o == 7'h49) ^ data_i[11];
		data_o[12] = (syndrome_o == 7'h31) ^ data_i[12];
		data_o[13] = (syndrome_o == 7'h51) ^ data_i[13];
		data_o[14] = (syndrome_o == 7'h61) ^ data_i[14];
		data_o[15] = (syndrome_o == 7'h0e) ^ data_i[15];
		data_o[16] = (syndrome_o == 7'h16) ^ data_i[16];
		data_o[17] = (syndrome_o == 7'h26) ^ data_i[17];
		data_o[18] = (syndrome_o == 7'h46) ^ data_i[18];
		data_o[19] = (syndrome_o == 7'h1a) ^ data_i[19];
		data_o[20] = (syndrome_o == 7'h2a) ^ data_i[20];
		data_o[21] = (syndrome_o == 7'h4a) ^ data_i[21];
		data_o[22] = (syndrome_o == 7'h32) ^ data_i[22];
		data_o[23] = (syndrome_o == 7'h52) ^ data_i[23];
		data_o[24] = (syndrome_o == 7'h62) ^ data_i[24];
		data_o[25] = (syndrome_o == 7'h1c) ^ data_i[25];
		data_o[26] = (syndrome_o == 7'h2c) ^ data_i[26];
		data_o[27] = (syndrome_o == 7'h4c) ^ data_i[27];
		data_o[28] = (syndrome_o == 7'h34) ^ data_i[28];
		data_o[29] = (syndrome_o == 7'h54) ^ data_i[29];
		data_o[30] = (syndrome_o == 7'h64) ^ data_i[30];
		data_o[31] = (syndrome_o == 7'h38) ^ data_i[31];
		data_o[32] = (syndrome_o == 7'h58) ^ data_i[32];
		data_o[33] = (syndrome_o == 7'h68) ^ data_i[33];
		data_o[34] = (syndrome_o == 7'h70) ^ data_i[34];
		data_o[35] = (syndrome_o == 7'h1f) ^ data_i[35];
		data_o[36] = (syndrome_o == 7'h2f) ^ data_i[36];
		data_o[37] = (syndrome_o == 7'h4f) ^ data_i[37];
		data_o[38] = (syndrome_o == 7'h37) ^ data_i[38];
		data_o[39] = (syndrome_o == 7'h57) ^ data_i[39];
		data_o[40] = (syndrome_o == 7'h67) ^ data_i[40];
		data_o[41] = (syndrome_o == 7'h3b) ^ data_i[41];
		data_o[42] = (syndrome_o == 7'h5b) ^ data_i[42];
		data_o[43] = (syndrome_o == 7'h6b) ^ data_i[43];
		data_o[44] = (syndrome_o == 7'h73) ^ data_i[44];
		data_o[45] = (syndrome_o == 7'h3d) ^ data_i[45];
		data_o[46] = (syndrome_o == 7'h5d) ^ data_i[46];
		data_o[47] = (syndrome_o == 7'h6d) ^ data_i[47];
		data_o[48] = (syndrome_o == 7'h75) ^ data_i[48];
		data_o[49] = (syndrome_o == 7'h79) ^ data_i[49];
		data_o[50] = (syndrome_o == 7'h3e) ^ data_i[50];
		data_o[51] = (syndrome_o == 7'h5e) ^ data_i[51];
		data_o[52] = (syndrome_o == 7'h6e) ^ data_i[52];
		data_o[53] = (syndrome_o == 7'h76) ^ data_i[53];
		data_o[54] = (syndrome_o == 7'h7a) ^ data_i[54];
		data_o[55] = (syndrome_o == 7'h7c) ^ data_i[55];
		data_o[56] = (syndrome_o == 7'h7f) ^ data_i[56];
		err_o[0] = ^syndrome_o;
		err_o[1] = ~err_o[0] & |syndrome_o;
	end
endmodule
module prim_secded_inv_64_57_enc (
	data_i,
	data_o
);
	input [56:0] data_i;
	output reg [63:0] data_o;
	function automatic [63:0] sv2v_cast_64;
		input reg [63:0] inp;
		sv2v_cast_64 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_64(data_i);
		data_o[57] = ^(data_o & 64'h0103fff800007fff);
		data_o[58] = ^(data_o & 64'h017c1ff801ff801f);
		data_o[59] = ^(data_o & 64'h01bde1f87e0781e1);
		data_o[60] = ^(data_o & 64'h01deee3b8e388e22);
		data_o[61] = ^(data_o & 64'h01ef76cdb2c93244);
		data_o[62] = ^(data_o & 64'h01f7bb56d5525488);
		data_o[63] = ^(data_o & 64'h01fbdda769a46910);
		data_o = data_o ^ 64'h5400000000000000;
	end
endmodule
module prim_secded_inv_72_64_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [71:0] data_i;
	output reg [63:0] data_o;
	output reg [7:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^((data_i ^ 72'haa0000000000000000) & 72'h01b9000000001fffff);
		syndrome_o[1] = ^((data_i ^ 72'haa0000000000000000) & 72'h025e00000fffe0003f);
		syndrome_o[2] = ^((data_i ^ 72'haa0000000000000000) & 72'h0467003ff003e007c1);
		syndrome_o[3] = ^((data_i ^ 72'haa0000000000000000) & 72'h08cd0fc0f03c207842);
		syndrome_o[4] = ^((data_i ^ 72'haa0000000000000000) & 72'h10b671c711c4438884);
		syndrome_o[5] = ^((data_i ^ 72'haa0000000000000000) & 72'h20b5b65926488c9108);
		syndrome_o[6] = ^((data_i ^ 72'haa0000000000000000) & 72'h40cbdaaa4a91152210);
		syndrome_o[7] = ^((data_i ^ 72'haa0000000000000000) & 72'h807aed348d221a4420);
		data_o[0] = (syndrome_o == 8'h07) ^ data_i[0];
		data_o[1] = (syndrome_o == 8'h0b) ^ data_i[1];
		data_o[2] = (syndrome_o == 8'h13) ^ data_i[2];
		data_o[3] = (syndrome_o == 8'h23) ^ data_i[3];
		data_o[4] = (syndrome_o == 8'h43) ^ data_i[4];
		data_o[5] = (syndrome_o == 8'h83) ^ data_i[5];
		data_o[6] = (syndrome_o == 8'h0d) ^ data_i[6];
		data_o[7] = (syndrome_o == 8'h15) ^ data_i[7];
		data_o[8] = (syndrome_o == 8'h25) ^ data_i[8];
		data_o[9] = (syndrome_o == 8'h45) ^ data_i[9];
		data_o[10] = (syndrome_o == 8'h85) ^ data_i[10];
		data_o[11] = (syndrome_o == 8'h19) ^ data_i[11];
		data_o[12] = (syndrome_o == 8'h29) ^ data_i[12];
		data_o[13] = (syndrome_o == 8'h49) ^ data_i[13];
		data_o[14] = (syndrome_o == 8'h89) ^ data_i[14];
		data_o[15] = (syndrome_o == 8'h31) ^ data_i[15];
		data_o[16] = (syndrome_o == 8'h51) ^ data_i[16];
		data_o[17] = (syndrome_o == 8'h91) ^ data_i[17];
		data_o[18] = (syndrome_o == 8'h61) ^ data_i[18];
		data_o[19] = (syndrome_o == 8'ha1) ^ data_i[19];
		data_o[20] = (syndrome_o == 8'hc1) ^ data_i[20];
		data_o[21] = (syndrome_o == 8'h0e) ^ data_i[21];
		data_o[22] = (syndrome_o == 8'h16) ^ data_i[22];
		data_o[23] = (syndrome_o == 8'h26) ^ data_i[23];
		data_o[24] = (syndrome_o == 8'h46) ^ data_i[24];
		data_o[25] = (syndrome_o == 8'h86) ^ data_i[25];
		data_o[26] = (syndrome_o == 8'h1a) ^ data_i[26];
		data_o[27] = (syndrome_o == 8'h2a) ^ data_i[27];
		data_o[28] = (syndrome_o == 8'h4a) ^ data_i[28];
		data_o[29] = (syndrome_o == 8'h8a) ^ data_i[29];
		data_o[30] = (syndrome_o == 8'h32) ^ data_i[30];
		data_o[31] = (syndrome_o == 8'h52) ^ data_i[31];
		data_o[32] = (syndrome_o == 8'h92) ^ data_i[32];
		data_o[33] = (syndrome_o == 8'h62) ^ data_i[33];
		data_o[34] = (syndrome_o == 8'ha2) ^ data_i[34];
		data_o[35] = (syndrome_o == 8'hc2) ^ data_i[35];
		data_o[36] = (syndrome_o == 8'h1c) ^ data_i[36];
		data_o[37] = (syndrome_o == 8'h2c) ^ data_i[37];
		data_o[38] = (syndrome_o == 8'h4c) ^ data_i[38];
		data_o[39] = (syndrome_o == 8'h8c) ^ data_i[39];
		data_o[40] = (syndrome_o == 8'h34) ^ data_i[40];
		data_o[41] = (syndrome_o == 8'h54) ^ data_i[41];
		data_o[42] = (syndrome_o == 8'h94) ^ data_i[42];
		data_o[43] = (syndrome_o == 8'h64) ^ data_i[43];
		data_o[44] = (syndrome_o == 8'ha4) ^ data_i[44];
		data_o[45] = (syndrome_o == 8'hc4) ^ data_i[45];
		data_o[46] = (syndrome_o == 8'h38) ^ data_i[46];
		data_o[47] = (syndrome_o == 8'h58) ^ data_i[47];
		data_o[48] = (syndrome_o == 8'h98) ^ data_i[48];
		data_o[49] = (syndrome_o == 8'h68) ^ data_i[49];
		data_o[50] = (syndrome_o == 8'ha8) ^ data_i[50];
		data_o[51] = (syndrome_o == 8'hc8) ^ data_i[51];
		data_o[52] = (syndrome_o == 8'h70) ^ data_i[52];
		data_o[53] = (syndrome_o == 8'hb0) ^ data_i[53];
		data_o[54] = (syndrome_o == 8'hd0) ^ data_i[54];
		data_o[55] = (syndrome_o == 8'he0) ^ data_i[55];
		data_o[56] = (syndrome_o == 8'h6d) ^ data_i[56];
		data_o[57] = (syndrome_o == 8'hd6) ^ data_i[57];
		data_o[58] = (syndrome_o == 8'h3e) ^ data_i[58];
		data_o[59] = (syndrome_o == 8'hcb) ^ data_i[59];
		data_o[60] = (syndrome_o == 8'hb3) ^ data_i[60];
		data_o[61] = (syndrome_o == 8'hb5) ^ data_i[61];
		data_o[62] = (syndrome_o == 8'hce) ^ data_i[62];
		data_o[63] = (syndrome_o == 8'h79) ^ data_i[63];
		err_o[0] = ^syndrome_o;
		err_o[1] = ~err_o[0] & |syndrome_o;
	end
endmodule
module prim_secded_inv_72_64_enc (
	data_i,
	data_o
);
	input [63:0] data_i;
	output reg [71:0] data_o;
	function automatic [71:0] sv2v_cast_72;
		input reg [71:0] inp;
		sv2v_cast_72 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_72(data_i);
		data_o[64] = ^(data_o & 72'h00b9000000001fffff);
		data_o[65] = ^(data_o & 72'h005e00000fffe0003f);
		data_o[66] = ^(data_o & 72'h0067003ff003e007c1);
		data_o[67] = ^(data_o & 72'h00cd0fc0f03c207842);
		data_o[68] = ^(data_o & 72'h00b671c711c4438884);
		data_o[69] = ^(data_o & 72'h00b5b65926488c9108);
		data_o[70] = ^(data_o & 72'h00cbdaaa4a91152210);
		data_o[71] = ^(data_o & 72'h007aed348d221a4420);
		data_o = data_o ^ 72'haa0000000000000000;
	end
endmodule
module prim_secded_inv_hamming_22_16_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [21:0] data_i;
	output reg [15:0] data_o;
	output reg [5:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^((data_i ^ 22'h2a0000) & 22'h01ad5b);
		syndrome_o[1] = ^((data_i ^ 22'h2a0000) & 22'h02366d);
		syndrome_o[2] = ^((data_i ^ 22'h2a0000) & 22'h04c78e);
		syndrome_o[3] = ^((data_i ^ 22'h2a0000) & 22'h0807f0);
		syndrome_o[4] = ^((data_i ^ 22'h2a0000) & 22'h10f800);
		syndrome_o[5] = ^((data_i ^ 22'h2a0000) & 22'h3fffff);
		data_o[0] = (syndrome_o == 6'h23) ^ data_i[0];
		data_o[1] = (syndrome_o == 6'h25) ^ data_i[1];
		data_o[2] = (syndrome_o == 6'h26) ^ data_i[2];
		data_o[3] = (syndrome_o == 6'h27) ^ data_i[3];
		data_o[4] = (syndrome_o == 6'h29) ^ data_i[4];
		data_o[5] = (syndrome_o == 6'h2a) ^ data_i[5];
		data_o[6] = (syndrome_o == 6'h2b) ^ data_i[6];
		data_o[7] = (syndrome_o == 6'h2c) ^ data_i[7];
		data_o[8] = (syndrome_o == 6'h2d) ^ data_i[8];
		data_o[9] = (syndrome_o == 6'h2e) ^ data_i[9];
		data_o[10] = (syndrome_o == 6'h2f) ^ data_i[10];
		data_o[11] = (syndrome_o == 6'h31) ^ data_i[11];
		data_o[12] = (syndrome_o == 6'h32) ^ data_i[12];
		data_o[13] = (syndrome_o == 6'h33) ^ data_i[13];
		data_o[14] = (syndrome_o == 6'h34) ^ data_i[14];
		data_o[15] = (syndrome_o == 6'h35) ^ data_i[15];
		err_o[0] = syndrome_o[5];
		err_o[1] = |syndrome_o[4:0] & ~syndrome_o[5];
	end
endmodule
module prim_secded_inv_hamming_22_16_enc (
	data_i,
	data_o
);
	input [15:0] data_i;
	output reg [21:0] data_o;
	function automatic [21:0] sv2v_cast_22;
		input reg [21:0] inp;
		sv2v_cast_22 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_22(data_i);
		data_o[16] = ^(data_o & 22'h00ad5b);
		data_o[17] = ^(data_o & 22'h00366d);
		data_o[18] = ^(data_o & 22'h00c78e);
		data_o[19] = ^(data_o & 22'h0007f0);
		data_o[20] = ^(data_o & 22'h00f800);
		data_o[21] = ^(data_o & 22'h1fffff);
		data_o = data_o ^ 22'h2a0000;
	end
endmodule
module prim_secded_inv_hamming_39_32_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [38:0] data_i;
	output reg [31:0] data_o;
	output reg [6:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^((data_i ^ 39'h2a00000000) & 39'h0156aaad5b);
		syndrome_o[1] = ^((data_i ^ 39'h2a00000000) & 39'h029b33366d);
		syndrome_o[2] = ^((data_i ^ 39'h2a00000000) & 39'h04e3c3c78e);
		syndrome_o[3] = ^((data_i ^ 39'h2a00000000) & 39'h0803fc07f0);
		syndrome_o[4] = ^((data_i ^ 39'h2a00000000) & 39'h1003fff800);
		syndrome_o[5] = ^((data_i ^ 39'h2a00000000) & 39'h20fc000000);
		syndrome_o[6] = ^((data_i ^ 39'h2a00000000) & 39'h7fffffffff);
		data_o[0] = (syndrome_o == 7'h43) ^ data_i[0];
		data_o[1] = (syndrome_o == 7'h45) ^ data_i[1];
		data_o[2] = (syndrome_o == 7'h46) ^ data_i[2];
		data_o[3] = (syndrome_o == 7'h47) ^ data_i[3];
		data_o[4] = (syndrome_o == 7'h49) ^ data_i[4];
		data_o[5] = (syndrome_o == 7'h4a) ^ data_i[5];
		data_o[6] = (syndrome_o == 7'h4b) ^ data_i[6];
		data_o[7] = (syndrome_o == 7'h4c) ^ data_i[7];
		data_o[8] = (syndrome_o == 7'h4d) ^ data_i[8];
		data_o[9] = (syndrome_o == 7'h4e) ^ data_i[9];
		data_o[10] = (syndrome_o == 7'h4f) ^ data_i[10];
		data_o[11] = (syndrome_o == 7'h51) ^ data_i[11];
		data_o[12] = (syndrome_o == 7'h52) ^ data_i[12];
		data_o[13] = (syndrome_o == 7'h53) ^ data_i[13];
		data_o[14] = (syndrome_o == 7'h54) ^ data_i[14];
		data_o[15] = (syndrome_o == 7'h55) ^ data_i[15];
		data_o[16] = (syndrome_o == 7'h56) ^ data_i[16];
		data_o[17] = (syndrome_o == 7'h57) ^ data_i[17];
		data_o[18] = (syndrome_o == 7'h58) ^ data_i[18];
		data_o[19] = (syndrome_o == 7'h59) ^ data_i[19];
		data_o[20] = (syndrome_o == 7'h5a) ^ data_i[20];
		data_o[21] = (syndrome_o == 7'h5b) ^ data_i[21];
		data_o[22] = (syndrome_o == 7'h5c) ^ data_i[22];
		data_o[23] = (syndrome_o == 7'h5d) ^ data_i[23];
		data_o[24] = (syndrome_o == 7'h5e) ^ data_i[24];
		data_o[25] = (syndrome_o == 7'h5f) ^ data_i[25];
		data_o[26] = (syndrome_o == 7'h61) ^ data_i[26];
		data_o[27] = (syndrome_o == 7'h62) ^ data_i[27];
		data_o[28] = (syndrome_o == 7'h63) ^ data_i[28];
		data_o[29] = (syndrome_o == 7'h64) ^ data_i[29];
		data_o[30] = (syndrome_o == 7'h65) ^ data_i[30];
		data_o[31] = (syndrome_o == 7'h66) ^ data_i[31];
		err_o[0] = syndrome_o[6];
		err_o[1] = |syndrome_o[5:0] & ~syndrome_o[6];
	end
endmodule
module prim_secded_inv_hamming_39_32_enc (
	data_i,
	data_o
);
	input [31:0] data_i;
	output reg [38:0] data_o;
	function automatic [38:0] sv2v_cast_39;
		input reg [38:0] inp;
		sv2v_cast_39 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_39(data_i);
		data_o[32] = ^(data_o & 39'h0056aaad5b);
		data_o[33] = ^(data_o & 39'h009b33366d);
		data_o[34] = ^(data_o & 39'h00e3c3c78e);
		data_o[35] = ^(data_o & 39'h0003fc07f0);
		data_o[36] = ^(data_o & 39'h0003fff800);
		data_o[37] = ^(data_o & 39'h00fc000000);
		data_o[38] = ^(data_o & 39'h3fffffffff);
		data_o = data_o ^ 39'h2a00000000;
	end
endmodule
module prim_secded_inv_hamming_72_64_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [71:0] data_i;
	output reg [63:0] data_o;
	output reg [7:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^((data_i ^ 72'haa0000000000000000) & 72'h01ab55555556aaad5b);
		syndrome_o[1] = ^((data_i ^ 72'haa0000000000000000) & 72'h02cd9999999b33366d);
		syndrome_o[2] = ^((data_i ^ 72'haa0000000000000000) & 72'h04f1e1e1e1e3c3c78e);
		syndrome_o[3] = ^((data_i ^ 72'haa0000000000000000) & 72'h0801fe01fe03fc07f0);
		syndrome_o[4] = ^((data_i ^ 72'haa0000000000000000) & 72'h1001fffe0003fff800);
		syndrome_o[5] = ^((data_i ^ 72'haa0000000000000000) & 72'h2001fffffffc000000);
		syndrome_o[6] = ^((data_i ^ 72'haa0000000000000000) & 72'h40fe00000000000000);
		syndrome_o[7] = ^((data_i ^ 72'haa0000000000000000) & 72'hffffffffffffffffff);
		data_o[0] = (syndrome_o == 8'h83) ^ data_i[0];
		data_o[1] = (syndrome_o == 8'h85) ^ data_i[1];
		data_o[2] = (syndrome_o == 8'h86) ^ data_i[2];
		data_o[3] = (syndrome_o == 8'h87) ^ data_i[3];
		data_o[4] = (syndrome_o == 8'h89) ^ data_i[4];
		data_o[5] = (syndrome_o == 8'h8a) ^ data_i[5];
		data_o[6] = (syndrome_o == 8'h8b) ^ data_i[6];
		data_o[7] = (syndrome_o == 8'h8c) ^ data_i[7];
		data_o[8] = (syndrome_o == 8'h8d) ^ data_i[8];
		data_o[9] = (syndrome_o == 8'h8e) ^ data_i[9];
		data_o[10] = (syndrome_o == 8'h8f) ^ data_i[10];
		data_o[11] = (syndrome_o == 8'h91) ^ data_i[11];
		data_o[12] = (syndrome_o == 8'h92) ^ data_i[12];
		data_o[13] = (syndrome_o == 8'h93) ^ data_i[13];
		data_o[14] = (syndrome_o == 8'h94) ^ data_i[14];
		data_o[15] = (syndrome_o == 8'h95) ^ data_i[15];
		data_o[16] = (syndrome_o == 8'h96) ^ data_i[16];
		data_o[17] = (syndrome_o == 8'h97) ^ data_i[17];
		data_o[18] = (syndrome_o == 8'h98) ^ data_i[18];
		data_o[19] = (syndrome_o == 8'h99) ^ data_i[19];
		data_o[20] = (syndrome_o == 8'h9a) ^ data_i[20];
		data_o[21] = (syndrome_o == 8'h9b) ^ data_i[21];
		data_o[22] = (syndrome_o == 8'h9c) ^ data_i[22];
		data_o[23] = (syndrome_o == 8'h9d) ^ data_i[23];
		data_o[24] = (syndrome_o == 8'h9e) ^ data_i[24];
		data_o[25] = (syndrome_o == 8'h9f) ^ data_i[25];
		data_o[26] = (syndrome_o == 8'ha1) ^ data_i[26];
		data_o[27] = (syndrome_o == 8'ha2) ^ data_i[27];
		data_o[28] = (syndrome_o == 8'ha3) ^ data_i[28];
		data_o[29] = (syndrome_o == 8'ha4) ^ data_i[29];
		data_o[30] = (syndrome_o == 8'ha5) ^ data_i[30];
		data_o[31] = (syndrome_o == 8'ha6) ^ data_i[31];
		data_o[32] = (syndrome_o == 8'ha7) ^ data_i[32];
		data_o[33] = (syndrome_o == 8'ha8) ^ data_i[33];
		data_o[34] = (syndrome_o == 8'ha9) ^ data_i[34];
		data_o[35] = (syndrome_o == 8'haa) ^ data_i[35];
		data_o[36] = (syndrome_o == 8'hab) ^ data_i[36];
		data_o[37] = (syndrome_o == 8'hac) ^ data_i[37];
		data_o[38] = (syndrome_o == 8'had) ^ data_i[38];
		data_o[39] = (syndrome_o == 8'hae) ^ data_i[39];
		data_o[40] = (syndrome_o == 8'haf) ^ data_i[40];
		data_o[41] = (syndrome_o == 8'hb0) ^ data_i[41];
		data_o[42] = (syndrome_o == 8'hb1) ^ data_i[42];
		data_o[43] = (syndrome_o == 8'hb2) ^ data_i[43];
		data_o[44] = (syndrome_o == 8'hb3) ^ data_i[44];
		data_o[45] = (syndrome_o == 8'hb4) ^ data_i[45];
		data_o[46] = (syndrome_o == 8'hb5) ^ data_i[46];
		data_o[47] = (syndrome_o == 8'hb6) ^ data_i[47];
		data_o[48] = (syndrome_o == 8'hb7) ^ data_i[48];
		data_o[49] = (syndrome_o == 8'hb8) ^ data_i[49];
		data_o[50] = (syndrome_o == 8'hb9) ^ data_i[50];
		data_o[51] = (syndrome_o == 8'hba) ^ data_i[51];
		data_o[52] = (syndrome_o == 8'hbb) ^ data_i[52];
		data_o[53] = (syndrome_o == 8'hbc) ^ data_i[53];
		data_o[54] = (syndrome_o == 8'hbd) ^ data_i[54];
		data_o[55] = (syndrome_o == 8'hbe) ^ data_i[55];
		data_o[56] = (syndrome_o == 8'hbf) ^ data_i[56];
		data_o[57] = (syndrome_o == 8'hc1) ^ data_i[57];
		data_o[58] = (syndrome_o == 8'hc2) ^ data_i[58];
		data_o[59] = (syndrome_o == 8'hc3) ^ data_i[59];
		data_o[60] = (syndrome_o == 8'hc4) ^ data_i[60];
		data_o[61] = (syndrome_o == 8'hc5) ^ data_i[61];
		data_o[62] = (syndrome_o == 8'hc6) ^ data_i[62];
		data_o[63] = (syndrome_o == 8'hc7) ^ data_i[63];
		err_o[0] = syndrome_o[7];
		err_o[1] = |syndrome_o[6:0] & ~syndrome_o[7];
	end
endmodule
module prim_secded_inv_hamming_72_64_enc (
	data_i,
	data_o
);
	input [63:0] data_i;
	output reg [71:0] data_o;
	function automatic [71:0] sv2v_cast_72;
		input reg [71:0] inp;
		sv2v_cast_72 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_72(data_i);
		data_o[64] = ^(data_o & 72'h00ab55555556aaad5b);
		data_o[65] = ^(data_o & 72'h00cd9999999b33366d);
		data_o[66] = ^(data_o & 72'h00f1e1e1e1e3c3c78e);
		data_o[67] = ^(data_o & 72'h0001fe01fe03fc07f0);
		data_o[68] = ^(data_o & 72'h0001fffe0003fff800);
		data_o[69] = ^(data_o & 72'h0001fffffffc000000);
		data_o[70] = ^(data_o & 72'h00fe00000000000000);
		data_o[71] = ^(data_o & 72'h7fffffffffffffffff);
		data_o = data_o ^ 72'haa0000000000000000;
	end
endmodule
module prim_secded_inv_hamming_76_68_dec (
	data_i,
	data_o,
	syndrome_o,
	err_o
);
	input [75:0] data_i;
	output reg [67:0] data_o;
	output reg [7:0] syndrome_o;
	output reg [1:0] err_o;
	always @(*) begin : p_encode
		syndrome_o[0] = ^((data_i ^ 76'haa00000000000000000) & 76'h01aab55555556aaad5b);
		syndrome_o[1] = ^((data_i ^ 76'haa00000000000000000) & 76'h02ccd9999999b33366d);
		syndrome_o[2] = ^((data_i ^ 76'haa00000000000000000) & 76'h040f1e1e1e1e3c3c78e);
		syndrome_o[3] = ^((data_i ^ 76'haa00000000000000000) & 76'h08f01fe01fe03fc07f0);
		syndrome_o[4] = ^((data_i ^ 76'haa00000000000000000) & 76'h10001fffe0003fff800);
		syndrome_o[5] = ^((data_i ^ 76'haa00000000000000000) & 76'h20001fffffffc000000);
		syndrome_o[6] = ^((data_i ^ 76'haa00000000000000000) & 76'h40ffe00000000000000);
		syndrome_o[7] = ^((data_i ^ 76'haa00000000000000000) & 76'hfffffffffffffffffff);
		data_o[0] = (syndrome_o == 8'h83) ^ data_i[0];
		data_o[1] = (syndrome_o == 8'h85) ^ data_i[1];
		data_o[2] = (syndrome_o == 8'h86) ^ data_i[2];
		data_o[3] = (syndrome_o == 8'h87) ^ data_i[3];
		data_o[4] = (syndrome_o == 8'h89) ^ data_i[4];
		data_o[5] = (syndrome_o == 8'h8a) ^ data_i[5];
		data_o[6] = (syndrome_o == 8'h8b) ^ data_i[6];
		data_o[7] = (syndrome_o == 8'h8c) ^ data_i[7];
		data_o[8] = (syndrome_o == 8'h8d) ^ data_i[8];
		data_o[9] = (syndrome_o == 8'h8e) ^ data_i[9];
		data_o[10] = (syndrome_o == 8'h8f) ^ data_i[10];
		data_o[11] = (syndrome_o == 8'h91) ^ data_i[11];
		data_o[12] = (syndrome_o == 8'h92) ^ data_i[12];
		data_o[13] = (syndrome_o == 8'h93) ^ data_i[13];
		data_o[14] = (syndrome_o == 8'h94) ^ data_i[14];
		data_o[15] = (syndrome_o == 8'h95) ^ data_i[15];
		data_o[16] = (syndrome_o == 8'h96) ^ data_i[16];
		data_o[17] = (syndrome_o == 8'h97) ^ data_i[17];
		data_o[18] = (syndrome_o == 8'h98) ^ data_i[18];
		data_o[19] = (syndrome_o == 8'h99) ^ data_i[19];
		data_o[20] = (syndrome_o == 8'h9a) ^ data_i[20];
		data_o[21] = (syndrome_o == 8'h9b) ^ data_i[21];
		data_o[22] = (syndrome_o == 8'h9c) ^ data_i[22];
		data_o[23] = (syndrome_o == 8'h9d) ^ data_i[23];
		data_o[24] = (syndrome_o == 8'h9e) ^ data_i[24];
		data_o[25] = (syndrome_o == 8'h9f) ^ data_i[25];
		data_o[26] = (syndrome_o == 8'ha1) ^ data_i[26];
		data_o[27] = (syndrome_o == 8'ha2) ^ data_i[27];
		data_o[28] = (syndrome_o == 8'ha3) ^ data_i[28];
		data_o[29] = (syndrome_o == 8'ha4) ^ data_i[29];
		data_o[30] = (syndrome_o == 8'ha5) ^ data_i[30];
		data_o[31] = (syndrome_o == 8'ha6) ^ data_i[31];
		data_o[32] = (syndrome_o == 8'ha7) ^ data_i[32];
		data_o[33] = (syndrome_o == 8'ha8) ^ data_i[33];
		data_o[34] = (syndrome_o == 8'ha9) ^ data_i[34];
		data_o[35] = (syndrome_o == 8'haa) ^ data_i[35];
		data_o[36] = (syndrome_o == 8'hab) ^ data_i[36];
		data_o[37] = (syndrome_o == 8'hac) ^ data_i[37];
		data_o[38] = (syndrome_o == 8'had) ^ data_i[38];
		data_o[39] = (syndrome_o == 8'hae) ^ data_i[39];
		data_o[40] = (syndrome_o == 8'haf) ^ data_i[40];
		data_o[41] = (syndrome_o == 8'hb0) ^ data_i[41];
		data_o[42] = (syndrome_o == 8'hb1) ^ data_i[42];
		data_o[43] = (syndrome_o == 8'hb2) ^ data_i[43];
		data_o[44] = (syndrome_o == 8'hb3) ^ data_i[44];
		data_o[45] = (syndrome_o == 8'hb4) ^ data_i[45];
		data_o[46] = (syndrome_o == 8'hb5) ^ data_i[46];
		data_o[47] = (syndrome_o == 8'hb6) ^ data_i[47];
		data_o[48] = (syndrome_o == 8'hb7) ^ data_i[48];
		data_o[49] = (syndrome_o == 8'hb8) ^ data_i[49];
		data_o[50] = (syndrome_o == 8'hb9) ^ data_i[50];
		data_o[51] = (syndrome_o == 8'hba) ^ data_i[51];
		data_o[52] = (syndrome_o == 8'hbb) ^ data_i[52];
		data_o[53] = (syndrome_o == 8'hbc) ^ data_i[53];
		data_o[54] = (syndrome_o == 8'hbd) ^ data_i[54];
		data_o[55] = (syndrome_o == 8'hbe) ^ data_i[55];
		data_o[56] = (syndrome_o == 8'hbf) ^ data_i[56];
		data_o[57] = (syndrome_o == 8'hc1) ^ data_i[57];
		data_o[58] = (syndrome_o == 8'hc2) ^ data_i[58];
		data_o[59] = (syndrome_o == 8'hc3) ^ data_i[59];
		data_o[60] = (syndrome_o == 8'hc4) ^ data_i[60];
		data_o[61] = (syndrome_o == 8'hc5) ^ data_i[61];
		data_o[62] = (syndrome_o == 8'hc6) ^ data_i[62];
		data_o[63] = (syndrome_o == 8'hc7) ^ data_i[63];
		data_o[64] = (syndrome_o == 8'hc8) ^ data_i[64];
		data_o[65] = (syndrome_o == 8'hc9) ^ data_i[65];
		data_o[66] = (syndrome_o == 8'hca) ^ data_i[66];
		data_o[67] = (syndrome_o == 8'hcb) ^ data_i[67];
		err_o[0] = syndrome_o[7];
		err_o[1] = |syndrome_o[6:0] & ~syndrome_o[7];
	end
endmodule
module prim_secded_inv_hamming_76_68_enc (
	data_i,
	data_o
);
	input [67:0] data_i;
	output reg [75:0] data_o;
	function automatic [75:0] sv2v_cast_76;
		input reg [75:0] inp;
		sv2v_cast_76 = inp;
	endfunction
	always @(*) begin : p_encode
		data_o = sv2v_cast_76(data_i);
		data_o[68] = ^(data_o & 76'h00aab55555556aaad5b);
		data_o[69] = ^(data_o & 76'h00ccd9999999b33366d);
		data_o[70] = ^(data_o & 76'h000f1e1e1e1e3c3c78e);
		data_o[71] = ^(data_o & 76'h00f01fe01fe03fc07f0);
		data_o[72] = ^(data_o & 76'h00001fffe0003fff800);
		data_o[73] = ^(data_o & 76'h00001fffffffc000000);
		data_o[74] = ^(data_o & 76'h00ffe00000000000000);
		data_o[75] = ^(data_o & 76'h7ffffffffffffffffff);
		data_o = data_o ^ 76'haa00000000000000000;
	end
endmodule
module prim_slicer (
	sel_i,
	data_i,
	data_o
);
	parameter signed [31:0] InW = 64;
	parameter signed [31:0] OutW = 8;
	parameter signed [31:0] IndexW = 4;
	input [IndexW - 1:0] sel_i;
	input [InW - 1:0] data_i;
	output wire [OutW - 1:0] data_o;
	localparam signed [31:0] UnrollW = OutW * (2 ** IndexW);
	wire [UnrollW - 1:0] unrolled_data;
	function automatic [UnrollW - 1:0] sv2v_cast_CF722;
		input reg [UnrollW - 1:0] inp;
		sv2v_cast_CF722 = inp;
	endfunction
	assign unrolled_data = sv2v_cast_CF722(data_i);
	assign data_o = unrolled_data[sel_i * OutW+:OutW];
endmodule
module prim_sparse_fsm_flop (
	clk_i,
	rst_ni,
	state_i,
	state_o
);
	parameter signed [31:0] Width = 1;
	parameter [Width - 1:0] ResetValue = 1'sb0;
	parameter [0:0] EnableAlertTriggerSVA = 1;
	input clk_i;
	input rst_ni;
	input wire [Width - 1:0] state_i;
	output wire [Width - 1:0] state_o;
	wire unused_err_o;
	wire [Width - 1:0] state_raw;
	prim_flop #(
		.Width(Width),
		.ResetValue(ResetValue)
	) u_state_flop(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(state_i),
		.q_o(state_raw)
	);
	assign state_o = state_raw;
	assign unused_err_o = 1'b0;
endmodule
module prim_sram_arbiter (
	clk_i,
	rst_ni,
	req_i,
	req_addr_i,
	req_write_i,
	req_wdata_i,
	req_wmask_i,
	gnt_o,
	rsp_rvalid_o,
	rsp_rdata_o,
	rsp_error_o,
	sram_req_o,
	sram_addr_o,
	sram_write_o,
	sram_wdata_o,
	sram_wmask_o,
	sram_rvalid_i,
	sram_rdata_i,
	sram_rerror_i
);
	parameter [31:0] N = 4;
	parameter [31:0] SramDw = 32;
	parameter [31:0] SramAw = 12;
	parameter ArbiterImpl = "PPC";
	parameter [0:0] EnMask = 1'b0;
	input clk_i;
	input rst_ni;
	input [N - 1:0] req_i;
	input [(N * SramAw) - 1:0] req_addr_i;
	input [N - 1:0] req_write_i;
	input [(N * SramDw) - 1:0] req_wdata_i;
	input [(N * SramDw) - 1:0] req_wmask_i;
	output wire [N - 1:0] gnt_o;
	output wire [N - 1:0] rsp_rvalid_o;
	output wire [(N * SramDw) - 1:0] rsp_rdata_o;
	output wire [(N * 2) - 1:0] rsp_error_o;
	output wire sram_req_o;
	output wire [SramAw - 1:0] sram_addr_o;
	output wire sram_write_o;
	output wire [SramDw - 1:0] sram_wdata_o;
	output wire [SramDw - 1:0] sram_wmask_o;
	input sram_rvalid_i;
	input [SramDw - 1:0] sram_rdata_i;
	input [1:0] sram_rerror_i;
	wire [(N * (((1 + SramAw) + SramDw) + SramDw)) - 1:0] req_packed;
	genvar i;
	generate
		for (i = 0; i < N; i = i + 1) begin : gen_reqs
			assign req_packed[((N - 1) - i) * (((1 + SramAw) + SramDw) + SramDw)+:((1 + SramAw) + SramDw) + SramDw] = {req_write_i[i], req_addr_i[((N - 1) - i) * SramAw+:SramAw], req_wdata_i[((N - 1) - i) * SramDw+:SramDw], (EnMask ? req_wmask_i[((N - 1) - i) * SramDw+:SramDw] : {SramDw {1'b1}})};
		end
	endgenerate
	localparam signed [31:0] ARB_DW = ((1 + SramAw) + SramDw) + SramDw;
	wire [(((1 + SramAw) + SramDw) + SramDw) - 1:0] sram_packed;
	assign sram_write_o = sram_packed[1 + (SramAw + (SramDw + (SramDw - 1)))];
	assign sram_addr_o = sram_packed[SramAw + (SramDw + (SramDw - 1))-:((SramAw + (SramDw + (SramDw - 1))) >= (SramDw + (SramDw + 0)) ? ((SramAw + (SramDw + (SramDw - 1))) - (SramDw + (SramDw + 0))) + 1 : ((SramDw + (SramDw + 0)) - (SramAw + (SramDw + (SramDw - 1)))) + 1)];
	assign sram_wdata_o = sram_packed[SramDw + (SramDw - 1)-:((SramDw + (SramDw - 1)) >= (SramDw + 0) ? ((SramDw + (SramDw - 1)) - (SramDw + 0)) + 1 : ((SramDw + 0) - (SramDw + (SramDw - 1))) + 1)];
	assign sram_wmask_o = (EnMask ? sram_packed[SramDw - 1-:SramDw] : {SramDw {1'b1}});
	generate
		if (EnMask == 1'b0) begin : g_unused
			reg unused_wmask;
			always @(*) begin
				unused_wmask = 1'b1;
				begin : sv2v_autoblock_1
					reg [31:0] i;
					for (i = 0; i < N; i = i + 1)
						unused_wmask = unused_wmask ^ ^req_wmask_i[((N - 1) - i) * SramDw+:SramDw];
				end
				unused_wmask = unused_wmask ^ ^sram_packed[SramDw - 1-:SramDw];
			end
		end
		if (ArbiterImpl == "PPC") begin : gen_arb_ppc
			prim_arbiter_ppc #(
				.N(N),
				.DW(ARB_DW)
			) u_reqarb(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_chk_i(1'b1),
				.req_i(req_i),
				.data_i(req_packed),
				.gnt_o(gnt_o),
				.valid_o(sram_req_o),
				.data_o(sram_packed),
				.ready_i(1'b1)
			);
		end
		else if (ArbiterImpl == "BINTREE") begin : gen_tree_arb
			prim_arbiter_tree #(
				.N(N),
				.DW(ARB_DW)
			) u_reqarb(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_chk_i(1'b1),
				.req_i(req_i),
				.data_i(req_packed),
				.gnt_o(gnt_o),
				.valid_o(sram_req_o),
				.data_o(sram_packed),
				.ready_i(1'b1)
			);
		end
	endgenerate
	wire [N - 1:0] steer;
	wire sram_ack;
	assign sram_ack = sram_rvalid_i & |steer;
	prim_fifo_sync #(
		.Width(N),
		.Pass(1'b0),
		.Depth(4)
	) u_req_fifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(1'b0),
		.wvalid_i(sram_req_o & ~sram_write_o),
		.wdata_i(gnt_o),
		.rready_i(sram_ack),
		.rdata_o(steer)
	);
	assign rsp_rvalid_o = steer & {N {sram_rvalid_i}};
	generate
		for (i = 0; i < N; i = i + 1) begin : gen_rsp
			assign rsp_rdata_o[((N - 1) - i) * SramDw+:SramDw] = sram_rdata_i;
			assign rsp_error_o[((N - 1) - i) * 2+:2] = sram_rerror_i;
		end
	endgenerate
endmodule
module prim_subreg (
	clk_i,
	rst_ni,
	we,
	wd,
	de,
	d,
	qe,
	q,
	ds,
	qs
);
	parameter signed [31:0] DW = 32;
	parameter [2:0] SwAccess = 3'd0;
	parameter [DW - 1:0] RESVAL = 1'sb0;
	input clk_i;
	input rst_ni;
	input we;
	input [DW - 1:0] wd;
	input de;
	input [DW - 1:0] d;
	output wire qe;
	output reg [DW - 1:0] q;
	output wire [DW - 1:0] ds;
	output wire [DW - 1:0] qs;
	wire wr_en;
	wire [DW - 1:0] wr_data;
	prim_subreg_arb #(
		.DW(DW),
		.SwAccess(SwAccess)
	) wr_en_data_arb(
		.we(we),
		.wd(wd),
		.de(de),
		.d(d),
		.q(q),
		.wr_en(wr_en),
		.wr_data(wr_data)
	);
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			q <= RESVAL;
		else if (wr_en)
			q <= wr_data;
	assign ds = (wr_en ? wr_data : qs);
	assign qe = wr_en;
	assign qs = q;
endmodule
module prim_subreg_ext (
	re,
	we,
	wd,
	d,
	qe,
	qre,
	q,
	ds,
	qs
);
	parameter [31:0] DW = 32;
	input re;
	input we;
	input [DW - 1:0] wd;
	input [DW - 1:0] d;
	output wire qe;
	output wire qre;
	output wire [DW - 1:0] q;
	output wire [DW - 1:0] ds;
	output wire [DW - 1:0] qs;
	assign ds = d;
	assign qs = d;
	assign q = wd;
	assign qe = we;
	assign qre = re;
endmodule
module prim_subreg_shadow (
	clk_i,
	rst_ni,
	rst_shadowed_ni,
	re,
	we,
	wd,
	de,
	d,
	qe,
	q,
	ds,
	qs,
	phase,
	err_update,
	err_storage
);
	parameter signed [31:0] DW = 32;
	parameter [2:0] SwAccess = 3'd0;
	parameter [DW - 1:0] RESVAL = 1'sb0;
	input clk_i;
	input rst_ni;
	input rst_shadowed_ni;
	input re;
	input we;
	input [DW - 1:0] wd;
	input de;
	input [DW - 1:0] d;
	output wire qe;
	output wire [DW - 1:0] q;
	output wire [DW - 1:0] ds;
	output wire [DW - 1:0] qs;
	output wire phase;
	output wire err_update;
	output wire err_storage;
	localparam [2:0] InvertedSwAccess = (SwAccess == 3'd4 ? 3'd5 : (SwAccess == 3'd5 ? 3'd4 : SwAccess));
	localparam [2:0] StagedSwAccess = (SwAccess == 3'd4 ? 3'd0 : (SwAccess == 3'd5 ? 3'd0 : SwAccess));
	wire phase_clear;
	reg phase_q;
	wire staged_we;
	wire shadow_we;
	wire committed_we;
	wire staged_de;
	wire shadow_de;
	wire committed_de;
	wire committed_qe;
	wire [DW - 1:0] staged_q;
	wire [DW - 1:0] shadow_q;
	wire [DW - 1:0] committed_q;
	wire [DW - 1:0] committed_qs;
	wire wr_en;
	wire [DW - 1:0] wr_data;
	prim_subreg_arb #(
		.DW(DW),
		.SwAccess(SwAccess)
	) wr_en_data_arb(
		.we(we),
		.wd(wd),
		.de(de),
		.d(d),
		.q(q),
		.wr_en(wr_en),
		.wr_data(wr_data)
	);
	assign phase_clear = (SwAccess == 3'd1 ? 1'b0 : re);
	always @(posedge clk_i or negedge rst_ni) begin : phase_reg
		if (!rst_ni)
			phase_q <= 1'b0;
		else if (wr_en && !err_storage)
			phase_q <= ~phase_q;
		else if (phase_clear || err_storage)
			phase_q <= 1'b0;
	end
	assign staged_we = (we & ~phase_q) & ~err_storage;
	assign staged_de = (de & ~phase_q) & ~err_storage;
	prim_subreg #(
		.DW(DW),
		.SwAccess(StagedSwAccess),
		.RESVAL(~RESVAL)
	) staged_reg(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(staged_we),
		.wd(~wr_data),
		.de(staged_de),
		.d(~d),
		.q(staged_q)
	);
	assign shadow_we = ((we & phase_q) & ~err_update) & ~err_storage;
	assign shadow_de = ((de & phase_q) & ~err_update) & ~err_storage;
	prim_subreg #(
		.DW(DW),
		.SwAccess(InvertedSwAccess),
		.RESVAL(~RESVAL)
	) shadow_reg(
		.clk_i(clk_i),
		.rst_ni(rst_shadowed_ni),
		.we(shadow_we),
		.wd(staged_q),
		.de(shadow_de),
		.d(staged_q),
		.q(shadow_q)
	);
	assign committed_we = shadow_we;
	assign committed_de = shadow_de;
	prim_subreg #(
		.DW(DW),
		.SwAccess(SwAccess),
		.RESVAL(RESVAL)
	) committed_reg(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(committed_we),
		.wd(wr_data),
		.de(committed_de),
		.d(d),
		.qe(committed_qe),
		.q(committed_q),
		.ds(ds),
		.qs(committed_qs)
	);
	assign phase = phase_q;
	assign err_update = (~staged_q != wr_data ? phase_q & wr_en : 1'b0);
	assign err_storage = ~shadow_q != committed_q;
	assign qe = committed_qe;
	assign q = committed_q;
	assign qs = committed_qs;
endmodule
module prim_subst_perm (
	data_i,
	key_i,
	data_o
);
	parameter signed [31:0] DataWidth = 64;
	parameter signed [31:0] NumRounds = 31;
	parameter [0:0] Decrypt = 0;
	input [DataWidth - 1:0] data_i;
	input [DataWidth - 1:0] key_i;
	output wire [DataWidth - 1:0] data_o;
	reg [(NumRounds >= 0 ? ((NumRounds + 1) * DataWidth) - 1 : ((1 - NumRounds) * DataWidth) + ((NumRounds * DataWidth) - 1)):(NumRounds >= 0 ? 0 : NumRounds * DataWidth)] data_state;
	wire [DataWidth * 1:1] sv2v_tmp_428CF;
	assign sv2v_tmp_428CF = data_i;
	always @(*) data_state[(NumRounds >= 0 ? 0 : NumRounds) * DataWidth+:DataWidth] = sv2v_tmp_428CF;
	genvar r;
	localparam [63:0] prim_cipher_pkg_PRESENT_SBOX4 = 64'h21748fe3da09b65c;
	localparam [63:0] prim_cipher_pkg_PRESENT_SBOX4_INV = 64'ha970364bd21c8fe5;
	generate
		for (r = 0; r < NumRounds; r = r + 1) begin : gen_round
			reg [DataWidth - 1:0] data_state_sbox;
			reg [DataWidth - 1:0] data_state_flipped;
			if (Decrypt) begin : gen_dec
				always @(*) begin : p_dec
					data_state_sbox = data_state[(NumRounds >= 0 ? r : NumRounds - r) * DataWidth+:DataWidth] ^ key_i;
					data_state_flipped = data_state_sbox;
					begin : sv2v_autoblock_1
						reg signed [31:0] k;
						for (k = 0; k < (DataWidth / 2); k = k + 1)
							begin
								data_state_flipped[k * 2] = data_state_sbox[k];
								data_state_flipped[(k * 2) + 1] = data_state_sbox[k + (DataWidth / 2)];
							end
					end
					begin : sv2v_autoblock_2
						reg signed [31:0] k;
						for (k = 0; k < DataWidth; k = k + 1)
							data_state_sbox[(DataWidth - 1) - k] = data_state_flipped[k];
					end
					begin : sv2v_autoblock_3
						reg signed [31:0] k;
						for (k = 0; k < (DataWidth / 4); k = k + 1)
							data_state_sbox[k * 4+:4] = prim_cipher_pkg_PRESENT_SBOX4_INV[data_state_sbox[k * 4+:4] * 4+:4];
					end
					data_state[(NumRounds >= 0 ? r + 1 : NumRounds - (r + 1)) * DataWidth+:DataWidth] = data_state_sbox;
				end
			end
			else begin : gen_enc
				always @(*) begin : p_enc
					data_state_sbox = data_state[(NumRounds >= 0 ? r : NumRounds - r) * DataWidth+:DataWidth] ^ key_i;
					begin : sv2v_autoblock_4
						reg signed [31:0] k;
						for (k = 0; k < (DataWidth / 4); k = k + 1)
							data_state_sbox[k * 4+:4] = prim_cipher_pkg_PRESENT_SBOX4[data_state_sbox[k * 4+:4] * 4+:4];
					end
					begin : sv2v_autoblock_5
						reg signed [31:0] k;
						for (k = 0; k < DataWidth; k = k + 1)
							data_state_flipped[(DataWidth - 1) - k] = data_state_sbox[k];
					end
					data_state_sbox = data_state_flipped;
					begin : sv2v_autoblock_6
						reg signed [31:0] k;
						for (k = 0; k < (DataWidth / 2); k = k + 1)
							begin
								data_state_sbox[k] = data_state_flipped[k * 2];
								data_state_sbox[k + (DataWidth / 2)] = data_state_flipped[(k * 2) + 1];
							end
					end
					data_state[(NumRounds >= 0 ? r + 1 : NumRounds - (r + 1)) * DataWidth+:DataWidth] = data_state_sbox;
				end
			end
		end
	endgenerate
	assign data_o = data_state[(NumRounds >= 0 ? NumRounds : NumRounds - NumRounds) * DataWidth+:DataWidth] ^ key_i;
endmodule
module prim_sync_reqack (
	clk_src_i,
	rst_src_ni,
	clk_dst_i,
	rst_dst_ni,
	req_chk_i,
	src_req_i,
	src_ack_o,
	dst_req_o,
	dst_ack_i
);
	parameter [0:0] EnRstChks = 1'b0;
	parameter [0:0] EnRzHs = 1'b0;
	input clk_src_i;
	input rst_src_ni;
	input clk_dst_i;
	input rst_dst_ni;
	input wire req_chk_i;
	input wire src_req_i;
	output reg src_ack_o;
	output reg dst_req_o;
	input wire dst_ack_i;
	wire unused_req_chk;
	assign unused_req_chk = req_chk_i;
	generate
		if (EnRzHs) begin : gen_rz_hs_protocol
			reg src_fsm_d;
			reg src_fsm_q;
			reg dst_fsm_d;
			reg dst_fsm_q;
			wire src_ack;
			reg dst_ack;
			reg src_req;
			wire dst_req;
			always @(*) begin : src_fsm
				src_fsm_d = src_fsm_q;
				src_ack_o = 1'b0;
				src_req = 1'b0;
				case (src_fsm_q)
					1'd0:
						if (!src_ack && src_req_i)
							src_fsm_d = 1'd1;
					1'd1: begin
						src_req = 1'b1;
						src_ack_o = src_ack;
						if (!src_req_i || src_ack)
							src_fsm_d = 1'd0;
					end
					default:
						;
				endcase
			end
			prim_flop_2sync #(.Width(1)) ack_sync(
				.clk_i(clk_src_i),
				.rst_ni(rst_src_ni),
				.d_i(dst_ack),
				.q_o(src_ack)
			);
			always @(posedge clk_src_i or negedge rst_src_ni)
				if (!rst_src_ni)
					src_fsm_q <= 1'd0;
				else
					src_fsm_q <= src_fsm_d;
			always @(*) begin : dst_fsm
				dst_fsm_d = dst_fsm_q;
				dst_req_o = 1'b0;
				dst_ack = 1'b0;
				case (dst_fsm_q)
					1'd0:
						if (dst_req) begin
							dst_req_o = 1'b1;
							if (dst_ack_i)
								dst_fsm_d = 1'd1;
						end
					1'd1: begin
						dst_ack = 1'b1;
						if (!dst_req)
							dst_fsm_d = 1'd0;
					end
					default:
						;
				endcase
			end
			prim_flop_2sync #(.Width(1)) req_sync(
				.clk_i(clk_dst_i),
				.rst_ni(rst_dst_ni),
				.d_i(src_req),
				.q_o(dst_req)
			);
			always @(posedge clk_dst_i or negedge rst_dst_ni)
				if (!rst_dst_ni)
					dst_fsm_q <= 1'd0;
				else
					dst_fsm_q <= dst_fsm_d;
		end
		else begin : gen_nrz_hs_protocol
			reg src_fsm_ns;
			reg src_fsm_cs;
			reg dst_fsm_ns;
			reg dst_fsm_cs;
			reg src_req_d;
			reg src_req_q;
			wire src_ack;
			reg dst_ack_d;
			reg dst_ack_q;
			wire dst_req;
			wire src_handshake;
			wire dst_handshake;
			assign src_handshake = src_req_i & src_ack_o;
			assign dst_handshake = dst_req_o & dst_ack_i;
			prim_flop_2sync #(.Width(1)) req_sync(
				.clk_i(clk_dst_i),
				.rst_ni(rst_dst_ni),
				.d_i(src_req_q),
				.q_o(dst_req)
			);
			prim_flop_2sync #(.Width(1)) ack_sync(
				.clk_i(clk_src_i),
				.rst_ni(rst_src_ni),
				.d_i(dst_ack_q),
				.q_o(src_ack)
			);
			always @(*) begin : src_fsm
				src_fsm_ns = src_fsm_cs;
				src_req_d = src_req_q;
				src_ack_o = 1'b0;
				case (src_fsm_cs)
					1'd0: begin
						src_req_d = src_req_i;
						src_ack_o = src_ack;
						if (src_handshake)
							src_fsm_ns = 1'd1;
					end
					1'd1: begin
						src_req_d = ~src_req_i;
						src_ack_o = ~src_ack;
						if (src_handshake)
							src_fsm_ns = 1'd0;
					end
					default:
						;
				endcase
			end
			always @(*) begin : dst_fsm
				dst_fsm_ns = dst_fsm_cs;
				dst_req_o = 1'b0;
				dst_ack_d = dst_ack_q;
				case (dst_fsm_cs)
					1'd0: begin
						dst_req_o = dst_req;
						dst_ack_d = dst_ack_i;
						if (dst_handshake)
							dst_fsm_ns = 1'd1;
					end
					1'd1: begin
						dst_req_o = ~dst_req;
						dst_ack_d = ~dst_ack_i;
						if (dst_handshake)
							dst_fsm_ns = 1'd0;
					end
					default:
						;
				endcase
			end
			always @(posedge clk_src_i or negedge rst_src_ni)
				if (!rst_src_ni) begin
					src_fsm_cs <= 1'd0;
					src_req_q <= 1'b0;
				end
				else begin
					src_fsm_cs <= src_fsm_ns;
					src_req_q <= src_req_d;
				end
			always @(posedge clk_dst_i or negedge rst_dst_ni)
				if (!rst_dst_ni) begin
					dst_fsm_cs <= 1'd0;
					dst_ack_q <= 1'b0;
				end
				else begin
					dst_fsm_cs <= dst_fsm_ns;
					dst_ack_q <= dst_ack_d;
				end
		end
	endgenerate
endmodule
module prim_sync_reqack_data (
	clk_src_i,
	rst_src_ni,
	clk_dst_i,
	rst_dst_ni,
	req_chk_i,
	src_req_i,
	src_ack_o,
	dst_req_o,
	dst_ack_i,
	data_i,
	data_o
);
	parameter [31:0] Width = 1;
	parameter [0:0] EnRstChks = 1'b0;
	parameter [0:0] DataSrc2Dst = 1'b1;
	parameter [0:0] DataReg = 1'b0;
	parameter [0:0] EnRzHs = 1'b0;
	input clk_src_i;
	input rst_src_ni;
	input clk_dst_i;
	input rst_dst_ni;
	input wire req_chk_i;
	input wire src_req_i;
	output wire src_ack_o;
	output wire dst_req_o;
	input wire dst_ack_i;
	input wire [Width - 1:0] data_i;
	output wire [Width - 1:0] data_o;
	prim_sync_reqack #(
		.EnRstChks(EnRstChks),
		.EnRzHs(EnRzHs)
	) u_prim_sync_reqack(
		.clk_src_i(clk_src_i),
		.rst_src_ni(rst_src_ni),
		.clk_dst_i(clk_dst_i),
		.rst_dst_ni(rst_dst_ni),
		.req_chk_i(req_chk_i),
		.src_req_i(src_req_i),
		.src_ack_o(src_ack_o),
		.dst_req_o(dst_req_o),
		.dst_ack_i(dst_ack_i)
	);
	generate
		if ((DataSrc2Dst == 1'b0) && (DataReg == 1'b1)) begin : gen_data_reg
			wire data_we;
			wire [Width - 1:0] data_d;
			reg [Width - 1:0] data_q;
			assign data_we = dst_req_o & dst_ack_i;
			assign data_d = data_i;
			always @(posedge clk_dst_i or negedge rst_dst_ni)
				if (!rst_dst_ni)
					data_q <= 1'sb0;
				else if (data_we)
					data_q <= data_d;
			assign data_o = data_q;
		end
		else begin : gen_no_data_reg
			assign data_o = data_i;
		end
	endgenerate
endmodule
module prim_sync_slow_fast (
	clk_slow_i,
	clk_fast_i,
	rst_fast_ni,
	wdata_i,
	rdata_o
);
	parameter [31:0] Width = 32;
	input wire clk_slow_i;
	input wire clk_fast_i;
	input wire rst_fast_ni;
	input wire [Width - 1:0] wdata_i;
	output wire [Width - 1:0] rdata_o;
	wire sync_clk_slow;
	reg sync_clk_slow_q;
	wire wdata_en;
	reg [Width - 1:0] wdata_q;
	prim_flop_2sync #(.Width(1)) sync_slow_clk(
		.clk_i(clk_fast_i),
		.rst_ni(rst_fast_ni),
		.d_i(clk_slow_i),
		.q_o(sync_clk_slow)
	);
	always @(posedge clk_fast_i or negedge rst_fast_ni)
		if (!rst_fast_ni)
			sync_clk_slow_q <= 1'b0;
		else
			sync_clk_slow_q <= sync_clk_slow;
	assign wdata_en = sync_clk_slow_q & !sync_clk_slow;
	always @(posedge clk_fast_i or negedge rst_fast_ni)
		if (!rst_fast_ni)
			wdata_q <= 1'sb0;
		else if (wdata_en)
			wdata_q <= wdata_i;
	assign rdata_o = wdata_q;
endmodule
(* DONT_TOUCH = "yes" *) module prim_xilinx_and2 (
	in0_i,
	in1_i,
	out_o
);
	parameter signed [31:0] Width = 1;
	input [Width - 1:0] in0_i;
	input [Width - 1:0] in1_i;
	output wire [Width - 1:0] out_o;
	assign out_o = in0_i & in1_i;
endmodule
(* DONT_TOUCH = "yes" *) module prim_xilinx_buf (
	in_i,
	out_o
);
	parameter signed [31:0] Width = 1;
	input [Width - 1:0] in_i;
	output wire [Width - 1:0] out_o;
	assign out_o = in_i;
endmodule
module prim_xilinx_clock_gating (
	clk_i,
	en_i,
	test_en_i,
	clk_o
);
	parameter [0:0] NoFpgaGate = 1'b0;
	parameter [0:0] FpgaBufGlobal = 1'b1;
	input clk_i;
	input en_i;
	input test_en_i;
	output wire clk_o;
	generate
		if (NoFpgaGate) begin : gen_no_gate
			assign clk_o = clk_i;
		end
		else begin : gen_gate
			if (FpgaBufGlobal) begin : gen_bufgce
				BUFGCE #(.SIM_DEVICE("7SERIES")) u_bufgce(
					.I(clk_i),
					.CE(en_i | test_en_i),
					.O(clk_o)
				);
			end
			else begin : gen_bufhce
				BUFHCE u_bufhce(
					.I(clk_i),
					.CE(en_i | test_en_i),
					.O(clk_o)
				);
			end
		end
	endgenerate
endmodule
module prim_xilinx_clock_mux2 (
	clk0_i,
	clk1_i,
	sel_i,
	clk_o
);
	parameter [0:0] NoFpgaBufG = 1'b0;
	input clk0_i;
	input clk1_i;
	input sel_i;
	output wire clk_o;
	generate
		if (NoFpgaBufG) begin : gen_no_bufg
			assign clk_o = (sel_i ? clk1_i : clk0_i);
		end
		else begin : gen_bufg
			BUFGMUX bufgmux_i(
				.S(sel_i),
				.I0(clk0_i),
				.I1(clk1_i),
				.O(clk_o)
			);
		end
	endgenerate
endmodule
(* DONT_TOUCH = "yes" *) module prim_xilinx_flop (
	clk_i,
	rst_ni,
	d_i,
	q_o
);
	parameter signed [31:0] Width = 1;
	parameter [Width - 1:0] ResetValue = 0;
	input clk_i;
	input rst_ni;
	input [Width - 1:0] d_i;
	output reg [Width - 1:0] q_o;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			q_o <= ResetValue;
		else
			q_o <= d_i;
endmodule
(* DONT_TOUCH = "yes" *) module prim_xilinx_flop_en (
	clk_i,
	rst_ni,
	en_i,
	d_i,
	q_o
);
	parameter signed [31:0] Width = 1;
	parameter [0:0] EnSecBuf = 0;
	parameter [Width - 1:0] ResetValue = 0;
	input clk_i;
	input rst_ni;
	input en_i;
	input [Width - 1:0] d_i;
	output reg [Width - 1:0] q_o;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			q_o <= ResetValue;
		else if (en_i)
			q_o <= d_i;
endmodule
(* DONT_TOUCH = "yes" *) module prim_xilinx_xor2 (
	in0_i,
	in1_i,
	out_o
);
	parameter signed [31:0] Width = 1;
	input [Width - 1:0] in0_i;
	input [Width - 1:0] in1_i;
	output wire [Width - 1:0] out_o;
	assign out_o = in0_i ^ in1_i;
endmodule
module prim_xnor2 (
	in0_i,
	in1_i,
	out_o
);
	parameter signed [31:0] Width = 1;
	input [Width - 1:0] in0_i;
	input [Width - 1:0] in1_i;
	output wire [Width - 1:0] out_o;
	generate
		if (1) begin : gen_generic
			prim_generic_xnor2 #(.Width(Width)) u_impl_generic(
				.in0_i(in0_i),
				.in1_i(in1_i),
				.out_o(out_o)
			);
		end
	endgenerate
endmodule
module prim_xor2 (
	in0_i,
	in1_i,
	out_o
);
	parameter signed [31:0] Width = 1;
	input [Width - 1:0] in0_i;
	input [Width - 1:0] in1_i;
	output wire [Width - 1:0] out_o;
	parameter integer Impl = 32'sd0;
	generate
		if (Impl == 32'sd2) begin : gen_xilinx
			prim_xilinx_xor2 #(.Width(Width)) u_impl_xilinx(
				.in0_i(in0_i),
				.in1_i(in1_i),
				.out_o(out_o)
			);
		end
		else begin : gen_generic
			prim_generic_xor2 #(.Width(Width)) u_impl_generic(
				.in0_i(in0_i),
				.in1_i(in1_i),
				.out_o(out_o)
			);
		end
	endgenerate
endmodule
module pwrmgr_reg_top (
	clk_i,
	rst_ni,
	clk_lc_i,
	rst_lc_ni,
	tl_i,
	tl_o,
	reg2hw,
	hw2reg,
	intg_err_o,
	devmode_i
);
	input clk_i;
	input rst_ni;
	input clk_lc_i;
	input rst_lc_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_i;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	output wire [36:0] reg2hw;
	input wire [38:0] hw2reg;
	output wire intg_err_o;
	input devmode_i;
	localparam signed [31:0] AW = 7;
	localparam signed [31:0] DW = 32;
	localparam signed [31:0] DBW = 4;
	wire reg_we;
	wire reg_re;
	wire [6:0] reg_addr;
	wire [31:0] reg_wdata;
	wire [3:0] reg_be;
	wire [31:0] reg_rdata;
	wire reg_error;
	wire addrmiss;
	reg wr_err;
	reg [31:0] reg_rdata_next;
	wire reg_busy;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_reg_h2d;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_reg_d2h;
	wire intg_err;
	tlul_cmd_intg_chk u_chk(
		.tl_i(tl_i),
		.err_o(intg_err)
	);
	wire reg_we_err;
	reg [16:0] reg_we_check;
	prim_reg_we_check #(.OneHotWidth(17)) u_prim_reg_we_check(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.oh_i(reg_we_check),
		.en_i(reg_we && !addrmiss),
		.err_o(reg_we_err)
	);
	reg err_q;
	always @(posedge clk_lc_i or negedge rst_lc_ni)
		if (!rst_lc_ni)
			err_q <= 1'sb0;
		else if (intg_err || reg_we_err)
			err_q <= 1'b1;
	assign intg_err_o = (err_q | intg_err) | reg_we_err;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o_pre;
	tlul_rsp_intg_gen #(
		.EnableRspIntgGen(1),
		.EnableDataIntgGen(1)
	) u_rsp_intg_gen(
		.tl_i(tl_o_pre),
		.tl_o(tl_o)
	);
	assign tl_reg_h2d = tl_i;
	assign tl_o_pre = tl_reg_d2h;
	function automatic [3:0] sv2v_cast_2253A;
		input reg [3:0] inp;
		sv2v_cast_2253A = inp;
	endfunction
	tlul_adapter_reg #(
		.RegAw(AW),
		.RegDw(DW),
		.EnableDataIntgGen(0)
	) u_reg_if(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_reg_h2d),
		.tl_o(tl_reg_d2h),
		.en_ifetch_i(sv2v_cast_2253A(4'h9)),
		.we_o(reg_we),
		.re_o(reg_re),
		.addr_o(reg_addr),
		.wdata_o(reg_wdata),
		.be_o(reg_be),
		.busy_i(reg_busy),
		.rdata_i(reg_rdata),
		.error_i(reg_error)
	);
	assign reg_rdata = reg_rdata_next;
	assign reg_error = ((devmode_i & addrmiss) | wr_err) | intg_err;
	wire intr_state_we;
	wire intr_state_qs;
	wire intr_state_wd;
	wire intr_enable_we;
	wire intr_enable_qs;
	wire intr_enable_wd;
	wire intr_test_we;
	wire intr_test_wd;
	wire alert_test_we;
	wire alert_test_wd;
	wire ctrl_cfg_regwen_re;
	wire ctrl_cfg_regwen_qs;
	wire control_we;
	wire control_low_power_hint_qs;
	wire control_low_power_hint_wd;
	wire control_core_clk_en_qs;
	wire control_core_clk_en_wd;
	wire control_io_clk_en_qs;
	wire control_io_clk_en_wd;
	wire control_usb_clk_en_lp_qs;
	wire control_usb_clk_en_lp_wd;
	wire control_usb_clk_en_active_qs;
	wire control_usb_clk_en_active_wd;
	wire control_main_pd_n_qs;
	wire control_main_pd_n_wd;
	wire cfg_cdc_sync_we;
	wire cfg_cdc_sync_qs;
	wire cfg_cdc_sync_wd;
	wire wakeup_en_regwen_we;
	wire wakeup_en_regwen_qs;
	wire wakeup_en_regwen_wd;
	wire wakeup_en_we;
	wire wakeup_en_en_0_qs;
	wire wakeup_en_en_0_wd;
	wire wakeup_en_en_1_qs;
	wire wakeup_en_en_1_wd;
	wire wakeup_en_en_2_qs;
	wire wakeup_en_en_2_wd;
	wire wakeup_en_en_3_qs;
	wire wakeup_en_en_3_wd;
	wire wakeup_en_en_4_qs;
	wire wakeup_en_en_4_wd;
	wire wakeup_en_en_5_qs;
	wire wakeup_en_en_5_wd;
	wire wake_status_val_0_qs;
	wire wake_status_val_1_qs;
	wire wake_status_val_2_qs;
	wire wake_status_val_3_qs;
	wire wake_status_val_4_qs;
	wire wake_status_val_5_qs;
	wire reset_en_regwen_we;
	wire reset_en_regwen_qs;
	wire reset_en_regwen_wd;
	wire reset_en_we;
	wire reset_en_en_0_qs;
	wire reset_en_en_0_wd;
	wire reset_en_en_1_qs;
	wire reset_en_en_1_wd;
	wire reset_status_val_0_qs;
	wire reset_status_val_1_qs;
	wire escalate_reset_status_qs;
	wire wake_info_capture_dis_we;
	wire wake_info_capture_dis_qs;
	wire wake_info_capture_dis_wd;
	wire wake_info_re;
	wire wake_info_we;
	wire [5:0] wake_info_reasons_qs;
	wire [5:0] wake_info_reasons_wd;
	wire wake_info_fall_through_qs;
	wire wake_info_fall_through_wd;
	wire wake_info_abort_qs;
	wire wake_info_abort_wd;
	wire fault_status_reg_intg_err_qs;
	wire fault_status_esc_timeout_qs;
	wire fault_status_main_pd_glitch_qs;
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_intr_state(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_state_we),
		.wd(intr_state_wd),
		.de(hw2reg[37]),
		.d(hw2reg[38]),
		.q(reg2hw[36]),
		.qs(intr_state_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_intr_enable(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(intr_enable_we),
		.wd(intr_enable_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[35]),
		.qs(intr_enable_qs)
	);
	wire intr_test_qe;
	wire [0:0] intr_test_flds_we;
	assign intr_test_qe = &intr_test_flds_we;
	prim_subreg_ext #(.DW(1)) u_intr_test(
		.re(1'b0),
		.we(intr_test_we),
		.wd(intr_test_wd),
		.d(1'sb0),
		.qe(intr_test_flds_we[0]),
		.q(reg2hw[34])
	);
	assign reg2hw[33] = intr_test_qe;
	wire alert_test_qe;
	wire [0:0] alert_test_flds_we;
	assign alert_test_qe = &alert_test_flds_we;
	prim_subreg_ext #(.DW(1)) u_alert_test(
		.re(1'b0),
		.we(alert_test_we),
		.wd(alert_test_wd),
		.d(1'sb0),
		.qe(alert_test_flds_we[0]),
		.q(reg2hw[32])
	);
	assign reg2hw[31] = alert_test_qe;
	prim_subreg_ext #(.DW(1)) u_ctrl_cfg_regwen(
		.re(ctrl_cfg_regwen_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[36]),
		.qs(ctrl_cfg_regwen_qs)
	);
	wire control_gated_we;
	assign control_gated_we = control_we & ctrl_cfg_regwen_qs;
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_control_low_power_hint(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(control_gated_we),
		.wd(control_low_power_hint_wd),
		.de(hw2reg[34]),
		.d(hw2reg[35]),
		.q(reg2hw[30]),
		.qs(control_low_power_hint_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_control_core_clk_en(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(control_gated_we),
		.wd(control_core_clk_en_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[29]),
		.qs(control_core_clk_en_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_control_io_clk_en(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(control_gated_we),
		.wd(control_io_clk_en_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[28]),
		.qs(control_io_clk_en_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_control_usb_clk_en_lp(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(control_gated_we),
		.wd(control_usb_clk_en_lp_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[27]),
		.qs(control_usb_clk_en_lp_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_control_usb_clk_en_active(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(control_gated_we),
		.wd(control_usb_clk_en_active_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[26]),
		.qs(control_usb_clk_en_active_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h1)
	) u_control_main_pd_n(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(control_gated_we),
		.wd(control_main_pd_n_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[25]),
		.qs(control_main_pd_n_qs)
	);
	wire cfg_cdc_sync_qe;
	wire [0:0] cfg_cdc_sync_flds_we;
	prim_flop #(
		.Width(1),
		.ResetValue(0)
	) u_cfg_cdc_sync0_qe(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i(&cfg_cdc_sync_flds_we),
		.q_o(cfg_cdc_sync_qe)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_cfg_cdc_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(cfg_cdc_sync_we),
		.wd(cfg_cdc_sync_wd),
		.de(hw2reg[32]),
		.d(hw2reg[33]),
		.qe(cfg_cdc_sync_flds_we[0]),
		.q(reg2hw[24]),
		.qs(cfg_cdc_sync_qs)
	);
	assign reg2hw[23] = cfg_cdc_sync_qe;
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_wakeup_en_regwen(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(wakeup_en_regwen_we),
		.wd(wakeup_en_regwen_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(wakeup_en_regwen_qs)
	);
	wire wakeup_en_gated_we;
	assign wakeup_en_gated_we = wakeup_en_we & wakeup_en_regwen_qs;
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_wakeup_en_en_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(wakeup_en_gated_we),
		.wd(wakeup_en_en_0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[17]),
		.qs(wakeup_en_en_0_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_wakeup_en_en_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(wakeup_en_gated_we),
		.wd(wakeup_en_en_1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[18]),
		.qs(wakeup_en_en_1_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_wakeup_en_en_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(wakeup_en_gated_we),
		.wd(wakeup_en_en_2_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[19]),
		.qs(wakeup_en_en_2_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_wakeup_en_en_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(wakeup_en_gated_we),
		.wd(wakeup_en_en_3_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[20]),
		.qs(wakeup_en_en_3_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_wakeup_en_en_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(wakeup_en_gated_we),
		.wd(wakeup_en_en_4_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[21]),
		.qs(wakeup_en_en_4_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_wakeup_en_en_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(wakeup_en_gated_we),
		.wd(wakeup_en_en_5_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[22]),
		.qs(wakeup_en_en_5_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd1),
		.RESVAL(1'h0)
	) u_wake_status_val_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(1'sb0),
		.de(hw2reg[20]),
		.d(hw2reg[21]),
		.qs(wake_status_val_0_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd1),
		.RESVAL(1'h0)
	) u_wake_status_val_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(1'sb0),
		.de(hw2reg[22]),
		.d(hw2reg[23]),
		.qs(wake_status_val_1_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd1),
		.RESVAL(1'h0)
	) u_wake_status_val_2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(1'sb0),
		.de(hw2reg[24]),
		.d(hw2reg[25]),
		.qs(wake_status_val_2_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd1),
		.RESVAL(1'h0)
	) u_wake_status_val_3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(1'sb0),
		.de(hw2reg[26]),
		.d(hw2reg[27]),
		.qs(wake_status_val_3_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd1),
		.RESVAL(1'h0)
	) u_wake_status_val_4(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(1'sb0),
		.de(hw2reg[28]),
		.d(hw2reg[29]),
		.qs(wake_status_val_4_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd1),
		.RESVAL(1'h0)
	) u_wake_status_val_5(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(1'sb0),
		.de(hw2reg[30]),
		.d(hw2reg[31]),
		.qs(wake_status_val_5_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_reset_en_regwen(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(reset_en_regwen_we),
		.wd(reset_en_regwen_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(reset_en_regwen_qs)
	);
	wire reset_en_gated_we;
	assign reset_en_gated_we = reset_en_we & reset_en_regwen_qs;
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_reset_en_en_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(reset_en_gated_we),
		.wd(reset_en_en_0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[15]),
		.qs(reset_en_en_0_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_reset_en_en_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(reset_en_gated_we),
		.wd(reset_en_en_1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[16]),
		.qs(reset_en_en_1_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd1),
		.RESVAL(1'h0)
	) u_reset_status_val_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(1'sb0),
		.de(hw2reg[16]),
		.d(hw2reg[17]),
		.qs(reset_status_val_0_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd1),
		.RESVAL(1'h0)
	) u_reset_status_val_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(1'sb0),
		.de(hw2reg[18]),
		.d(hw2reg[19]),
		.qs(reset_status_val_1_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd1),
		.RESVAL(1'h0)
	) u_escalate_reset_status(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(1'b0),
		.wd(1'sb0),
		.de(hw2reg[14]),
		.d(hw2reg[15]),
		.qs(escalate_reset_status_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_wake_info_capture_dis(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(wake_info_capture_dis_we),
		.wd(wake_info_capture_dis_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[14]),
		.qs(wake_info_capture_dis_qs)
	);
	wire wake_info_qe;
	wire [2:0] wake_info_flds_we;
	assign wake_info_qe = &wake_info_flds_we;
	prim_subreg_ext #(.DW(6)) u_wake_info_reasons(
		.re(wake_info_re),
		.we(wake_info_we),
		.wd(wake_info_reasons_wd),
		.d(hw2reg[13-:6]),
		.qe(wake_info_flds_we[0]),
		.q(reg2hw[13-:6]),
		.qs(wake_info_reasons_qs)
	);
	assign reg2hw[7] = wake_info_qe;
	prim_subreg_ext #(.DW(1)) u_wake_info_fall_through(
		.re(wake_info_re),
		.we(wake_info_we),
		.wd(wake_info_fall_through_wd),
		.d(hw2reg[7]),
		.qe(wake_info_flds_we[1]),
		.q(reg2hw[6]),
		.qs(wake_info_fall_through_qs)
	);
	assign reg2hw[5] = wake_info_qe;
	prim_subreg_ext #(.DW(1)) u_wake_info_abort(
		.re(wake_info_re),
		.we(wake_info_we),
		.wd(wake_info_abort_wd),
		.d(hw2reg[6]),
		.qe(wake_info_flds_we[2]),
		.q(reg2hw[4]),
		.qs(wake_info_abort_qs)
	);
	assign reg2hw[3] = wake_info_qe;
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd1),
		.RESVAL(1'h0)
	) u_fault_status_reg_intg_err(
		.clk_i(clk_lc_i),
		.rst_ni(rst_lc_ni),
		.we(1'b0),
		.wd(1'sb0),
		.de(hw2reg[4]),
		.d(hw2reg[5]),
		.q(reg2hw[2]),
		.qs(fault_status_reg_intg_err_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd1),
		.RESVAL(1'h0)
	) u_fault_status_esc_timeout(
		.clk_i(clk_lc_i),
		.rst_ni(rst_lc_ni),
		.we(1'b0),
		.wd(1'sb0),
		.de(hw2reg[2]),
		.d(hw2reg[3]),
		.q(reg2hw[1]),
		.qs(fault_status_esc_timeout_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd1),
		.RESVAL(1'h0)
	) u_fault_status_main_pd_glitch(
		.clk_i(clk_lc_i),
		.rst_ni(rst_lc_ni),
		.we(1'b0),
		.wd(1'sb0),
		.de(hw2reg[0]),
		.d(hw2reg[1]),
		.q(reg2hw[0]),
		.qs(fault_status_main_pd_glitch_qs)
	);
	reg [16:0] addr_hit;
	localparam signed [31:0] pwrmgr_reg_pkg_BlockAw = 7;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_ALERT_TEST_OFFSET = 7'h0c;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_CFG_CDC_SYNC_OFFSET = 7'h18;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_CONTROL_OFFSET = 7'h14;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_CTRL_CFG_REGWEN_OFFSET = 7'h10;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_ESCALATE_RESET_STATUS_OFFSET = 7'h34;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_FAULT_STATUS_OFFSET = 7'h40;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_INTR_ENABLE_OFFSET = 7'h04;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_INTR_STATE_OFFSET = 7'h00;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_INTR_TEST_OFFSET = 7'h08;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_RESET_EN_OFFSET = 7'h2c;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_RESET_EN_REGWEN_OFFSET = 7'h28;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_RESET_STATUS_OFFSET = 7'h30;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_WAKEUP_EN_OFFSET = 7'h20;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_WAKEUP_EN_REGWEN_OFFSET = 7'h1c;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_WAKE_INFO_CAPTURE_DIS_OFFSET = 7'h38;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_WAKE_INFO_OFFSET = 7'h3c;
	localparam [6:0] pwrmgr_reg_pkg_PWRMGR_WAKE_STATUS_OFFSET = 7'h24;
	always @(*) begin
		addr_hit = 1'sb0;
		addr_hit[0] = reg_addr == pwrmgr_reg_pkg_PWRMGR_INTR_STATE_OFFSET;
		addr_hit[1] = reg_addr == pwrmgr_reg_pkg_PWRMGR_INTR_ENABLE_OFFSET;
		addr_hit[2] = reg_addr == pwrmgr_reg_pkg_PWRMGR_INTR_TEST_OFFSET;
		addr_hit[3] = reg_addr == pwrmgr_reg_pkg_PWRMGR_ALERT_TEST_OFFSET;
		addr_hit[4] = reg_addr == pwrmgr_reg_pkg_PWRMGR_CTRL_CFG_REGWEN_OFFSET;
		addr_hit[5] = reg_addr == pwrmgr_reg_pkg_PWRMGR_CONTROL_OFFSET;
		addr_hit[6] = reg_addr == pwrmgr_reg_pkg_PWRMGR_CFG_CDC_SYNC_OFFSET;
		addr_hit[7] = reg_addr == pwrmgr_reg_pkg_PWRMGR_WAKEUP_EN_REGWEN_OFFSET;
		addr_hit[8] = reg_addr == pwrmgr_reg_pkg_PWRMGR_WAKEUP_EN_OFFSET;
		addr_hit[9] = reg_addr == pwrmgr_reg_pkg_PWRMGR_WAKE_STATUS_OFFSET;
		addr_hit[10] = reg_addr == pwrmgr_reg_pkg_PWRMGR_RESET_EN_REGWEN_OFFSET;
		addr_hit[11] = reg_addr == pwrmgr_reg_pkg_PWRMGR_RESET_EN_OFFSET;
		addr_hit[12] = reg_addr == pwrmgr_reg_pkg_PWRMGR_RESET_STATUS_OFFSET;
		addr_hit[13] = reg_addr == pwrmgr_reg_pkg_PWRMGR_ESCALATE_RESET_STATUS_OFFSET;
		addr_hit[14] = reg_addr == pwrmgr_reg_pkg_PWRMGR_WAKE_INFO_CAPTURE_DIS_OFFSET;
		addr_hit[15] = reg_addr == pwrmgr_reg_pkg_PWRMGR_WAKE_INFO_OFFSET;
		addr_hit[16] = reg_addr == pwrmgr_reg_pkg_PWRMGR_FAULT_STATUS_OFFSET;
	end
	assign addrmiss = (reg_re || reg_we ? ~|addr_hit : 1'b0);
	localparam [67:0] pwrmgr_reg_pkg_PWRMGR_PERMIT = 68'b00010001000100010001001100010001000100010001000100010001000100010001;
	always @(*) wr_err = reg_we & (((((((((((((((((addr_hit[0] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[64+:4] & ~reg_be)) | (addr_hit[1] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[60+:4] & ~reg_be))) | (addr_hit[2] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[56+:4] & ~reg_be))) | (addr_hit[3] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[52+:4] & ~reg_be))) | (addr_hit[4] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[48+:4] & ~reg_be))) | (addr_hit[5] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[44+:4] & ~reg_be))) | (addr_hit[6] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[40+:4] & ~reg_be))) | (addr_hit[7] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[36+:4] & ~reg_be))) | (addr_hit[8] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[32+:4] & ~reg_be))) | (addr_hit[9] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[28+:4] & ~reg_be))) | (addr_hit[10] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[24+:4] & ~reg_be))) | (addr_hit[11] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[20+:4] & ~reg_be))) | (addr_hit[12] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[16+:4] & ~reg_be))) | (addr_hit[13] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[12+:4] & ~reg_be))) | (addr_hit[14] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[8+:4] & ~reg_be))) | (addr_hit[15] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[4+:4] & ~reg_be))) | (addr_hit[16] & |(pwrmgr_reg_pkg_PWRMGR_PERMIT[0+:4] & ~reg_be)));
	assign intr_state_we = (addr_hit[0] & reg_we) & !reg_error;
	assign intr_state_wd = reg_wdata[0];
	assign intr_enable_we = (addr_hit[1] & reg_we) & !reg_error;
	assign intr_enable_wd = reg_wdata[0];
	assign intr_test_we = (addr_hit[2] & reg_we) & !reg_error;
	assign intr_test_wd = reg_wdata[0];
	assign alert_test_we = (addr_hit[3] & reg_we) & !reg_error;
	assign alert_test_wd = reg_wdata[0];
	assign ctrl_cfg_regwen_re = (addr_hit[4] & reg_re) & !reg_error;
	assign control_we = (addr_hit[5] & reg_we) & !reg_error;
	assign control_low_power_hint_wd = reg_wdata[0];
	assign control_core_clk_en_wd = reg_wdata[4];
	assign control_io_clk_en_wd = reg_wdata[5];
	assign control_usb_clk_en_lp_wd = reg_wdata[6];
	assign control_usb_clk_en_active_wd = reg_wdata[7];
	assign control_main_pd_n_wd = reg_wdata[8];
	assign cfg_cdc_sync_we = (addr_hit[6] & reg_we) & !reg_error;
	assign cfg_cdc_sync_wd = reg_wdata[0];
	assign wakeup_en_regwen_we = (addr_hit[7] & reg_we) & !reg_error;
	assign wakeup_en_regwen_wd = reg_wdata[0];
	assign wakeup_en_we = (addr_hit[8] & reg_we) & !reg_error;
	assign wakeup_en_en_0_wd = reg_wdata[0];
	assign wakeup_en_en_1_wd = reg_wdata[1];
	assign wakeup_en_en_2_wd = reg_wdata[2];
	assign wakeup_en_en_3_wd = reg_wdata[3];
	assign wakeup_en_en_4_wd = reg_wdata[4];
	assign wakeup_en_en_5_wd = reg_wdata[5];
	assign reset_en_regwen_we = (addr_hit[10] & reg_we) & !reg_error;
	assign reset_en_regwen_wd = reg_wdata[0];
	assign reset_en_we = (addr_hit[11] & reg_we) & !reg_error;
	assign reset_en_en_0_wd = reg_wdata[0];
	assign reset_en_en_1_wd = reg_wdata[1];
	assign wake_info_capture_dis_we = (addr_hit[14] & reg_we) & !reg_error;
	assign wake_info_capture_dis_wd = reg_wdata[0];
	assign wake_info_re = (addr_hit[15] & reg_re) & !reg_error;
	assign wake_info_we = (addr_hit[15] & reg_we) & !reg_error;
	assign wake_info_reasons_wd = reg_wdata[5:0];
	assign wake_info_fall_through_wd = reg_wdata[6];
	assign wake_info_abort_wd = reg_wdata[7];
	always @(*) begin
		reg_we_check = 1'sb0;
		reg_we_check[0] = intr_state_we;
		reg_we_check[1] = intr_enable_we;
		reg_we_check[2] = intr_test_we;
		reg_we_check[3] = alert_test_we;
		reg_we_check[4] = 1'b0;
		reg_we_check[5] = control_gated_we;
		reg_we_check[6] = cfg_cdc_sync_we;
		reg_we_check[7] = wakeup_en_regwen_we;
		reg_we_check[8] = wakeup_en_gated_we;
		reg_we_check[9] = 1'b0;
		reg_we_check[10] = reset_en_regwen_we;
		reg_we_check[11] = reset_en_gated_we;
		reg_we_check[12] = 1'b0;
		reg_we_check[13] = 1'b0;
		reg_we_check[14] = wake_info_capture_dis_we;
		reg_we_check[15] = wake_info_we;
		reg_we_check[16] = 1'b0;
	end
	always @(*) begin
		reg_rdata_next = 1'sb0;
		case (1'b1)
			addr_hit[0]: reg_rdata_next[0] = intr_state_qs;
			addr_hit[1]: reg_rdata_next[0] = intr_enable_qs;
			addr_hit[2]: reg_rdata_next[0] = 1'sb0;
			addr_hit[3]: reg_rdata_next[0] = 1'sb0;
			addr_hit[4]: reg_rdata_next[0] = ctrl_cfg_regwen_qs;
			addr_hit[5]: begin
				reg_rdata_next[0] = control_low_power_hint_qs;
				reg_rdata_next[4] = control_core_clk_en_qs;
				reg_rdata_next[5] = control_io_clk_en_qs;
				reg_rdata_next[6] = control_usb_clk_en_lp_qs;
				reg_rdata_next[7] = control_usb_clk_en_active_qs;
				reg_rdata_next[8] = control_main_pd_n_qs;
			end
			addr_hit[6]: reg_rdata_next[0] = cfg_cdc_sync_qs;
			addr_hit[7]: reg_rdata_next[0] = wakeup_en_regwen_qs;
			addr_hit[8]: begin
				reg_rdata_next[0] = wakeup_en_en_0_qs;
				reg_rdata_next[1] = wakeup_en_en_1_qs;
				reg_rdata_next[2] = wakeup_en_en_2_qs;
				reg_rdata_next[3] = wakeup_en_en_3_qs;
				reg_rdata_next[4] = wakeup_en_en_4_qs;
				reg_rdata_next[5] = wakeup_en_en_5_qs;
			end
			addr_hit[9]: begin
				reg_rdata_next[0] = wake_status_val_0_qs;
				reg_rdata_next[1] = wake_status_val_1_qs;
				reg_rdata_next[2] = wake_status_val_2_qs;
				reg_rdata_next[3] = wake_status_val_3_qs;
				reg_rdata_next[4] = wake_status_val_4_qs;
				reg_rdata_next[5] = wake_status_val_5_qs;
			end
			addr_hit[10]: reg_rdata_next[0] = reset_en_regwen_qs;
			addr_hit[11]: begin
				reg_rdata_next[0] = reset_en_en_0_qs;
				reg_rdata_next[1] = reset_en_en_1_qs;
			end
			addr_hit[12]: begin
				reg_rdata_next[0] = reset_status_val_0_qs;
				reg_rdata_next[1] = reset_status_val_1_qs;
			end
			addr_hit[13]: reg_rdata_next[0] = escalate_reset_status_qs;
			addr_hit[14]: reg_rdata_next[0] = wake_info_capture_dis_qs;
			addr_hit[15]: begin
				reg_rdata_next[5:0] = wake_info_reasons_qs;
				reg_rdata_next[6] = wake_info_fall_through_qs;
				reg_rdata_next[7] = wake_info_abort_qs;
			end
			addr_hit[16]: begin
				reg_rdata_next[0] = fault_status_reg_intg_err_qs;
				reg_rdata_next[1] = fault_status_esc_timeout_qs;
				reg_rdata_next[2] = fault_status_main_pd_glitch_qs;
			end
			default: reg_rdata_next = 1'sb1;
		endcase
	end
	wire shadow_busy;
	assign shadow_busy = 1'b0;
	assign reg_busy = shadow_busy;
	wire unused_wdata;
	wire unused_be;
	assign unused_wdata = ^reg_wdata;
	assign unused_be = ^reg_be;
endmodule
module rv_core_addr_trans (
	clk_i,
	rst_ni,
	region_cfg_i,
	addr_i,
	addr_o
);
	parameter signed [31:0] AddrWidth = 32;
	parameter signed [31:0] NumRegions = 2;
	input wire clk_i;
	input wire rst_ni;
	input wire [(NumRegions * 65) - 1:0] region_cfg_i;
	input wire [AddrWidth - 1:0] addr_i;
	output wire [AddrWidth - 1:0] addr_o;
	wire [(NumRegions * (AddrWidth + AddrWidth)) - 1:0] region_ctrls;
	wire [(NumRegions * AddrWidth) - 1:0] input_masks;
	genvar i;
	generate
		for (i = 0; i < NumRegions; i = i + 1) begin : gen_region_ctrls
			assign input_masks[i * AddrWidth] = 1'b0;
			genvar j;
			for (j = 1; j < AddrWidth; j = j + 1) begin : gen_addr_masks_lower_bits
				assign input_masks[(i * AddrWidth) + j] = ~&region_cfg_i[(i * 65) + ((31 + j) >= 32 ? 31 + j : ((31 + j) + ((31 + j) >= 32 ? (31 + j) - 31 : 33 - (31 + j))) - 1)-:((31 + j) >= 32 ? (31 + j) - 31 : 33 - (31 + j))];
			end
			assign region_ctrls[(((NumRegions - 1) - i) * (AddrWidth + AddrWidth)) + (AddrWidth + (AddrWidth - 1))-:((AddrWidth + (AddrWidth - 1)) >= (AddrWidth + 0) ? ((AddrWidth + (AddrWidth - 1)) - (AddrWidth + 0)) + 1 : ((AddrWidth + 0) - (AddrWidth + (AddrWidth - 1))) + 1)] = ~input_masks[i * AddrWidth+:AddrWidth];
			assign region_ctrls[(((NumRegions - 1) - i) * (AddrWidth + AddrWidth)) + (AddrWidth - 1)-:AddrWidth] = region_cfg_i[(i * 65) + 31-:32];
		end
	endgenerate
	wire [NumRegions - 1:0] all_matches;
	generate
		for (i = 0; i < NumRegions; i = i + 1) begin : gen_region_matches
			assign all_matches[i] = region_cfg_i[(i * 65) + 64] & ((region_cfg_i[(i * 65) + 63-:32] & input_masks[i * AddrWidth+:AddrWidth]) == (addr_i & input_masks[i * AddrWidth+:AddrWidth]));
		end
	endgenerate
	wire sel_match;
	wire [(AddrWidth + AddrWidth) - 1:0] sel_region;
	prim_arbiter_fixed #(
		.N(NumRegions),
		.DW(AddrWidth + AddrWidth),
		.EnDataPort(1)
	) u_sel_region(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.req_i(all_matches),
		.data_i(region_ctrls),
		.valid_o(sel_match),
		.data_o(sel_region),
		.ready_i(1'b1)
	);
	assign addr_o = (sel_match ? (addr_i & sel_region[AddrWidth + (AddrWidth - 1)-:((AddrWidth + (AddrWidth - 1)) >= (AddrWidth + 0) ? ((AddrWidth + (AddrWidth - 1)) - (AddrWidth + 0)) + 1 : ((AddrWidth + 0) - (AddrWidth + (AddrWidth - 1))) + 1)]) | sel_region[AddrWidth - 1-:AddrWidth] : addr_i);
	wire unused_clk;
	wire unused_rst_n;
	assign unused_clk = clk_i;
	assign unused_rst_n = rst_ni;
endmodule
module rv_core_ibex_cfg_reg_top (
	clk_i,
	rst_ni,
	tl_i,
	tl_o,
	tl_win_o,
	tl_win_i,
	reg2hw,
	hw2reg,
	intg_err_o,
	devmode_i
);
	input clk_i;
	input rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_i;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_win_o;
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_win_i;
	output wire [312:0] reg2hw;
	input wire [82:0] hw2reg;
	output wire intg_err_o;
	input devmode_i;
	localparam signed [31:0] AW = 8;
	localparam signed [31:0] DW = 32;
	localparam signed [31:0] DBW = 4;
	wire reg_we;
	wire reg_re;
	wire [7:0] reg_addr;
	wire [31:0] reg_wdata;
	wire [3:0] reg_be;
	wire [31:0] reg_rdata;
	wire reg_error;
	wire addrmiss;
	reg wr_err;
	reg [31:0] reg_rdata_next;
	wire reg_busy;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_reg_h2d;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_reg_d2h;
	wire intg_err;
	tlul_cmd_intg_chk u_chk(
		.tl_i(tl_i),
		.err_o(intg_err)
	);
	wire reg_we_err;
	reg [24:0] reg_we_check;
	prim_reg_we_check #(.OneHotWidth(25)) u_prim_reg_we_check(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.oh_i(reg_we_check),
		.en_i(reg_we && !addrmiss),
		.err_o(reg_we_err)
	);
	reg err_q;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			err_q <= 1'sb0;
		else if (intg_err || reg_we_err)
			err_q <= 1'b1;
	assign intg_err_o = (err_q | intg_err) | reg_we_err;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o_pre;
	tlul_rsp_intg_gen #(
		.EnableRspIntgGen(1),
		.EnableDataIntgGen(1)
	) u_rsp_intg_gen(
		.tl_i(tl_o_pre),
		.tl_o(tl_o)
	);
	wire [(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (2 * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24)) - 1 : (2 * (1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 22)):(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23)] tl_socket_h2d;
	wire [((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (2 * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2)) - 1 : (2 * (1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1))) + ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 0)):((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1)] tl_socket_d2h;
	reg [0:0] reg_steer;
	assign tl_reg_h2d = tl_socket_h2d[(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) + 0+:(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))];
	assign tl_socket_d2h[((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1) + 0+:((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1))] = tl_reg_d2h;
	assign tl_win_o = tl_socket_h2d[(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))+:(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))];
	assign tl_socket_d2h[((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1) + ((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1))+:((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1))] = tl_win_i;
	tlul_socket_1n #(
		.N(2),
		.HReqPass(1'b1),
		.HRspPass(1'b1),
		.DReqPass({2 {1'b1}}),
		.DRspPass({2 {1'b1}}),
		.HReqDepth(4'h0),
		.HRspDepth(4'h0),
		.DReqDepth({2 {4'h0}}),
		.DRspDepth({2 {4'h0}}),
		.ExplicitErrs(1'b0)
	) u_socket(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_h_i(tl_i),
		.tl_h_o(tl_o_pre),
		.tl_d_o(tl_socket_h2d),
		.tl_d_i(tl_socket_d2h),
		.dev_select_i(reg_steer)
	);
	always @(*) begin
		reg_steer = ((128 <= tl_i[(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - 24:(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - 31]) && (159 >= tl_i[(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - 24:(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - 31]) ? 1'd0 : 1'd1);
		if (intg_err)
			reg_steer = 1'd1;
	end
	function automatic [3:0] sv2v_cast_E79FB;
		input reg [3:0] inp;
		sv2v_cast_E79FB = inp;
	endfunction
	tlul_adapter_reg #(
		.RegAw(AW),
		.RegDw(DW),
		.EnableDataIntgGen(0)
	) u_reg_if(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_reg_h2d),
		.tl_o(tl_reg_d2h),
		.en_ifetch_i(sv2v_cast_E79FB(4'h9)),
		.we_o(reg_we),
		.re_o(reg_re),
		.addr_o(reg_addr),
		.wdata_o(reg_wdata),
		.be_o(reg_be),
		.busy_i(reg_busy),
		.rdata_i(reg_rdata),
		.error_i(reg_error)
	);
	assign reg_rdata = reg_rdata_next;
	assign reg_error = ((devmode_i & addrmiss) | wr_err) | intg_err;
	wire alert_test_we;
	wire alert_test_fatal_sw_err_wd;
	wire alert_test_recov_sw_err_wd;
	wire alert_test_fatal_hw_err_wd;
	wire alert_test_recov_hw_err_wd;
	wire sw_recov_err_we;
	wire [3:0] sw_recov_err_qs;
	wire [3:0] sw_recov_err_wd;
	wire sw_fatal_err_we;
	wire [3:0] sw_fatal_err_qs;
	wire [3:0] sw_fatal_err_wd;
	wire ibus_regwen_0_we;
	wire ibus_regwen_0_qs;
	wire ibus_regwen_0_wd;
	wire ibus_regwen_1_we;
	wire ibus_regwen_1_qs;
	wire ibus_regwen_1_wd;
	wire ibus_addr_en_0_we;
	wire ibus_addr_en_0_qs;
	wire ibus_addr_en_0_wd;
	wire ibus_addr_en_1_we;
	wire ibus_addr_en_1_qs;
	wire ibus_addr_en_1_wd;
	wire ibus_addr_matching_0_we;
	wire [31:0] ibus_addr_matching_0_qs;
	wire [31:0] ibus_addr_matching_0_wd;
	wire ibus_addr_matching_1_we;
	wire [31:0] ibus_addr_matching_1_qs;
	wire [31:0] ibus_addr_matching_1_wd;
	wire ibus_remap_addr_0_we;
	wire [31:0] ibus_remap_addr_0_qs;
	wire [31:0] ibus_remap_addr_0_wd;
	wire ibus_remap_addr_1_we;
	wire [31:0] ibus_remap_addr_1_qs;
	wire [31:0] ibus_remap_addr_1_wd;
	wire dbus_regwen_0_we;
	wire dbus_regwen_0_qs;
	wire dbus_regwen_0_wd;
	wire dbus_regwen_1_we;
	wire dbus_regwen_1_qs;
	wire dbus_regwen_1_wd;
	wire dbus_addr_en_0_we;
	wire dbus_addr_en_0_qs;
	wire dbus_addr_en_0_wd;
	wire dbus_addr_en_1_we;
	wire dbus_addr_en_1_qs;
	wire dbus_addr_en_1_wd;
	wire dbus_addr_matching_0_we;
	wire [31:0] dbus_addr_matching_0_qs;
	wire [31:0] dbus_addr_matching_0_wd;
	wire dbus_addr_matching_1_we;
	wire [31:0] dbus_addr_matching_1_qs;
	wire [31:0] dbus_addr_matching_1_wd;
	wire dbus_remap_addr_0_we;
	wire [31:0] dbus_remap_addr_0_qs;
	wire [31:0] dbus_remap_addr_0_wd;
	wire dbus_remap_addr_1_we;
	wire [31:0] dbus_remap_addr_1_qs;
	wire [31:0] dbus_remap_addr_1_wd;
	wire nmi_enable_we;
	wire nmi_enable_alert_en_qs;
	wire nmi_enable_alert_en_wd;
	wire nmi_enable_wdog_en_qs;
	wire nmi_enable_wdog_en_wd;
	wire nmi_state_we;
	wire nmi_state_alert_qs;
	wire nmi_state_alert_wd;
	wire nmi_state_wdog_qs;
	wire nmi_state_wdog_wd;
	wire err_status_we;
	wire err_status_reg_intg_err_qs;
	wire err_status_reg_intg_err_wd;
	wire err_status_fatal_intg_err_qs;
	wire err_status_fatal_intg_err_wd;
	wire err_status_fatal_core_err_qs;
	wire err_status_fatal_core_err_wd;
	wire err_status_recov_core_err_qs;
	wire err_status_recov_core_err_wd;
	wire rnd_data_re;
	wire [31:0] rnd_data_qs;
	wire rnd_status_re;
	wire rnd_status_rnd_data_valid_qs;
	wire rnd_status_rnd_data_fips_qs;
	wire fpga_info_re;
	wire [31:0] fpga_info_qs;
	wire alert_test_qe;
	wire [3:0] alert_test_flds_we;
	assign alert_test_qe = &alert_test_flds_we;
	prim_subreg_ext #(.DW(1)) u_alert_test_fatal_sw_err(
		.re(1'b0),
		.we(alert_test_we),
		.wd(alert_test_fatal_sw_err_wd),
		.d(1'sb0),
		.qe(alert_test_flds_we[0]),
		.q(reg2hw[312])
	);
	assign reg2hw[311] = alert_test_qe;
	prim_subreg_ext #(.DW(1)) u_alert_test_recov_sw_err(
		.re(1'b0),
		.we(alert_test_we),
		.wd(alert_test_recov_sw_err_wd),
		.d(1'sb0),
		.qe(alert_test_flds_we[1]),
		.q(reg2hw[310])
	);
	assign reg2hw[309] = alert_test_qe;
	prim_subreg_ext #(.DW(1)) u_alert_test_fatal_hw_err(
		.re(1'b0),
		.we(alert_test_we),
		.wd(alert_test_fatal_hw_err_wd),
		.d(1'sb0),
		.qe(alert_test_flds_we[2]),
		.q(reg2hw[308])
	);
	assign reg2hw[307] = alert_test_qe;
	prim_subreg_ext #(.DW(1)) u_alert_test_recov_hw_err(
		.re(1'b0),
		.we(alert_test_we),
		.wd(alert_test_recov_hw_err_wd),
		.d(1'sb0),
		.qe(alert_test_flds_we[3]),
		.q(reg2hw[306])
	);
	assign reg2hw[305] = alert_test_qe;
	prim_subreg #(
		.DW(4),
		.SwAccess(3'd0),
		.RESVAL(4'h9)
	) u_sw_recov_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(sw_recov_err_we),
		.wd(sw_recov_err_wd),
		.de(hw2reg[78]),
		.d(hw2reg[82-:4]),
		.q(reg2hw[304-:4]),
		.qs(sw_recov_err_qs)
	);
	prim_subreg #(
		.DW(4),
		.SwAccess(3'd5),
		.RESVAL(4'h9)
	) u_sw_fatal_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(sw_fatal_err_we),
		.wd(sw_fatal_err_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[300-:4]),
		.qs(sw_fatal_err_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_ibus_regwen_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ibus_regwen_0_we),
		.wd(ibus_regwen_0_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(ibus_regwen_0_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_ibus_regwen_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ibus_regwen_1_we),
		.wd(ibus_regwen_1_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(ibus_regwen_1_qs)
	);
	wire ibus_addr_en_0_gated_we;
	assign ibus_addr_en_0_gated_we = ibus_addr_en_0_we & ibus_regwen_0_qs;
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_ibus_addr_en_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ibus_addr_en_0_gated_we),
		.wd(ibus_addr_en_0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[295]),
		.qs(ibus_addr_en_0_qs)
	);
	wire ibus_addr_en_1_gated_we;
	assign ibus_addr_en_1_gated_we = ibus_addr_en_1_we & ibus_regwen_1_qs;
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_ibus_addr_en_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ibus_addr_en_1_gated_we),
		.wd(ibus_addr_en_1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[296]),
		.qs(ibus_addr_en_1_qs)
	);
	wire ibus_addr_matching_0_gated_we;
	assign ibus_addr_matching_0_gated_we = ibus_addr_matching_0_we & ibus_regwen_0_qs;
	prim_subreg #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_ibus_addr_matching_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ibus_addr_matching_0_gated_we),
		.wd(ibus_addr_matching_0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[262-:32]),
		.qs(ibus_addr_matching_0_qs)
	);
	wire ibus_addr_matching_1_gated_we;
	assign ibus_addr_matching_1_gated_we = ibus_addr_matching_1_we & ibus_regwen_1_qs;
	prim_subreg #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_ibus_addr_matching_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ibus_addr_matching_1_gated_we),
		.wd(ibus_addr_matching_1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[294-:32]),
		.qs(ibus_addr_matching_1_qs)
	);
	wire ibus_remap_addr_0_gated_we;
	assign ibus_remap_addr_0_gated_we = ibus_remap_addr_0_we & ibus_regwen_0_qs;
	prim_subreg #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_ibus_remap_addr_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ibus_remap_addr_0_gated_we),
		.wd(ibus_remap_addr_0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[198-:32]),
		.qs(ibus_remap_addr_0_qs)
	);
	wire ibus_remap_addr_1_gated_we;
	assign ibus_remap_addr_1_gated_we = ibus_remap_addr_1_we & ibus_regwen_1_qs;
	prim_subreg #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_ibus_remap_addr_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(ibus_remap_addr_1_gated_we),
		.wd(ibus_remap_addr_1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[230-:32]),
		.qs(ibus_remap_addr_1_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_dbus_regwen_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(dbus_regwen_0_we),
		.wd(dbus_regwen_0_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(dbus_regwen_0_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd5),
		.RESVAL(1'h1)
	) u_dbus_regwen_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(dbus_regwen_1_we),
		.wd(dbus_regwen_1_wd),
		.de(1'b0),
		.d(1'sb0),
		.qs(dbus_regwen_1_qs)
	);
	wire dbus_addr_en_0_gated_we;
	assign dbus_addr_en_0_gated_we = dbus_addr_en_0_we & dbus_regwen_0_qs;
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_dbus_addr_en_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(dbus_addr_en_0_gated_we),
		.wd(dbus_addr_en_0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[165]),
		.qs(dbus_addr_en_0_qs)
	);
	wire dbus_addr_en_1_gated_we;
	assign dbus_addr_en_1_gated_we = dbus_addr_en_1_we & dbus_regwen_1_qs;
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd0),
		.RESVAL(1'h0)
	) u_dbus_addr_en_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(dbus_addr_en_1_gated_we),
		.wd(dbus_addr_en_1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[166]),
		.qs(dbus_addr_en_1_qs)
	);
	wire dbus_addr_matching_0_gated_we;
	assign dbus_addr_matching_0_gated_we = dbus_addr_matching_0_we & dbus_regwen_0_qs;
	prim_subreg #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_dbus_addr_matching_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(dbus_addr_matching_0_gated_we),
		.wd(dbus_addr_matching_0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[132-:32]),
		.qs(dbus_addr_matching_0_qs)
	);
	wire dbus_addr_matching_1_gated_we;
	assign dbus_addr_matching_1_gated_we = dbus_addr_matching_1_we & dbus_regwen_1_qs;
	prim_subreg #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_dbus_addr_matching_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(dbus_addr_matching_1_gated_we),
		.wd(dbus_addr_matching_1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[164-:32]),
		.qs(dbus_addr_matching_1_qs)
	);
	wire dbus_remap_addr_0_gated_we;
	assign dbus_remap_addr_0_gated_we = dbus_remap_addr_0_we & dbus_regwen_0_qs;
	prim_subreg #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_dbus_remap_addr_0(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(dbus_remap_addr_0_gated_we),
		.wd(dbus_remap_addr_0_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[68-:32]),
		.qs(dbus_remap_addr_0_qs)
	);
	wire dbus_remap_addr_1_gated_we;
	assign dbus_remap_addr_1_gated_we = dbus_remap_addr_1_we & dbus_regwen_1_qs;
	prim_subreg #(
		.DW(32),
		.SwAccess(3'd0),
		.RESVAL(32'h00000000)
	) u_dbus_remap_addr_1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(dbus_remap_addr_1_gated_we),
		.wd(dbus_remap_addr_1_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[100-:32]),
		.qs(dbus_remap_addr_1_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd4),
		.RESVAL(1'h0)
	) u_nmi_enable_alert_en(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(nmi_enable_we),
		.wd(nmi_enable_alert_en_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[36]),
		.qs(nmi_enable_alert_en_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd4),
		.RESVAL(1'h0)
	) u_nmi_enable_wdog_en(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(nmi_enable_we),
		.wd(nmi_enable_wdog_en_wd),
		.de(1'b0),
		.d(1'sb0),
		.q(reg2hw[35]),
		.qs(nmi_enable_wdog_en_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_nmi_state_alert(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(nmi_state_we),
		.wd(nmi_state_alert_wd),
		.de(hw2reg[76]),
		.d(hw2reg[77]),
		.q(reg2hw[34]),
		.qs(nmi_state_alert_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_nmi_state_wdog(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(nmi_state_we),
		.wd(nmi_state_wdog_wd),
		.de(hw2reg[74]),
		.d(hw2reg[75]),
		.q(reg2hw[33]),
		.qs(nmi_state_wdog_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_err_status_reg_intg_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(err_status_we),
		.wd(err_status_reg_intg_err_wd),
		.de(hw2reg[72]),
		.d(hw2reg[73]),
		.qs(err_status_reg_intg_err_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_err_status_fatal_intg_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(err_status_we),
		.wd(err_status_fatal_intg_err_wd),
		.de(hw2reg[70]),
		.d(hw2reg[71]),
		.qs(err_status_fatal_intg_err_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_err_status_fatal_core_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(err_status_we),
		.wd(err_status_fatal_core_err_wd),
		.de(hw2reg[68]),
		.d(hw2reg[69]),
		.qs(err_status_fatal_core_err_qs)
	);
	prim_subreg #(
		.DW(1),
		.SwAccess(3'd3),
		.RESVAL(1'h0)
	) u_err_status_recov_core_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.we(err_status_we),
		.wd(err_status_recov_core_err_wd),
		.de(hw2reg[66]),
		.d(hw2reg[67]),
		.qs(err_status_recov_core_err_qs)
	);
	prim_subreg_ext #(.DW(32)) u_rnd_data(
		.re(rnd_data_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[65-:32]),
		.qre(reg2hw[0]),
		.q(reg2hw[32-:32]),
		.qs(rnd_data_qs)
	);
	prim_subreg_ext #(.DW(1)) u_rnd_status_rnd_data_valid(
		.re(rnd_status_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[33]),
		.qs(rnd_status_rnd_data_valid_qs)
	);
	prim_subreg_ext #(.DW(1)) u_rnd_status_rnd_data_fips(
		.re(rnd_status_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[32]),
		.qs(rnd_status_rnd_data_fips_qs)
	);
	prim_subreg_ext #(.DW(32)) u_fpga_info(
		.re(fpga_info_re),
		.we(1'b0),
		.wd(1'sb0),
		.d(hw2reg[31-:32]),
		.qs(fpga_info_qs)
	);
	reg [24:0] addr_hit;
	localparam signed [31:0] rv_core_ibex_reg_pkg_CfgAw = 8;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_ALERT_TEST_OFFSET = 8'h00;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_DBUS_ADDR_EN_0_OFFSET = 8'h34;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_DBUS_ADDR_EN_1_OFFSET = 8'h38;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_DBUS_ADDR_MATCHING_0_OFFSET = 8'h3c;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_DBUS_ADDR_MATCHING_1_OFFSET = 8'h40;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_DBUS_REGWEN_0_OFFSET = 8'h2c;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_DBUS_REGWEN_1_OFFSET = 8'h30;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_DBUS_REMAP_ADDR_0_OFFSET = 8'h44;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_DBUS_REMAP_ADDR_1_OFFSET = 8'h48;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_ERR_STATUS_OFFSET = 8'h54;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_FPGA_INFO_OFFSET = 8'h60;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_IBUS_ADDR_EN_0_OFFSET = 8'h14;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_IBUS_ADDR_EN_1_OFFSET = 8'h18;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_IBUS_ADDR_MATCHING_0_OFFSET = 8'h1c;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_IBUS_ADDR_MATCHING_1_OFFSET = 8'h20;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_IBUS_REGWEN_0_OFFSET = 8'h0c;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_IBUS_REGWEN_1_OFFSET = 8'h10;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_IBUS_REMAP_ADDR_0_OFFSET = 8'h24;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_IBUS_REMAP_ADDR_1_OFFSET = 8'h28;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_NMI_ENABLE_OFFSET = 8'h4c;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_NMI_STATE_OFFSET = 8'h50;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_RND_DATA_OFFSET = 8'h58;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_RND_STATUS_OFFSET = 8'h5c;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_SW_FATAL_ERR_OFFSET = 8'h08;
	localparam [7:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_SW_RECOV_ERR_OFFSET = 8'h04;
	always @(*) begin
		addr_hit = 1'sb0;
		addr_hit[0] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_ALERT_TEST_OFFSET;
		addr_hit[1] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_SW_RECOV_ERR_OFFSET;
		addr_hit[2] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_SW_FATAL_ERR_OFFSET;
		addr_hit[3] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_IBUS_REGWEN_0_OFFSET;
		addr_hit[4] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_IBUS_REGWEN_1_OFFSET;
		addr_hit[5] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_IBUS_ADDR_EN_0_OFFSET;
		addr_hit[6] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_IBUS_ADDR_EN_1_OFFSET;
		addr_hit[7] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_IBUS_ADDR_MATCHING_0_OFFSET;
		addr_hit[8] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_IBUS_ADDR_MATCHING_1_OFFSET;
		addr_hit[9] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_IBUS_REMAP_ADDR_0_OFFSET;
		addr_hit[10] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_IBUS_REMAP_ADDR_1_OFFSET;
		addr_hit[11] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_DBUS_REGWEN_0_OFFSET;
		addr_hit[12] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_DBUS_REGWEN_1_OFFSET;
		addr_hit[13] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_DBUS_ADDR_EN_0_OFFSET;
		addr_hit[14] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_DBUS_ADDR_EN_1_OFFSET;
		addr_hit[15] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_DBUS_ADDR_MATCHING_0_OFFSET;
		addr_hit[16] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_DBUS_ADDR_MATCHING_1_OFFSET;
		addr_hit[17] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_DBUS_REMAP_ADDR_0_OFFSET;
		addr_hit[18] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_DBUS_REMAP_ADDR_1_OFFSET;
		addr_hit[19] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_NMI_ENABLE_OFFSET;
		addr_hit[20] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_NMI_STATE_OFFSET;
		addr_hit[21] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_ERR_STATUS_OFFSET;
		addr_hit[22] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_RND_DATA_OFFSET;
		addr_hit[23] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_RND_STATUS_OFFSET;
		addr_hit[24] = reg_addr == rv_core_ibex_reg_pkg_RV_CORE_IBEX_FPGA_INFO_OFFSET;
	end
	assign addrmiss = (reg_re || reg_we ? ~|addr_hit : 1'b0);
	localparam [99:0] rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT = 100'b0001000100010001000100010001111111111111111100010001000100011111111111111111000100010011111100011111;
	always @(*) wr_err = reg_we & (((((((((((((((((((((((((addr_hit[0] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[96+:4] & ~reg_be)) | (addr_hit[1] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[92+:4] & ~reg_be))) | (addr_hit[2] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[88+:4] & ~reg_be))) | (addr_hit[3] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[84+:4] & ~reg_be))) | (addr_hit[4] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[80+:4] & ~reg_be))) | (addr_hit[5] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[76+:4] & ~reg_be))) | (addr_hit[6] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[72+:4] & ~reg_be))) | (addr_hit[7] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[68+:4] & ~reg_be))) | (addr_hit[8] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[64+:4] & ~reg_be))) | (addr_hit[9] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[60+:4] & ~reg_be))) | (addr_hit[10] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[56+:4] & ~reg_be))) | (addr_hit[11] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[52+:4] & ~reg_be))) | (addr_hit[12] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[48+:4] & ~reg_be))) | (addr_hit[13] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[44+:4] & ~reg_be))) | (addr_hit[14] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[40+:4] & ~reg_be))) | (addr_hit[15] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[36+:4] & ~reg_be))) | (addr_hit[16] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[32+:4] & ~reg_be))) | (addr_hit[17] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[28+:4] & ~reg_be))) | (addr_hit[18] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[24+:4] & ~reg_be))) | (addr_hit[19] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[20+:4] & ~reg_be))) | (addr_hit[20] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[16+:4] & ~reg_be))) | (addr_hit[21] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[12+:4] & ~reg_be))) | (addr_hit[22] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[8+:4] & ~reg_be))) | (addr_hit[23] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[4+:4] & ~reg_be))) | (addr_hit[24] & |(rv_core_ibex_reg_pkg_RV_CORE_IBEX_CFG_PERMIT[0+:4] & ~reg_be)));
	assign alert_test_we = (addr_hit[0] & reg_we) & !reg_error;
	assign alert_test_fatal_sw_err_wd = reg_wdata[0];
	assign alert_test_recov_sw_err_wd = reg_wdata[1];
	assign alert_test_fatal_hw_err_wd = reg_wdata[2];
	assign alert_test_recov_hw_err_wd = reg_wdata[3];
	assign sw_recov_err_we = (addr_hit[1] & reg_we) & !reg_error;
	assign sw_recov_err_wd = reg_wdata[3:0];
	assign sw_fatal_err_we = (addr_hit[2] & reg_we) & !reg_error;
	assign sw_fatal_err_wd = reg_wdata[3:0];
	assign ibus_regwen_0_we = (addr_hit[3] & reg_we) & !reg_error;
	assign ibus_regwen_0_wd = reg_wdata[0];
	assign ibus_regwen_1_we = (addr_hit[4] & reg_we) & !reg_error;
	assign ibus_regwen_1_wd = reg_wdata[0];
	assign ibus_addr_en_0_we = (addr_hit[5] & reg_we) & !reg_error;
	assign ibus_addr_en_0_wd = reg_wdata[0];
	assign ibus_addr_en_1_we = (addr_hit[6] & reg_we) & !reg_error;
	assign ibus_addr_en_1_wd = reg_wdata[0];
	assign ibus_addr_matching_0_we = (addr_hit[7] & reg_we) & !reg_error;
	assign ibus_addr_matching_0_wd = reg_wdata[31:0];
	assign ibus_addr_matching_1_we = (addr_hit[8] & reg_we) & !reg_error;
	assign ibus_addr_matching_1_wd = reg_wdata[31:0];
	assign ibus_remap_addr_0_we = (addr_hit[9] & reg_we) & !reg_error;
	assign ibus_remap_addr_0_wd = reg_wdata[31:0];
	assign ibus_remap_addr_1_we = (addr_hit[10] & reg_we) & !reg_error;
	assign ibus_remap_addr_1_wd = reg_wdata[31:0];
	assign dbus_regwen_0_we = (addr_hit[11] & reg_we) & !reg_error;
	assign dbus_regwen_0_wd = reg_wdata[0];
	assign dbus_regwen_1_we = (addr_hit[12] & reg_we) & !reg_error;
	assign dbus_regwen_1_wd = reg_wdata[0];
	assign dbus_addr_en_0_we = (addr_hit[13] & reg_we) & !reg_error;
	assign dbus_addr_en_0_wd = reg_wdata[0];
	assign dbus_addr_en_1_we = (addr_hit[14] & reg_we) & !reg_error;
	assign dbus_addr_en_1_wd = reg_wdata[0];
	assign dbus_addr_matching_0_we = (addr_hit[15] & reg_we) & !reg_error;
	assign dbus_addr_matching_0_wd = reg_wdata[31:0];
	assign dbus_addr_matching_1_we = (addr_hit[16] & reg_we) & !reg_error;
	assign dbus_addr_matching_1_wd = reg_wdata[31:0];
	assign dbus_remap_addr_0_we = (addr_hit[17] & reg_we) & !reg_error;
	assign dbus_remap_addr_0_wd = reg_wdata[31:0];
	assign dbus_remap_addr_1_we = (addr_hit[18] & reg_we) & !reg_error;
	assign dbus_remap_addr_1_wd = reg_wdata[31:0];
	assign nmi_enable_we = (addr_hit[19] & reg_we) & !reg_error;
	assign nmi_enable_alert_en_wd = reg_wdata[0];
	assign nmi_enable_wdog_en_wd = reg_wdata[1];
	assign nmi_state_we = (addr_hit[20] & reg_we) & !reg_error;
	assign nmi_state_alert_wd = reg_wdata[0];
	assign nmi_state_wdog_wd = reg_wdata[1];
	assign err_status_we = (addr_hit[21] & reg_we) & !reg_error;
	assign err_status_reg_intg_err_wd = reg_wdata[0];
	assign err_status_fatal_intg_err_wd = reg_wdata[8];
	assign err_status_fatal_core_err_wd = reg_wdata[9];
	assign err_status_recov_core_err_wd = reg_wdata[10];
	assign rnd_data_re = (addr_hit[22] & reg_re) & !reg_error;
	assign rnd_status_re = (addr_hit[23] & reg_re) & !reg_error;
	assign fpga_info_re = (addr_hit[24] & reg_re) & !reg_error;
	always @(*) begin
		reg_we_check = 1'sb0;
		reg_we_check[0] = alert_test_we;
		reg_we_check[1] = sw_recov_err_we;
		reg_we_check[2] = sw_fatal_err_we;
		reg_we_check[3] = ibus_regwen_0_we;
		reg_we_check[4] = ibus_regwen_1_we;
		reg_we_check[5] = ibus_addr_en_0_gated_we;
		reg_we_check[6] = ibus_addr_en_1_gated_we;
		reg_we_check[7] = ibus_addr_matching_0_gated_we;
		reg_we_check[8] = ibus_addr_matching_1_gated_we;
		reg_we_check[9] = ibus_remap_addr_0_gated_we;
		reg_we_check[10] = ibus_remap_addr_1_gated_we;
		reg_we_check[11] = dbus_regwen_0_we;
		reg_we_check[12] = dbus_regwen_1_we;
		reg_we_check[13] = dbus_addr_en_0_gated_we;
		reg_we_check[14] = dbus_addr_en_1_gated_we;
		reg_we_check[15] = dbus_addr_matching_0_gated_we;
		reg_we_check[16] = dbus_addr_matching_1_gated_we;
		reg_we_check[17] = dbus_remap_addr_0_gated_we;
		reg_we_check[18] = dbus_remap_addr_1_gated_we;
		reg_we_check[19] = nmi_enable_we;
		reg_we_check[20] = nmi_state_we;
		reg_we_check[21] = err_status_we;
		reg_we_check[22] = 1'b0;
		reg_we_check[23] = 1'b0;
		reg_we_check[24] = 1'b0;
	end
	always @(*) begin
		reg_rdata_next = 1'sb0;
		case (1'b1)
			addr_hit[0]: begin
				reg_rdata_next[0] = 1'sb0;
				reg_rdata_next[1] = 1'sb0;
				reg_rdata_next[2] = 1'sb0;
				reg_rdata_next[3] = 1'sb0;
			end
			addr_hit[1]: reg_rdata_next[3:0] = sw_recov_err_qs;
			addr_hit[2]: reg_rdata_next[3:0] = sw_fatal_err_qs;
			addr_hit[3]: reg_rdata_next[0] = ibus_regwen_0_qs;
			addr_hit[4]: reg_rdata_next[0] = ibus_regwen_1_qs;
			addr_hit[5]: reg_rdata_next[0] = ibus_addr_en_0_qs;
			addr_hit[6]: reg_rdata_next[0] = ibus_addr_en_1_qs;
			addr_hit[7]: reg_rdata_next[31:0] = ibus_addr_matching_0_qs;
			addr_hit[8]: reg_rdata_next[31:0] = ibus_addr_matching_1_qs;
			addr_hit[9]: reg_rdata_next[31:0] = ibus_remap_addr_0_qs;
			addr_hit[10]: reg_rdata_next[31:0] = ibus_remap_addr_1_qs;
			addr_hit[11]: reg_rdata_next[0] = dbus_regwen_0_qs;
			addr_hit[12]: reg_rdata_next[0] = dbus_regwen_1_qs;
			addr_hit[13]: reg_rdata_next[0] = dbus_addr_en_0_qs;
			addr_hit[14]: reg_rdata_next[0] = dbus_addr_en_1_qs;
			addr_hit[15]: reg_rdata_next[31:0] = dbus_addr_matching_0_qs;
			addr_hit[16]: reg_rdata_next[31:0] = dbus_addr_matching_1_qs;
			addr_hit[17]: reg_rdata_next[31:0] = dbus_remap_addr_0_qs;
			addr_hit[18]: reg_rdata_next[31:0] = dbus_remap_addr_1_qs;
			addr_hit[19]: begin
				reg_rdata_next[0] = nmi_enable_alert_en_qs;
				reg_rdata_next[1] = nmi_enable_wdog_en_qs;
			end
			addr_hit[20]: begin
				reg_rdata_next[0] = nmi_state_alert_qs;
				reg_rdata_next[1] = nmi_state_wdog_qs;
			end
			addr_hit[21]: begin
				reg_rdata_next[0] = err_status_reg_intg_err_qs;
				reg_rdata_next[8] = err_status_fatal_intg_err_qs;
				reg_rdata_next[9] = err_status_fatal_core_err_qs;
				reg_rdata_next[10] = err_status_recov_core_err_qs;
			end
			addr_hit[22]: reg_rdata_next[31:0] = rnd_data_qs;
			addr_hit[23]: begin
				reg_rdata_next[0] = rnd_status_rnd_data_valid_qs;
				reg_rdata_next[1] = rnd_status_rnd_data_fips_qs;
			end
			addr_hit[24]: reg_rdata_next[31:0] = fpga_info_qs;
			default: reg_rdata_next = 1'sb1;
		endcase
	end
	wire shadow_busy;
	assign shadow_busy = 1'b0;
	assign reg_busy = shadow_busy;
	wire unused_wdata;
	wire unused_be;
	assign unused_wdata = ^reg_wdata;
	assign unused_be = ^reg_be;
endmodule
module sram2tlul (
	clk_i,
	rst_ni,
	tl_o,
	tl_i,
	mem_req_i,
	mem_write_i,
	mem_addr_i,
	mem_wdata_i,
	mem_rvalid_o,
	mem_rdata_o,
	mem_error_o
);
	parameter signed [31:0] SramAw = 12;
	parameter signed [31:0] SramDw = 32;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	parameter [31:0] TlBaseAddr = 'h0;
	input clk_i;
	input rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_o;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_i;
	input mem_req_i;
	input mem_write_i;
	input [SramAw - 1:0] mem_addr_i;
	input [SramDw - 1:0] mem_wdata_i;
	output wire mem_rvalid_o;
	output wire [SramDw - 1:0] mem_rdata_o;
	output wire [1:0] mem_error_o;
	localparam [31:0] SRAM_DWB = $clog2(SramDw / 8);
	assign tl_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] = mem_req_i;
	assign tl_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] = (mem_write_i ? 3'h0 : 3'h4);
	assign tl_o[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] = 1'sb0;
	function automatic [top_pkg_TL_SZW - 1:0] sv2v_cast_53D14;
		input reg [top_pkg_TL_SZW - 1:0] inp;
		sv2v_cast_53D14 = inp;
	endfunction
	assign tl_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)] = sv2v_cast_53D14(SRAM_DWB);
	assign tl_o[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) >= (32'sd32 + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 56)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1)] = 1'sb0;
	assign tl_o[top_pkg_TL_AW + (top_pkg_TL_DBW + 55)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)] = TlBaseAddr | {{(top_pkg_TL_AW - SramAw) - SRAM_DWB {1'b0}}, mem_addr_i, {SRAM_DWB {1'b0}}};
	assign tl_o[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))] = 1'sb1;
	assign tl_o[55-:32] = mem_wdata_i;
	assign tl_o[23-:23] = 1'sb0;
	assign tl_o[0] = 1'b1;
	assign mem_rvalid_o = tl_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] && (tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)] == 3'h1);
	assign mem_rdata_o = tl_i[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)];
	assign mem_error_o = {2 {tl_i[1]}};
endmodule
module tlul_adapter_host (
	clk_i,
	rst_ni,
	req_i,
	gnt_o,
	addr_i,
	we_i,
	wdata_i,
	wdata_intg_i,
	be_i,
	instr_type_i,
	valid_o,
	rdata_o,
	rdata_intg_o,
	err_o,
	intg_err_o,
	tl_o,
	tl_i
);
	parameter [31:0] MAX_REQS = 2;
	parameter [0:0] EnableDataIntgGen = 0;
	parameter [0:0] EnableRspDataIntgCheck = 0;
	input clk_i;
	input rst_ni;
	input req_i;
	output wire gnt_o;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	input wire [31:0] addr_i;
	input wire we_i;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	input wire [31:0] wdata_i;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	input wire [6:0] wdata_intg_i;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	input wire [top_pkg_TL_DBW - 1:0] be_i;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	input wire [3:0] instr_type_i;
	output wire valid_o;
	output wire [31:0] rdata_o;
	output wire [6:0] rdata_intg_o;
	output wire err_o;
	output wire intg_err_o;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_o;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_i;
	localparam signed [31:0] WordSize = $clog2(top_pkg_TL_DBW);
	wire [7:0] tl_source;
	wire [top_pkg_TL_DBW - 1:0] tl_be;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_out;
	function automatic [7:0] sv2v_cast_8;
		input reg [7:0] inp;
		sv2v_cast_8 = inp;
	endfunction
	generate
		if (MAX_REQS == 1) begin : g_single_req
			assign tl_source = 1'sb0;
		end
		else begin : g_multiple_reqs
			localparam signed [31:0] ReqNumW = $clog2(MAX_REQS);
			localparam [31:0] MaxSource = MAX_REQS - 1;
			reg [ReqNumW - 1:0] source_d;
			reg [ReqNumW - 1:0] source_q;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					source_q <= 1'sb0;
				else
					source_q <= source_d;
			always @(*) begin
				source_d = source_q;
				if (req_i && gnt_o)
					if (source_q == MaxSource[ReqNumW - 1:0])
						source_d = 1'sb0;
					else
						source_d = source_q + 1;
			end
			assign tl_source = sv2v_cast_8(source_q);
		end
	endgenerate
	assign tl_be = (~we_i ? {top_pkg_TL_DBW {1'b1}} : be_i);
	function automatic signed [top_pkg_TL_SZW - 1:0] sv2v_cast_53D14_signed;
		input reg signed [top_pkg_TL_SZW - 1:0] inp;
		sv2v_cast_53D14_signed = inp;
	endfunction
	function automatic [6:0] sv2v_cast_6BD77;
		input reg [6:0] inp;
		sv2v_cast_6BD77 = inp;
	endfunction
	function automatic [top_pkg_TL_SZW - 1:0] sv2v_cast_87CE4;
		input reg [top_pkg_TL_SZW - 1:0] inp;
		sv2v_cast_87CE4 = inp;
	endfunction
	function automatic [7:0] sv2v_cast_DE545;
		input reg [7:0] inp;
		sv2v_cast_DE545 = inp;
	endfunction
	function automatic [31:0] sv2v_cast_4B555;
		input reg [31:0] inp;
		sv2v_cast_4B555 = inp;
	endfunction
	function automatic [31:0] sv2v_cast_B57C0;
		input reg [31:0] inp;
		sv2v_cast_B57C0 = inp;
	endfunction
	function automatic [22:0] sv2v_cast_CEE27;
		input reg [22:0] inp;
		sv2v_cast_CEE27 = inp;
	endfunction
	assign tl_out = {req_i, (~we_i ? 3'h4 : (&be_i ? 3'h0 : 3'h1)), 3'h0, sv2v_cast_87CE4(sv2v_cast_53D14_signed(WordSize)), sv2v_cast_DE545(tl_source), sv2v_cast_4B555({addr_i[31:WordSize], {WordSize {1'b0}}}), tl_be, sv2v_cast_B57C0(wdata_i), sv2v_cast_CEE27({5'b00000, instr_type_i, sv2v_cast_6BD77(1'sb0), wdata_intg_i}), 1'b1};
	tlul_cmd_intg_gen #(.EnableDataIntgGen(EnableDataIntgGen)) u_cmd_intg_gen(
		.tl_i(tl_out),
		.tl_o(tl_o)
	);
	assign gnt_o = tl_i[0];
	assign valid_o = tl_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))];
	assign rdata_o = tl_i[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)];
	assign rdata_intg_o = tl_i[((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 7)-:tlul_pkg_DataIntgWidth];
	wire intg_err;
	tlul_rsp_intg_chk #(.EnableRspDataIntgCheck(EnableRspDataIntgCheck)) u_rsp_chk(
		.tl_i(tl_i),
		.err_o(intg_err)
	);
	reg intg_err_q;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			intg_err_q <= 1'sb0;
		else if (intg_err)
			intg_err_q <= 1'b1;
	assign err_o = tl_i[1] | intg_err;
	assign intg_err_o = intg_err_q | intg_err;
	wire unused_addr_bottom_bits;
	assign unused_addr_bottom_bits = ^addr_i[WordSize - 1:0];
	wire unused_tl_i_fields;
	assign unused_tl_i_fields = ^{tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)], tl_i[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)], tl_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)], tl_i[top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))-:((32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))) >= ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) + 1 : ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) + 1)], tl_i[top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))-:(((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)) >= (32'sd32 + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) + 1 : ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) + 1)], tl_i[(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1-:(((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) >= 2 ? (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 0 : 3 - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))]};
endmodule
module tlul_adapter_reg (
	clk_i,
	rst_ni,
	tl_i,
	tl_o,
	en_ifetch_i,
	intg_error_o,
	re_o,
	we_o,
	addr_o,
	wdata_o,
	be_o,
	busy_i,
	rdata_i,
	error_i
);
	parameter [0:0] CmdIntgCheck = 0;
	parameter [0:0] EnableRspIntgGen = 0;
	parameter [0:0] EnableDataIntgGen = 0;
	parameter signed [31:0] RegAw = 8;
	parameter signed [31:0] RegDw = 32;
	parameter signed [31:0] AccessLatency = 0;
	localparam signed [31:0] RegBw = RegDw / 8;
	input clk_i;
	input rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_i;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	input wire [3:0] en_ifetch_i;
	output wire intg_error_o;
	output wire re_o;
	output wire we_o;
	output wire [RegAw - 1:0] addr_o;
	output wire [RegDw - 1:0] wdata_o;
	output wire [RegBw - 1:0] be_o;
	input busy_i;
	input [RegDw - 1:0] rdata_i;
	input error_i;
	localparam signed [31:0] IW = top_pkg_TL_AIW;
	localparam signed [31:0] SZW = top_pkg_TL_SZW;
	reg outstanding_q;
	wire a_ack;
	wire d_ack;
	wire [RegDw - 1:0] rdata;
	reg [RegDw - 1:0] rdata_q;
	reg error_q;
	wire error;
	wire err_internal;
	wire instr_error;
	wire intg_error;
	reg addr_align_err;
	wire malformed_meta_err;
	wire tl_err;
	reg [7:0] reqid_q;
	reg [SZW - 1:0] reqsz_q;
	reg [2:0] rspop_q;
	wire rd_req;
	wire wr_req;
	assign a_ack = tl_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & tl_o[0];
	assign d_ack = tl_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] & tl_i[0];
	assign wr_req = a_ack & ((tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h0) | (tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h1));
	assign rd_req = a_ack & (tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h4);
	assign we_o = wr_req & ~err_internal;
	assign re_o = rd_req & ~err_internal;
	assign wdata_o = tl_i[55-:32];
	assign be_o = tl_i[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))];
	generate
		if (RegAw <= 2) begin : gen_only_one_reg
			assign addr_o = 1'sb0;
		end
		else begin : gen_more_regs
			assign addr_o = {tl_i[(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (32 - RegAw):(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - 29], 2'b00};
		end
	endgenerate
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			outstanding_q <= 1'b0;
		else if (a_ack)
			outstanding_q <= 1'b1;
		else if (d_ack)
			outstanding_q <= 1'b0;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			reqid_q <= 1'sb0;
			reqsz_q <= 1'sb0;
			rspop_q <= 3'h0;
		end
		else if (a_ack) begin
			reqid_q <= tl_i[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) >= (32'sd32 + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 56)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1)];
			reqsz_q <= tl_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)];
			rspop_q <= (rd_req ? 3'h1 : 3'h0);
		end
	generate
		if (AccessLatency == 1) begin : gen_access_latency1
			reg wr_req_q;
			reg rd_req_q;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni) begin
					rdata_q <= 1'sb0;
					error_q <= 1'b0;
					wr_req_q <= 1'b0;
					rd_req_q <= 1'b0;
				end
				else begin
					rd_req_q <= rd_req;
					wr_req_q <= wr_req;
					if (a_ack)
						error_q <= err_internal;
					else begin
						error_q <= error;
						rdata_q <= rdata;
					end
				end
			assign rdata = ((error_i || error_q) || wr_req_q ? {RegDw {1'sb1}} : (rd_req_q ? rdata_i : rdata_q));
			assign error = (rd_req_q || wr_req_q ? error_q || error_i : error_q);
		end
		else begin : gen_access_latency0
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni) begin
					rdata_q <= 1'sb0;
					error_q <= 1'b0;
				end
				else if (a_ack) begin
					rdata_q <= ((error_i || err_internal) || wr_req ? {RegDw {1'sb1}} : rdata_i);
					error_q <= error_i || err_internal;
				end
			assign rdata = rdata_q;
			assign error = error_q;
		end
	endgenerate
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o_pre;
	function automatic [top_pkg_TL_SZW - 1:0] sv2v_cast_9E41F;
		input reg [top_pkg_TL_SZW - 1:0] inp;
		sv2v_cast_9E41F = inp;
	endfunction
	function automatic [7:0] sv2v_cast_5359E;
		input reg [7:0] inp;
		sv2v_cast_5359E = inp;
	endfunction
	function automatic [0:0] sv2v_cast_8A6A9;
		input reg [0:0] inp;
		sv2v_cast_8A6A9 = inp;
	endfunction
	function automatic [31:0] sv2v_cast_D64A5;
		input reg [31:0] inp;
		sv2v_cast_D64A5 = inp;
	endfunction
	function automatic [(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 1:0] sv2v_cast_F43C7;
		input reg [(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 1:0] inp;
		sv2v_cast_F43C7 = inp;
	endfunction
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	assign tl_o_pre = {outstanding_q, rspop_q, 3'b000, sv2v_cast_9E41F(reqsz_q), sv2v_cast_5359E(reqid_q), sv2v_cast_8A6A9(1'sb0), sv2v_cast_D64A5(rdata), sv2v_cast_F43C7(1'sb0), error, sv2v_cast_1(~(outstanding_q | (tl_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & busy_i)))};
	tlul_rsp_intg_gen #(
		.EnableRspIntgGen(EnableRspIntgGen),
		.EnableDataIntgGen(EnableDataIntgGen)
	) u_rsp_intg_gen(
		.tl_i(tl_o_pre),
		.tl_o(tl_o)
	);
	generate
		if (CmdIntgCheck) begin : gen_cmd_intg_check
			reg intg_error_q;
			tlul_cmd_intg_chk u_cmd_intg_chk(
				.tl_i(tl_i),
				.err_o(intg_error)
			);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					intg_error_q <= 1'b0;
				else if (intg_error)
					intg_error_q <= 1'b1;
			assign intg_error_o = intg_error_q;
		end
		else begin : gen_no_cmd_intg_check
			assign intg_error = 1'b0;
			assign intg_error_o = 1'b0;
		end
	endgenerate
	function automatic [3:0] sv2v_cast_70B14;
		input reg [3:0] inp;
		sv2v_cast_70B14 = inp;
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_false_loose;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_false_loose = sv2v_cast_70B14(4'h6) != val;
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_invalid;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_invalid = ~(|{((sv2v_cast_70B14(4'h6) ^ (val ^ val)) === (val ^ (sv2v_cast_70B14(4'h6) ^ sv2v_cast_70B14(4'h6)))) & ((((val ^ val) ^ (sv2v_cast_70B14(4'h6) ^ sv2v_cast_70B14(4'h6))) === (sv2v_cast_70B14(4'h6) ^ sv2v_cast_70B14(4'h6))) | 1'bx), ((sv2v_cast_70B14(4'h9) ^ (val ^ val)) === (val ^ (sv2v_cast_70B14(4'h9) ^ sv2v_cast_70B14(4'h9)))) & ((((val ^ val) ^ (sv2v_cast_70B14(4'h9) ^ sv2v_cast_70B14(4'h9))) === (sv2v_cast_70B14(4'h9) ^ sv2v_cast_70B14(4'h9))) | 1'bx)});
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_true_strict;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_true_strict = sv2v_cast_70B14(4'h6) == val;
	endfunction
	assign instr_error = prim_mubi_pkg_mubi4_test_invalid(tl_i[18-:4]) | (prim_mubi_pkg_mubi4_test_true_strict(tl_i[18-:4]) & prim_mubi_pkg_mubi4_test_false_loose(en_ifetch_i));
	assign err_internal = (((addr_align_err | malformed_meta_err) | tl_err) | instr_error) | intg_error;
	function automatic tlul_pkg_tl_a_user_chk;
		input reg [22:0] user;
		reg malformed_err;
		reg unused_user;
		begin
			unused_user = |user;
			malformed_err = prim_mubi_pkg_mubi4_test_invalid(user[17-:4]);
			tlul_pkg_tl_a_user_chk = malformed_err;
		end
	endfunction
	assign malformed_meta_err = tlul_pkg_tl_a_user_chk(tl_i[23-:23]);
	always @(*)
		if (wr_req)
			addr_align_err = |tl_i[(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - 30:(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - 31];
		else
			addr_align_err = 1'b0;
	tlul_err u_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_i),
		.err_o(tl_err)
	);
endmodule
module tlul_adapter_sram (
	clk_i,
	rst_ni,
	tl_i,
	tl_o,
	en_ifetch_i,
	req_o,
	req_type_o,
	gnt_i,
	we_o,
	addr_o,
	wdata_o,
	wmask_o,
	intg_error_o,
	rdata_i,
	rvalid_i,
	rerror_i
);
	parameter signed [31:0] SramAw = 12;
	parameter signed [31:0] SramDw = 32;
	parameter signed [31:0] Outstanding = 1;
	parameter [0:0] ByteAccess = 1;
	parameter [0:0] ErrOnWrite = 0;
	parameter [0:0] ErrOnRead = 0;
	parameter [0:0] CmdIntgCheck = 0;
	parameter [0:0] EnableRspIntgGen = 0;
	parameter [0:0] EnableDataIntgGen = 0;
	parameter [0:0] EnableDataIntgPt = 0;
	parameter [0:0] SecFifoPtr = 0;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] WidthMult = SramDw / top_pkg_TL_DW;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] IntgWidth = tlul_pkg_DataIntgWidth * WidthMult;
	localparam signed [31:0] DataOutW = (EnableDataIntgPt ? SramDw + IntgWidth : SramDw);
	input clk_i;
	input rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_i;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	input wire [3:0] en_ifetch_i;
	output wire req_o;
	output wire [3:0] req_type_o;
	input gnt_i;
	output wire we_o;
	output wire [SramAw - 1:0] addr_o;
	output wire [DataOutW - 1:0] wdata_o;
	output wire [DataOutW - 1:0] wmask_o;
	output wire intg_error_o;
	input [DataOutW - 1:0] rdata_i;
	input rvalid_i;
	input [1:0] rerror_i;
	localparam signed [31:0] SramByte = SramDw / 8;
	function automatic integer prim_util_pkg_vbits;
		input integer value;
		prim_util_pkg_vbits = (value == 1 ? 1 : $clog2(value));
	endfunction
	localparam signed [31:0] DataBitWidth = prim_util_pkg_vbits(SramByte);
	localparam signed [31:0] WoffsetWidth = (SramByte == top_pkg_TL_DBW ? 1 : DataBitWidth - prim_util_pkg_vbits(top_pkg_TL_DBW));
	wire error_det;
	wire error_internal;
	wire wr_attr_error;
	wire instr_error;
	wire wr_vld_error;
	wire rd_vld_error;
	wire rsp_fifo_error;
	wire intg_error;
	wire tlul_error;
	generate
		if (CmdIntgCheck) begin : gen_cmd_intg_check
			tlul_cmd_intg_chk u_cmd_intg_chk(
				.tl_i(tl_i),
				.err_o(intg_error)
			);
		end
		else begin : gen_no_cmd_intg_check
			assign intg_error = 1'sb0;
		end
	endgenerate
	reg intg_error_q;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			intg_error_q <= 1'sb0;
		else if (intg_error || rsp_fifo_error)
			intg_error_q <= 1'b1;
	assign intg_error_o = (intg_error | rsp_fifo_error) | intg_error_q;
	assign wr_attr_error = ((tl_i[6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) - (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))))) + 1 : ((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) - (6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))))) + 1)] == 3'h0) || (tl_i[6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) - (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))))) + 1 : ((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) - (6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))))) + 1)] == 3'h1) ? (ByteAccess == 0 ? (tl_i[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))] != {((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55)) * 1 {1'sb1}}) || (tl_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)] != 2'h2) : 1'b0) : 1'b0);
	function automatic [3:0] sv2v_cast_84290;
		input reg [3:0] inp;
		sv2v_cast_84290 = inp;
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_false_loose;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_false_loose = sv2v_cast_84290(4'h6) != val;
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_invalid;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_invalid = ~(|{((sv2v_cast_84290(4'h6) ^ (val ^ val)) === (val ^ (sv2v_cast_84290(4'h6) ^ sv2v_cast_84290(4'h6)))) & ((((val ^ val) ^ (sv2v_cast_84290(4'h6) ^ sv2v_cast_84290(4'h6))) === (sv2v_cast_84290(4'h6) ^ sv2v_cast_84290(4'h6))) | 1'bx), ((sv2v_cast_84290(4'h9) ^ (val ^ val)) === (val ^ (sv2v_cast_84290(4'h9) ^ sv2v_cast_84290(4'h9)))) & ((((val ^ val) ^ (sv2v_cast_84290(4'h9) ^ sv2v_cast_84290(4'h9))) === (sv2v_cast_84290(4'h9) ^ sv2v_cast_84290(4'h9))) | 1'bx)});
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_true_strict;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_true_strict = sv2v_cast_84290(4'h6) == val;
	endfunction
	assign instr_error = prim_mubi_pkg_mubi4_test_invalid(tl_i[18-:4]) | (prim_mubi_pkg_mubi4_test_true_strict(tl_i[18-:4]) & prim_mubi_pkg_mubi4_test_false_loose(en_ifetch_i));
	generate
		if (ErrOnWrite == 1) begin : gen_no_writes
			assign wr_vld_error = tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] != 3'h4;
		end
		else begin : gen_writes_allowed
			assign wr_vld_error = 1'b0;
		end
		if (ErrOnRead == 1) begin : gen_no_reads
			assign rd_vld_error = tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h4;
		end
		else begin : gen_reads_allowed
			assign rd_vld_error = 1'b0;
		end
	endgenerate
	tlul_err u_err(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_i),
		.err_o(tlul_error)
	);
	assign error_det = ((((wr_attr_error | wr_vld_error) | rd_vld_error) | instr_error) | tlul_error) | intg_error;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_i_int;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o_int;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_out;
	wire unused_tl_i_int;
	assign unused_tl_i_int = ^tl_i_int;
	tlul_rsp_intg_gen #(
		.EnableRspIntgGen(EnableRspIntgGen),
		.EnableDataIntgGen(EnableDataIntgGen)
	) u_rsp_gen(
		.tl_i(tl_out),
		.tl_o(tl_o)
	);
	tlul_sram_byte #(
		.EnableIntg((ByteAccess & EnableDataIntgPt) & !ErrOnWrite),
		.Outstanding(Outstanding)
	) u_sram_byte(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_i(tl_i),
		.tl_o(tl_out),
		.tl_sram_o(tl_i_int),
		.tl_sram_i(tl_o_int),
		.error_i(error_det),
		.error_o(error_internal)
	);
	localparam signed [31:0] SramReqFifoWidth = top_pkg_TL_DBW + WoffsetWidth;
	localparam signed [31:0] ReqFifoWidth = (7 + top_pkg_TL_SZW) + top_pkg_TL_AIW;
	localparam signed [31:0] RspFifoWidth = (((top_pkg_TL_DW + tlul_pkg_DataIntgWidth) + 0) >= 0 ? (top_pkg_TL_DW + tlul_pkg_DataIntgWidth) + 1 : 1 - ((top_pkg_TL_DW + tlul_pkg_DataIntgWidth) + 0));
	wire reqfifo_wvalid;
	wire reqfifo_wready;
	wire reqfifo_rvalid;
	wire reqfifo_rready;
	wire [((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) - 1:0] reqfifo_wdata;
	wire [((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) - 1:0] reqfifo_rdata;
	wire sramreqfifo_wvalid;
	wire sramreqfifo_wready;
	wire sramreqfifo_rready;
	wire [(top_pkg_TL_DBW + WoffsetWidth) - 1:0] sramreqfifo_wdata;
	wire [(top_pkg_TL_DBW + WoffsetWidth) - 1:0] sramreqfifo_rdata;
	wire rspfifo_wvalid;
	wire rspfifo_wready;
	wire rspfifo_rvalid;
	wire rspfifo_rready;
	wire [(top_pkg_TL_DW + tlul_pkg_DataIntgWidth) + 0:0] rspfifo_wdata;
	wire [(top_pkg_TL_DW + tlul_pkg_DataIntgWidth) + 0:0] rspfifo_rdata;
	wire a_ack;
	wire d_ack;
	wire sram_ack;
	assign a_ack = tl_i_int[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & tl_o_int[0];
	assign d_ack = tl_o_int[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] & tl_i_int[0];
	assign sram_ack = req_o & gnt_i;
	reg d_valid;
	reg d_error;
	always @(*) begin
		d_valid = 1'b0;
		if (reqfifo_rvalid) begin
			if (reqfifo_rdata[1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))])
				d_valid = 1'b1;
			else if (reqfifo_rdata[3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))-:((7 + (top_pkg_TL_SZW + 7)) >= (5 + (top_pkg_TL_SZW + 8)) ? ((3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))) - (1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 8)))) + 1 : ((1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 8))) - (3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)))) + 1)] == 2'd1)
				d_valid = rspfifo_rvalid;
			else
				d_valid = 1'b1;
		end
		else
			d_valid = 1'b0;
	end
	always @(*) begin
		d_error = 1'b0;
		if (reqfifo_rvalid) begin
			if (reqfifo_rdata[3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))-:((7 + (top_pkg_TL_SZW + 7)) >= (5 + (top_pkg_TL_SZW + 8)) ? ((3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))) - (1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 8)))) + 1 : ((1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 8))) - (3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)))) + 1)] == 2'd1)
				d_error = rspfifo_rdata[0] | reqfifo_rdata[1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))];
			else
				d_error = reqfifo_rdata[1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))];
		end
		else
			d_error = 1'b0;
	end
	wire vld_rd_rsp;
	assign vld_rd_rsp = ((d_valid & reqfifo_rvalid) & rspfifo_rvalid) & (reqfifo_rdata[3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))-:((7 + (top_pkg_TL_SZW + 7)) >= (5 + (top_pkg_TL_SZW + 8)) ? ((3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))) - (1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 8)))) + 1 : ((1 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 8))) - (3 + (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)))) + 1)] == 2'd1);
	wire [31:0] error_blanking_data;
	localparam [31:0] tlul_pkg_DataWhenError = {top_pkg_TL_DW {1'b1}};
	localparam [31:0] tlul_pkg_DataWhenInstrError = 1'sb0;
	assign error_blanking_data = (prim_mubi_pkg_mubi4_test_true_strict(reqfifo_rdata[prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)-:((prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)) >= (top_pkg_TL_SZW + 8) ? ((prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)) - (top_pkg_TL_SZW + 8)) + 1 : ((top_pkg_TL_SZW + 8) - (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))) + 1)]) ? tlul_pkg_DataWhenInstrError : tlul_pkg_DataWhenError);
	wire [31:0] unused_instr;
	wire [31:0] unused_data;
	wire [6:0] error_instr_integ;
	wire [6:0] error_data_integ;
	localparam signed [31:0] tlul_pkg_DataMaxWidth = 32;
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	tlul_data_integ_enc u_tlul_data_integ_enc_instr(
		.data_i(sv2v_cast_32(tlul_pkg_DataWhenInstrError)),
		.data_intg_o({error_instr_integ, unused_instr})
	);
	tlul_data_integ_enc u_tlul_data_integ_enc_data(
		.data_i(sv2v_cast_32(tlul_pkg_DataWhenError)),
		.data_intg_o({error_data_integ, unused_data})
	);
	wire [6:0] error_blanking_integ;
	assign error_blanking_integ = (prim_mubi_pkg_mubi4_test_true_strict(reqfifo_rdata[prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)-:((prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)) >= (top_pkg_TL_SZW + 8) ? ((prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7)) - (top_pkg_TL_SZW + 8)) + 1 : ((top_pkg_TL_SZW + 8) - (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_SZW + 7))) + 1)]) ? error_instr_integ : error_data_integ);
	wire [31:0] d_data;
	assign d_data = (vld_rd_rsp & ~d_error ? rspfifo_rdata[39-:32] : error_blanking_data);
	wire [6:0] data_intg;
	localparam [6:0] prim_secded_pkg_SecdedInv3932ZeroEcc = 7'h2a;
	assign data_intg = (vld_rd_rsp && reqfifo_rdata[5 + (top_pkg_TL_SZW + 7)] ? error_blanking_integ : (vld_rd_rsp ? rspfifo_rdata[7-:7] : prim_secded_pkg_SecdedInv3932ZeroEcc));
	function automatic [6:0] sv2v_cast_360E7;
		input reg [6:0] inp;
		sv2v_cast_360E7 = inp;
	endfunction
	function automatic [top_pkg_TL_SZW - 1:0] sv2v_cast_9AB5F;
		input reg [top_pkg_TL_SZW - 1:0] inp;
		sv2v_cast_9AB5F = inp;
	endfunction
	function automatic [7:0] sv2v_cast_81C02;
		input reg [7:0] inp;
		sv2v_cast_81C02 = inp;
	endfunction
	function automatic [0:0] sv2v_cast_ACC85;
		input reg [0:0] inp;
		sv2v_cast_ACC85 = inp;
	endfunction
	function automatic [31:0] sv2v_cast_1B895;
		input reg [31:0] inp;
		sv2v_cast_1B895 = inp;
	endfunction
	function automatic [(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 1:0] sv2v_cast_42B55;
		input reg [(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 1:0] inp;
		sv2v_cast_42B55 = inp;
	endfunction
	assign tl_o_int = {d_valid, (d_valid && (reqfifo_rdata[7 + (top_pkg_TL_SZW + 7)-:((7 + (top_pkg_TL_SZW + 7)) >= (5 + (top_pkg_TL_SZW + 8)) ? ((7 + (top_pkg_TL_SZW + 7)) - (5 + (top_pkg_TL_SZW + 8))) + 1 : ((5 + (top_pkg_TL_SZW + 8)) - (7 + (top_pkg_TL_SZW + 7))) + 1)] != 2'd1) ? 3'h0 : 3'h1), 3'b000, sv2v_cast_9AB5F((d_valid ? reqfifo_rdata[top_pkg_TL_SZW + 7-:((top_pkg_TL_SZW + 7) >= 8 ? top_pkg_TL_SZW : 9 - (top_pkg_TL_SZW + 7))] : {((top_pkg_TL_SZW + 7) >= 8 ? top_pkg_TL_SZW : 9 - (top_pkg_TL_SZW + 7)) * 1 {1'sb0}})), sv2v_cast_81C02((d_valid ? reqfifo_rdata[7-:top_pkg_TL_AIW] : {8 {1'sb0}})), sv2v_cast_ACC85(1'b0), sv2v_cast_1B895(d_data), sv2v_cast_42B55({sv2v_cast_360E7(1'sb0), data_intg}), d_valid && d_error, ((gnt_i | error_internal) & reqfifo_wready) & sramreqfifo_wready};
	assign req_o = (tl_i_int[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & reqfifo_wready) & ~error_internal;
	assign req_type_o = tl_i_int[18-:4];
	assign we_o = tl_i_int[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & |{tl_i_int[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h0, tl_i_int[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h1};
	assign addr_o = (tl_i_int[7 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))] ? tl_i_int[(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (31 - DataBitWidth)+:SramAw] : {SramAw {1'sb0}});
	wire [WoffsetWidth - 1:0] woffset;
	generate
		if (top_pkg_TL_DW != SramDw) begin : gen_wordwidthadapt
			assign woffset = tl_i_int[(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (32 - DataBitWidth):(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (31 - prim_util_pkg_vbits(top_pkg_TL_DBW))];
		end
		else begin : gen_no_wordwidthadapt
			assign woffset = 1'sb0;
		end
	endgenerate
	localparam signed [31:0] DataWidth = (EnableDataIntgPt ? top_pkg_TL_DW + tlul_pkg_DataIntgWidth : top_pkg_TL_DW);
	wire [(WidthMult * DataWidth) - 1:0] wmask_combined;
	wire [(WidthMult * DataWidth) - 1:0] wdata_combined;
	reg [(WidthMult * top_pkg_TL_DW) - 1:0] wmask_int;
	reg [(WidthMult * top_pkg_TL_DW) - 1:0] wdata_int;
	reg [(WidthMult * tlul_pkg_DataIntgWidth) - 1:0] wmask_intg;
	reg [(WidthMult * tlul_pkg_DataIntgWidth) - 1:0] wdata_intg;
	always @(*) begin
		wmask_int = 1'sb0;
		wdata_int = 1'sb0;
		if (tl_i_int[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))]) begin : sv2v_autoblock_1
			reg signed [31:0] i;
			for (i = 0; i < 4; i = i + 1)
				begin
					wmask_int[(woffset * top_pkg_TL_DW) + (8 * i)+:8] = {8 {tl_i_int[(top_pkg_TL_DBW + 55) - ((top_pkg_TL_DBW - 1) - i)]}};
					wdata_int[(woffset * top_pkg_TL_DW) + (8 * i)+:8] = (tl_i_int[(top_pkg_TL_DBW + 55) - ((top_pkg_TL_DBW - 1) - i)] && we_o ? tl_i_int[24 + (8 * i)+:8] : {8 {1'sb0}});
				end
		end
	end
	always @(*) begin
		wmask_intg = 1'sb0;
		wdata_intg = 1'sb0;
		if (tl_i_int[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))]) begin
			wmask_intg[woffset * tlul_pkg_DataIntgWidth+:tlul_pkg_DataIntgWidth] = {tlul_pkg_DataIntgWidth {1'b1}};
			wdata_intg[woffset * tlul_pkg_DataIntgWidth+:tlul_pkg_DataIntgWidth] = tl_i_int[7-:tlul_pkg_DataIntgWidth];
		end
	end
	genvar i;
	generate
		for (i = 0; i < WidthMult; i = i + 1) begin : gen_write_output
			if (EnableDataIntgPt) begin : gen_combined_output
				assign wmask_combined[i * DataWidth+:DataWidth] = {wmask_intg[i * tlul_pkg_DataIntgWidth+:tlul_pkg_DataIntgWidth], wmask_int[i * top_pkg_TL_DW+:top_pkg_TL_DW]};
				assign wdata_combined[i * DataWidth+:DataWidth] = {wdata_intg[i * tlul_pkg_DataIntgWidth+:tlul_pkg_DataIntgWidth], wdata_int[i * top_pkg_TL_DW+:top_pkg_TL_DW]};
			end
			else begin : gen_ft_output
				wire unused_w;
				assign wmask_combined[i * DataWidth+:DataWidth] = wmask_int[i * top_pkg_TL_DW+:top_pkg_TL_DW];
				assign wdata_combined[i * DataWidth+:DataWidth] = wdata_int[i * top_pkg_TL_DW+:top_pkg_TL_DW];
				assign unused_w = |wmask_intg & |wdata_intg;
			end
		end
	endgenerate
	assign wmask_o = wmask_combined;
	assign wdata_o = wdata_combined;
	assign reqfifo_wvalid = a_ack;
	assign reqfifo_wdata = {(tl_i_int[6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) - (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))))) + 1 : ((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) - (6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))))) + 1)] != 3'h4 ? 2'd0 : 2'd1), error_internal, sv2v_cast_84290(tl_i_int[18-:4]), tl_i_int[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)], tl_i_int[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) >= (32'sd32 + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 56)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1)]};
	assign reqfifo_rready = d_ack;
	assign sramreqfifo_wdata = {tl_i_int[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))], woffset};
	assign sramreqfifo_wvalid = sram_ack & ~we_o;
	assign sramreqfifo_rready = rspfifo_wvalid;
	assign rspfifo_wvalid = rvalid_i & reqfifo_rvalid;
	wire [(WidthMult * DataWidth) - 1:0] rdata_reshaped;
	reg [DataWidth - 1:0] rdata_tlword;
	assign rdata_reshaped = rdata_i;
	localparam [38:0] prim_secded_pkg_SecdedInv3932ZeroWord = 39'h2a00000000;
	generate
		if (EnableDataIntgPt) begin : gen_no_rmask
			always @(*) begin
				rdata_tlword = prim_secded_pkg_SecdedInv3932ZeroWord;
				if (|sramreqfifo_rdata[top_pkg_TL_DBW + (WoffsetWidth - 1)-:((top_pkg_TL_DBW + (WoffsetWidth - 1)) >= (WoffsetWidth + 0) ? ((top_pkg_TL_DBW + (WoffsetWidth - 1)) - (WoffsetWidth + 0)) + 1 : ((WoffsetWidth + 0) - (top_pkg_TL_DBW + (WoffsetWidth - 1))) + 1)])
					rdata_tlword = rdata_reshaped[sramreqfifo_rdata[WoffsetWidth - 1-:WoffsetWidth] * DataWidth+:DataWidth];
			end
		end
		else begin : gen_rmask
			reg [DataWidth - 1:0] rmask;
			always @(*) begin
				rmask = 1'sb0;
				begin : sv2v_autoblock_2
					reg signed [31:0] i;
					for (i = 0; i < 4; i = i + 1)
						rmask[8 * i+:8] = {8 {sramreqfifo_rdata[(top_pkg_TL_DBW + (WoffsetWidth - 1)) - ((top_pkg_TL_DBW - 1) - i)]}};
				end
			end
			wire [DataWidth:1] sv2v_tmp_64F5A;
			assign sv2v_tmp_64F5A = rdata_reshaped[sramreqfifo_rdata[WoffsetWidth - 1-:WoffsetWidth] * DataWidth+:DataWidth] & rmask;
			always @(*) rdata_tlword = sv2v_tmp_64F5A;
		end
	endgenerate
	function automatic [6:0] sv2v_cast_CDF18;
		input reg [6:0] inp;
		sv2v_cast_CDF18 = inp;
	endfunction
	assign rspfifo_wdata = {sv2v_cast_1B895(rdata_tlword[31:0]), sv2v_cast_CDF18((EnableDataIntgPt ? rdata_tlword[DataWidth - 1-:tlul_pkg_DataIntgWidth] : {7 {1'sb0}})), rerror_i[1]};
	assign rspfifo_rready = ((reqfifo_rdata[7 + (top_pkg_TL_SZW + 7)-:((7 + (top_pkg_TL_SZW + 7)) >= (5 + (top_pkg_TL_SZW + 8)) ? ((7 + (top_pkg_TL_SZW + 7)) - (5 + (top_pkg_TL_SZW + 8))) + 1 : ((5 + (top_pkg_TL_SZW + 8)) - (7 + (top_pkg_TL_SZW + 7))) + 1)] == 2'd1) & ~reqfifo_rdata[5 + (top_pkg_TL_SZW + 7)] ? reqfifo_rready : 1'b0);
	wire unused_rerror;
	assign unused_rerror = rerror_i[0];
	prim_fifo_sync #(
		.Width(ReqFifoWidth),
		.Pass(1'b0),
		.Depth(Outstanding)
	) u_reqfifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(1'b0),
		.wvalid_i(reqfifo_wvalid),
		.wready_o(reqfifo_wready),
		.wdata_i(reqfifo_wdata),
		.rvalid_o(reqfifo_rvalid),
		.rready_i(reqfifo_rready),
		.rdata_o(reqfifo_rdata)
	);
	prim_fifo_sync #(
		.Width(SramReqFifoWidth),
		.Pass(1'b0),
		.Depth(Outstanding)
	) u_sramreqfifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(1'b0),
		.wvalid_i(sramreqfifo_wvalid),
		.wready_o(sramreqfifo_wready),
		.wdata_i(sramreqfifo_wdata),
		.rready_i(sramreqfifo_rready),
		.rdata_o(sramreqfifo_rdata)
	);
	prim_fifo_sync #(
		.Width(RspFifoWidth),
		.Pass(1'b1),
		.Depth(Outstanding),
		.Secure(SecFifoPtr)
	) u_rspfifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(1'b0),
		.wvalid_i(rspfifo_wvalid),
		.wready_o(rspfifo_wready),
		.wdata_i(rspfifo_wdata),
		.rvalid_o(rspfifo_rvalid),
		.rready_i(rspfifo_rready),
		.rdata_o(rspfifo_rdata),
		.err_o(rsp_fifo_error)
	);
endmodule
module tlul_assert (
	clk_i,
	rst_ni,
	h2d,
	d2h
);
	parameter EndpointType = "Device";
	input clk_i;
	input rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] h2d;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] d2h;
endmodule
module tlul_assert_multiple (
	clk_i,
	rst_ni,
	h2d,
	d2h
);
	parameter [31:0] N = 2;
	parameter EndpointType = "Device";
	input clk_i;
	input rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (N * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24)) - 1 : (N * (1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 22)):(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23)] h2d;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	input wire [((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (N * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2)) - 1 : (N * (1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1))) + ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 0)):((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1)] d2h;
	genvar ii;
	generate
		for (ii = 0; ii < N; ii = ii + 1) begin : gen_assert
			tlul_assert #(.EndpointType(EndpointType)) tlul_assert(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.h2d(h2d[(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) + (((N - 1) - ii) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23)))+:(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))]),
				.d2h(d2h[((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1) + (((N - 1) - ii) * ((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1)))+:((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1))])
			);
		end
	endgenerate
endmodule
module tlul_cmd_intg_chk (
	tl_i,
	err_o
);
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_i;
	output wire err_o;
	wire [1:0] err;
	wire data_err;
	wire [(((prim_mubi_pkg_MuBi4Width + top_pkg_TL_AW) + 3) + top_pkg_TL_DBW) - 1:0] cmd;
	function automatic [(((prim_mubi_pkg_MuBi4Width + top_pkg_TL_AW) + 3) + top_pkg_TL_DBW) - 1:0] tlul_pkg_extract_h2d_cmd_intg;
		input reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl;
		reg [(((prim_mubi_pkg_MuBi4Width + top_pkg_TL_AW) + 3) + top_pkg_TL_DBW) - 1:0] payload;
		reg unused_tlul;
		begin
			unused_tlul = ^tl;
			payload[top_pkg_TL_AW + (top_pkg_TL_DBW + 2)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 2)) >= (3 + (top_pkg_TL_DBW + 0)) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 2)) - (3 + (top_pkg_TL_DBW + 0))) + 1 : ((3 + (top_pkg_TL_DBW + 0)) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 2))) + 1)] = tl[top_pkg_TL_AW + (top_pkg_TL_DBW + 55)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)];
			payload[top_pkg_TL_DBW + 2-:((top_pkg_TL_DBW + 2) >= (top_pkg_TL_DBW + 0) ? ((top_pkg_TL_DBW + 2) - (top_pkg_TL_DBW + 0)) + 1 : ((top_pkg_TL_DBW + 0) - (top_pkg_TL_DBW + 2)) + 1)] = tl[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)];
			payload[top_pkg_TL_DBW - 1-:top_pkg_TL_DBW] = tl[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))];
			payload[prim_mubi_pkg_MuBi4Width + (top_pkg_TL_AW + (top_pkg_TL_DBW + 2))-:(((32'sd4 + 32'sd32) + (top_pkg_TL_DBW + 2)) >= (35 + (top_pkg_TL_DBW + 0)) ? ((prim_mubi_pkg_MuBi4Width + (top_pkg_TL_AW + (top_pkg_TL_DBW + 2))) - (top_pkg_TL_AW + (3 + (top_pkg_TL_DBW + 0)))) + 1 : ((top_pkg_TL_AW + (3 + (top_pkg_TL_DBW + 0))) - (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_AW + (top_pkg_TL_DBW + 2)))) + 1)] = tl[18-:4];
			tlul_pkg_extract_h2d_cmd_intg = payload;
		end
	endfunction
	assign cmd = tlul_pkg_extract_h2d_cmd_intg(tl_i);
	localparam signed [31:0] tlul_pkg_H2DCmdMaxWidth = 57;
	function automatic [56:0] sv2v_cast_57;
		input reg [56:0] inp;
		sv2v_cast_57 = inp;
	endfunction
	prim_secded_inv_64_57_dec u_chk(
		.data_i({tl_i[14-:7], sv2v_cast_57(cmd)}),
		.err_o(err)
	);
	localparam signed [31:0] tlul_pkg_DataMaxWidth = 32;
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	tlul_data_integ_dec u_tlul_data_integ_dec(
		.data_intg_i({tl_i[7-:tlul_pkg_DataIntgWidth], sv2v_cast_32(tl_i[55-:32])}),
		.data_err_o(data_err)
	);
	assign err_o = tl_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & (|err | |data_err);
	wire unused_tl;
	assign unused_tl = |tl_i;
endmodule
module tlul_cmd_intg_gen (
	tl_i,
	tl_o
);
	parameter [0:0] EnableDataIntgGen = 1'b1;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_i;
	output reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_o;
	wire [(((prim_mubi_pkg_MuBi4Width + top_pkg_TL_AW) + 3) + top_pkg_TL_DBW) - 1:0] cmd;
	function automatic [(((prim_mubi_pkg_MuBi4Width + top_pkg_TL_AW) + 3) + top_pkg_TL_DBW) - 1:0] tlul_pkg_extract_h2d_cmd_intg;
		input reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl;
		reg [(((prim_mubi_pkg_MuBi4Width + top_pkg_TL_AW) + 3) + top_pkg_TL_DBW) - 1:0] payload;
		reg unused_tlul;
		begin
			unused_tlul = ^tl;
			payload[top_pkg_TL_AW + (top_pkg_TL_DBW + 2)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 2)) >= (3 + (top_pkg_TL_DBW + 0)) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 2)) - (3 + (top_pkg_TL_DBW + 0))) + 1 : ((3 + (top_pkg_TL_DBW + 0)) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 2))) + 1)] = tl[top_pkg_TL_AW + (top_pkg_TL_DBW + 55)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)];
			payload[top_pkg_TL_DBW + 2-:((top_pkg_TL_DBW + 2) >= (top_pkg_TL_DBW + 0) ? ((top_pkg_TL_DBW + 2) - (top_pkg_TL_DBW + 0)) + 1 : ((top_pkg_TL_DBW + 0) - (top_pkg_TL_DBW + 2)) + 1)] = tl[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)];
			payload[top_pkg_TL_DBW - 1-:top_pkg_TL_DBW] = tl[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))];
			payload[prim_mubi_pkg_MuBi4Width + (top_pkg_TL_AW + (top_pkg_TL_DBW + 2))-:(((32'sd4 + 32'sd32) + (top_pkg_TL_DBW + 2)) >= (35 + (top_pkg_TL_DBW + 0)) ? ((prim_mubi_pkg_MuBi4Width + (top_pkg_TL_AW + (top_pkg_TL_DBW + 2))) - (top_pkg_TL_AW + (3 + (top_pkg_TL_DBW + 0)))) + 1 : ((top_pkg_TL_AW + (3 + (top_pkg_TL_DBW + 0))) - (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_AW + (top_pkg_TL_DBW + 2)))) + 1)] = tl[18-:4];
			tlul_pkg_extract_h2d_cmd_intg = payload;
		end
	endfunction
	assign cmd = tlul_pkg_extract_h2d_cmd_intg(tl_i);
	localparam signed [31:0] tlul_pkg_H2DCmdMaxWidth = 57;
	wire [56:0] unused_cmd_payload;
	wire [6:0] cmd_intg;
	function automatic [56:0] sv2v_cast_57;
		input reg [56:0] inp;
		sv2v_cast_57 = inp;
	endfunction
	prim_secded_inv_64_57_enc u_cmd_gen(
		.data_i(sv2v_cast_57(cmd)),
		.data_o({cmd_intg, unused_cmd_payload})
	);
	wire [31:0] data_final;
	wire [6:0] data_intg;
	localparam signed [31:0] tlul_pkg_DataMaxWidth = 32;
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	generate
		if (EnableDataIntgGen) begin : gen_data_intg
			assign data_final = tl_i[55-:32];
			wire [31:0] unused_data;
			prim_secded_inv_39_32_enc u_data_gen(
				.data_i(sv2v_cast_32(data_final)),
				.data_o({data_intg, unused_data})
			);
		end
		else begin : gen_passthrough_data_intg
			assign data_final = tl_i[55-:32];
			assign data_intg = tl_i[7-:tlul_pkg_DataIntgWidth];
		end
	endgenerate
	always @(*) begin
		tl_o = tl_i;
		tl_o[55-:32] = data_final;
		tl_o[14-:7] = cmd_intg;
		tl_o[7-:tlul_pkg_DataIntgWidth] = data_intg;
	end
	wire unused_tl;
	assign unused_tl = ^tl_i;
endmodule
module tlul_data_integ_dec (
	data_intg_i,
	data_err_o
);
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_DataMaxWidth = 32;
	input [(tlul_pkg_DataMaxWidth + tlul_pkg_DataIntgWidth) - 1:0] data_intg_i;
	output wire data_err_o;
	wire [1:0] data_err;
	prim_secded_inv_39_32_dec u_data_chk(
		.data_i(data_intg_i),
		.err_o(data_err)
	);
	assign data_err_o = |data_err;
endmodule
module tlul_data_integ_enc (
	data_i,
	data_intg_o
);
	localparam signed [31:0] tlul_pkg_DataMaxWidth = 32;
	input [31:0] data_i;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	output wire [(tlul_pkg_DataMaxWidth + tlul_pkg_DataIntgWidth) - 1:0] data_intg_o;
	prim_secded_inv_39_32_enc u_data_gen(
		.data_i(data_i),
		.data_o(data_intg_o)
	);
endmodule
module tlul_err (
	clk_i,
	rst_ni,
	tl_i,
	err_o
);
	input clk_i;
	input rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_i;
	output wire err_o;
	localparam signed [31:0] IW = top_pkg_TL_AIW;
	localparam signed [31:0] SZW = top_pkg_TL_SZW;
	localparam signed [31:0] DW = top_pkg_TL_DW;
	localparam signed [31:0] MW = top_pkg_TL_DBW;
	localparam signed [31:0] SubAW = 2;
	wire opcode_allowed;
	wire a_config_allowed;
	wire op_full;
	wire op_partial;
	wire op_get;
	assign op_full = tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h0;
	assign op_partial = tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h1;
	assign op_get = tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h4;
	wire instr_wr_err;
	function automatic [3:0] sv2v_cast_D5347;
		input reg [3:0] inp;
		sv2v_cast_D5347 = inp;
	endfunction
	function automatic prim_mubi_pkg_mubi4_test_true_strict;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_true_strict = sv2v_cast_D5347(4'h6) == val;
	endfunction
	assign instr_wr_err = prim_mubi_pkg_mubi4_test_true_strict(tl_i[18-:4]) & (op_full | op_partial);
	wire instr_type_err;
	function automatic prim_mubi_pkg_mubi4_test_invalid;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_invalid = ~(|{((sv2v_cast_D5347(4'h6) ^ (val ^ val)) === (val ^ (sv2v_cast_D5347(4'h6) ^ sv2v_cast_D5347(4'h6)))) & ((((val ^ val) ^ (sv2v_cast_D5347(4'h6) ^ sv2v_cast_D5347(4'h6))) === (sv2v_cast_D5347(4'h6) ^ sv2v_cast_D5347(4'h6))) | 1'bx), ((sv2v_cast_D5347(4'h9) ^ (val ^ val)) === (val ^ (sv2v_cast_D5347(4'h9) ^ sv2v_cast_D5347(4'h9)))) & ((((val ^ val) ^ (sv2v_cast_D5347(4'h9) ^ sv2v_cast_D5347(4'h9))) === (sv2v_cast_D5347(4'h9) ^ sv2v_cast_D5347(4'h9))) | 1'bx)});
	endfunction
	assign instr_type_err = prim_mubi_pkg_mubi4_test_invalid(tl_i[18-:4]);
	assign err_o = (~(opcode_allowed & a_config_allowed) | instr_wr_err) | instr_type_err;
	assign opcode_allowed = ((tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h0) | (tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h1)) | (tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h4);
	reg addr_sz_chk;
	reg mask_chk;
	reg fulldata_chk;
	wire [MW - 1:0] mask;
	assign mask = 1 << tl_i[(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - 30:(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - 31];
	always @(*) begin
		addr_sz_chk = 1'b0;
		mask_chk = 1'b0;
		fulldata_chk = 1'b0;
		if (tl_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))])
			case (tl_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)])
				'h0: begin
					addr_sz_chk = 1'b1;
					mask_chk = ~|(tl_i[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))] & ~mask);
					fulldata_chk = |(tl_i[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))] & mask);
				end
				'h1: begin
					addr_sz_chk = ~tl_i[(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - 31];
					mask_chk = (tl_i[(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - 30] ? ~|(tl_i[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))] & 4'b0011) : ~|(tl_i[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))] & 4'b1100));
					fulldata_chk = (tl_i[(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - 30] ? &tl_i[(top_pkg_TL_DBW + 55) - (top_pkg_TL_DBW - 4):(top_pkg_TL_DBW + 55) - (top_pkg_TL_DBW - 3)] : &tl_i[(top_pkg_TL_DBW + 55) - (top_pkg_TL_DBW - 2):(top_pkg_TL_DBW + 55) - (top_pkg_TL_DBW - 1)]);
				end
				'h2: begin
					addr_sz_chk = ~|tl_i[(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - 30:(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - 31];
					mask_chk = 1'b1;
					fulldata_chk = &tl_i[(top_pkg_TL_DBW + 55) - (top_pkg_TL_DBW - 4):(top_pkg_TL_DBW + 55) - (top_pkg_TL_DBW - 1)];
				end
				default: begin
					addr_sz_chk = 1'b0;
					mask_chk = 1'b0;
					fulldata_chk = 1'b0;
				end
			endcase
		else begin
			addr_sz_chk = 1'b0;
			mask_chk = 1'b0;
			fulldata_chk = 1'b0;
		end
	end
	assign a_config_allowed = (addr_sz_chk & mask_chk) & ((op_get | op_partial) | fulldata_chk);
endmodule
module tlul_err_resp (
	clk_i,
	rst_ni,
	tl_h_i,
	tl_h_o
);
	input clk_i;
	input rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_h_i;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_h_o;
	reg [2:0] err_opcode;
	reg [7:0] err_source;
	reg [top_pkg_TL_SZW - 1:0] err_size;
	reg err_req_pending;
	reg err_rsp_pending;
	reg [3:0] err_instr_type;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_h_o_int;
	tlul_rsp_intg_gen #(
		.EnableRspIntgGen(1),
		.EnableDataIntgGen(1)
	) u_intg_gen(
		.tl_i(tl_h_o_int),
		.tl_o(tl_h_o)
	);
	function automatic [3:0] sv2v_cast_210BB;
		input reg [3:0] inp;
		sv2v_cast_210BB = inp;
	endfunction
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			err_req_pending <= 1'b0;
			err_source <= {top_pkg_TL_AIW {1'b0}};
			err_opcode <= 3'h4;
			err_size <= 1'sb0;
			err_instr_type <= sv2v_cast_210BB(4'h9);
		end
		else if (tl_h_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] && tl_h_o_int[0]) begin
			err_req_pending <= 1'b1;
			err_source <= tl_h_i[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) >= (32'sd32 + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 56)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1)];
			err_opcode <= tl_h_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)];
			err_size <= tl_h_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)];
			err_instr_type <= tl_h_i[18-:4];
		end
		else if (!err_rsp_pending)
			err_req_pending <= 1'b0;
	assign tl_h_o_int[0] = ~err_rsp_pending & ~(err_req_pending & ~tl_h_i[0]);
	assign tl_h_o_int[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] = err_req_pending | err_rsp_pending;
	function automatic prim_mubi_pkg_mubi4_test_true_strict;
		input reg [3:0] val;
		prim_mubi_pkg_mubi4_test_true_strict = sv2v_cast_210BB(4'h6) == val;
	endfunction
	localparam [31:0] tlul_pkg_DataWhenError = {top_pkg_TL_DW {1'b1}};
	localparam [31:0] tlul_pkg_DataWhenInstrError = 1'sb0;
	assign tl_h_o_int[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)] = (prim_mubi_pkg_mubi4_test_true_strict(err_instr_type) ? tlul_pkg_DataWhenInstrError : tlul_pkg_DataWhenError);
	assign tl_h_o_int[top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))-:((32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))) >= ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) + 1 : ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) + 1)] = err_source;
	assign tl_h_o_int[top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))-:(((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)) >= (32'sd32 + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) + 1 : ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) + 1)] = 1'sb0;
	assign tl_h_o_int[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)] = 1'sb0;
	assign tl_h_o_int[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)] = err_size;
	assign tl_h_o_int[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)] = (err_opcode == 3'h4 ? 3'h1 : 3'h0);
	assign tl_h_o_int[(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1-:(((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) >= 2 ? (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 0 : 3 - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))] = 1'sb0;
	assign tl_h_o_int[1] = 1'b1;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			err_rsp_pending <= 1'b0;
		else if ((err_req_pending || err_rsp_pending) && !tl_h_i[0])
			err_rsp_pending <= 1'b1;
		else
			err_rsp_pending <= 1'b0;
	wire unused_tl_h;
	assign unused_tl_h = ^tl_h_i;
endmodule
module tlul_fifo_async (
	clk_h_i,
	rst_h_ni,
	clk_d_i,
	rst_d_ni,
	tl_h_i,
	tl_h_o,
	tl_d_o,
	tl_d_i
);
	parameter [31:0] ReqDepth = 3;
	parameter [31:0] RspDepth = 3;
	input clk_h_i;
	input rst_h_ni;
	input clk_d_i;
	input rst_d_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_h_i;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_h_o;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_d_o;
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_d_i;
	localparam [31:0] REQFIFO_WIDTH = (1 * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24)) - 2;
	prim_fifo_async #(
		.Width(REQFIFO_WIDTH),
		.Depth(ReqDepth),
		.OutputZeroIfInvalid(1)
	) reqfifo(
		.clk_wr_i(clk_h_i),
		.rst_wr_ni(rst_h_ni),
		.clk_rd_i(clk_d_i),
		.rst_rd_ni(rst_d_ni),
		.wvalid_i(tl_h_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))]),
		.wready_o(tl_h_o[0]),
		.wdata_i({tl_h_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)], tl_h_i[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)], tl_h_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)], tl_h_i[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) >= (32'sd32 + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 56)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1)], tl_h_i[top_pkg_TL_AW + (top_pkg_TL_DBW + 55)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)], tl_h_i[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))], tl_h_i[55-:32], tl_h_i[23-:23]}),
		.rvalid_o(tl_d_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))]),
		.rready_i(tl_d_i[0]),
		.rdata_o({tl_d_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)], tl_d_o[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)], tl_d_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)], tl_d_o[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) >= (32'sd32 + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 56)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1)], tl_d_o[top_pkg_TL_AW + (top_pkg_TL_DBW + 55)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)], tl_d_o[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))], tl_d_o[55-:32], tl_d_o[23-:23]})
	);
	localparam [31:0] RSPFIFO_WIDTH = (1 * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2)) - 2;
	prim_fifo_async #(
		.Width(RSPFIFO_WIDTH),
		.Depth(RspDepth),
		.OutputZeroIfInvalid(1)
	) rspfifo(
		.clk_wr_i(clk_d_i),
		.rst_wr_ni(rst_d_ni),
		.clk_rd_i(clk_h_i),
		.rst_rd_ni(rst_h_ni),
		.wvalid_i(tl_d_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))]),
		.wready_o(tl_d_o[0]),
		.wdata_i({tl_d_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)], tl_d_i[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)], tl_d_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)], tl_d_i[top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))-:((32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))) >= ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) + 1 : ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) + 1)], tl_d_i[top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))-:(((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)) >= (32'sd32 + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) + 1 : ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) + 1)], tl_d_i[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)], tl_d_i[(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1-:(((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) >= 2 ? (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 0 : 3 - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))], tl_d_i[1]}),
		.rvalid_o(tl_h_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))]),
		.rready_i(tl_h_i[0]),
		.rdata_o({tl_h_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)], tl_h_o[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)], tl_h_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)], tl_h_o[top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))-:((32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))) >= ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) + 1 : ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) + 1)], tl_h_o[top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))-:(((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)) >= (32'sd32 + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) + 1 : ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) + 1)], tl_h_o[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)], tl_h_o[(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1-:(((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) >= 2 ? (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 0 : 3 - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))], tl_h_o[1]})
	);
endmodule
module tlul_fifo_sync (
	clk_i,
	rst_ni,
	tl_h_i,
	tl_h_o,
	tl_d_o,
	tl_d_i,
	spare_req_i,
	spare_req_o,
	spare_rsp_i,
	spare_rsp_o
);
	parameter [0:0] ReqPass = 1'b1;
	parameter [0:0] RspPass = 1'b1;
	parameter [31:0] ReqDepth = 2;
	parameter [31:0] RspDepth = 2;
	parameter [31:0] SpareReqW = 1;
	parameter [31:0] SpareRspW = 1;
	input clk_i;
	input rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_h_i;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_h_o;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_d_o;
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_d_i;
	input [SpareReqW - 1:0] spare_req_i;
	output wire [SpareReqW - 1:0] spare_req_o;
	input [SpareRspW - 1:0] spare_rsp_i;
	output wire [SpareRspW - 1:0] spare_rsp_o;
	localparam [31:0] REQFIFO_WIDTH = ((1 * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24)) - 2) + SpareReqW;
	prim_fifo_sync #(
		.Width(REQFIFO_WIDTH),
		.Pass(ReqPass),
		.Depth(ReqDepth)
	) reqfifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(1'b0),
		.wvalid_i(tl_h_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))]),
		.wready_o(tl_h_o[0]),
		.wdata_i({tl_h_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)], tl_h_i[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)], tl_h_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)], tl_h_i[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) >= (32'sd32 + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 56)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1)], tl_h_i[top_pkg_TL_AW + (top_pkg_TL_DBW + 55)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)], tl_h_i[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))], tl_h_i[55-:32], tl_h_i[23-:23], spare_req_i}),
		.rvalid_o(tl_d_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))]),
		.rready_i(tl_d_i[0]),
		.rdata_o({tl_d_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)], tl_d_o[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)], tl_d_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)], tl_d_o[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) >= (32'sd32 + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 56)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1)], tl_d_o[top_pkg_TL_AW + (top_pkg_TL_DBW + 55)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)], tl_d_o[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))], tl_d_o[55-:32], tl_d_o[23-:23], spare_req_o})
	);
	localparam [31:0] RSPFIFO_WIDTH = ((1 * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2)) - 2) + SpareRspW;
	prim_fifo_sync #(
		.Width(RSPFIFO_WIDTH),
		.Pass(RspPass),
		.Depth(RspDepth)
	) rspfifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_i(1'b0),
		.wvalid_i(tl_d_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))]),
		.wready_o(tl_d_o[0]),
		.wdata_i({tl_d_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)], tl_d_i[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)], tl_d_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)], tl_d_i[top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))-:((32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))) >= ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) + 1 : ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) + 1)], tl_d_i[top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))-:(((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)) >= (32'sd32 + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) + 1 : ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) + 1)], (tl_d_i[6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) - (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))))) + 1 : ((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) - (6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))))) + 1)] == 3'h1 ? tl_d_i[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)] : {top_pkg_TL_DW {1'b0}}), tl_d_i[(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1-:(((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) >= 2 ? (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 0 : 3 - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))], tl_d_i[1], spare_rsp_i}),
		.rvalid_o(tl_h_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))]),
		.rready_i(tl_h_i[0]),
		.rdata_o({tl_h_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)], tl_h_o[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)], tl_h_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)], tl_h_o[top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))-:((32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))) >= ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) + 1 : ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) + 1)], tl_h_o[top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))-:(((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)) >= (32'sd32 + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) + 1 : ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) + 1)], tl_h_o[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)], tl_h_o[(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1-:(((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) >= 2 ? (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 0 : 3 - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))], tl_h_o[1], spare_rsp_o})
	);
endmodule
module tlul_lc_gate (
	clk_i,
	rst_ni,
	tl_h2d_i,
	tl_d2h_o,
	tl_h2d_o,
	tl_d2h_i,
	flush_req_i,
	flush_ack_o,
	resp_pending_o,
	lc_en_i,
	err_o
);
	parameter signed [31:0] NumGatesPerDirection = 2;
	input clk_i;
	input rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_h2d_i;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	output reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_d2h_o;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_h2d_o;
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_d2h_i;
	input flush_req_i;
	output reg flush_ack_o;
	output reg resp_pending_o;
	localparam signed [31:0] lc_ctrl_pkg_TxWidth = 4;
	input wire [3:0] lc_en_i;
	output reg err_o;
	reg [3:0] err_en;
	wire [(NumGatesPerDirection * lc_ctrl_pkg_TxWidth) - 1:0] err_en_buf;
	prim_lc_sync #(
		.NumCopies(NumGatesPerDirection),
		.AsyncOn(0)
	) u_err_en_sync(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.lc_en_i(err_en),
		.lc_en_o(err_en_buf)
	);
	reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_h2d_int [0:NumGatesPerDirection + 0];
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_d2h_int [0:NumGatesPerDirection + 0];
	genvar k;
	function automatic [3:0] sv2v_cast_4BF1C;
		input reg [3:0] inp;
		sv2v_cast_4BF1C = inp;
	endfunction
	function automatic lc_ctrl_pkg_lc_tx_test_false_strict;
		input reg [3:0] val;
		lc_ctrl_pkg_lc_tx_test_false_strict = sv2v_cast_4BF1C(4'b1010) == val;
	endfunction
	generate
		for (k = 0; k < NumGatesPerDirection; k = k + 1) begin : gen_lc_gating_muxes
			wire [(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23)):1] sv2v_tmp_u_prim_blanker_h2d_out_o;
			always @(*) tl_h2d_int[k + 1] = sv2v_tmp_u_prim_blanker_h2d_out_o;
			prim_blanker #(.Width(1 * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24))) u_prim_blanker_h2d(
				.in_i(tl_h2d_int[k]),
				.en_i(lc_ctrl_pkg_lc_tx_test_false_strict(err_en_buf[k * lc_ctrl_pkg_TxWidth+:lc_ctrl_pkg_TxWidth])),
				.out_o(sv2v_tmp_u_prim_blanker_h2d_out_o)
			);
			prim_blanker #(.Width(1 * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2))) u_prim_blanker_d2h(
				.in_i(tl_d2h_int[k + 1]),
				.en_i(lc_ctrl_pkg_lc_tx_test_false_strict(err_en_buf[k * lc_ctrl_pkg_TxWidth+:lc_ctrl_pkg_TxWidth])),
				.out_o(tl_d2h_int[k])
			);
		end
	endgenerate
	assign tl_h2d_o = tl_h2d_int[NumGatesPerDirection];
	assign tl_d2h_int[NumGatesPerDirection] = tl_d2h_i;
	localparam signed [31:0] StateWidth = 9;
	reg [8:0] state_d;
	wire [8:0] state_q;
	function automatic [8:0] sv2v_cast_84C2F;
		input reg [8:0] inp;
		sv2v_cast_84C2F = inp;
	endfunction
	prim_sparse_fsm_flop_378FE_346F8 #(
		.StateEnumT_StateWidth(StateWidth),
		.Width(StateWidth),
		.ResetValue(sv2v_cast_84C2F(9'b010111010)),
		.EnableAlertTriggerSVA(1)
	) u_state_regs(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.state_i(state_d),
		.state_o(state_q)
	);
	reg [1:0] outstanding_txn;
	wire a_ack;
	wire d_ack;
	assign a_ack = tl_h2d_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & tl_d2h_o[0];
	assign d_ack = tl_h2d_i[0] & tl_d2h_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))];
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			outstanding_txn <= 1'sb0;
		else if (a_ack && !d_ack)
			outstanding_txn <= outstanding_txn + 1'b1;
		else if (d_ack && !a_ack)
			outstanding_txn <= outstanding_txn - 1'b1;
	reg block_cmd;
	function automatic lc_ctrl_pkg_lc_tx_test_false_loose;
		input reg [3:0] val;
		lc_ctrl_pkg_lc_tx_test_false_loose = sv2v_cast_4BF1C(4'b0101) != val;
	endfunction
	function automatic lc_ctrl_pkg_lc_tx_test_true_strict;
		input reg [3:0] val;
		lc_ctrl_pkg_lc_tx_test_true_strict = sv2v_cast_4BF1C(4'b0101) == val;
	endfunction
	always @(*) begin
		block_cmd = 1'sb0;
		state_d = state_q;
		err_en = sv2v_cast_4BF1C(4'b1010);
		err_o = 1'sb0;
		flush_ack_o = 1'sb0;
		resp_pending_o = 1'b0;
		case (state_q)
			sv2v_cast_84C2F(9'b100100001): begin
				if (lc_ctrl_pkg_lc_tx_test_false_loose(lc_en_i) || flush_req_i)
					state_d = sv2v_cast_84C2F(9'b011100111);
				if (outstanding_txn != {2 {1'sb0}})
					resp_pending_o = 1'b1;
			end
			sv2v_cast_84C2F(9'b011100111): begin
				block_cmd = 1'b1;
				if (outstanding_txn == {2 {1'sb0}})
					state_d = (lc_ctrl_pkg_lc_tx_test_false_loose(lc_en_i) ? sv2v_cast_84C2F(9'b010111010) : sv2v_cast_84C2F(9'b001001100));
				else
					resp_pending_o = 1'b1;
			end
			sv2v_cast_84C2F(9'b001001100): begin
				block_cmd = 1'b1;
				flush_ack_o = 1'b1;
				if (lc_ctrl_pkg_lc_tx_test_false_loose(lc_en_i))
					state_d = sv2v_cast_84C2F(9'b010111010);
				else if (!flush_req_i)
					state_d = sv2v_cast_84C2F(9'b100100001);
			end
			sv2v_cast_84C2F(9'b010111010): begin
				err_en = sv2v_cast_4BF1C(4'b0101);
				if (lc_ctrl_pkg_lc_tx_test_true_strict(lc_en_i))
					state_d = sv2v_cast_84C2F(9'b100010110);
			end
			sv2v_cast_84C2F(9'b100010110): begin
				err_en = sv2v_cast_4BF1C(4'b0101);
				block_cmd = 1'b1;
				if (outstanding_txn == {2 {1'sb0}})
					state_d = sv2v_cast_84C2F(9'b100100001);
			end
			default: begin
				err_o = 1'b1;
				err_en = sv2v_cast_4BF1C(4'b0101);
			end
		endcase
	end
	reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_h2d_error;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_d2h_error;
	function automatic lc_ctrl_pkg_lc_tx_test_true_loose;
		input reg [3:0] val;
		lc_ctrl_pkg_lc_tx_test_true_loose = sv2v_cast_4BF1C(4'b1010) != val;
	endfunction
	always @(*) begin
		tl_h2d_int[0] = tl_h2d_i;
		tl_d2h_o = tl_d2h_int[0];
		tl_h2d_error = 1'sb0;
		if (lc_ctrl_pkg_lc_tx_test_true_loose(err_en)) begin
			tl_h2d_error = tl_h2d_i;
			tl_d2h_o = tl_d2h_error;
		end
		if (block_cmd) begin
			tl_d2h_o[0] = 1'b0;
			tl_h2d_int[0][7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] = 1'b0;
			tl_h2d_error[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] = 1'b0;
		end
	end
	tlul_err_resp u_tlul_err_resp(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_h_i(tl_h2d_error),
		.tl_h_o(tl_d2h_error)
	);
endmodule
module tlul_rsp_intg_chk (
	tl_i,
	err_o
);
	parameter [0:0] EnableRspDataIntgCheck = 0;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_i;
	output wire err_o;
	wire [1:0] rsp_err;
	wire [(3 + top_pkg_TL_SZW) + 0:0] rsp;
	function automatic [(3 + top_pkg_TL_SZW) + 0:0] tlul_pkg_extract_d2h_rsp_intg;
		input reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl;
		reg [(3 + top_pkg_TL_SZW) + 0:0] payload;
		reg unused_tlul;
		begin
			unused_tlul = ^tl;
			payload[3 + (top_pkg_TL_SZW + 0)-:((3 + (top_pkg_TL_SZW + 0)) >= (top_pkg_TL_SZW + 1) ? ((3 + (top_pkg_TL_SZW + 0)) - (top_pkg_TL_SZW + 1)) + 1 : ((top_pkg_TL_SZW + 1) - (3 + (top_pkg_TL_SZW + 0))) + 1)] = tl[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)];
			payload[top_pkg_TL_SZW + 0-:((top_pkg_TL_SZW + 0) >= 1 ? top_pkg_TL_SZW + 0 : 2 - (top_pkg_TL_SZW + 0))] = tl[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)];
			payload[0] = tl[1];
			tlul_pkg_extract_d2h_rsp_intg = payload;
		end
	endfunction
	assign rsp = tlul_pkg_extract_d2h_rsp_intg(tl_i);
	localparam signed [31:0] tlul_pkg_D2HRspMaxWidth = 57;
	function automatic [56:0] sv2v_cast_57;
		input reg [56:0] inp;
		sv2v_cast_57 = inp;
	endfunction
	prim_secded_inv_64_57_dec u_chk(
		.data_i({tl_i[((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 14)-:7], sv2v_cast_57(rsp)}),
		.err_o(rsp_err)
	);
	wire rsp_data_err;
	localparam signed [31:0] tlul_pkg_DataMaxWidth = 32;
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	generate
		if (EnableRspDataIntgCheck) begin : gen_rsp_data_intg_check
			tlul_data_integ_dec u_tlul_data_integ_dec(
				.data_intg_i({tl_i[((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 7)-:tlul_pkg_DataIntgWidth], sv2v_cast_32(tl_i[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)])}),
				.data_err_o(rsp_data_err)
			);
		end
		else begin : gen_no_rsp_data_intg_check
			assign rsp_data_err = 1'b0;
		end
	endgenerate
	assign err_o = tl_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] & (|rsp_err | rsp_data_err);
	wire unused_tl;
	assign unused_tl = |tl_i;
endmodule
module tlul_rsp_intg_gen (
	tl_i,
	tl_o
);
	parameter [0:0] EnableRspIntgGen = 1'b1;
	parameter [0:0] EnableDataIntgGen = 1'b1;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_i;
	output reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	wire [6:0] rsp_intg;
	localparam signed [31:0] tlul_pkg_D2HRspMaxWidth = 57;
	function automatic [(3 + top_pkg_TL_SZW) + 0:0] tlul_pkg_extract_d2h_rsp_intg;
		input reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl;
		reg [(3 + top_pkg_TL_SZW) + 0:0] payload;
		reg unused_tlul;
		begin
			unused_tlul = ^tl;
			payload[3 + (top_pkg_TL_SZW + 0)-:((3 + (top_pkg_TL_SZW + 0)) >= (top_pkg_TL_SZW + 1) ? ((3 + (top_pkg_TL_SZW + 0)) - (top_pkg_TL_SZW + 1)) + 1 : ((top_pkg_TL_SZW + 1) - (3 + (top_pkg_TL_SZW + 0))) + 1)] = tl[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)];
			payload[top_pkg_TL_SZW + 0-:((top_pkg_TL_SZW + 0) >= 1 ? top_pkg_TL_SZW + 0 : 2 - (top_pkg_TL_SZW + 0))] = tl[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)];
			payload[0] = tl[1];
			tlul_pkg_extract_d2h_rsp_intg = payload;
		end
	endfunction
	function automatic [56:0] sv2v_cast_57;
		input reg [56:0] inp;
		sv2v_cast_57 = inp;
	endfunction
	generate
		if (EnableRspIntgGen) begin : gen_rsp_intg
			wire [(3 + top_pkg_TL_SZW) + 0:0] rsp;
			wire [56:0] unused_payload;
			assign rsp = tlul_pkg_extract_d2h_rsp_intg(tl_i);
			prim_secded_inv_64_57_enc u_rsp_gen(
				.data_i(sv2v_cast_57(rsp)),
				.data_o({rsp_intg, unused_payload})
			);
		end
		else begin : gen_passthrough_rsp_intg
			assign rsp_intg = tl_i[((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 14)-:7];
		end
	endgenerate
	wire [6:0] data_intg;
	localparam signed [31:0] tlul_pkg_DataMaxWidth = 32;
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	generate
		if (EnableDataIntgGen) begin : gen_data_intg
			wire [31:0] unused_data;
			tlul_data_integ_enc u_tlul_data_integ_enc(
				.data_i(sv2v_cast_32(tl_i[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)])),
				.data_intg_o({data_intg, unused_data})
			);
		end
		else begin : gen_passthrough_data_intg
			assign data_intg = tl_i[((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 7)-:tlul_pkg_DataIntgWidth];
		end
	endgenerate
	always @(*) begin
		tl_o = tl_i;
		tl_o[((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 14)-:7] = rsp_intg;
		tl_o[((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 7)-:tlul_pkg_DataIntgWidth] = data_intg;
	end
	wire unused_tl;
	assign unused_tl = ^tl_i;
endmodule
module tlul_socket_1n (
	clk_i,
	rst_ni,
	tl_h_i,
	tl_h_o,
	tl_d_o,
	tl_d_i,
	dev_select_i
);
	parameter [31:0] N = 4;
	parameter [0:0] HReqPass = 1'b1;
	parameter [0:0] HRspPass = 1'b1;
	parameter [N - 1:0] DReqPass = {N {1'b1}};
	parameter [N - 1:0] DRspPass = {N {1'b1}};
	parameter [3:0] HReqDepth = 4'h1;
	parameter [3:0] HRspDepth = 4'h1;
	parameter [(N * 4) - 1:0] DReqDepth = {N {4'h1}};
	parameter [(N * 4) - 1:0] DRspDepth = {N {4'h1}};
	parameter [0:0] ExplicitErrs = 1'b1;
	localparam [31:0] NWD = $clog2((ExplicitErrs ? N + 1 : N));
	input clk_i;
	input rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_h_i;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_h_o;
	output wire [(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (N * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24)) - 1 : (N * (1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 22)):(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23)] tl_d_o;
	input wire [((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (N * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2)) - 1 : (N * (1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1))) + ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 0)):((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1)] tl_d_i;
	input [NWD - 1:0] dev_select_i;
	wire [NWD - 1:0] dev_select_t;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_t_o;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_t_i;
	tlul_fifo_sync #(
		.ReqPass(HReqPass),
		.RspPass(HRspPass),
		.ReqDepth(HReqDepth),
		.RspDepth(HRspDepth),
		.SpareReqW(NWD)
	) fifo_h(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_h_i(tl_h_i),
		.tl_h_o(tl_h_o),
		.tl_d_o(tl_t_o),
		.tl_d_i(tl_t_i),
		.spare_req_i(dev_select_i),
		.spare_req_o(dev_select_t),
		.spare_rsp_i(1'b0)
	);
	localparam signed [31:0] MaxOutstanding = 256;
	localparam signed [31:0] OutstandingW = 9;
	reg [8:0] num_req_outstanding;
	reg [NWD - 1:0] dev_select_outstanding;
	wire hold_all_requests;
	wire accept_t_req;
	wire accept_t_rsp;
	assign accept_t_req = tl_t_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & tl_t_i[0];
	assign accept_t_rsp = tl_t_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] & tl_t_o[0];
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			num_req_outstanding <= 1'sb0;
			dev_select_outstanding <= 1'sb0;
		end
		else if (accept_t_req) begin
			if (!accept_t_rsp)
				num_req_outstanding <= num_req_outstanding + 1'b1;
			dev_select_outstanding <= dev_select_t;
		end
		else if (accept_t_rsp)
			num_req_outstanding <= num_req_outstanding - 1'b1;
	assign hold_all_requests = (num_req_outstanding != {9 {1'sb0}}) & (dev_select_t != dev_select_outstanding);
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_u_o [0:N + 0];
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_u_i [0:N + 0];
	wire [22:0] blanked_auser;
	localparam [31:0] tlul_pkg_BlankedAData = {top_pkg_TL_DW {1'b1}};
	function automatic [63:0] sv2v_cast_64;
		input reg [63:0] inp;
		sv2v_cast_64 = inp;
	endfunction
	function automatic [63:0] prim_secded_pkg_prim_secded_inv_64_57_enc;
		input reg [56:0] data_i;
		reg [63:0] data_o;
		begin
			data_o = sv2v_cast_64(data_i);
			data_o[57] = ^(data_o & 64'h0103fff800007fff);
			data_o[58] = ^(data_o & 64'h017c1ff801ff801f);
			data_o[59] = ^(data_o & 64'h01bde1f87e0781e1);
			data_o[60] = ^(data_o & 64'h01deee3b8e388e22);
			data_o[61] = ^(data_o & 64'h01ef76cdb2c93244);
			data_o[62] = ^(data_o & 64'h01f7bb56d5525488);
			data_o[63] = ^(data_o & 64'h01fbdda769a46910);
			data_o = data_o ^ 64'h5400000000000000;
			prim_secded_pkg_prim_secded_inv_64_57_enc = data_o;
		end
	endfunction
	localparam signed [31:0] tlul_pkg_H2DCmdMaxWidth = 57;
	function automatic [(((prim_mubi_pkg_MuBi4Width + top_pkg_TL_AW) + 3) + top_pkg_TL_DBW) - 1:0] tlul_pkg_extract_h2d_cmd_intg;
		input reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl;
		reg [(((prim_mubi_pkg_MuBi4Width + top_pkg_TL_AW) + 3) + top_pkg_TL_DBW) - 1:0] payload;
		reg unused_tlul;
		begin
			unused_tlul = ^tl;
			payload[top_pkg_TL_AW + (top_pkg_TL_DBW + 2)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 2)) >= (3 + (top_pkg_TL_DBW + 0)) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 2)) - (3 + (top_pkg_TL_DBW + 0))) + 1 : ((3 + (top_pkg_TL_DBW + 0)) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 2))) + 1)] = tl[top_pkg_TL_AW + (top_pkg_TL_DBW + 55)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)];
			payload[top_pkg_TL_DBW + 2-:((top_pkg_TL_DBW + 2) >= (top_pkg_TL_DBW + 0) ? ((top_pkg_TL_DBW + 2) - (top_pkg_TL_DBW + 0)) + 1 : ((top_pkg_TL_DBW + 0) - (top_pkg_TL_DBW + 2)) + 1)] = tl[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)];
			payload[top_pkg_TL_DBW - 1-:top_pkg_TL_DBW] = tl[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))];
			payload[prim_mubi_pkg_MuBi4Width + (top_pkg_TL_AW + (top_pkg_TL_DBW + 2))-:(((32'sd4 + 32'sd32) + (top_pkg_TL_DBW + 2)) >= (35 + (top_pkg_TL_DBW + 0)) ? ((prim_mubi_pkg_MuBi4Width + (top_pkg_TL_AW + (top_pkg_TL_DBW + 2))) - (top_pkg_TL_AW + (3 + (top_pkg_TL_DBW + 0)))) + 1 : ((top_pkg_TL_AW + (3 + (top_pkg_TL_DBW + 0))) - (prim_mubi_pkg_MuBi4Width + (top_pkg_TL_AW + (top_pkg_TL_DBW + 2)))) + 1)] = tl[18-:4];
			tlul_pkg_extract_h2d_cmd_intg = payload;
		end
	endfunction
	function automatic [56:0] sv2v_cast_57;
		input reg [56:0] inp;
		sv2v_cast_57 = inp;
	endfunction
	function automatic [6:0] tlul_pkg_get_cmd_intg;
		input reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl;
		reg [6:0] cmd_intg;
		reg [56:0] unused_cmd_payload;
		reg [(((prim_mubi_pkg_MuBi4Width + top_pkg_TL_AW) + 3) + top_pkg_TL_DBW) - 1:0] cmd;
		begin
			cmd = tlul_pkg_extract_h2d_cmd_intg(tl);
			{cmd_intg, unused_cmd_payload} = prim_secded_pkg_prim_secded_inv_64_57_enc(sv2v_cast_57(cmd));
			tlul_pkg_get_cmd_intg = cmd_intg;
		end
	endfunction
	function automatic [6:0] tlul_pkg_get_bad_cmd_intg;
		input reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl;
		reg [6:0] cmd_intg;
		begin
			cmd_intg = tlul_pkg_get_cmd_intg(tl);
			tlul_pkg_get_bad_cmd_intg = ~cmd_intg;
		end
	endfunction
	function automatic [38:0] sv2v_cast_39;
		input reg [38:0] inp;
		sv2v_cast_39 = inp;
	endfunction
	function automatic [38:0] prim_secded_pkg_prim_secded_inv_39_32_enc;
		input reg [31:0] data_i;
		reg [38:0] data_o;
		begin
			data_o = sv2v_cast_39(data_i);
			data_o[32] = ^(data_o & 39'h002606bd25);
			data_o[33] = ^(data_o & 39'h00deba8050);
			data_o[34] = ^(data_o & 39'h00413d89aa);
			data_o[35] = ^(data_o & 39'h0031234ed1);
			data_o[36] = ^(data_o & 39'h00c2c1323b);
			data_o[37] = ^(data_o & 39'h002dcc624c);
			data_o[38] = ^(data_o & 39'h0098505586);
			data_o = data_o ^ 39'h2a00000000;
			prim_secded_pkg_prim_secded_inv_39_32_enc = data_o;
		end
	endfunction
	function automatic [6:0] tlul_pkg_get_data_intg;
		input reg [31:0] data;
		reg [6:0] data_intg;
		reg [31:0] unused_data;
		reg [(tlul_pkg_DataIntgWidth + top_pkg_TL_DW) - 1:0] enc_data;
		begin
			enc_data = prim_secded_pkg_prim_secded_inv_39_32_enc(data);
			data_intg = enc_data[(tlul_pkg_DataIntgWidth + top_pkg_TL_DW) - 1:top_pkg_TL_DW];
			unused_data = enc_data[31:0];
			tlul_pkg_get_data_intg = data_intg;
		end
	endfunction
	function automatic [6:0] tlul_pkg_get_bad_data_intg;
		input reg [31:0] data;
		reg [6:0] data_intg;
		begin
			data_intg = tlul_pkg_get_data_intg(data);
			tlul_pkg_get_bad_data_intg = ~data_intg;
		end
	endfunction
	function automatic [4:0] sv2v_cast_5;
		input reg [4:0] inp;
		sv2v_cast_5 = inp;
	endfunction
	function automatic [3:0] sv2v_cast_51AC7;
		input reg [3:0] inp;
		sv2v_cast_51AC7 = inp;
	endfunction
	function automatic [6:0] sv2v_cast_D1AC3;
		input reg [6:0] inp;
		sv2v_cast_D1AC3 = inp;
	endfunction
	assign blanked_auser = {sv2v_cast_5(tl_t_o[23-:5]), sv2v_cast_51AC7(tl_t_o[18-:4]), tlul_pkg_get_bad_cmd_intg(tl_t_o), sv2v_cast_D1AC3(tlul_pkg_get_bad_data_intg(tlul_pkg_BlankedAData))};
	genvar i;
	function automatic signed [NWD - 1:0] sv2v_cast_28286_signed;
		input reg signed [NWD - 1:0] inp;
		sv2v_cast_28286_signed = inp;
	endfunction
	generate
		for (i = 0; i < N; i = i + 1) begin : gen_u_o
			wire dev_select;
			assign dev_select = (dev_select_t == sv2v_cast_28286_signed(i)) & ~hold_all_requests;
			assign tl_u_o[i][7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] = tl_t_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & dev_select;
			assign tl_u_o[i][6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] = tl_t_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)];
			assign tl_u_o[i][3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] = tl_t_o[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)];
			assign tl_u_o[i][top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)] = tl_t_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)];
			assign tl_u_o[i][top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) >= (32'sd32 + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 56)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1)] = tl_t_o[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) >= (32'sd32 + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 56)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1)];
			assign tl_u_o[i][top_pkg_TL_AW + (top_pkg_TL_DBW + 55)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)] = tl_t_o[top_pkg_TL_AW + (top_pkg_TL_DBW + 55)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)];
			assign tl_u_o[i][top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))] = tl_t_o[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))];
			assign tl_u_o[i][55-:32] = (dev_select ? tl_t_o[55-:32] : tlul_pkg_BlankedAData);
			assign tl_u_o[i][23-:23] = (dev_select ? tl_t_o[23-:23] : blanked_auser);
			assign tl_u_o[i][0] = tl_t_o[0];
		end
	endgenerate
	reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_t_p;
	reg hfifo_reqready;
	always @(*) begin
		hfifo_reqready = tl_u_i[N][0];
		begin : sv2v_autoblock_1
			reg signed [31:0] idx;
			for (idx = 0; idx < N; idx = idx + 1)
				if (dev_select_t == sv2v_cast_28286_signed(idx))
					hfifo_reqready = tl_u_i[idx][0];
		end
		if (hold_all_requests)
			hfifo_reqready = 1'b0;
	end
	assign tl_t_i[0] = tl_t_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & hfifo_reqready;
	always @(*) begin
		tl_t_p = tl_u_i[N];
		begin : sv2v_autoblock_2
			reg signed [31:0] idx;
			for (idx = 0; idx < N; idx = idx + 1)
				if (dev_select_outstanding == sv2v_cast_28286_signed(idx))
					tl_t_p = tl_u_i[idx];
		end
	end
	assign tl_t_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] = tl_t_p[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))];
	assign tl_t_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)] = tl_t_p[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)];
	assign tl_t_i[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)] = tl_t_p[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)];
	assign tl_t_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)] = tl_t_p[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)];
	assign tl_t_i[top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))-:((32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))) >= ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) + 1 : ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) + 1)] = tl_t_p[top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))-:((32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))) >= ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) + 1 : ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) + 1)];
	assign tl_t_i[top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))-:(((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)) >= (32'sd32 + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) + 1 : ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) + 1)] = tl_t_p[top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))-:(((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)) >= (32'sd32 + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) + 1 : ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) + 1)];
	assign tl_t_i[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)] = tl_t_p[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)];
	assign tl_t_i[(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1-:(((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) >= 2 ? (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 0 : 3 - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))] = tl_t_p[(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1-:(((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) >= 2 ? (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 0 : 3 - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))];
	assign tl_t_i[1] = tl_t_p[1];
	generate
		for (i = 0; i < N; i = i + 1) begin : gen_dfifo
			tlul_fifo_sync #(
				.ReqPass(DReqPass[i]),
				.RspPass(DRspPass[i]),
				.ReqDepth(DReqDepth[i * 4+:4]),
				.RspDepth(DRspDepth[i * 4+:4])
			) fifo_d(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.tl_h_i(tl_u_o[i]),
				.tl_h_o(tl_u_i[i]),
				.tl_d_o(tl_d_o[(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) + (((N - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23)))+:(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))]),
				.tl_d_i(tl_d_i[((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1) + (((N - 1) - i) * ((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1)))+:((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1))]),
				.spare_req_i(1'b0),
				.spare_rsp_i(1'b0)
			);
		end
	endgenerate
	function automatic [NWD - 1:0] sv2v_cast_28286;
		input reg [NWD - 1:0] inp;
		sv2v_cast_28286 = inp;
	endfunction
	generate
		if ($clog2(N + 1) <= NWD) begin : gen_err_resp
			assign tl_u_o[N][0] = tl_t_o[0];
			assign tl_u_o[N][7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] = (tl_t_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & (dev_select_t >= sv2v_cast_28286(N))) & ~hold_all_requests;
			assign tl_u_o[N][6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] = tl_t_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)];
			assign tl_u_o[N][3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] = tl_t_o[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)];
			assign tl_u_o[N][top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)] = tl_t_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)];
			assign tl_u_o[N][top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) >= (32'sd32 + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 56)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1)] = tl_t_o[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) >= (32'sd32 + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 56)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1)];
			assign tl_u_o[N][top_pkg_TL_AW + (top_pkg_TL_DBW + 55)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)] = tl_t_o[top_pkg_TL_AW + (top_pkg_TL_DBW + 55)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)];
			assign tl_u_o[N][top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))] = tl_t_o[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))];
			assign tl_u_o[N][55-:32] = tl_t_o[55-:32];
			assign tl_u_o[N][23-:23] = tl_t_o[23-:23];
			tlul_err_resp err_resp(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.tl_h_i(tl_u_o[N]),
				.tl_h_o(tl_u_i[N])
			);
		end
		else begin : gen_no_err_resp
			assign tl_u_o[N] = 1'sb0;
			assign tl_u_i[N] = 1'sb0;
			wire unused_sig;
			assign unused_sig = ^tl_u_o[N];
		end
	endgenerate
endmodule
module tlul_socket_m1 (
	clk_i,
	rst_ni,
	tl_h_i,
	tl_h_o,
	tl_d_o,
	tl_d_i
);
	parameter [31:0] M = 4;
	parameter [M - 1:0] HReqPass = {M {1'b1}};
	parameter [M - 1:0] HRspPass = {M {1'b1}};
	parameter [(M * 4) - 1:0] HReqDepth = {M {4'h1}};
	parameter [(M * 4) - 1:0] HRspDepth = {M {4'h1}};
	parameter [0:0] DReqPass = 1'b1;
	parameter [0:0] DRspPass = 1'b1;
	parameter [3:0] DReqDepth = 4'h1;
	parameter [3:0] DRspDepth = 4'h1;
	input clk_i;
	input rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (M * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24)) - 1 : (M * (1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 22)):(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23)] tl_h_i;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	output wire [((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (M * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2)) - 1 : (M * (1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1))) + ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 0)):((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1)] tl_h_o;
	output wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_d_o;
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_d_i;
	localparam [31:0] IDW = top_pkg_TL_AIW;
	localparam [31:0] STIDW = $clog2(M);
	wire [(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (M * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24)) - 1 : (M * (1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 22)):(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23)] hreq_fifo_o;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] hrsp_fifo_i [0:M - 1];
	wire [M - 1:0] hrequest;
	wire [M - 1:0] hgrant;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] dreq_fifo_i;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] drsp_fifo_o;
	wire arb_valid;
	wire arb_ready;
	wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] arb_data;
	genvar i;
	function automatic [2:0] sv2v_cast_3;
		input reg [2:0] inp;
		sv2v_cast_3 = inp;
	endfunction
	function automatic [top_pkg_TL_SZW - 1:0] sv2v_cast_F164F;
		input reg [top_pkg_TL_SZW - 1:0] inp;
		sv2v_cast_F164F = inp;
	endfunction
	function automatic [7:0] sv2v_cast_5656E;
		input reg [7:0] inp;
		sv2v_cast_5656E = inp;
	endfunction
	function automatic [31:0] sv2v_cast_AEF98;
		input reg [31:0] inp;
		sv2v_cast_AEF98 = inp;
	endfunction
	function automatic [top_pkg_TL_DBW - 1:0] sv2v_cast_895D2;
		input reg [top_pkg_TL_DBW - 1:0] inp;
		sv2v_cast_895D2 = inp;
	endfunction
	function automatic [31:0] sv2v_cast_19205;
		input reg [31:0] inp;
		sv2v_cast_19205 = inp;
	endfunction
	function automatic [22:0] sv2v_cast_6B624;
		input reg [22:0] inp;
		sv2v_cast_6B624 = inp;
	endfunction
	generate
		for (i = 0; i < M; i = i + 1) begin : gen_host_fifo
			wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] hreq_fifo_i;
			wire [STIDW - 1:0] reqid_sub;
			wire [7:0] shifted_id;
			assign reqid_sub = i;
			assign shifted_id = {tl_h_i[(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - 7 : ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) - ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - 7)) : (((((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - 7 : ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) - ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - 7))) - (IDW - STIDW)) + 1)+:IDW - STIDW], reqid_sub};
			wire [7:IDW - STIDW] unused_tl_h_source;
			assign unused_tl_h_source = tl_h_i[(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) : ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) : (((((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) : ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + STIDW) - 1)-:STIDW];
			assign hreq_fifo_i = {tl_h_i[(((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) : ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) - (7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))))], sv2v_cast_3(tl_h_i[(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) : ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) : (((((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) : ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))))) + ((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)) - 1)-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)]), sv2v_cast_3(tl_h_i[(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) : ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) : (((((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) : ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))))) + ((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)) - 1)-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)]), sv2v_cast_F164F(tl_h_i[(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) : ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) : (((((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) : ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + ((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)) - 1)-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)]), sv2v_cast_5656E(shifted_id), sv2v_cast_AEF98(tl_h_i[(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? top_pkg_TL_AW + (top_pkg_TL_DBW + 55) : ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) : (((((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? top_pkg_TL_AW + (top_pkg_TL_DBW + 55) : ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)) - 1)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)]), sv2v_cast_895D2(tl_h_i[(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? top_pkg_TL_DBW + 55 : ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) - (top_pkg_TL_DBW + 55)) : (((((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? top_pkg_TL_DBW + 55 : ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) - (top_pkg_TL_DBW + 55))) + ((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))) - 1)-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))]), sv2v_cast_19205(tl_h_i[(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 55 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) - 32) : ((((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 55 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) - 32)) + 31)-:32]), sv2v_cast_6B624(tl_h_i[(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 23 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 0) : ((((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 23 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 0)) + 22)-:23]), tl_h_i[(((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23)]};
			tlul_fifo_sync #(
				.ReqPass(HReqPass[i]),
				.RspPass(HRspPass[i]),
				.ReqDepth(HReqDepth[i * 4+:4]),
				.RspDepth(HRspDepth[i * 4+:4]),
				.SpareReqW(1)
			) u_hostfifo(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.tl_h_i(hreq_fifo_i),
				.tl_h_o(tl_h_o[((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1) + (((M - 1) - i) * ((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1)))+:((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1))]),
				.tl_d_o(hreq_fifo_o[(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) + (((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23)))+:(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))]),
				.tl_d_i(hrsp_fifo_i[i]),
				.spare_req_i(1'b0),
				.spare_rsp_i(1'b0)
			);
		end
	endgenerate
	tlul_fifo_sync #(
		.ReqPass(DReqPass),
		.RspPass(DRspPass),
		.ReqDepth(DReqDepth),
		.RspDepth(DRspDepth),
		.SpareReqW(1)
	) u_devicefifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.tl_h_i(dreq_fifo_i),
		.tl_h_o(drsp_fifo_o),
		.tl_d_o(tl_d_o),
		.tl_d_i(tl_d_i),
		.spare_req_i(1'b0),
		.spare_rsp_i(1'b0)
	);
	generate
		for (i = 0; i < M; i = i + 1) begin : gen_arbreqgnt
			assign hrequest[i] = hreq_fifo_o[(((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) : ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23) - (7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))))];
		end
	endgenerate
	assign arb_ready = drsp_fifo_o[0];
	localparam tlul_pkg_ArbiterImpl = "PPC";
	generate
		if (tlul_pkg_ArbiterImpl == "PPC") begin : gen_arb_ppc
			prim_arbiter_ppc #(
				.N(M),
				.DW(1 * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24))
			) u_reqarb(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_chk_i(1'b0),
				.req_i(hrequest),
				.data_i(hreq_fifo_o),
				.gnt_o(hgrant),
				.valid_o(arb_valid),
				.data_o(arb_data),
				.ready_i(arb_ready)
			);
		end
		else if (tlul_pkg_ArbiterImpl == "BINTREE") begin : gen_tree_arb
			prim_arbiter_tree #(
				.N(M),
				.DW(1 * ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24))
			) u_reqarb(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_chk_i(1'b0),
				.req_i(hrequest),
				.data_i(hreq_fifo_o),
				.gnt_o(hgrant),
				.valid_o(arb_valid),
				.data_o(arb_data),
				.ready_i(arb_ready)
			);
		end
	endgenerate
	wire [M - 1:0] hfifo_rspvalid;
	wire [M - 1:0] dfifo_rspready;
	wire [7:0] hfifo_rspid;
	wire dfifo_rspready_merged;
	assign dfifo_rspready_merged = |dfifo_rspready;
	assign dreq_fifo_i = {arb_valid, sv2v_cast_3(arb_data[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)]), sv2v_cast_3(arb_data[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)]), sv2v_cast_F164F(arb_data[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)]), sv2v_cast_5656E(arb_data[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) >= (32'sd32 + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 56)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1)]), sv2v_cast_AEF98(arb_data[top_pkg_TL_AW + (top_pkg_TL_DBW + 55)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)]), sv2v_cast_895D2(arb_data[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))]), sv2v_cast_19205(arb_data[55-:32]), sv2v_cast_6B624(arb_data[23-:23]), dfifo_rspready_merged};
	assign hfifo_rspid = {{STIDW {1'b0}}, drsp_fifo_o[top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))):(top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - (7 - STIDW)]};
	function automatic [0:0] sv2v_cast_9DEED;
		input reg [0:0] inp;
		sv2v_cast_9DEED = inp;
	endfunction
	function automatic [(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 1:0] sv2v_cast_1E00F;
		input reg [(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) - 1:0] inp;
		sv2v_cast_1E00F = inp;
	endfunction
	generate
		for (i = 0; i < M; i = i + 1) begin : gen_idrouting
			assign hfifo_rspvalid[i] = drsp_fifo_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] & (drsp_fifo_o[(top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - 7+:STIDW] == i);
			assign dfifo_rspready[i] = (hreq_fifo_o[(((M - 1) - i) * (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23))) + (((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? 0 : (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23)] & (drsp_fifo_o[(top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) - 7+:STIDW] == i)) & drsp_fifo_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))];
			assign hrsp_fifo_i[i] = {hfifo_rspvalid[i], sv2v_cast_3(drsp_fifo_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((6 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)]), sv2v_cast_3(drsp_fifo_o[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))-:((3 + (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1))))) >= (top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2)))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))))) + 1)]), sv2v_cast_F164F(drsp_fifo_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)]), sv2v_cast_5656E(hfifo_rspid), sv2v_cast_9DEED(drsp_fifo_o[top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))-:(((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)) >= (32'sd32 + ((32'sd7 + 32'sd7) + 2)) ? ((top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))) + 1 : ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) - (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))) + 1)]), sv2v_cast_19205(drsp_fifo_o[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)]), sv2v_cast_1E00F(drsp_fifo_o[(tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1-:(((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1) >= 2 ? (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 0 : 3 - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))]), drsp_fifo_o[1], hgrant[i]};
		end
	endgenerate
endmodule
module tlul_sram_byte (
	clk_i,
	rst_ni,
	tl_i,
	tl_o,
	tl_sram_o,
	tl_sram_i,
	error_i,
	error_o
);
	parameter [0:0] EnableIntg = 0;
	parameter signed [31:0] Outstanding = 1;
	input clk_i;
	input rst_ni;
	localparam signed [31:0] prim_mubi_pkg_MuBi4Width = 4;
	localparam signed [31:0] tlul_pkg_DataIntgWidth = 7;
	localparam signed [31:0] tlul_pkg_H2DCmdIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_AIW = 8;
	localparam signed [31:0] top_pkg_TL_AW = 32;
	localparam signed [31:0] top_pkg_TL_DW = 32;
	localparam signed [31:0] top_pkg_TL_DBW = top_pkg_TL_DW >> 3;
	localparam signed [31:0] top_pkg_TL_SZW = $clog2($clog2(top_pkg_TL_DBW) + 1);
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_i;
	localparam signed [31:0] tlul_pkg_D2HRspIntgWidth = 7;
	localparam signed [31:0] top_pkg_TL_DIW = 1;
	output reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_o;
	output reg [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23:0] tl_sram_o;
	input wire [(((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1:0] tl_sram_i;
	input error_i;
	output wire error_o;
	function automatic integer prim_util_pkg_vbits;
		input integer value;
		prim_util_pkg_vbits = (value == 1 ? 1 : $clog2(value));
	endfunction
	function automatic signed [tlul_sram_byte.prim_util_pkg_vbits(Outstanding + 1) - 1:0] sv2v_cast_C8BB0_signed;
		input reg signed [tlul_sram_byte.prim_util_pkg_vbits(Outstanding + 1) - 1:0] inp;
		sv2v_cast_C8BB0_signed = inp;
	endfunction
	function automatic [top_pkg_TL_SZW - 1:0] sv2v_cast_53D14;
		input reg [top_pkg_TL_SZW - 1:0] inp;
		sv2v_cast_53D14 = inp;
	endfunction
	function automatic [2:0] sv2v_cast_3;
		input reg [2:0] inp;
		sv2v_cast_3 = inp;
	endfunction
	function automatic [top_pkg_TL_SZW - 1:0] sv2v_cast_BFA8D;
		input reg [top_pkg_TL_SZW - 1:0] inp;
		sv2v_cast_BFA8D = inp;
	endfunction
	function automatic [7:0] sv2v_cast_3FC4C;
		input reg [7:0] inp;
		sv2v_cast_3FC4C = inp;
	endfunction
	function automatic [31:0] sv2v_cast_B3982;
		input reg [31:0] inp;
		sv2v_cast_B3982 = inp;
	endfunction
	function automatic [top_pkg_TL_DBW - 1:0] sv2v_cast_10924;
		input reg [top_pkg_TL_DBW - 1:0] inp;
		sv2v_cast_10924 = inp;
	endfunction
	function automatic [31:0] sv2v_cast_F9BF7;
		input reg [31:0] inp;
		sv2v_cast_F9BF7 = inp;
	endfunction
	function automatic [22:0] sv2v_cast_BC556;
		input reg [22:0] inp;
		sv2v_cast_BC556 = inp;
	endfunction
	generate
		if (EnableIntg) begin : gen_integ_handling
			reg stall_host;
			reg rd_phase;
			reg rd_wait;
			reg wr_phase;
			reg [1:0] state_d;
			reg [1:0] state_q;
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					state_q <= 2'd0;
				else
					state_q <= state_d;
			wire a_ack;
			wire d_ack;
			wire sram_a_ack;
			wire sram_d_ack;
			wire wr_txn;
			wire byte_wr_txn;
			wire byte_req_ack;
			wire [prim_util_pkg_vbits(Outstanding + 1) - 1:0] pending_txn_cnt;
			assign a_ack = tl_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & tl_o[0];
			assign d_ack = tl_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] & tl_i[0];
			assign sram_a_ack = tl_sram_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & tl_sram_i[0];
			assign sram_d_ack = tl_sram_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] & tl_sram_o[0];
			assign wr_txn = (tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h0) | (tl_i[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] == 3'h1);
			assign byte_req_ack = (byte_wr_txn & a_ack) & ~error_i;
			assign byte_wr_txn = (tl_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & ~&tl_i[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))]) & wr_txn;
			always @(*) begin
				rd_wait = 1'b0;
				stall_host = 1'b0;
				wr_phase = 1'b0;
				rd_phase = 1'b0;
				state_d = state_q;
				case (state_q)
					2'd0:
						if (byte_wr_txn) begin
							rd_phase = 1'b1;
							if (byte_req_ack)
								state_d = 2'd1;
						end
					2'd1: begin
						rd_phase = 1'b1;
						stall_host = 1'b1;
						if (pending_txn_cnt == sv2v_cast_C8BB0_signed(1)) begin
							rd_wait = 1'b1;
							if (sram_d_ack)
								state_d = 2'd2;
						end
					end
					2'd2: begin
						stall_host = 1'b1;
						wr_phase = 1'b1;
						if (sram_a_ack)
							state_d = 2'd0;
					end
					default:
						;
				endcase
			end
			wire [(((((3 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 22:0] txn_data;
			wire [(((((3 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 22:0] held_data;
			wire fifo_rdy;
			localparam signed [31:0] TxnDataWidth = 1 * ((((((3 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23);
			wire [top_pkg_TL_SZW - 1:0] a_size;
			assign txn_data = {sv2v_cast_3(tl_i[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)]), sv2v_cast_BFA8D(tl_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)]), sv2v_cast_3FC4C(tl_i[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) >= (32'sd32 + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 56)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1)]), sv2v_cast_B3982(tl_i[top_pkg_TL_AW + (top_pkg_TL_DBW + 55)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)]), sv2v_cast_10924(tl_i[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))]), sv2v_cast_F9BF7(tl_i[55-:32]), sv2v_cast_BC556(tl_i[23-:23])};
			prim_fifo_sync #(
				.Width(TxnDataWidth),
				.Pass(1'b0),
				.Depth(1),
				.OutputZeroIfEmpty(1'b0)
			) u_sync_fifo(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.clr_i(1'b0),
				.wvalid_i(byte_req_ack),
				.wready_o(fifo_rdy),
				.wdata_i(txn_data),
				.rready_i(sram_a_ack),
				.rdata_o(held_data)
			);
			reg [31:0] rsp_data;
			always @(posedge clk_i)
				if (sram_d_ack && rd_wait)
					rsp_data <= tl_sram_i[top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)-:((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) >= ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) ? ((top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)) - ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)) + 1 : (((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2) - (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))) + 1)];
			reg [31:0] combined_data;
			wire [31:0] unused_data;
			always @(*) begin : sv2v_autoblock_1
				reg signed [31:0] i;
				for (i = 0; i < top_pkg_TL_DBW; i = i + 1)
					combined_data[i * 8+:8] = (held_data[(top_pkg_TL_DBW + 54) - ((top_pkg_TL_DBW - 1) - i)] ? held_data[23 + (i * 8)+:8] : rsp_data[i * 8+:8]);
			end
			wire [6:0] data_intg;
			tlul_data_integ_enc u_tlul_data_integ_enc(
				.data_i(combined_data),
				.data_intg_o({data_intg, unused_data})
			);
			reg [22:0] combined_user;
			always @(*) begin
				combined_user = held_data[22-:23];
				combined_user[6-:tlul_pkg_DataIntgWidth] = data_intg;
			end
			localparam [31:0] AccessSize = $clog2(top_pkg_TL_DBW);
			always @(*) begin
				tl_sram_o = tl_i;
				tl_sram_o[0] = tl_i[0] | rd_wait;
				if (wr_phase) begin
					tl_sram_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] = 1'b1;
					tl_sram_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] = 3'h0;
					tl_sram_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)] = sv2v_cast_53D14(AccessSize);
					tl_sram_o[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))] = {top_pkg_TL_DBW {1'b1}};
					tl_sram_o[top_pkg_TL_AW + (top_pkg_TL_DBW + 55)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) >= (top_pkg_TL_DBW + 56) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_DBW + 56)) + 1 : ((top_pkg_TL_DBW + 56) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1)] = held_data[top_pkg_TL_AW + (top_pkg_TL_DBW + 54)-:((top_pkg_TL_AW + (top_pkg_TL_DBW + 54)) >= (top_pkg_TL_DBW + 55) ? ((top_pkg_TL_AW + (top_pkg_TL_DBW + 54)) - (top_pkg_TL_DBW + 55)) + 1 : ((top_pkg_TL_DBW + 55) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) + 1)];
					tl_sram_o[(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (32 - AccessSize):(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - 31] = 1'sb0;
					tl_sram_o[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) >= (32'sd32 + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 56)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1)] = held_data[top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))-:(((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)) >= (32'sd32 + (top_pkg_TL_DBW + 55)) ? ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))) - (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) + 1 : ((top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) + 1)];
					tl_sram_o[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] = held_data[3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))-:((3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54)))) >= (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) ? ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1 : ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))))) + 1)];
					tl_sram_o[55-:32] = combined_data;
					tl_sram_o[23-:23] = combined_user;
				end
				else if (rd_phase) begin
					tl_sram_o[(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - (32 - AccessSize):(top_pkg_TL_AW + (top_pkg_TL_DBW + 55)) - 31] = 1'sb0;
					if (!error_i || stall_host) begin
						tl_sram_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)] = sv2v_cast_53D14(AccessSize);
						tl_sram_o[top_pkg_TL_DBW + 55-:((top_pkg_TL_DBW + 55) >= 56 ? top_pkg_TL_DBW : 57 - (top_pkg_TL_DBW + 55))] = {top_pkg_TL_DBW {1'b1}};
						tl_sram_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] = tl_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))] & ~stall_host;
						tl_sram_o[6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))-:((6 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)))) >= (3 + (top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)))) ? ((6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) - (3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))))) + 1 : ((3 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))))) - (6 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))))) + 1)] = 3'h4;
					end
				end
			end
			wire unused_held_data;
			assign unused_held_data = ^{held_data[(top_pkg_TL_AW + (top_pkg_TL_DBW + 54)) - (32 - AccessSize):(top_pkg_TL_AW + (top_pkg_TL_DBW + 54)) - 31], held_data[6-:tlul_pkg_DataIntgWidth], held_data[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 54))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 54))))) + 1)]};
			assign error_o = error_i & ~stall_host;
			wire size_fifo_rdy;
			prim_fifo_sync #(
				.Width(top_pkg_TL_SZW),
				.Pass(1'b0),
				.Depth(Outstanding),
				.OutputZeroIfEmpty(1'b1)
			) u_sync_fifo_a_size(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.clr_i(1'b0),
				.wvalid_i(a_ack),
				.wready_o(size_fifo_rdy),
				.wdata_i(tl_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))-:((top_pkg_TL_SZW + ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 55))) >= ((32'sd8 + 32'sd32) + (top_pkg_TL_DBW + 56)) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55)))) - (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56)))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 56))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_AW + (top_pkg_TL_DBW + 55))))) + 1)]),
				.rready_i(d_ack),
				.rdata_o(a_size),
				.depth_o(pending_txn_cnt)
			);
			always @(*) begin
				tl_o = tl_sram_i;
				tl_o[0] = ((tl_sram_i[0] & ~stall_host) & fifo_rdy) & size_fifo_rdy;
				tl_o[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] = tl_sram_i[7 + (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))] & ~rd_wait;
				tl_o[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)] = a_size;
			end
			wire unused_tl;
			assign unused_tl = |tl_sram_i[top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))-:((top_pkg_TL_SZW + (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 1)))) >= (32'sd8 + ((32'sd1 + 32'sd32) + ((32'sd7 + 32'sd7) + 2))) ? ((top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1))))) - (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2))))) + 1 : ((top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 2)))) - (top_pkg_TL_SZW + (top_pkg_TL_AIW + (top_pkg_TL_DIW + (top_pkg_TL_DW + ((tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth) + 1)))))) + 1)];
		end
		else begin : gen_no_integ_handling
			wire [(((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd32)) + top_pkg_TL_DBW) + 55) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 24 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_AW) + top_pkg_TL_DBW) + top_pkg_TL_DW) + 23)):1] sv2v_tmp_3382F;
			assign sv2v_tmp_3382F = tl_i;
			always @(*) tl_sram_o = sv2v_tmp_3382F;
			wire [((((((7 + top_pkg_TL_SZW) + (32'sd8 + 32'sd1)) + 32'sd32) + (32'sd7 + 32'sd7)) + 1) >= 0 ? (((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 2 : 1 - ((((((7 + top_pkg_TL_SZW) + top_pkg_TL_AIW) + top_pkg_TL_DIW) + top_pkg_TL_DW) + (tlul_pkg_D2HRspIntgWidth + tlul_pkg_DataIntgWidth)) + 1)):1] sv2v_tmp_1F073;
			assign sv2v_tmp_1F073 = tl_sram_i;
			always @(*) tl_o = sv2v_tmp_1F073;
			assign error_o = error_i;
		end
	endgenerate
endmodule
