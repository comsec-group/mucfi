`include "formal/assumptions/ibex_top_di_asm.sv"
`include "formal/assumptions/ibex_top_ti_asm.sv"
