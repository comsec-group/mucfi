bit gen_rs1_uc_orig;

assign gen_rs1_uc_orig =

((($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h10), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h11), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h14), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h15), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h18), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h19), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1c), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1d), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h12) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h13)), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h16) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h17)), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1a) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1b)), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1e) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1f)) }) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h18), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h19), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1c), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1d), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1a) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1b)), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1e) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1f)) }) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1c), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1d), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1e) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1f)) }) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | (((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1e) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1f)) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1f) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [31])))) | ((~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1f)) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [30])))))) | ((~ ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1e) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1f))) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1d) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [29])))) | ((~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1d)) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [28])))))))) | ((~ (| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1c), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1d), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1e) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1f)) })) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | (((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1a) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1b)) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1b) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [27])))) | ((~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1b)) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [26])))))) | ((~ ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1a) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1b))) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h19) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [25])))) | ((~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h19)) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [24])))))))))) | ((~ (| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h18), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h19), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1c), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1d), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1a) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1b)), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1e) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1f)) })) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h14), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h15), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h16) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h17)) }) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | (((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h16) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h17)) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h17) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [23])))) | ((~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h17)) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [22])))))) | ((~ ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h16) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h17))) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h15) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [21])))) | ((~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h15)) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [20])))))))) | ((~ (| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h14), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h15), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h16) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h17)) })) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | (((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h12) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h13)) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h13) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [19])))) | ((~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h13)) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [18])))))) | ((~ ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h12) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h13))) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h11) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [17])))) | ((~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h11)) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [16])))))))))))) | ((~ (| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h10), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h11), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h14), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h15), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h18), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h19), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1c), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1d), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h12) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h13)), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h16) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h17)), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1a) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1b)), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1e) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h1f)) })) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h08), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h09), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0c), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0d), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0a) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0b)), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0e) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0f)) }) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0c), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0d), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0e) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0f)) }) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | (((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0e) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0f)) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0f) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [15])))) | ((~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0f)) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [14])))))) | ((~ ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0e) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0f))) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0d) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [13])))) | ((~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0d)) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [12])))))))) | ((~ (| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0c), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0d), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0e) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0f)) })) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | (((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0a) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0b)) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0b) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [11])))) | ((~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0b)) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [10])))))) | ((~ ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0a) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0b))) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h09) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [9])))) | ((~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h09)) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [8])))))))))) | ((~ (| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h08), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h09), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0c), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0d), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0a) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0b)), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0e) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h0f)) })) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h04), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h05), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h06) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h07)) }) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | (((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h06) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h07)) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h07) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [7])))) | ((~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h07)) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [6])))))) | ((~ ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h06) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h07))) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h05) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [5])))) | ((~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h05)) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [4])))))))) | ((~ (| { (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h04), (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h05), ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h06) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h07)) })) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | (((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h02) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h03)) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h03) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [3])))) | ((~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h03)) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [2])))))) | ((~ ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h02) | (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h03))) & (($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | ((u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h01) & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__gen_wren_check__u_prim_buf__gen_generic__u_impl_generic__in_i [1])))) | ((~ (u_ibex_core__id_stage_i__controller_i__instr_i [19:15] ==  5'h01)) & ($past(((~ rst_ni) | u_ibex_core__if_stage_i__if_id_pipe_reg_we )) | (gen_regfile_ff__register_file_i__dummy_instr_id_i  & $past(((~ rst_ni) | gen_regfile_ff__register_file_i__g_dummy_r0__we_r0_dummy )))))))))))))));

