
bit[31:0] op1_CSRRS_t0;
assign op1_CSRRS_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_CSRRC_t0;
assign op1_CSRRC_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_FENCE_t0;
assign op1_FENCE_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_CSRRWI_t0;
assign op1_CSRRWI_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_FENCE_I_t0;
assign op1_FENCE_I_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_CSRRSI_t0;
assign op1_CSRRSI_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_CSRRW_t0;
assign op1_CSRRW_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_EBREAK_t0;
assign op1_EBREAK_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_CSRRCI_t0;
assign op1_CSRRCI_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_ECALL_t0;
assign op1_ECALL_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_ADD_t0;
assign op1_ADD_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_ADD_t0;
assign op2_ADD_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_ADDI_t0;
assign op1_ADDI_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_AND_t0;
assign op1_AND_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_AND_t0;
assign op2_AND_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_ANDI_t0;
assign op1_ANDI_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_BEQ_t0;
assign op1_BEQ_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_BEQ_t0;
assign op2_BEQ_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_BGE_t0;
assign op1_BGE_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_BGE_t0;
assign op2_BGE_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_BGEU_t0;
assign op1_BGEU_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_BGEU_t0;
assign op2_BGEU_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_BLT_t0;
assign op1_BLT_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_BLT_t0;
assign op2_BLT_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_BLTU_t0;
assign op1_BLTU_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_BLTU_t0;
assign op2_BLTU_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_BNE_t0;
assign op1_BNE_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_BNE_t0;
assign op2_BNE_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_DIV_t0;
assign op1_DIV_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_DIV_t0;
assign op2_DIV_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_DIVU_t0;
assign op1_DIVU_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_DIVU_t0;
assign op2_DIVU_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_JALR_t0;
assign op1_JALR_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_LB_t0;
assign op1_LB_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_LBU_t0;
assign op1_LBU_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_LH_t0;
assign op1_LH_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_LHU_t0;
assign op1_LHU_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_LW_t0;
assign op1_LW_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_MUL_t0;
assign op1_MUL_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_MUL_t0;
assign op2_MUL_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_MULH_t0;
assign op1_MULH_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_MULH_t0;
assign op2_MULH_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_MULHSU_t0;
assign op1_MULHSU_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_MULHSU_t0;
assign op2_MULHSU_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_MULHU_t0;
assign op1_MULHU_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_MULHU_t0;
assign op2_MULHU_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_OR_t0;
assign op1_OR_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_OR_t0;
assign op2_OR_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_ORI_t0;
assign op1_ORI_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_REM_t0;
assign op1_REM_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_REM_t0;
assign op2_REM_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_REMU_t0;
assign op1_REMU_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_REMU_t0;
assign op2_REMU_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SB_t0;
assign op1_SB_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_SH_t0;
assign op1_SH_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_SLL_t0;
assign op1_SLL_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_SLL_t0;
assign op2_SLL_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SLLI_t0;
assign op1_SLLI_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_SLT_t0;
assign op1_SLT_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_SLT_t0;
assign op2_SLT_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SLTI_t0;
assign op1_SLTI_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_SLTIU_t0;
assign op1_SLTIU_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_SLTU_t0;
assign op1_SLTU_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_SLTU_t0;
assign op2_SLTU_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SRA_t0;
assign op1_SRA_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_SRA_t0;
assign op2_SRA_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SRAI_t0;
assign op1_SRAI_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_SRL_t0;
assign op1_SRL_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_SRL_t0;
assign op2_SRL_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SRLI_t0;
assign op1_SRLI_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_SUB_t0;
assign op1_SUB_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_SUB_t0;
assign op2_SUB_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SW_t0;
assign op1_SW_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_XOR_t0;
assign op1_XOR_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_XOR_t0;
assign op2_XOR_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_XORI_t0;
assign op1_XORI_t0 = i_pipeline__i_gprs__rs1_data_t0;

// Generated by gen_checker_inst.py


bit[31:0] op1_SHA512SIG1L_t0;
assign op1_SHA512SIG1L_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_SHA512SIG1L_t0;
assign op2_SHA512SIG1L_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_AES32DSI_t0;
assign op1_AES32DSI_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_AES32DSI_t0;
assign op2_AES32DSI_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SM4ED_t0;
assign op1_SM4ED_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_SM4ED_t0;
assign op2_SM4ED_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SHA512SUM1_t0;
assign op1_SHA512SUM1_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_AES32ESI_t0;
assign op1_AES32ESI_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_AES32ESI_t0;
assign op2_AES32ESI_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SHA512SUM1R_t0;
assign op1_SHA512SUM1R_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_SHA512SUM1R_t0;
assign op2_SHA512SUM1R_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SHA512SIG0L_t0;
assign op1_SHA512SIG0L_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_SHA512SIG0L_t0;
assign op2_SHA512SIG0L_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SM3P1_t0;
assign op1_SM3P1_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_SM3P0_t0;
assign op1_SM3P0_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_AES64ES_t0;
assign op1_AES64ES_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_AES64ES_t0;
assign op2_AES64ES_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SHA256SIG1_t0;
assign op1_SHA256SIG1_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_AES64IM_t0;
assign op1_AES64IM_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_SHA512SUM0R_t0;
assign op1_SHA512SUM0R_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_SHA512SUM0R_t0;
assign op2_SHA512SUM0R_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_AES32DSMI_t0;
assign op1_AES32DSMI_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_AES32DSMI_t0;
assign op2_AES32DSMI_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SHA512SUM0_t0;
assign op1_SHA512SUM0_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_SHA512SIG0_t0;
assign op1_SHA512SIG0_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_AES64ESM_t0;
assign op1_AES64ESM_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_AES64ESM_t0;
assign op2_AES64ESM_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_AES64KS1I_t0;
assign op1_AES64KS1I_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_AES64KS2_t0;
assign op1_AES64KS2_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_AES64KS2_t0;
assign op2_AES64KS2_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SHA256SIG0_t0;
assign op1_SHA256SIG0_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_AES64DSM_t0;
assign op1_AES64DSM_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_AES64DSM_t0;
assign op2_AES64DSM_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_AES64DS_t0;
assign op1_AES64DS_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_AES64DS_t0;
assign op2_AES64DS_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SHA512SIG0H_t0;
assign op1_SHA512SIG0H_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_SHA512SIG0H_t0;
assign op2_SHA512SIG0H_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SHA256SUM0_t0;
assign op1_SHA256SUM0_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_SHA512SIG1H_t0;
assign op1_SHA512SIG1H_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_SHA512SIG1H_t0;
assign op2_SHA512SIG1H_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SHA512SIG1_t0;
assign op1_SHA512SIG1_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_SM4KS_t0;
assign op1_SM4KS_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_SM4KS_t0;
assign op2_SM4KS_t0 = i_pipeline__i_gprs__rs2_data_t0;

bit[31:0] op1_SHA256SUM1_t0;
assign op1_SHA256SUM1_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op1_AES32ESMI_t0;
assign op1_AES32ESMI_t0 = i_pipeline__i_gprs__rs1_data_t0;

bit[31:0] op2_AES32ESMI_t0;
assign op2_AES32ESMI_t0 = i_pipeline__i_gprs__rs2_data_t0;


