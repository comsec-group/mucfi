module \$paramod$038d6e761af5e8bbfc2ed9b8473abfd849408d7b\ibex_id_stage (clk_i, rst_ni, ctrl_busy_o, illegal_insn_o, instr_valid_i, instr_rdata_i, instr_rdata_alu_i, instr_rdata_c_i, instr_is_compressed_i, instr_bp_taken_i, instr_req_o, instr_first_cycle_id_o, instr_valid_clear_o, id_in_ready_o, instr_exec_i, icache_inval_o, branch_decision_i, pc_set_o, pc_mux_o, nt_branch_mispredict_o, nt_branch_addr_o
, exc_pc_mux_o, exc_cause_o, illegal_c_insn_i, instr_fetch_err_i, instr_fetch_err_plus2_i, pc_id_i, ex_valid_i, lsu_resp_valid_i, alu_operator_ex_o, alu_operand_a_ex_o, alu_operand_b_ex_o, imd_val_we_ex_i, imd_val_d_ex_i, imd_val_q_ex_o, bt_a_operand_o, bt_b_operand_o, mult_en_ex_o, div_en_ex_o, mult_sel_ex_o, div_sel_ex_o, multdiv_operator_ex_o
, multdiv_signed_mode_ex_o, multdiv_operand_a_ex_o, multdiv_operand_b_ex_o, multdiv_ready_id_o, csr_access_o, csr_op_o, csr_op_en_o, csr_save_if_o, csr_save_id_o, csr_save_wb_o, csr_restore_mret_id_o, csr_restore_dret_id_o, csr_save_cause_o, csr_mtval_o, priv_mode_i, csr_mstatus_tw_i, illegal_csr_insn_i, data_ind_timing_i, lsu_req_o, lsu_we_o, lsu_type_o
, lsu_sign_ext_o, lsu_wdata_o, lsu_req_done_i, lsu_addr_incr_req_i, lsu_addr_last_i, csr_mstatus_mie_i, irq_pending_i, irqs_i, irq_nm_i, nmi_mode_o, lsu_load_err_i, lsu_load_resp_intg_err_i, lsu_store_err_i, lsu_store_resp_intg_err_i, debug_mode_o, debug_mode_entering_o, debug_cause_o, debug_csr_save_o, debug_req_i, debug_single_step_i, debug_ebreakm_i
, debug_ebreaku_i, trigger_match_i, result_ex_i, csr_rdata_i, rf_raddr_a_o, rf_rdata_a_i, rf_raddr_b_o, rf_rdata_b_i, rf_ren_a_o, rf_ren_b_o, rf_waddr_id_o, rf_wdata_id_o, rf_we_id_o, rf_rd_a_wb_match_o, rf_rd_b_wb_match_o, rf_waddr_wb_i, rf_wdata_fwd_wb_i, rf_write_wb_i, en_wb_o, instr_type_wb_o, instr_perf_count_id_o
, ready_wb_i, outstanding_load_wb_i, outstanding_store_wb_i, perf_jump_o, perf_branch_o, perf_tbranch_o, perf_dside_wait_o, perf_mul_wait_o, perf_div_wait_o, instr_id_done_o, trigger_match_i_t0, debug_cause_o_t0, debug_csr_save_o_t0, debug_ebreakm_i_t0, debug_ebreaku_i_t0, debug_mode_entering_o_t0, debug_mode_o_t0, debug_req_i_t0, debug_single_step_i_t0, exc_cause_o_t0, exc_pc_mux_o_t0
, id_in_ready_o_t0, instr_bp_taken_i_t0, instr_exec_i_t0, instr_fetch_err_i_t0, instr_fetch_err_plus2_i_t0, instr_is_compressed_i_t0, instr_valid_clear_o_t0, instr_valid_i_t0, irq_pending_i_t0, irqs_i_t0, lsu_addr_last_i_t0, nmi_mode_o_t0, nt_branch_mispredict_o_t0, pc_id_i_t0, pc_mux_o_t0, pc_set_o_t0, perf_jump_o_t0, csr_mstatus_mie_i_t0, perf_tbranch_o_t0, priv_mode_i_t0, csr_mtval_o_t0
, ready_wb_i_t0, csr_restore_dret_id_o_t0, csr_restore_mret_id_o_t0, csr_save_cause_o_t0, csr_save_id_o_t0, csr_save_if_o_t0, csr_save_wb_o_t0, ctrl_busy_o_t0, alu_operand_a_ex_o_t0, alu_operand_b_ex_o_t0, alu_operator_ex_o_t0, branch_decision_i_t0, bt_a_operand_o_t0, bt_b_operand_o_t0, csr_mstatus_tw_i_t0, csr_op_en_o_t0, csr_rdata_i_t0, data_ind_timing_i_t0, div_en_ex_o_t0, div_sel_ex_o_t0, en_wb_o_t0
, ex_valid_i_t0, illegal_csr_insn_i_t0, imd_val_d_ex_i_t0, imd_val_q_ex_o_t0, imd_val_we_ex_i_t0, instr_first_cycle_id_o_t0, instr_id_done_o_t0, instr_perf_count_id_o_t0, instr_rdata_c_i_t0, instr_type_wb_o_t0, irq_nm_i_t0, lsu_addr_incr_req_i_t0, lsu_load_err_i_t0, lsu_load_resp_intg_err_i_t0, lsu_req_done_i_t0, lsu_req_o_t0, lsu_resp_valid_i_t0, lsu_sign_ext_o_t0, lsu_store_err_i_t0, lsu_store_resp_intg_err_i_t0, lsu_type_o_t0
, lsu_wdata_o_t0, lsu_we_o_t0, mult_en_ex_o_t0, mult_sel_ex_o_t0, multdiv_operand_a_ex_o_t0, multdiv_operand_b_ex_o_t0, multdiv_operator_ex_o_t0, multdiv_ready_id_o_t0, multdiv_signed_mode_ex_o_t0, nt_branch_addr_o_t0, outstanding_load_wb_i_t0, outstanding_store_wb_i_t0, perf_branch_o_t0, perf_div_wait_o_t0, perf_dside_wait_o_t0, perf_mul_wait_o_t0, result_ex_i_t0, rf_rd_a_wb_match_o_t0, rf_rd_b_wb_match_o_t0, rf_rdata_a_i_t0, rf_rdata_b_i_t0
, rf_waddr_id_o_t0, rf_waddr_wb_i_t0, rf_wdata_fwd_wb_i_t0, rf_wdata_id_o_t0, rf_we_id_o_t0, rf_write_wb_i_t0, rf_ren_b_o_t0, rf_ren_a_o_t0, rf_raddr_b_o_t0, rf_raddr_a_o_t0, instr_rdata_alu_i_t0, illegal_insn_o_t0, illegal_c_insn_i_t0, icache_inval_o_t0, csr_op_o_t0, csr_access_o_t0, instr_req_o_t0, instr_rdata_i_t0);
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0001_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0003_;
/* src = "generated/sv2v_out.v:17539.2-17548.5" */
wire _0004_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0005_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0007_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0008_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0009_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0010_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0011_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0013_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0015_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0016_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0017_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0018_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0019_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0021_;
/* src = "generated/sv2v_out.v:17539.2-17548.5" */
wire _0022_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0023_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0024_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0025_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0026_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0027_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0028_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0029_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0030_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0031_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0032_;
/* src = "generated/sv2v_out.v:17539.2-17548.5" */
wire _0033_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0034_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0035_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0036_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0037_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0038_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0039_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0040_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0041_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0042_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0043_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0044_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0045_;
/* src = "generated/sv2v_out.v:17693.2-17752.5" */
wire _0046_;
/* src = "generated/sv2v_out.v:17359.22-17359.56" */
wire _0047_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17359.22-17359.56" */
wire _0048_;
/* src = "generated/sv2v_out.v:17359.21-17359.75" */
wire _0049_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17359.21-17359.75" */
wire _0050_;
/* src = "generated/sv2v_out.v:17474.23-17474.50" */
wire _0051_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17474.23-17474.50" */
wire _0052_;
/* src = "generated/sv2v_out.v:17550.73-17550.104" */
wire _0053_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17550.73-17550.104" */
wire _0054_;
/* src = "generated/sv2v_out.v:17625.38-17625.68" */
wire _0055_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17625.38-17625.68" */
wire _0056_;
/* src = "generated/sv2v_out.v:17633.24-17633.54" */
wire _0057_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17633.24-17633.54" */
wire _0058_;
/* src = "generated/sv2v_out.v:17741.19-17741.41" */
wire _0059_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17741.19-17741.41" */
wire _0060_;
/* src = "generated/sv2v_out.v:17742.10-17742.38" */
wire _0061_;
/* src = "generated/sv2v_out.v:17755.23-17755.44" */
wire _0062_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17755.23-17755.44" */
wire _0063_;
/* src = "generated/sv2v_out.v:17770.35-17770.88" */
wire _0064_;
/* src = "generated/sv2v_out.v:17771.31-17771.58" */
wire _0065_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17771.31-17771.58" */
wire _0066_;
/* src = "generated/sv2v_out.v:17771.30-17771.74" */
wire _0067_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17771.30-17771.74" */
wire _0068_;
/* src = "generated/sv2v_out.v:17772.69-17772.98" */
wire _0069_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17772.69-17772.98" */
wire _0070_;
/* src = "generated/sv2v_out.v:17779.29-17779.61" */
wire _0071_;
/* src = "generated/sv2v_out.v:17780.29-17780.61" */
wire _0072_;
/* src = "generated/sv2v_out.v:17820.36-17820.64" */
wire _0073_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17820.36-17820.64" */
wire _0074_;
/* src = "generated/sv2v_out.v:17820.35-17820.85" */
wire _0075_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17820.35-17820.85" */
wire _0076_;
/* src = "generated/sv2v_out.v:17820.34-17820.108" */
wire _0077_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17820.34-17820.108" */
wire _0078_;
wire [31:0] _0079_;
wire _0080_;
wire _0081_;
wire _0082_;
wire [31:0] _0083_;
wire [31:0] _0084_;
wire [31:0] _0085_;
wire [31:0] _0086_;
wire [31:0] _0087_;
wire _0088_;
wire [31:0] _0089_;
wire [31:0] _0090_;
wire [31:0] _0091_;
wire [31:0] _0092_;
wire _0093_;
wire _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire [31:0] _0101_;
wire [31:0] _0102_;
wire [31:0] _0103_;
wire [31:0] _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire _0109_;
wire _0110_;
wire _0111_;
wire _0112_;
wire _0113_;
wire _0114_;
wire _0115_;
wire _0116_;
wire _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire _0139_;
wire _0140_;
wire _0141_;
wire _0142_;
wire _0143_;
wire [31:0] _0144_;
wire [31:0] _0145_;
wire _0146_;
wire _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
wire _0152_;
wire _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire _0186_;
wire _0187_;
wire _0188_;
wire _0189_;
wire _0190_;
wire _0191_;
wire _0192_;
wire _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire _0199_;
wire _0200_;
wire _0201_;
wire _0202_;
wire _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
wire _0221_;
wire _0222_;
wire _0223_;
wire _0224_;
wire _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire _0241_;
wire _0242_;
wire _0243_;
wire _0244_;
wire _0245_;
wire _0246_;
wire _0247_;
wire [33:0] _0248_;
wire [33:0] _0249_;
wire [33:0] _0250_;
wire [33:0] _0251_;
wire _0252_;
wire [31:0] _0253_;
wire [31:0] _0254_;
wire [31:0] _0255_;
wire [31:0] _0256_;
wire [31:0] _0257_;
wire [31:0] _0258_;
wire [31:0] _0259_;
wire [31:0] _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire [31:0] _0264_;
wire [31:0] _0265_;
wire [31:0] _0266_;
wire [31:0] _0267_;
wire [31:0] _0268_;
wire [31:0] _0269_;
wire [31:0] _0270_;
wire [31:0] _0271_;
wire _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire _0276_;
wire _0277_;
wire _0278_;
wire _0279_;
wire _0280_;
wire _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire _0285_;
wire _0286_;
wire _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire _0294_;
wire _0295_;
wire _0296_;
wire _0297_;
wire _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire _0324_;
wire _0325_;
wire _0326_;
wire _0327_;
wire _0328_;
wire _0329_;
wire _0330_;
wire _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire _0335_;
wire _0336_;
wire _0337_;
wire _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire _0344_;
wire _0345_;
wire _0346_;
wire [31:0] _0347_;
wire [31:0] _0348_;
wire [31:0] _0349_;
wire [31:0] _0350_;
wire [31:0] _0351_;
wire [31:0] _0352_;
wire [31:0] _0353_;
wire _0354_;
wire _0355_;
wire _0356_;
wire _0357_;
wire _0358_;
wire _0359_;
wire _0360_;
wire _0361_;
wire _0362_;
wire _0363_;
wire _0364_;
wire _0365_;
wire _0366_;
wire _0367_;
wire _0368_;
wire _0369_;
wire _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire _0376_;
wire _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire _0382_;
wire _0383_;
wire _0384_;
wire _0385_;
wire _0386_;
wire _0387_;
wire _0388_;
wire [33:0] _0389_;
wire [33:0] _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire _0398_;
wire _0399_;
wire _0400_;
wire _0401_;
wire _0402_;
wire _0403_;
wire _0404_;
wire _0405_;
wire _0406_;
wire _0407_;
wire _0408_;
wire _0409_;
wire _0410_;
wire _0411_;
wire _0412_;
wire _0413_;
wire [31:0] _0414_;
wire [31:0] _0415_;
wire [31:0] _0416_;
wire [31:0] _0417_;
/* cellift = 32'd1 */
wire [31:0] _0418_;
wire [31:0] _0419_;
/* cellift = 32'd1 */
wire [31:0] _0420_;
wire [31:0] _0421_;
/* cellift = 32'd1 */
wire [31:0] _0422_;
wire [31:0] _0423_;
/* cellift = 32'd1 */
wire [31:0] _0424_;
wire [31:0] _0425_;
/* cellift = 32'd1 */
wire [31:0] _0426_;
wire [31:0] _0427_;
/* cellift = 32'd1 */
wire [31:0] _0428_;
wire [31:0] _0429_;
/* cellift = 32'd1 */
wire [31:0] _0430_;
/* src = "generated/sv2v_out.v:17541.34-17541.50" */
wire _0431_;
/* src = "generated/sv2v_out.v:17541.56-17541.72" */
wire _0432_;
/* src = "generated/sv2v_out.v:17542.11-17542.42" */
wire _0433_;
/* src = "generated/sv2v_out.v:17542.48-17542.79" */
wire _0434_;
/* src = "generated/sv2v_out.v:17542.86-17542.117" */
wire _0435_;
/* src = "generated/sv2v_out.v:17542.124-17542.153" */
wire _0436_;
/* src = "generated/sv2v_out.v:17546.11-17546.42" */
wire _0437_;
/* src = "generated/sv2v_out.v:17546.48-17546.79" */
wire _0438_;
/* src = "generated/sv2v_out.v:17546.86-17546.117" */
wire _0439_;
/* src = "generated/sv2v_out.v:17546.124-17546.155" */
wire _0440_;
/* src = "generated/sv2v_out.v:17773.31-17773.60" */
wire _0441_;
/* src = "generated/sv2v_out.v:17774.31-17774.60" */
wire _0442_;
/* src = "generated/sv2v_out.v:17541.7-17541.74" */
wire _0443_;
/* src = "generated/sv2v_out.v:17545.12-17545.55" */
wire _0444_;
/* src = "generated/sv2v_out.v:17541.33-17541.73" */
wire _0445_;
/* src = "generated/sv2v_out.v:17542.10-17542.80" */
wire _0446_;
/* src = "generated/sv2v_out.v:17542.9-17542.118" */
wire _0447_;
/* src = "generated/sv2v_out.v:17542.8-17542.154" */
wire _0448_;
/* src = "generated/sv2v_out.v:17546.10-17546.80" */
wire _0449_;
/* src = "generated/sv2v_out.v:17546.9-17546.118" */
wire _0450_;
/* src = "generated/sv2v_out.v:17546.8-17546.156" */
wire _0451_;
/* src = "generated/sv2v_out.v:17720.20-17720.80" */
wire _0452_;
/* src = "generated/sv2v_out.v:17545.38-17545.54" */
wire _0453_;
/* src = "generated/sv2v_out.v:17550.31-17550.51" */
wire _0454_;
/* src = "generated/sv2v_out.v:17359.60-17359.75" */
wire _0455_;
/* src = "generated/sv2v_out.v:17549.45-17549.58" */
wire _0456_;
/* src = "generated/sv2v_out.v:17657.95-17657.115" */
wire _0457_;
/* src = "generated/sv2v_out.v:17755.23-17755.32" */
wire _0458_;
/* src = "generated/sv2v_out.v:17755.35-17755.44" */
wire _0459_;
/* src = "generated/sv2v_out.v:17767.90-17767.107" */
wire _0460_;
/* src = "generated/sv2v_out.v:17769.78-17769.93" */
wire _0461_;
/* src = "generated/sv2v_out.v:17771.47-17771.58" */
wire _0462_;
/* src = "generated/sv2v_out.v:17784.32-17784.43" */
wire _0463_;
/* src = "generated/sv2v_out.v:17820.36-17820.46" */
wire _0464_;
/* src = "generated/sv2v_out.v:17820.49-17820.64" */
wire _0465_;
/* src = "generated/sv2v_out.v:17550.56-17550.105" */
wire _0466_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17550.56-17550.105" */
wire _0467_;
/* src = "generated/sv2v_out.v:17551.45-17551.82" */
wire _0468_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17551.45-17551.82" */
wire _0469_;
/* src = "generated/sv2v_out.v:17551.44-17551.103" */
wire _0470_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17551.44-17551.103" */
wire _0471_;
/* src = "generated/sv2v_out.v:17551.43-17551.125" */
wire _0472_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17551.43-17551.125" */
wire _0473_;
/* src = "generated/sv2v_out.v:17657.36-17657.65" */
wire _0474_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17657.36-17657.65" */
wire _0475_;
/* src = "generated/sv2v_out.v:17657.35-17657.91" */
wire _0476_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17657.35-17657.91" */
wire _0477_;
/* src = "generated/sv2v_out.v:17721.23-17721.81" */
wire _0478_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17721.23-17721.81" */
wire _0479_;
/* src = "generated/sv2v_out.v:17754.24-17754.47" */
wire _0480_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17754.24-17754.47" */
wire _0481_;
/* src = "generated/sv2v_out.v:17754.23-17754.64" */
wire _0482_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17754.23-17754.64" */
wire _0483_;
/* src = "generated/sv2v_out.v:17754.22-17754.78" */
wire _0484_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17754.22-17754.78" */
wire _0485_;
/* src = "generated/sv2v_out.v:17754.21-17754.94" */
wire _0486_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17754.21-17754.94" */
wire _0487_;
/* src = "generated/sv2v_out.v:17767.40-17767.86" */
wire _0488_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17767.40-17767.86" */
wire _0489_;
/* src = "generated/sv2v_out.v:17769.26-17769.58" */
wire _0490_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17769.26-17769.58" */
wire _0491_;
/* src = "generated/sv2v_out.v:17769.25-17769.74" */
wire _0492_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17769.25-17769.74" */
wire _0493_;
/* src = "generated/sv2v_out.v:17772.40-17772.99" */
wire _0494_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17772.40-17772.99" */
wire _0495_;
/* src = "generated/sv2v_out.v:17781.50-17781.73" */
wire _0496_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17781.50-17781.73" */
wire _0497_;
/* src = "generated/sv2v_out.v:17785.64-17785.103" */
wire _0498_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17785.64-17785.103" */
wire _0499_;
wire _0500_;
wire _0501_;
wire _0502_;
wire _0503_;
wire _0504_;
wire _0505_;
wire _0506_;
wire _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
/* cellift = 32'd1 */
wire _0514_;
wire _0515_;
/* cellift = 32'd1 */
wire _0516_;
wire _0517_;
/* cellift = 32'd1 */
wire _0518_;
wire _0519_;
/* cellift = 32'd1 */
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
/* cellift = 32'd1 */
wire _0525_;
wire _0526_;
/* cellift = 32'd1 */
wire _0527_;
wire _0528_;
wire _0529_;
/* cellift = 32'd1 */
wire _0530_;
wire _0531_;
/* cellift = 32'd1 */
wire _0532_;
wire _0533_;
/* cellift = 32'd1 */
wire _0534_;
wire _0535_;
/* cellift = 32'd1 */
wire _0536_;
wire _0537_;
/* cellift = 32'd1 */
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0542_;
wire _0543_;
/* src = "generated/sv2v_out.v:17773.64-17773.77" */
wire _0544_;
/* src = "generated/sv2v_out.v:17774.64-17774.77" */
wire _0545_;
/* src = "generated/sv2v_out.v:17720.20-17720.94" */
wire _0546_;
/* src = "generated/sv2v_out.v:17782.53-17782.73" */
wire [1:0] _0547_;
/* src = "generated/sv2v_out.v:17370.7-17370.25" */
wire alu_multicycle_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17370.7-17370.25" */
/* unused_bits = "0" */
wire alu_multicycle_dec_t0;
/* src = "generated/sv2v_out.v:17366.13-17366.29" */
wire [1:0] alu_op_a_mux_sel;
/* src = "generated/sv2v_out.v:17367.13-17367.33" */
wire [1:0] alu_op_a_mux_sel_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17367.13-17367.33" */
/* unused_bits = "0 1" */
wire [1:0] alu_op_a_mux_sel_dec_t0;
/* src = "generated/sv2v_out.v:17368.7-17368.23" */
wire alu_op_b_mux_sel;
/* src = "generated/sv2v_out.v:17369.7-17369.27" */
wire alu_op_b_mux_sel_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17369.7-17369.27" */
/* unused_bits = "0" */
wire alu_op_b_mux_sel_dec_t0;
/* src = "generated/sv2v_out.v:17222.21-17222.39" */
output [31:0] alu_operand_a_ex_o;
wire [31:0] alu_operand_a_ex_o;
/* cellift = 32'd1 */
output [31:0] alu_operand_a_ex_o_t0;
wire [31:0] alu_operand_a_ex_o_t0;
/* src = "generated/sv2v_out.v:17223.21-17223.39" */
output [31:0] alu_operand_b_ex_o;
wire [31:0] alu_operand_b_ex_o;
/* cellift = 32'd1 */
output [31:0] alu_operand_b_ex_o_t0;
wire [31:0] alu_operand_b_ex_o_t0;
/* src = "generated/sv2v_out.v:17221.20-17221.37" */
output [6:0] alu_operator_ex_o;
wire [6:0] alu_operator_ex_o;
/* cellift = 32'd1 */
output [6:0] alu_operator_ex_o_t0;
wire [6:0] alu_operator_ex_o_t0;
/* src = "generated/sv2v_out.v:17208.13-17208.30" */
input branch_decision_i;
wire branch_decision_i;
/* cellift = 32'd1 */
input branch_decision_i_t0;
wire branch_decision_i_t0;
/* src = "generated/sv2v_out.v:17317.7-17317.20" */
wire branch_in_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17317.7-17317.20" */
wire branch_in_dec_t0;
/* src = "generated/sv2v_out.v:17322.7-17322.29" */
wire branch_jump_set_done_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17322.7-17322.29" */
wire branch_jump_set_done_d_t0;
/* src = "generated/sv2v_out.v:17321.6-17321.28" */
reg branch_jump_set_done_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17321.6-17321.28" */
reg branch_jump_set_done_q_t0;
/* src = "generated/sv2v_out.v:17323.6-17323.20" */
wire branch_not_set;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17323.6-17323.20" */
wire branch_not_set_t0;
/* src = "generated/sv2v_out.v:17318.7-17318.17" */
wire branch_set;
/* src = "generated/sv2v_out.v:17319.7-17319.21" */
reg branch_set_raw;
/* src = "generated/sv2v_out.v:17320.6-17320.22" */
wire branch_set_raw_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17320.6-17320.22" */
wire branch_set_raw_d_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17319.7-17319.21" */
reg branch_set_raw_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17318.7-17318.17" */
wire branch_set_t0;
/* src = "generated/sv2v_out.v:17324.7-17324.19" */
wire branch_taken;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17324.7-17324.19" */
wire branch_taken_t0;
/* src = "generated/sv2v_out.v:17373.13-17373.25" */
/* unused_bits = "0 1" */
wire [1:0] bt_a_mux_sel;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17373.13-17373.25" */
/* unused_bits = "0 1" */
wire [1:0] bt_a_mux_sel_t0;
/* src = "generated/sv2v_out.v:17227.20-17227.34" */
output [31:0] bt_a_operand_o;
wire [31:0] bt_a_operand_o;
/* cellift = 32'd1 */
output [31:0] bt_a_operand_o_t0;
wire [31:0] bt_a_operand_o_t0;
/* src = "generated/sv2v_out.v:17374.13-17374.25" */
/* unused_bits = "0 1 2" */
wire [2:0] bt_b_mux_sel;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17374.13-17374.25" */
/* unused_bits = "0 1 2" */
wire [2:0] bt_b_mux_sel_t0;
/* src = "generated/sv2v_out.v:17228.20-17228.34" */
output [31:0] bt_b_operand_o;
wire [31:0] bt_b_operand_o;
/* cellift = 32'd1 */
output [31:0] bt_b_operand_o_t0;
wire [31:0] bt_b_operand_o_t0;
/* src = "generated/sv2v_out.v:17192.13-17192.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:17333.7-17333.21" */
wire controller_run;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17333.7-17333.21" */
wire controller_run_t0;
/* src = "generated/sv2v_out.v:17238.14-17238.26" */
output csr_access_o;
wire csr_access_o;
/* cellift = 32'd1 */
output csr_access_o_t0;
wire csr_access_o_t0;
/* src = "generated/sv2v_out.v:17260.13-17260.30" */
input csr_mstatus_mie_i;
wire csr_mstatus_mie_i;
/* cellift = 32'd1 */
input csr_mstatus_mie_i_t0;
wire csr_mstatus_mie_i_t0;
/* src = "generated/sv2v_out.v:17249.13-17249.29" */
input csr_mstatus_tw_i;
wire csr_mstatus_tw_i;
/* cellift = 32'd1 */
input csr_mstatus_tw_i_t0;
wire csr_mstatus_tw_i_t0;
/* src = "generated/sv2v_out.v:17247.21-17247.32" */
output [31:0] csr_mtval_o;
wire [31:0] csr_mtval_o;
/* cellift = 32'd1 */
output [31:0] csr_mtval_o_t0;
wire [31:0] csr_mtval_o_t0;
/* src = "generated/sv2v_out.v:17240.14-17240.25" */
output csr_op_en_o;
wire csr_op_en_o;
/* cellift = 32'd1 */
output csr_op_en_o_t0;
wire csr_op_en_o_t0;
/* src = "generated/sv2v_out.v:17239.20-17239.28" */
output [1:0] csr_op_o;
wire [1:0] csr_op_o;
/* cellift = 32'd1 */
output [1:0] csr_op_o_t0;
wire [1:0] csr_op_o_t0;
/* src = "generated/sv2v_out.v:17391.6-17391.20" */
wire csr_pipe_flush;
/* src = "generated/sv2v_out.v:17279.20-17279.31" */
input [31:0] csr_rdata_i;
wire [31:0] csr_rdata_i;
/* cellift = 32'd1 */
input [31:0] csr_rdata_i_t0;
wire [31:0] csr_rdata_i_t0;
/* src = "generated/sv2v_out.v:17245.14-17245.35" */
output csr_restore_dret_id_o;
wire csr_restore_dret_id_o;
/* cellift = 32'd1 */
output csr_restore_dret_id_o_t0;
wire csr_restore_dret_id_o_t0;
/* src = "generated/sv2v_out.v:17244.14-17244.35" */
output csr_restore_mret_id_o;
wire csr_restore_mret_id_o;
/* cellift = 32'd1 */
output csr_restore_mret_id_o_t0;
wire csr_restore_mret_id_o_t0;
/* src = "generated/sv2v_out.v:17246.14-17246.30" */
output csr_save_cause_o;
wire csr_save_cause_o;
/* cellift = 32'd1 */
output csr_save_cause_o_t0;
wire csr_save_cause_o_t0;
/* src = "generated/sv2v_out.v:17242.14-17242.27" */
output csr_save_id_o;
wire csr_save_id_o;
/* cellift = 32'd1 */
output csr_save_id_o_t0;
wire csr_save_id_o_t0;
/* src = "generated/sv2v_out.v:17241.14-17241.27" */
output csr_save_if_o;
wire csr_save_if_o;
/* cellift = 32'd1 */
output csr_save_if_o_t0;
wire csr_save_if_o_t0;
/* src = "generated/sv2v_out.v:17243.14-17243.27" */
output csr_save_wb_o;
wire csr_save_wb_o;
/* cellift = 32'd1 */
output csr_save_wb_o_t0;
wire csr_save_wb_o_t0;
/* src = "generated/sv2v_out.v:17194.14-17194.25" */
output ctrl_busy_o;
wire ctrl_busy_o;
/* cellift = 32'd1 */
output ctrl_busy_o_t0;
wire ctrl_busy_o_t0;
/* src = "generated/sv2v_out.v:17251.13-17251.30" */
input data_ind_timing_i;
wire data_ind_timing_i;
/* cellift = 32'd1 */
input data_ind_timing_i_t0;
wire data_ind_timing_i_t0;
/* src = "generated/sv2v_out.v:17390.7-17390.23" */
wire data_req_allowed;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17390.7-17390.23" */
wire data_req_allowed_t0;
/* src = "generated/sv2v_out.v:17271.20-17271.33" */
output [2:0] debug_cause_o;
wire [2:0] debug_cause_o;
/* cellift = 32'd1 */
output [2:0] debug_cause_o_t0;
wire [2:0] debug_cause_o_t0;
/* src = "generated/sv2v_out.v:17272.14-17272.30" */
output debug_csr_save_o;
wire debug_csr_save_o;
/* cellift = 32'd1 */
output debug_csr_save_o_t0;
wire debug_csr_save_o_t0;
/* src = "generated/sv2v_out.v:17275.13-17275.28" */
input debug_ebreakm_i;
wire debug_ebreakm_i;
/* cellift = 32'd1 */
input debug_ebreakm_i_t0;
wire debug_ebreakm_i_t0;
/* src = "generated/sv2v_out.v:17276.13-17276.28" */
input debug_ebreaku_i;
wire debug_ebreaku_i;
/* cellift = 32'd1 */
input debug_ebreaku_i_t0;
wire debug_ebreaku_i_t0;
/* src = "generated/sv2v_out.v:17270.14-17270.35" */
output debug_mode_entering_o;
wire debug_mode_entering_o;
/* cellift = 32'd1 */
output debug_mode_entering_o_t0;
wire debug_mode_entering_o_t0;
/* src = "generated/sv2v_out.v:17269.14-17269.26" */
output debug_mode_o;
wire debug_mode_o;
/* cellift = 32'd1 */
output debug_mode_o_t0;
wire debug_mode_o_t0;
/* src = "generated/sv2v_out.v:17273.13-17273.24" */
input debug_req_i;
wire debug_req_i;
/* cellift = 32'd1 */
input debug_req_i_t0;
wire debug_req_i_t0;
/* src = "generated/sv2v_out.v:17274.13-17274.32" */
input debug_single_step_i;
wire debug_single_step_i;
/* cellift = 32'd1 */
input debug_single_step_i_t0;
wire debug_single_step_i_t0;
/* src = "generated/sv2v_out.v:17381.7-17381.17" */
wire div_en_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17381.7-17381.17" */
wire div_en_dec_t0;
/* src = "generated/sv2v_out.v:17230.14-17230.25" */
output div_en_ex_o;
wire div_en_ex_o;
/* cellift = 32'd1 */
output div_en_ex_o_t0;
wire div_en_ex_o_t0;
/* src = "generated/sv2v_out.v:17232.14-17232.26" */
output div_sel_ex_o;
wire div_sel_ex_o;
/* cellift = 32'd1 */
output div_sel_ex_o_t0;
wire div_sel_ex_o_t0;
/* src = "generated/sv2v_out.v:17312.7-17312.20" */
wire dret_insn_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17312.7-17312.20" */
wire dret_insn_dec_t0;
/* src = "generated/sv2v_out.v:17310.7-17310.16" */
wire ebrk_insn;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17310.7-17310.16" */
wire ebrk_insn_t0;
/* src = "generated/sv2v_out.v:17313.7-17313.21" */
wire ecall_insn_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17313.7-17313.21" */
wire ecall_insn_dec_t0;
/* src = "generated/sv2v_out.v:17294.14-17294.21" */
output en_wb_o;
wire en_wb_o;
/* cellift = 32'd1 */
output en_wb_o_t0;
wire en_wb_o_t0;
/* src = "generated/sv2v_out.v:17219.13-17219.23" */
input ex_valid_i;
wire ex_valid_i;
/* cellift = 32'd1 */
input ex_valid_i_t0;
wire ex_valid_i_t0;
/* src = "generated/sv2v_out.v:17214.20-17214.31" */
output [6:0] exc_cause_o;
wire [6:0] exc_cause_o;
/* cellift = 32'd1 */
output [6:0] exc_cause_o_t0;
wire [6:0] exc_cause_o_t0;
/* src = "generated/sv2v_out.v:17213.20-17213.32" */
output [1:0] exc_pc_mux_o;
wire [1:0] exc_pc_mux_o;
/* cellift = 32'd1 */
output [1:0] exc_pc_mux_o_t0;
wire [1:0] exc_pc_mux_o_t0;
/* src = "generated/sv2v_out.v:17341.7-17341.15" */
wire flush_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17341.7-17341.15" */
wire flush_id_t0;
/* src = "generated/sv2v_out.v:17667.8-17667.22" */
reg \g_sec_branch_taken.branch_taken_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17667.8-17667.22" */
reg \g_sec_branch_taken.branch_taken_q_t0 ;
/* src = "generated/sv2v_out.v:17765.9-17765.19" */
wire \gen_stall_mem.instr_kill ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17765.9-17765.19" */
wire \gen_stall_mem.instr_kill_t0 ;
/* src = "generated/sv2v_out.v:17764.9-17764.34" */
wire \gen_stall_mem.outstanding_memory_access ;
/* src = "generated/sv2v_out.v:17762.9-17762.19" */
wire \gen_stall_mem.rf_rd_a_hz ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17762.9-17762.19" */
wire \gen_stall_mem.rf_rd_a_hz_t0 ;
/* src = "generated/sv2v_out.v:17763.9-17763.19" */
wire \gen_stall_mem.rf_rd_b_hz ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17763.9-17763.19" */
wire \gen_stall_mem.rf_rd_b_hz_t0 ;
/* src = "generated/sv2v_out.v:17207.14-17207.28" */
output icache_inval_o;
wire icache_inval_o;
/* cellift = 32'd1 */
output icache_inval_o_t0;
wire icache_inval_o_t0;
/* src = "generated/sv2v_out.v:17316.7-17316.19" */
wire id_exception;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17316.7-17316.19" */
wire id_exception_t0;
/* src = "generated/sv2v_out.v:17685.6-17685.14" */
reg id_fsm_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17685.6-17685.14" */
reg id_fsm_q_t0;
/* src = "generated/sv2v_out.v:17205.14-17205.27" */
output id_in_ready_o;
wire id_in_ready_o;
/* cellift = 32'd1 */
output id_in_ready_o_t0;
wire id_in_ready_o_t0;
/* src = "generated/sv2v_out.v:17215.13-17215.29" */
input illegal_c_insn_i;
wire illegal_c_insn_i;
/* cellift = 32'd1 */
input illegal_c_insn_i_t0;
wire illegal_c_insn_i_t0;
/* src = "generated/sv2v_out.v:17250.13-17250.31" */
input illegal_csr_insn_i;
wire illegal_csr_insn_i;
/* cellift = 32'd1 */
input illegal_csr_insn_i_t0;
wire illegal_csr_insn_i_t0;
/* src = "generated/sv2v_out.v:17308.7-17308.24" */
wire illegal_dret_insn;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17308.7-17308.24" */
wire illegal_dret_insn_t0;
/* src = "generated/sv2v_out.v:17307.7-17307.23" */
wire illegal_insn_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17307.7-17307.23" */
wire illegal_insn_dec_t0;
/* src = "generated/sv2v_out.v:17195.14-17195.28" */
output illegal_insn_o;
wire illegal_insn_o;
/* cellift = 32'd1 */
output illegal_insn_o_t0;
wire illegal_insn_o_t0;
/* src = "generated/sv2v_out.v:17309.7-17309.25" */
wire illegal_umode_insn;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17309.7-17309.25" */
wire illegal_umode_insn_t0;
/* src = "generated/sv2v_out.v:17225.20-17225.34" */
input [67:0] imd_val_d_ex_i;
wire [67:0] imd_val_d_ex_i;
/* cellift = 32'd1 */
input [67:0] imd_val_d_ex_i_t0;
wire [67:0] imd_val_d_ex_i_t0;
/* src = "generated/sv2v_out.v:17226.21-17226.35" */
output [67:0] imd_val_q_ex_o;
reg [67:0] imd_val_q_ex_o;
/* cellift = 32'd1 */
output [67:0] imd_val_q_ex_o_t0;
reg [67:0] imd_val_q_ex_o_t0;
/* src = "generated/sv2v_out.v:17224.19-17224.34" */
input [1:0] imd_val_we_ex_i;
wire [1:0] imd_val_we_ex_i;
/* cellift = 32'd1 */
input [1:0] imd_val_we_ex_i_t0;
wire [1:0] imd_val_we_ex_i_t0;
/* src = "generated/sv2v_out.v:17350.14-17350.19" */
wire [31:0] imm_a;
/* src = "generated/sv2v_out.v:17375.7-17375.20" */
wire imm_a_mux_sel;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17375.7-17375.20" */
/* unused_bits = "0" */
wire imm_a_mux_sel_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17350.14-17350.19" */
wire [31:0] imm_a_t0;
/* src = "generated/sv2v_out.v:17351.13-17351.18" */
wire [31:0] imm_b;
/* src = "generated/sv2v_out.v:17376.13-17376.26" */
wire [2:0] imm_b_mux_sel;
/* src = "generated/sv2v_out.v:17377.13-17377.30" */
wire [2:0] imm_b_mux_sel_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17377.13-17377.30" */
/* unused_bits = "0 1 2" */
wire [2:0] imm_b_mux_sel_dec_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17351.13-17351.18" */
wire [31:0] imm_b_t0;
/* src = "generated/sv2v_out.v:17346.14-17346.24" */
wire [31:0] imm_b_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17346.14-17346.24" */
wire [31:0] imm_b_type_t0;
/* src = "generated/sv2v_out.v:17344.14-17344.24" */
wire [31:0] imm_i_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17344.14-17344.24" */
wire [31:0] imm_i_type_t0;
/* src = "generated/sv2v_out.v:17348.14-17348.24" */
wire [31:0] imm_j_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17348.14-17348.24" */
wire [31:0] imm_j_type_t0;
/* src = "generated/sv2v_out.v:17345.14-17345.24" */
wire [31:0] imm_s_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17345.14-17345.24" */
wire [31:0] imm_s_type_t0;
/* src = "generated/sv2v_out.v:17347.14-17347.24" */
wire [31:0] imm_u_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17347.14-17347.24" */
wire [31:0] imm_u_type_t0;
/* src = "generated/sv2v_out.v:17201.13-17201.29" */
input instr_bp_taken_i;
wire instr_bp_taken_i;
/* cellift = 32'd1 */
input instr_bp_taken_i_t0;
wire instr_bp_taken_i_t0;
/* src = "generated/sv2v_out.v:17206.13-17206.25" */
input instr_exec_i;
wire instr_exec_i;
/* cellift = 32'd1 */
input instr_exec_i_t0;
wire instr_exec_i_t0;
/* src = "generated/sv2v_out.v:17331.7-17331.22" */
wire instr_executing;
/* src = "generated/sv2v_out.v:17330.7-17330.27" */
wire instr_executing_spec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17331.7-17331.22" */
wire instr_executing_t0;
/* src = "generated/sv2v_out.v:17216.13-17216.30" */
input instr_fetch_err_i;
wire instr_fetch_err_i;
/* cellift = 32'd1 */
input instr_fetch_err_i_t0;
wire instr_fetch_err_i_t0;
/* src = "generated/sv2v_out.v:17217.13-17217.36" */
input instr_fetch_err_plus2_i;
wire instr_fetch_err_plus2_i;
/* cellift = 32'd1 */
input instr_fetch_err_plus2_i_t0;
wire instr_fetch_err_plus2_i_t0;
/* src = "generated/sv2v_out.v:17203.14-17203.36" */
output instr_first_cycle_id_o;
wire instr_first_cycle_id_o;
/* cellift = 32'd1 */
output instr_first_cycle_id_o_t0;
wire instr_first_cycle_id_o_t0;
/* src = "generated/sv2v_out.v:17306.14-17306.29" */
output instr_id_done_o;
wire instr_id_done_o;
/* cellift = 32'd1 */
output instr_id_done_o_t0;
wire instr_id_done_o_t0;
/* src = "generated/sv2v_out.v:17200.13-17200.34" */
input instr_is_compressed_i;
wire instr_is_compressed_i;
/* cellift = 32'd1 */
input instr_is_compressed_i_t0;
wire instr_is_compressed_i_t0;
/* src = "generated/sv2v_out.v:17296.14-17296.35" */
output instr_perf_count_id_o;
wire instr_perf_count_id_o;
/* cellift = 32'd1 */
output instr_perf_count_id_o_t0;
wire instr_perf_count_id_o_t0;
/* src = "generated/sv2v_out.v:17198.20-17198.37" */
input [31:0] instr_rdata_alu_i;
wire [31:0] instr_rdata_alu_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_alu_i_t0;
wire [31:0] instr_rdata_alu_i_t0;
/* src = "generated/sv2v_out.v:17199.20-17199.35" */
input [15:0] instr_rdata_c_i;
wire [15:0] instr_rdata_c_i;
/* cellift = 32'd1 */
input [15:0] instr_rdata_c_i_t0;
wire [15:0] instr_rdata_c_i_t0;
/* src = "generated/sv2v_out.v:17197.20-17197.33" */
input [31:0] instr_rdata_i;
wire [31:0] instr_rdata_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_i_t0;
wire [31:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:17202.14-17202.25" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:17295.20-17295.35" */
output [1:0] instr_type_wb_o;
wire [1:0] instr_type_wb_o;
/* cellift = 32'd1 */
output [1:0] instr_type_wb_o_t0;
wire [1:0] instr_type_wb_o_t0;
/* src = "generated/sv2v_out.v:17204.14-17204.33" */
output instr_valid_clear_o;
wire instr_valid_clear_o;
/* cellift = 32'd1 */
output instr_valid_clear_o_t0;
wire instr_valid_clear_o_t0;
/* src = "generated/sv2v_out.v:17196.13-17196.26" */
input instr_valid_i;
wire instr_valid_i;
/* cellift = 32'd1 */
input instr_valid_i_t0;
wire instr_valid_i_t0;
/* src = "generated/sv2v_out.v:17263.13-17263.21" */
input irq_nm_i;
wire irq_nm_i;
/* cellift = 32'd1 */
input irq_nm_i_t0;
wire irq_nm_i_t0;
/* src = "generated/sv2v_out.v:17261.13-17261.26" */
input irq_pending_i;
wire irq_pending_i;
/* cellift = 32'd1 */
input irq_pending_i_t0;
wire irq_pending_i_t0;
/* src = "generated/sv2v_out.v:17262.20-17262.26" */
input [17:0] irqs_i;
wire [17:0] irqs_i;
/* cellift = 32'd1 */
input [17:0] irqs_i_t0;
wire [17:0] irqs_i_t0;
/* src = "generated/sv2v_out.v:17325.7-17325.18" */
wire jump_in_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17325.7-17325.18" */
wire jump_in_dec_t0;
/* src = "generated/sv2v_out.v:17327.7-17327.15" */
wire jump_set;
/* src = "generated/sv2v_out.v:17326.7-17326.19" */
wire jump_set_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17326.7-17326.19" */
wire jump_set_dec_t0;
/* src = "generated/sv2v_out.v:17328.6-17328.18" */
wire jump_set_raw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17328.6-17328.18" */
wire jump_set_raw_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17327.7-17327.15" */
wire jump_set_t0;
/* src = "generated/sv2v_out.v:17258.13-17258.32" */
input lsu_addr_incr_req_i;
wire lsu_addr_incr_req_i;
/* cellift = 32'd1 */
input lsu_addr_incr_req_i_t0;
wire lsu_addr_incr_req_i_t0;
/* src = "generated/sv2v_out.v:17259.20-17259.35" */
input [31:0] lsu_addr_last_i;
wire [31:0] lsu_addr_last_i;
/* cellift = 32'd1 */
input [31:0] lsu_addr_last_i_t0;
wire [31:0] lsu_addr_last_i_t0;
/* src = "generated/sv2v_out.v:17265.13-17265.27" */
input lsu_load_err_i;
wire lsu_load_err_i;
/* cellift = 32'd1 */
input lsu_load_err_i_t0;
wire lsu_load_err_i_t0;
/* src = "generated/sv2v_out.v:17266.13-17266.37" */
input lsu_load_resp_intg_err_i;
wire lsu_load_resp_intg_err_i;
/* cellift = 32'd1 */
input lsu_load_resp_intg_err_i_t0;
wire lsu_load_resp_intg_err_i_t0;
/* src = "generated/sv2v_out.v:17389.7-17389.18" */
wire lsu_req_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17389.7-17389.18" */
wire lsu_req_dec_t0;
/* src = "generated/sv2v_out.v:17257.13-17257.27" */
input lsu_req_done_i;
wire lsu_req_done_i;
/* cellift = 32'd1 */
input lsu_req_done_i_t0;
wire lsu_req_done_i_t0;
/* src = "generated/sv2v_out.v:17252.14-17252.23" */
output lsu_req_o;
wire lsu_req_o;
/* cellift = 32'd1 */
output lsu_req_o_t0;
wire lsu_req_o_t0;
/* src = "generated/sv2v_out.v:17220.13-17220.29" */
input lsu_resp_valid_i;
wire lsu_resp_valid_i;
/* cellift = 32'd1 */
input lsu_resp_valid_i_t0;
wire lsu_resp_valid_i_t0;
/* src = "generated/sv2v_out.v:17255.14-17255.28" */
output lsu_sign_ext_o;
wire lsu_sign_ext_o;
/* cellift = 32'd1 */
output lsu_sign_ext_o_t0;
wire lsu_sign_ext_o_t0;
/* src = "generated/sv2v_out.v:17267.13-17267.28" */
input lsu_store_err_i;
wire lsu_store_err_i;
/* cellift = 32'd1 */
input lsu_store_err_i_t0;
wire lsu_store_err_i_t0;
/* src = "generated/sv2v_out.v:17268.13-17268.38" */
input lsu_store_resp_intg_err_i;
wire lsu_store_resp_intg_err_i;
/* cellift = 32'd1 */
input lsu_store_resp_intg_err_i_t0;
wire lsu_store_resp_intg_err_i_t0;
/* src = "generated/sv2v_out.v:17254.20-17254.30" */
output [1:0] lsu_type_o;
wire [1:0] lsu_type_o;
/* cellift = 32'd1 */
output [1:0] lsu_type_o_t0;
wire [1:0] lsu_type_o_t0;
/* src = "generated/sv2v_out.v:17256.21-17256.32" */
output [31:0] lsu_wdata_o;
wire [31:0] lsu_wdata_o;
/* cellift = 32'd1 */
output [31:0] lsu_wdata_o_t0;
wire [31:0] lsu_wdata_o_t0;
/* src = "generated/sv2v_out.v:17253.14-17253.22" */
output lsu_we_o;
wire lsu_we_o;
/* cellift = 32'd1 */
output lsu_we_o_t0;
wire lsu_we_o_t0;
/* src = "generated/sv2v_out.v:17343.7-17343.24" */
wire mem_resp_intg_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17343.7-17343.24" */
wire mem_resp_intg_err_t0;
/* src = "generated/sv2v_out.v:17311.7-17311.20" */
wire mret_insn_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17311.7-17311.20" */
wire mret_insn_dec_t0;
/* src = "generated/sv2v_out.v:17379.7-17379.18" */
wire mult_en_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17379.7-17379.18" */
wire mult_en_dec_t0;
/* src = "generated/sv2v_out.v:17229.14-17229.26" */
output mult_en_ex_o;
wire mult_en_ex_o;
/* cellift = 32'd1 */
output mult_en_ex_o_t0;
wire mult_en_ex_o_t0;
/* src = "generated/sv2v_out.v:17231.14-17231.27" */
output mult_sel_ex_o;
wire mult_sel_ex_o;
/* cellift = 32'd1 */
output mult_sel_ex_o_t0;
wire mult_sel_ex_o_t0;
/* src = "generated/sv2v_out.v:17382.7-17382.21" */
wire multdiv_en_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17382.7-17382.21" */
wire multdiv_en_dec_t0;
/* src = "generated/sv2v_out.v:17235.21-17235.43" */
output [31:0] multdiv_operand_a_ex_o;
wire [31:0] multdiv_operand_a_ex_o;
/* cellift = 32'd1 */
output [31:0] multdiv_operand_a_ex_o_t0;
wire [31:0] multdiv_operand_a_ex_o_t0;
/* src = "generated/sv2v_out.v:17236.21-17236.43" */
output [31:0] multdiv_operand_b_ex_o;
wire [31:0] multdiv_operand_b_ex_o;
/* cellift = 32'd1 */
output [31:0] multdiv_operand_b_ex_o_t0;
wire [31:0] multdiv_operand_b_ex_o_t0;
/* src = "generated/sv2v_out.v:17233.20-17233.41" */
output [1:0] multdiv_operator_ex_o;
wire [1:0] multdiv_operator_ex_o;
/* cellift = 32'd1 */
output [1:0] multdiv_operator_ex_o_t0;
wire [1:0] multdiv_operator_ex_o_t0;
/* src = "generated/sv2v_out.v:17237.14-17237.32" */
output multdiv_ready_id_o;
wire multdiv_ready_id_o;
/* cellift = 32'd1 */
output multdiv_ready_id_o_t0;
wire multdiv_ready_id_o_t0;
/* src = "generated/sv2v_out.v:17234.20-17234.44" */
output [1:0] multdiv_signed_mode_ex_o;
wire [1:0] multdiv_signed_mode_ex_o;
/* cellift = 32'd1 */
output [1:0] multdiv_signed_mode_ex_o_t0;
wire [1:0] multdiv_signed_mode_ex_o_t0;
/* src = "generated/sv2v_out.v:17342.7-17342.22" */
wire multicycle_done;
/* src = "generated/sv2v_out.v:17264.14-17264.24" */
output nmi_mode_o;
wire nmi_mode_o;
/* cellift = 32'd1 */
output nmi_mode_o_t0;
wire nmi_mode_o_t0;
/* src = "generated/sv2v_out.v:17212.21-17212.37" */
output [31:0] nt_branch_addr_o;
wire [31:0] nt_branch_addr_o;
/* cellift = 32'd1 */
output [31:0] nt_branch_addr_o_t0;
wire [31:0] nt_branch_addr_o_t0;
/* src = "generated/sv2v_out.v:17211.14-17211.36" */
output nt_branch_mispredict_o;
wire nt_branch_mispredict_o;
/* cellift = 32'd1 */
output nt_branch_mispredict_o_t0;
wire nt_branch_mispredict_o_t0;
/* src = "generated/sv2v_out.v:17298.13-17298.34" */
input outstanding_load_wb_i;
wire outstanding_load_wb_i;
/* cellift = 32'd1 */
input outstanding_load_wb_i_t0;
wire outstanding_load_wb_i_t0;
/* src = "generated/sv2v_out.v:17299.13-17299.35" */
input outstanding_store_wb_i;
wire outstanding_store_wb_i;
/* cellift = 32'd1 */
input outstanding_store_wb_i_t0;
wire outstanding_store_wb_i_t0;
/* src = "generated/sv2v_out.v:17218.20-17218.27" */
input [31:0] pc_id_i;
wire [31:0] pc_id_i;
/* cellift = 32'd1 */
input [31:0] pc_id_i_t0;
wire [31:0] pc_id_i_t0;
/* src = "generated/sv2v_out.v:17210.20-17210.28" */
output [2:0] pc_mux_o;
wire [2:0] pc_mux_o;
/* cellift = 32'd1 */
output [2:0] pc_mux_o_t0;
wire [2:0] pc_mux_o_t0;
/* src = "generated/sv2v_out.v:17209.14-17209.22" */
output pc_set_o;
wire pc_set_o;
/* cellift = 32'd1 */
output pc_set_o_t0;
wire pc_set_o_t0;
/* src = "generated/sv2v_out.v:17301.13-17301.26" */
output perf_branch_o;
wire perf_branch_o;
/* cellift = 32'd1 */
output perf_branch_o_t0;
wire perf_branch_o_t0;
/* src = "generated/sv2v_out.v:17305.14-17305.29" */
output perf_div_wait_o;
wire perf_div_wait_o;
/* cellift = 32'd1 */
output perf_div_wait_o_t0;
wire perf_div_wait_o_t0;
/* src = "generated/sv2v_out.v:17303.14-17303.31" */
output perf_dside_wait_o;
wire perf_dside_wait_o;
/* cellift = 32'd1 */
output perf_dside_wait_o_t0;
wire perf_dside_wait_o_t0;
/* src = "generated/sv2v_out.v:17300.14-17300.25" */
output perf_jump_o;
wire perf_jump_o;
/* cellift = 32'd1 */
output perf_jump_o_t0;
wire perf_jump_o_t0;
/* src = "generated/sv2v_out.v:17304.14-17304.29" */
output perf_mul_wait_o;
wire perf_mul_wait_o;
/* cellift = 32'd1 */
output perf_mul_wait_o_t0;
wire perf_mul_wait_o_t0;
/* src = "generated/sv2v_out.v:17302.14-17302.28" */
output perf_tbranch_o;
wire perf_tbranch_o;
/* cellift = 32'd1 */
output perf_tbranch_o_t0;
wire perf_tbranch_o_t0;
/* src = "generated/sv2v_out.v:17248.19-17248.30" */
input [1:0] priv_mode_i;
wire [1:0] priv_mode_i;
/* cellift = 32'd1 */
input [1:0] priv_mode_i_t0;
wire [1:0] priv_mode_i_t0;
/* src = "generated/sv2v_out.v:17297.13-17297.23" */
input ready_wb_i;
wire ready_wb_i;
/* cellift = 32'd1 */
input ready_wb_i_t0;
wire ready_wb_i_t0;
/* src = "generated/sv2v_out.v:17278.20-17278.31" */
input [31:0] result_ex_i;
wire [31:0] result_ex_i;
/* cellift = 32'd1 */
input [31:0] result_ex_i_t0;
wire [31:0] result_ex_i_t0;
/* src = "generated/sv2v_out.v:17280.20-17280.32" */
output [4:0] rf_raddr_a_o;
wire [4:0] rf_raddr_a_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_a_o_t0;
wire [4:0] rf_raddr_a_o_t0;
/* src = "generated/sv2v_out.v:17282.20-17282.32" */
output [4:0] rf_raddr_b_o;
wire [4:0] rf_raddr_b_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_b_o_t0;
wire [4:0] rf_raddr_b_o_t0;
/* src = "generated/sv2v_out.v:17289.14-17289.32" */
output rf_rd_a_wb_match_o;
wire rf_rd_a_wb_match_o;
/* cellift = 32'd1 */
output rf_rd_a_wb_match_o_t0;
wire rf_rd_a_wb_match_o_t0;
/* src = "generated/sv2v_out.v:17290.14-17290.32" */
output rf_rd_b_wb_match_o;
wire rf_rd_b_wb_match_o;
/* cellift = 32'd1 */
output rf_rd_b_wb_match_o_t0;
wire rf_rd_b_wb_match_o_t0;
/* src = "generated/sv2v_out.v:17281.20-17281.32" */
input [31:0] rf_rdata_a_i;
wire [31:0] rf_rdata_a_i;
/* cellift = 32'd1 */
input [31:0] rf_rdata_a_i_t0;
wire [31:0] rf_rdata_a_i_t0;
/* src = "generated/sv2v_out.v:17283.20-17283.32" */
input [31:0] rf_rdata_b_i;
wire [31:0] rf_rdata_b_i;
/* cellift = 32'd1 */
input [31:0] rf_rdata_b_i_t0;
wire [31:0] rf_rdata_b_i_t0;
/* src = "generated/sv2v_out.v:17357.7-17357.19" */
wire rf_ren_a_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17357.7-17357.19" */
wire rf_ren_a_dec_t0;
/* src = "generated/sv2v_out.v:17284.14-17284.24" */
output rf_ren_a_o;
wire rf_ren_a_o;
/* cellift = 32'd1 */
output rf_ren_a_o_t0;
wire rf_ren_a_o_t0;
/* src = "generated/sv2v_out.v:17358.7-17358.19" */
wire rf_ren_b_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17358.7-17358.19" */
wire rf_ren_b_dec_t0;
/* src = "generated/sv2v_out.v:17285.14-17285.24" */
output rf_ren_b_o;
wire rf_ren_b_o;
/* cellift = 32'd1 */
output rf_ren_b_o_t0;
wire rf_ren_b_o_t0;
/* src = "generated/sv2v_out.v:17286.20-17286.33" */
output [4:0] rf_waddr_id_o;
wire [4:0] rf_waddr_id_o;
/* cellift = 32'd1 */
output [4:0] rf_waddr_id_o_t0;
wire [4:0] rf_waddr_id_o_t0;
/* src = "generated/sv2v_out.v:17291.19-17291.32" */
input [4:0] rf_waddr_wb_i;
wire [4:0] rf_waddr_wb_i;
/* cellift = 32'd1 */
input [4:0] rf_waddr_wb_i_t0;
wire [4:0] rf_waddr_wb_i_t0;
/* src = "generated/sv2v_out.v:17292.20-17292.37" */
input [31:0] rf_wdata_fwd_wb_i;
wire [31:0] rf_wdata_fwd_wb_i;
/* cellift = 32'd1 */
input [31:0] rf_wdata_fwd_wb_i_t0;
wire [31:0] rf_wdata_fwd_wb_i_t0;
/* src = "generated/sv2v_out.v:17287.20-17287.33" */
output [31:0] rf_wdata_id_o;
wire [31:0] rf_wdata_id_o;
/* cellift = 32'd1 */
output [31:0] rf_wdata_id_o_t0;
wire [31:0] rf_wdata_id_o_t0;
/* src = "generated/sv2v_out.v:17352.7-17352.19" */
wire rf_wdata_sel;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17352.7-17352.19" */
/* unused_bits = "0" */
wire rf_wdata_sel_t0;
/* src = "generated/sv2v_out.v:17353.7-17353.16" */
wire rf_we_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17353.7-17353.16" */
wire rf_we_dec_t0;
/* src = "generated/sv2v_out.v:17288.14-17288.24" */
output rf_we_id_o;
wire rf_we_id_o;
/* cellift = 32'd1 */
output rf_we_id_o_t0;
wire rf_we_id_o_t0;
/* src = "generated/sv2v_out.v:17354.6-17354.15" */
wire rf_we_raw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17354.6-17354.15" */
wire rf_we_raw_t0;
/* src = "generated/sv2v_out.v:17293.13-17293.26" */
input rf_write_wb_i;
wire rf_write_wb_i;
/* cellift = 32'd1 */
input rf_write_wb_i_t0;
wire rf_write_wb_i_t0;
/* src = "generated/sv2v_out.v:17193.13-17193.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:17371.6-17371.15" */
wire stall_alu;
/* src = "generated/sv2v_out.v:17337.6-17337.18" */
wire stall_branch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17337.6-17337.18" */
wire stall_branch_t0;
/* src = "generated/sv2v_out.v:17339.7-17339.15" */
wire stall_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17339.7-17339.15" */
wire stall_id_t0;
/* src = "generated/sv2v_out.v:17338.6-17338.16" */
wire stall_jump;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17338.6-17338.16" */
wire stall_jump_t0;
/* src = "generated/sv2v_out.v:17334.7-17334.18" */
wire stall_ld_hz;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17334.7-17334.18" */
wire stall_ld_hz_t0;
/* src = "generated/sv2v_out.v:17335.7-17335.16" */
wire stall_mem;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17335.7-17335.16" */
wire stall_mem_t0;
/* src = "generated/sv2v_out.v:17336.6-17336.19" */
wire stall_multdiv;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17336.6-17336.19" */
wire stall_multdiv_t0;
/* src = "generated/sv2v_out.v:17340.7-17340.15" */
wire stall_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17340.7-17340.15" */
wire stall_wb_t0;
/* src = "generated/sv2v_out.v:17277.13-17277.28" */
input trigger_match_i;
wire trigger_match_i;
/* cellift = 32'd1 */
input trigger_match_i_t0;
wire trigger_match_i_t0;
/* src = "generated/sv2v_out.v:17315.7-17315.19" */
wire wb_exception;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17315.7-17315.19" */
wire wb_exception_t0;
/* src = "generated/sv2v_out.v:17314.7-17314.19" */
wire wfi_insn_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17314.7-17314.19" */
wire wfi_insn_dec_t0;
/* src = "generated/sv2v_out.v:17349.14-17349.27" */
wire [31:0] zimm_rs1_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17349.14-17349.27" */
wire [31:0] zimm_rs1_type_t0;
assign nt_branch_addr_o = pc_id_i + /* src = "generated/sv2v_out.v:17679.30-17679.79" */ _0145_;
assign rf_ren_a_o = _0049_ & /* src = "generated/sv2v_out.v:17359.20-17359.91" */ rf_ren_a_dec;
assign _0049_ = _0047_ & /* src = "generated/sv2v_out.v:17360.21-17360.75" */ _0455_;
assign rf_ren_b_o = _0049_ & /* src = "generated/sv2v_out.v:17360.20-17360.91" */ rf_ren_b_dec;
assign _0051_ = rf_we_raw & /* src = "generated/sv2v_out.v:17474.23-17474.50" */ instr_executing;
assign rf_we_id_o = _0051_ & /* src = "generated/sv2v_out.v:17474.22-17474.73" */ _0123_;
assign illegal_dret_insn = dret_insn_dec & /* src = "generated/sv2v_out.v:17549.29-17549.58" */ _0456_;
assign _0053_ = csr_mstatus_tw_i & /* src = "generated/sv2v_out.v:17550.73-17550.104" */ wfi_insn_dec;
assign illegal_umode_insn = _0454_ & /* src = "generated/sv2v_out.v:17550.30-17550.106" */ _0466_;
assign illegal_insn_o = instr_valid_i & /* src = "generated/sv2v_out.v:17551.26-17551.126" */ _0472_;
assign _0055_ = data_req_allowed & /* src = "generated/sv2v_out.v:17625.38-17625.68" */ lsu_req_dec;
assign _0057_ = csr_access_o & /* src = "generated/sv2v_out.v:17633.24-17633.54" */ instr_executing;
assign csr_op_en_o = _0057_ & /* src = "generated/sv2v_out.v:17633.23-17633.73" */ instr_id_done_o;
assign branch_jump_set_done_d = _0476_ & /* src = "generated/sv2v_out.v:17657.34-17657.115" */ _0457_;
assign jump_set = jump_set_raw & /* src = "generated/sv2v_out.v:17663.20-17663.58" */ _0129_;
assign branch_set = branch_set_raw & /* src = "generated/sv2v_out.v:17664.22-17664.62" */ _0129_;
assign _0059_ = rf_we_dec & /* src = "generated/sv2v_out.v:17741.19-17741.41" */ ex_valid_i;
assign _0061_ = multicycle_done & /* src = "generated/sv2v_out.v:17742.10-17742.38" */ ready_wb_i;
assign _0062_ = _0458_ & /* src = "generated/sv2v_out.v:17755.23-17755.44" */ _0459_;
assign en_wb_o = _0062_ & /* src = "generated/sv2v_out.v:17755.22-17755.63" */ instr_executing;
assign instr_first_cycle_id_o = instr_valid_i & /* src = "generated/sv2v_out.v:17756.29-17756.63" */ _0088_;
assign \gen_stall_mem.outstanding_memory_access  = _0488_ & /* src = "generated/sv2v_out.v:17767.39-17767.107" */ _0460_;
assign _0047_ = instr_valid_i & /* src = "generated/sv2v_out.v:17770.36-17770.70" */ _0118_;
assign _0064_ = _0047_ & /* src = "generated/sv2v_out.v:17770.35-17770.88" */ controller_run;
assign instr_executing_spec = _0064_ & /* src = "generated/sv2v_out.v:17770.34-17770.104" */ _0113_;
assign _0067_ = _0065_ & /* src = "generated/sv2v_out.v:17771.30-17771.74" */ _0113_;
assign instr_executing = _0067_ & /* src = "generated/sv2v_out.v:17771.29-17771.104" */ data_req_allowed;
assign _0069_ = lsu_req_dec & /* src = "generated/sv2v_out.v:17772.69-17772.98" */ _0095_;
assign stall_mem = instr_valid_i & /* src = "generated/sv2v_out.v:17772.23-17772.100" */ _0494_;
assign rf_rd_a_wb_match_o = _0441_ & /* src = "generated/sv2v_out.v:17773.30-17773.77" */ _0544_;
assign rf_rd_b_wb_match_o = _0442_ & /* src = "generated/sv2v_out.v:17774.30-17774.77" */ _0545_;
assign \gen_stall_mem.rf_rd_a_hz  = rf_rd_a_wb_match_o & /* src = "generated/sv2v_out.v:17777.24-17777.51" */ rf_ren_a_o;
assign \gen_stall_mem.rf_rd_b_hz  = rf_rd_b_wb_match_o & /* src = "generated/sv2v_out.v:17778.24-17778.51" */ rf_ren_b_o;
assign _0071_ = rf_rd_a_wb_match_o & /* src = "generated/sv2v_out.v:17779.29-17779.61" */ rf_write_wb_i;
assign _0072_ = rf_rd_b_wb_match_o & /* src = "generated/sv2v_out.v:17780.29-17780.61" */ rf_write_wb_i;
assign stall_ld_hz = outstanding_load_wb_i & /* src = "generated/sv2v_out.v:17781.25-17781.74" */ _0496_;
assign instr_id_done_o = en_wb_o & /* src = "generated/sv2v_out.v:17783.29-17783.49" */ ready_wb_i;
assign stall_wb = en_wb_o & /* src = "generated/sv2v_out.v:17784.22-17784.43" */ _0463_;
assign _0065_ = instr_valid_i & /* src = "generated/sv2v_out.v:17785.32-17785.59" */ _0462_;
assign perf_dside_wait_o = _0065_ & /* src = "generated/sv2v_out.v:17785.31-17785.104" */ _0498_;
assign _0073_ = _0464_ & /* src = "generated/sv2v_out.v:17820.36-17820.64" */ _0465_;
assign _0075_ = _0073_ & /* src = "generated/sv2v_out.v:17820.35-17820.85" */ _0106_;
assign _0077_ = _0075_ & /* src = "generated/sv2v_out.v:17820.34-17820.108" */ _0123_;
assign instr_perf_count_id_o = _0077_ & /* src = "generated/sv2v_out.v:17820.33-17820.130" */ _0118_;
assign perf_mul_wait_o = stall_multdiv & /* src = "generated/sv2v_out.v:17822.27-17822.54" */ mult_en_dec;
assign perf_div_wait_o = stall_multdiv & /* src = "generated/sv2v_out.v:17823.27-17823.53" */ div_en_dec;
assign _0079_ = ~ pc_id_i_t0;
assign _0144_ = pc_id_i & _0079_;
assign _0415_ = _0144_ + _0145_;
assign _0353_ = pc_id_i | pc_id_i_t0;
assign _0416_ = _0353_ + _0145_;
assign _0414_ = _0415_ ^ _0416_;
assign nt_branch_addr_o_t0 = _0414_ | pc_id_i_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$038d6e761af5e8bbfc2ed9b8473abfd849408d7b\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME \g_sec_branch_taken.branch_taken_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_sec_branch_taken.branch_taken_q_t0  <= 1'h0;
else \g_sec_branch_taken.branch_taken_q_t0  <= branch_decision_i_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$038d6e761af5e8bbfc2ed9b8473abfd849408d7b\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME branch_set_raw_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_set_raw_t0 <= 1'h0;
else branch_set_raw_t0 <= branch_set_raw_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$038d6e761af5e8bbfc2ed9b8473abfd849408d7b\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME branch_jump_set_done_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_jump_set_done_q_t0 <= 1'h0;
else branch_jump_set_done_q_t0 <= branch_jump_set_done_d_t0;
assign _0080_ = ~ imd_val_we_ex_i[1];
assign _0081_ = ~ imd_val_we_ex_i[0];
assign _0082_ = ~ _0143_;
assign _0248_ = { imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1] } & imd_val_d_ex_i_t0[33:0];
assign _0250_ = { imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0] } & imd_val_d_ex_i_t0[67:34];
assign _0249_ = { _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_ } & imd_val_q_ex_o_t0[33:0];
assign _0251_ = { _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_, _0081_ } & imd_val_q_ex_o_t0[67:34];
assign _0252_ = _0082_ & id_fsm_q_t0;
assign _0389_ = _0248_ | _0249_;
assign _0390_ = _0250_ | _0251_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$038d6e761af5e8bbfc2ed9b8473abfd849408d7b\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME imd_val_q_ex_o_t0[33:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) imd_val_q_ex_o_t0[33:0] <= 34'h000000000;
else imd_val_q_ex_o_t0[33:0] <= _0389_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$038d6e761af5e8bbfc2ed9b8473abfd849408d7b\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME imd_val_q_ex_o_t0[67:34] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) imd_val_q_ex_o_t0[67:34] <= 34'h000000000;
else imd_val_q_ex_o_t0[67:34] <= _0390_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$038d6e761af5e8bbfc2ed9b8473abfd849408d7b\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME id_fsm_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) id_fsm_q_t0 <= 1'h0;
else id_fsm_q_t0 <= _0252_;
assign _0146_ = _0050_ & rf_ren_a_dec;
assign _0149_ = _0048_ & _0455_;
assign _0152_ = _0050_ & rf_ren_b_dec;
assign _0155_ = rf_we_raw_t0 & instr_executing;
assign _0158_ = _0052_ & _0123_;
assign _0161_ = dret_insn_dec_t0 & _0456_;
assign _0164_ = csr_mstatus_tw_i_t0 & wfi_insn_dec;
assign _0167_ = instr_valid_i_t0 & _0472_;
assign _0170_ = data_req_allowed_t0 & lsu_req_dec;
assign _0173_ = csr_access_o_t0 & instr_executing;
assign _0176_ = _0058_ & instr_id_done_o;
assign _0179_ = _0477_ & _0457_;
assign _0182_ = jump_set_raw_t0 & _0129_;
assign _0185_ = branch_set_raw_t0 & _0129_;
assign _0036_ = rf_we_dec_t0 & ex_valid_i;
assign _0190_ = stall_id_t0 & _0459_;
assign _0193_ = _0063_ & instr_executing;
assign _0196_ = instr_valid_i_t0 & _0088_;
assign _0199_ = _0489_ & _0460_;
assign _0202_ = instr_valid_i_t0 & _0118_;
assign _0205_ = _0066_ & _0113_;
assign _0208_ = _0068_ & data_req_allowed;
assign _0211_ = lsu_req_dec_t0 & _0095_;
assign _0214_ = instr_valid_i_t0 & _0494_;
assign _0217_ = outstanding_load_wb_i_t0 & _0496_;
assign _0220_ = en_wb_o_t0 & ready_wb_i;
assign _0223_ = en_wb_o_t0 & _0463_;
assign _0224_ = instr_valid_i_t0 & _0462_;
assign _0227_ = _0066_ & _0498_;
assign _0230_ = ebrk_insn_t0 & _0465_;
assign _0233_ = _0074_ & _0106_;
assign _0236_ = _0076_ & _0123_;
assign _0239_ = _0078_ & _0118_;
assign _0242_ = stall_multdiv_t0 & mult_en_dec;
assign _0245_ = stall_multdiv_t0 & div_en_dec;
assign _0147_ = rf_ren_a_dec_t0 & _0049_;
assign _0150_ = illegal_insn_o_t0 & _0047_;
assign _0153_ = rf_ren_b_dec_t0 & _0049_;
assign _0156_ = instr_executing_t0 & rf_we_raw;
assign _0159_ = illegal_csr_insn_i_t0 & _0051_;
assign _0162_ = debug_mode_o_t0 & dret_insn_dec;
assign _0165_ = wfi_insn_dec_t0 & csr_mstatus_tw_i;
assign illegal_umode_insn_t0 = _0467_ & _0454_;
assign _0168_ = _0473_ & instr_valid_i;
assign _0171_ = lsu_req_dec_t0 & data_req_allowed;
assign _0174_ = instr_executing_t0 & csr_access_o;
assign _0177_ = instr_id_done_o_t0 & _0057_;
assign _0180_ = instr_valid_clear_o_t0 & _0476_;
assign _0183_ = branch_jump_set_done_q_t0 & jump_set_raw;
assign _0186_ = branch_jump_set_done_q_t0 & branch_set_raw;
assign _0188_ = ex_valid_i_t0 & rf_we_dec;
assign _0191_ = flush_id_t0 & _0458_;
assign _0194_ = instr_executing_t0 & _0062_;
assign _0197_ = id_fsm_q_t0 & instr_valid_i;
assign _0200_ = lsu_resp_valid_i_t0 & _0488_;
assign _0203_ = instr_fetch_err_i_t0 & instr_valid_i;
assign _0206_ = stall_ld_hz_t0 & _0065_;
assign _0209_ = data_req_allowed_t0 & _0067_;
assign _0212_ = lsu_req_done_i_t0 & lsu_req_dec;
assign _0215_ = _0495_ & instr_valid_i;
assign \gen_stall_mem.rf_rd_a_hz_t0  = rf_ren_a_o_t0 & rf_rd_a_wb_match_o;
assign \gen_stall_mem.rf_rd_b_hz_t0  = rf_ren_b_o_t0 & rf_rd_b_wb_match_o;
assign _0218_ = _0497_ & outstanding_load_wb_i;
assign _0221_ = ready_wb_i_t0 & en_wb_o;
assign _0225_ = \gen_stall_mem.instr_kill_t0  & instr_valid_i;
assign _0228_ = _0499_ & _0065_;
assign _0231_ = ecall_insn_dec_t0 & _0464_;
assign _0234_ = illegal_insn_dec_t0 & _0073_;
assign _0237_ = illegal_csr_insn_i_t0 & _0075_;
assign _0240_ = instr_fetch_err_i_t0 & _0077_;
assign _0243_ = mult_en_dec_t0 & stall_multdiv;
assign _0246_ = div_en_dec_t0 & stall_multdiv;
assign _0148_ = _0050_ & rf_ren_a_dec_t0;
assign _0151_ = _0048_ & illegal_insn_o_t0;
assign _0154_ = _0050_ & rf_ren_b_dec_t0;
assign _0157_ = rf_we_raw_t0 & instr_executing_t0;
assign _0160_ = _0052_ & illegal_csr_insn_i_t0;
assign _0163_ = dret_insn_dec_t0 & debug_mode_o_t0;
assign _0166_ = csr_mstatus_tw_i_t0 & wfi_insn_dec_t0;
assign _0169_ = instr_valid_i_t0 & _0473_;
assign _0172_ = data_req_allowed_t0 & lsu_req_dec_t0;
assign _0175_ = csr_access_o_t0 & instr_executing_t0;
assign _0178_ = _0058_ & instr_id_done_o_t0;
assign _0181_ = _0477_ & instr_valid_clear_o_t0;
assign _0184_ = jump_set_raw_t0 & branch_jump_set_done_q_t0;
assign _0187_ = branch_set_raw_t0 & branch_jump_set_done_q_t0;
assign _0189_ = rf_we_dec_t0 & ex_valid_i_t0;
assign _0192_ = stall_id_t0 & flush_id_t0;
assign _0195_ = _0063_ & instr_executing_t0;
assign _0198_ = instr_valid_i_t0 & id_fsm_q_t0;
assign _0201_ = _0489_ & lsu_resp_valid_i_t0;
assign _0204_ = instr_valid_i_t0 & instr_fetch_err_i_t0;
assign _0207_ = _0066_ & stall_ld_hz_t0;
assign _0210_ = _0068_ & data_req_allowed_t0;
assign _0213_ = lsu_req_dec_t0 & lsu_req_done_i_t0;
assign _0216_ = instr_valid_i_t0 & _0495_;
assign _0219_ = outstanding_load_wb_i_t0 & _0497_;
assign _0222_ = en_wb_o_t0 & ready_wb_i_t0;
assign _0226_ = instr_valid_i_t0 & \gen_stall_mem.instr_kill_t0 ;
assign _0229_ = _0066_ & _0499_;
assign _0232_ = ebrk_insn_t0 & ecall_insn_dec_t0;
assign _0235_ = _0074_ & illegal_insn_dec_t0;
assign _0238_ = _0076_ & illegal_csr_insn_i_t0;
assign _0241_ = _0078_ & instr_fetch_err_i_t0;
assign _0244_ = stall_multdiv_t0 & mult_en_dec_t0;
assign _0247_ = stall_multdiv_t0 & div_en_dec_t0;
assign _0354_ = _0146_ | _0147_;
assign _0355_ = _0149_ | _0150_;
assign _0356_ = _0152_ | _0153_;
assign _0357_ = _0155_ | _0156_;
assign _0358_ = _0158_ | _0159_;
assign _0359_ = _0161_ | _0162_;
assign _0360_ = _0164_ | _0165_;
assign _0361_ = _0167_ | _0168_;
assign _0362_ = _0170_ | _0171_;
assign _0363_ = _0173_ | _0174_;
assign _0364_ = _0176_ | _0177_;
assign _0365_ = _0179_ | _0180_;
assign _0366_ = _0182_ | _0183_;
assign _0367_ = _0185_ | _0186_;
assign _0368_ = _0036_ | _0188_;
assign _0369_ = _0190_ | _0191_;
assign _0370_ = _0193_ | _0194_;
assign _0371_ = _0196_ | _0197_;
assign _0372_ = _0199_ | _0200_;
assign _0373_ = _0202_ | _0203_;
assign _0374_ = _0205_ | _0206_;
assign _0375_ = _0208_ | _0209_;
assign _0376_ = _0211_ | _0212_;
assign _0377_ = _0214_ | _0215_;
assign _0378_ = _0217_ | _0218_;
assign _0379_ = _0220_ | _0221_;
assign _0380_ = _0223_ | _0221_;
assign _0381_ = _0224_ | _0225_;
assign _0382_ = _0227_ | _0228_;
assign _0383_ = _0230_ | _0231_;
assign _0384_ = _0233_ | _0234_;
assign _0385_ = _0236_ | _0237_;
assign _0386_ = _0239_ | _0240_;
assign _0387_ = _0242_ | _0243_;
assign _0388_ = _0245_ | _0246_;
assign rf_ren_a_o_t0 = _0354_ | _0148_;
assign _0050_ = _0355_ | _0151_;
assign rf_ren_b_o_t0 = _0356_ | _0154_;
assign _0052_ = _0357_ | _0157_;
assign rf_we_id_o_t0 = _0358_ | _0160_;
assign illegal_dret_insn_t0 = _0359_ | _0163_;
assign _0054_ = _0360_ | _0166_;
assign illegal_insn_o_t0 = _0361_ | _0169_;
assign _0056_ = _0362_ | _0172_;
assign _0058_ = _0363_ | _0175_;
assign csr_op_en_o_t0 = _0364_ | _0178_;
assign branch_jump_set_done_d_t0 = _0365_ | _0181_;
assign jump_set_t0 = _0366_ | _0184_;
assign branch_set_t0 = _0367_ | _0187_;
assign _0060_ = _0368_ | _0189_;
assign _0063_ = _0369_ | _0192_;
assign en_wb_o_t0 = _0370_ | _0195_;
assign instr_first_cycle_id_o_t0 = _0371_ | _0198_;
assign data_req_allowed_t0 = _0372_ | _0201_;
assign _0048_ = _0373_ | _0204_;
assign _0068_ = _0374_ | _0207_;
assign instr_executing_t0 = _0375_ | _0210_;
assign _0070_ = _0376_ | _0213_;
assign stall_mem_t0 = _0377_ | _0216_;
assign stall_ld_hz_t0 = _0378_ | _0219_;
assign instr_id_done_o_t0 = _0379_ | _0222_;
assign stall_wb_t0 = _0380_ | _0222_;
assign _0066_ = _0381_ | _0226_;
assign perf_dside_wait_o_t0 = _0382_ | _0229_;
assign _0074_ = _0383_ | _0232_;
assign _0076_ = _0384_ | _0235_;
assign _0078_ = _0385_ | _0238_;
assign instr_perf_count_id_o_t0 = _0386_ | _0241_;
assign perf_mul_wait_o_t0 = _0387_ | _0244_;
assign perf_div_wait_o_t0 = _0388_ | _0247_;
/* src = "generated/sv2v_out.v:17465.4-17470.7" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$038d6e761af5e8bbfc2ed9b8473abfd849408d7b\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME imd_val_q_ex_o[33:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) imd_val_q_ex_o[33:0] <= 34'h000000000;
else if (imd_val_we_ex_i[1]) imd_val_q_ex_o[33:0] <= imd_val_d_ex_i[33:0];
/* src = "generated/sv2v_out.v:17465.4-17470.7" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$038d6e761af5e8bbfc2ed9b8473abfd849408d7b\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME imd_val_q_ex_o[67:34] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) imd_val_q_ex_o[67:34] <= 34'h000000000;
else if (imd_val_we_ex_i[0]) imd_val_q_ex_o[67:34] <= imd_val_d_ex_i[67:34];
/* src = "generated/sv2v_out.v:17687.2-17692.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$038d6e761af5e8bbfc2ed9b8473abfd849408d7b\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME id_fsm_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) id_fsm_q <= 1'h0;
else if (_0143_) id_fsm_q <= _0005_;
assign _0083_ = ~ { _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_ };
assign _0084_ = ~ { _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_ };
assign _0085_ = ~ { _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_ };
assign _0086_ = ~ { _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_ };
assign _0087_ = ~ { _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_ };
assign _0088_ = ~ id_fsm_q;
assign _0089_ = ~ { rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel };
assign _0090_ = ~ { _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_ };
assign _0091_ = ~ { _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_ };
assign _0092_ = ~ { _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_ };
assign _0093_ = ~ _0061_;
assign _0094_ = ~ multdiv_en_dec;
assign _0095_ = ~ lsu_req_done_i;
assign _0096_ = ~ jump_in_dec;
assign _0097_ = ~ branch_in_dec;
assign _0098_ = ~ lsu_req_dec;
assign _0099_ = ~ alu_multicycle_dec;
assign _0100_ = ~ instr_executing_spec;
assign _0101_ = ~ { imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel };
assign _0102_ = ~ { alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel };
assign _0103_ = ~ { _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_ };
assign _0104_ = ~ { _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_ };
assign _0253_ = _0083_ & imm_u_type_t0;
assign _0420_ = _0084_ & _0418_;
assign _0255_ = _0085_ & imm_s_type_t0;
assign _0257_ = _0086_ & _0424_;
assign _0259_ = _0087_ & _0426_;
assign _0261_ = _0088_ & _0028_;
assign _0003_ = _0088_ & _0021_;
assign _0007_ = _0088_ & _0025_;
assign _0001_ = _0088_ & _0019_;
assign _0264_ = _0089_ & result_ex_i_t0;
assign _0266_ = _0090_ & pc_id_i_t0;
assign _0268_ = _0091_ & multdiv_operand_a_ex_o_t0;
assign _0270_ = _0092_ & _0430_;
assign _0040_ = _0093_ & jump_in_dec_t0;
assign _0038_ = _0093_ & branch_in_dec_t0;
assign _0045_ = _0093_ & multdiv_en_dec_t0;
assign _0335_ = _0094_ & rf_we_dec_t0;
assign _0514_ = _0099_ & rf_we_dec_t0;
assign _0337_ = _0096_ & _0514_;
assign _0339_ = _0097_ & _0516_;
assign _0341_ = _0094_ & _0518_;
assign _0343_ = _0098_ & _0520_;
assign _0527_ = _0094_ & _0525_;
assign _0532_ = _0097_ & _0530_;
assign _0534_ = _0094_ & _0532_;
assign _0025_ = _0098_ & _0534_;
assign _0538_ = _0094_ & _0536_;
assign _0019_ = _0098_ & _0538_;
assign _0021_ = _0098_ & _0527_;
assign _0345_ = _0100_ & rf_we_dec_t0;
assign imm_a_t0 = _0101_ & zimm_rs1_type_t0;
assign _0347_ = _0102_ & lsu_wdata_o_t0;
assign _0349_ = _0103_ & rf_rdata_a_i_t0;
assign _0351_ = _0104_ & rf_rdata_b_i_t0;
assign _0254_ = { _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_, _0501_ } & imm_j_type_t0;
assign _0256_ = { _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_ } & imm_b_type_t0;
assign _0424_ = { _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_ } & imm_i_type_t0;
assign _0258_ = { _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_, _0412_ } & _0422_;
assign _0260_ = { _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_, _0142_ } & _0420_;
assign _0262_ = id_fsm_q & _0043_;
assign _0015_ = id_fsm_q & _0040_;
assign _0263_ = id_fsm_q & _0038_;
assign _0017_ = id_fsm_q & _0045_;
assign _0265_ = { rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel } & csr_rdata_i_t0;
assign _0267_ = { _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_ } & imm_a_t0;
assign _0269_ = { _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_ } & lsu_addr_last_i_t0;
assign _0271_ = { _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_, _0413_ } & _0428_;
assign _0336_ = multdiv_en_dec & _0060_;
assign _0338_ = jump_in_dec & rf_we_dec_t0;
assign _0340_ = branch_in_dec & rf_we_dec_t0;
assign _0342_ = multdiv_en_dec & _0036_;
assign _0344_ = lsu_req_dec & rf_we_dec_t0;
assign _0525_ = branch_in_dec & _0479_;
assign _0530_ = jump_in_dec & jump_set_dec_t0;
assign _0536_ = branch_in_dec & branch_decision_i_t0;
assign _0346_ = instr_executing_spec & _0010_;
assign stall_jump_t0 = instr_executing_spec & _0015_;
assign stall_branch_t0 = instr_executing_spec & _0013_;
assign stall_multdiv_t0 = instr_executing_spec & _0017_;
assign jump_set_raw_t0 = instr_executing_spec & _0007_;
assign branch_not_set_t0 = instr_executing_spec & _0001_;
assign branch_set_raw_d_t0 = instr_executing_spec & _0003_;
assign _0348_ = { alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel } & imm_b_t0;
assign lsu_req_o_t0 = instr_executing & _0056_;
assign mult_en_ex_o_t0 = instr_executing & mult_en_dec_t0;
assign div_en_ex_o_t0 = instr_executing & div_en_dec_t0;
assign _0350_ = { _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_, _0071_ } & rf_wdata_fwd_wb_i_t0;
assign _0352_ = { _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_ } & rf_wdata_fwd_wb_i_t0;
assign _0418_ = _0253_ | _0254_;
assign _0422_ = _0255_ | _0256_;
assign _0426_ = _0257_ | _0258_;
assign imm_b_t0 = _0259_ | _0260_;
assign _0010_ = _0261_ | _0262_;
assign _0013_ = _0003_ | _0263_;
assign rf_wdata_id_o_t0 = _0264_ | _0265_;
assign _0428_ = _0266_ | _0267_;
assign _0430_ = _0268_ | _0269_;
assign alu_operand_a_ex_o_t0 = _0270_ | _0271_;
assign _0043_ = _0335_ | _0336_;
assign _0516_ = _0337_ | _0338_;
assign _0518_ = _0339_ | _0340_;
assign _0520_ = _0341_ | _0342_;
assign _0028_ = _0343_ | _0344_;
assign rf_we_raw_t0 = _0345_ | _0346_;
assign alu_operand_b_ex_o_t0 = _0347_ | _0348_;
assign multdiv_operand_a_ex_o_t0 = _0349_ | _0350_;
assign lsu_wdata_o_t0 = _0351_ | _0352_;
assign _0143_ = & { instr_executing, instr_executing_spec };
assign _0105_ = ~ mret_insn_dec;
assign _0106_ = ~ illegal_insn_dec;
assign _0107_ = ~ _0468_;
assign _0108_ = ~ _0470_;
assign _0109_ = ~ lsu_load_resp_intg_err_i;
assign _0110_ = ~ mult_en_dec;
assign _0111_ = ~ branch_set_raw;
assign _0112_ = ~ _0474_;
assign _0032_ = ~ branch_decision_i;
assign _0113_ = ~ stall_ld_hz;
assign _0114_ = ~ _0480_;
assign _0115_ = ~ _0482_;
assign _0116_ = ~ _0484_;
assign _0117_ = ~ outstanding_load_wb_i;
assign _0118_ = ~ instr_fetch_err_i;
assign _0119_ = ~ _0490_;
assign _0120_ = ~ _0492_;
assign data_req_allowed = ~ \gen_stall_mem.outstanding_memory_access ;
assign _0121_ = ~ \gen_stall_mem.rf_rd_a_hz ;
assign _0122_ = ~ _0053_;
assign _0123_ = ~ illegal_csr_insn_i;
assign _0124_ = ~ illegal_dret_insn;
assign _0125_ = ~ illegal_umode_insn;
assign _0126_ = ~ lsu_store_resp_intg_err_i;
assign _0127_ = ~ div_en_dec;
assign _0128_ = ~ jump_set_raw;
assign _0129_ = ~ branch_jump_set_done_q;
assign _0130_ = ~ \g_sec_branch_taken.branch_taken_q ;
assign _0131_ = ~ data_ind_timing_i;
assign _0132_ = ~ stall_mem;
assign _0133_ = ~ stall_multdiv;
assign _0134_ = ~ stall_jump;
assign _0135_ = ~ stall_branch;
assign _0136_ = ~ stall_alu;
assign _0137_ = ~ outstanding_store_wb_i;
assign _0138_ = ~ wb_exception;
assign _0139_ = ~ id_exception;
assign _0140_ = ~ _0069_;
assign _0141_ = ~ \gen_stall_mem.rf_rd_b_hz ;
assign _0272_ = mret_insn_dec_t0 & _0122_;
assign _0275_ = illegal_insn_dec_t0 & _0123_;
assign _0278_ = _0469_ & _0124_;
assign _0281_ = _0471_ & _0125_;
assign _0284_ = lsu_load_resp_intg_err_i_t0 & _0126_;
assign _0287_ = mult_en_dec_t0 & _0127_;
assign _0290_ = branch_set_raw_t0 & _0128_;
assign _0293_ = _0475_ & _0129_;
assign _0296_ = data_ind_timing_i_t0 & _0130_;
assign _0299_ = branch_decision_i_t0 & _0131_;
assign _0302_ = stall_ld_hz_t0 & _0132_;
assign _0305_ = _0481_ & _0133_;
assign _0308_ = _0483_ & _0134_;
assign _0311_ = _0485_ & _0135_;
assign stall_id_t0 = _0487_ & _0136_;
assign _0314_ = outstanding_load_wb_i_t0 & _0137_;
assign _0317_ = instr_fetch_err_i_t0 & _0138_;
assign _0320_ = _0491_ & _0139_;
assign _0323_ = _0493_ & controller_run;
assign _0326_ = data_req_allowed_t0 & _0140_;
assign _0329_ = \gen_stall_mem.rf_rd_a_hz_t0  & _0141_;
assign _0332_ = data_req_allowed_t0 & _0113_;
assign _0273_ = _0054_ & _0105_;
assign _0276_ = illegal_csr_insn_i_t0 & _0106_;
assign _0279_ = illegal_dret_insn_t0 & _0107_;
assign _0282_ = illegal_umode_insn_t0 & _0108_;
assign _0285_ = lsu_store_resp_intg_err_i_t0 & _0109_;
assign _0288_ = div_en_dec_t0 & _0110_;
assign _0291_ = jump_set_raw_t0 & _0111_;
assign _0294_ = branch_jump_set_done_q_t0 & _0112_;
assign _0297_ = \g_sec_branch_taken.branch_taken_q_t0  & data_ind_timing_i;
assign _0300_ = data_ind_timing_i_t0 & _0032_;
assign _0303_ = stall_mem_t0 & _0113_;
assign _0306_ = stall_multdiv_t0 & _0114_;
assign _0309_ = stall_jump_t0 & _0115_;
assign _0312_ = stall_branch_t0 & _0116_;
assign _0315_ = outstanding_store_wb_i_t0 & _0117_;
assign _0318_ = wb_exception_t0 & _0118_;
assign _0321_ = id_exception_t0 & _0119_;
assign _0324_ = controller_run_t0 & _0120_;
assign _0327_ = _0070_ & data_req_allowed;
assign _0330_ = \gen_stall_mem.rf_rd_b_hz_t0  & _0121_;
assign _0333_ = stall_ld_hz_t0 & data_req_allowed;
assign _0274_ = mret_insn_dec_t0 & _0054_;
assign _0277_ = illegal_insn_dec_t0 & illegal_csr_insn_i_t0;
assign _0280_ = _0469_ & illegal_dret_insn_t0;
assign _0283_ = _0471_ & illegal_umode_insn_t0;
assign _0286_ = lsu_load_resp_intg_err_i_t0 & lsu_store_resp_intg_err_i_t0;
assign _0289_ = mult_en_dec_t0 & div_en_dec_t0;
assign _0292_ = branch_set_raw_t0 & jump_set_raw_t0;
assign _0295_ = _0475_ & branch_jump_set_done_q_t0;
assign _0298_ = data_ind_timing_i_t0 & \g_sec_branch_taken.branch_taken_q_t0 ;
assign _0301_ = branch_decision_i_t0 & data_ind_timing_i_t0;
assign _0304_ = stall_ld_hz_t0 & stall_mem_t0;
assign _0307_ = _0481_ & stall_multdiv_t0;
assign _0310_ = _0483_ & stall_jump_t0;
assign _0313_ = _0485_ & stall_branch_t0;
assign _0316_ = outstanding_load_wb_i_t0 & outstanding_store_wb_i_t0;
assign _0319_ = instr_fetch_err_i_t0 & wb_exception_t0;
assign _0322_ = _0491_ & id_exception_t0;
assign _0325_ = _0493_ & controller_run_t0;
assign _0328_ = data_req_allowed_t0 & _0070_;
assign _0331_ = \gen_stall_mem.rf_rd_a_hz_t0  & \gen_stall_mem.rf_rd_b_hz_t0 ;
assign _0334_ = data_req_allowed_t0 & stall_ld_hz_t0;
assign _0391_ = _0272_ | _0273_;
assign _0392_ = _0275_ | _0276_;
assign _0393_ = _0278_ | _0279_;
assign _0394_ = _0281_ | _0282_;
assign _0395_ = _0284_ | _0285_;
assign _0396_ = _0287_ | _0288_;
assign _0397_ = _0290_ | _0291_;
assign _0398_ = _0293_ | _0294_;
assign _0399_ = _0296_ | _0297_;
assign _0400_ = _0299_ | _0300_;
assign _0401_ = _0302_ | _0303_;
assign _0402_ = _0305_ | _0306_;
assign _0403_ = _0308_ | _0309_;
assign _0404_ = _0311_ | _0312_;
assign _0405_ = _0314_ | _0315_;
assign _0406_ = _0317_ | _0318_;
assign _0407_ = _0320_ | _0321_;
assign _0408_ = _0323_ | _0324_;
assign _0409_ = _0326_ | _0327_;
assign _0410_ = _0329_ | _0330_;
assign _0411_ = _0332_ | _0333_;
assign _0467_ = _0391_ | _0274_;
assign _0469_ = _0392_ | _0277_;
assign _0471_ = _0393_ | _0280_;
assign _0473_ = _0394_ | _0283_;
assign mem_resp_intg_err_t0 = _0395_ | _0286_;
assign multdiv_en_dec_t0 = _0396_ | _0289_;
assign _0475_ = _0397_ | _0292_;
assign _0477_ = _0398_ | _0295_;
assign branch_taken_t0 = _0399_ | _0298_;
assign _0479_ = _0400_ | _0301_;
assign _0481_ = _0401_ | _0304_;
assign _0483_ = _0402_ | _0307_;
assign _0485_ = _0403_ | _0310_;
assign _0487_ = _0404_ | _0313_;
assign _0489_ = _0405_ | _0316_;
assign _0491_ = _0406_ | _0319_;
assign _0493_ = _0407_ | _0322_;
assign \gen_stall_mem.instr_kill_t0  = _0408_ | _0325_;
assign _0495_ = _0409_ | _0328_;
assign _0497_ = _0410_ | _0331_;
assign _0499_ = _0411_ | _0334_;
assign _0412_ = _0504_ | _0503_;
assign _0413_ = _0542_ | _0541_;
assign _0142_ = | { _0502_, _0501_, _0500_ };
assign _0417_ = _0501_ ? imm_j_type : imm_u_type;
assign _0419_ = _0500_ ? _0145_ : _0417_;
assign _0421_ = _0503_ ? imm_b_type : imm_s_type;
assign _0423_ = _0505_ ? imm_i_type : 32'd4;
assign _0425_ = _0412_ ? _0421_ : _0423_;
assign imm_b = _0142_ ? _0419_ : _0425_;
assign _0005_ = id_fsm_q ? _0046_ : _0023_;
assign _0011_ = id_fsm_q ? 1'h0 : _0029_;
assign _0009_ = id_fsm_q ? _0042_ : _0027_;
assign _0014_ = id_fsm_q ? _0039_ : _0030_;
assign _0012_ = id_fsm_q ? _0037_ : _0020_;
assign _0016_ = id_fsm_q ? _0044_ : _0031_;
assign _0006_ = id_fsm_q ? 1'h0 : _0024_;
assign _0000_ = id_fsm_q ? 1'h0 : _0018_;
assign _0002_ = id_fsm_q ? 1'h0 : _0020_;
assign _0008_ = id_fsm_q ? 1'h0 : _0026_;
assign rf_wdata_id_o = rf_wdata_sel ? csr_rdata_i : result_ex_i;
assign _0427_ = _0541_ ? imm_a : pc_id_i;
assign _0429_ = _0543_ ? lsu_addr_last_i : multdiv_operand_a_ex_o;
assign alu_operand_a_ex_o = _0413_ ? _0427_ : _0429_;
assign _0431_ = csr_op_o == /* src = "generated/sv2v_out.v:17541.34-17541.50" */ 2'h1;
assign _0432_ = csr_op_o == /* src = "generated/sv2v_out.v:17541.56-17541.72" */ 2'h2;
assign _0433_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17542.11-17542.42" */ 12'h300;
assign _0434_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17542.48-17542.79" */ 12'h304;
assign _0435_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17542.86-17542.117" */ 12'h747;
assign _0436_ = instr_rdata_i[31:25] == /* src = "generated/sv2v_out.v:17542.124-17542.153" */ 7'h1d;
assign _0437_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17546.11-17546.42" */ 12'h7b0;
assign _0438_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17546.48-17546.79" */ 12'h7b1;
assign _0439_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17546.86-17546.117" */ 12'h7b2;
assign _0440_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17546.124-17546.155" */ 12'h7b3;
assign _0441_ = rf_waddr_wb_i == /* src = "generated/sv2v_out.v:17773.31-17773.60" */ rf_raddr_a_o;
assign _0442_ = rf_waddr_wb_i == /* src = "generated/sv2v_out.v:17774.31-17774.60" */ rf_raddr_b_o;
assign _0443_ = csr_op_en_o && /* src = "generated/sv2v_out.v:17541.7-17541.74" */ _0445_;
assign _0444_ = csr_op_en_o && /* src = "generated/sv2v_out.v:17545.12-17545.55" */ _0453_;
assign _0445_ = _0431_ || /* src = "generated/sv2v_out.v:17541.33-17541.73" */ _0432_;
assign _0446_ = _0433_ || /* src = "generated/sv2v_out.v:17542.10-17542.80" */ _0434_;
assign _0447_ = _0446_ || /* src = "generated/sv2v_out.v:17542.9-17542.118" */ _0435_;
assign _0448_ = _0447_ || /* src = "generated/sv2v_out.v:17542.8-17542.154" */ _0436_;
assign _0449_ = _0437_ || /* src = "generated/sv2v_out.v:17546.10-17546.80" */ _0438_;
assign _0450_ = _0449_ || /* src = "generated/sv2v_out.v:17546.9-17546.118" */ _0439_;
assign _0451_ = _0450_ || /* src = "generated/sv2v_out.v:17546.8-17546.156" */ _0440_;
assign _0452_ = data_ind_timing_i || /* src = "generated/sv2v_out.v:17720.20-17720.80" */ branch_decision_i;
assign _0453_ = | /* src = "generated/sv2v_out.v:17545.38-17545.54" */ csr_op_o;
assign _0454_ = priv_mode_i != /* src = "generated/sv2v_out.v:17550.31-17550.51" */ 2'h3;
assign _0455_ = ~ /* src = "generated/sv2v_out.v:17360.60-17360.75" */ illegal_insn_o;
assign _0456_ = ~ /* src = "generated/sv2v_out.v:17549.45-17549.58" */ debug_mode_o;
assign _0457_ = ~ /* src = "generated/sv2v_out.v:17657.95-17657.115" */ instr_valid_clear_o;
assign _0458_ = ~ /* src = "generated/sv2v_out.v:17755.23-17755.32" */ stall_id;
assign _0459_ = ~ /* src = "generated/sv2v_out.v:17755.35-17755.44" */ flush_id;
assign _0460_ = ~ /* src = "generated/sv2v_out.v:17767.90-17767.107" */ lsu_resp_valid_i;
assign _0461_ = ~ /* src = "generated/sv2v_out.v:17769.78-17769.93" */ controller_run;
assign _0463_ = ~ /* src = "generated/sv2v_out.v:17784.32-17784.43" */ ready_wb_i;
assign _0462_ = ~ /* src = "generated/sv2v_out.v:17785.48-17785.59" */ \gen_stall_mem.instr_kill ;
assign _0464_ = ~ /* src = "generated/sv2v_out.v:17820.36-17820.46" */ ebrk_insn;
assign _0465_ = ~ /* src = "generated/sv2v_out.v:17820.49-17820.64" */ ecall_insn_dec;
assign _0466_ = mret_insn_dec | /* src = "generated/sv2v_out.v:17550.56-17550.105" */ _0053_;
assign _0468_ = illegal_insn_dec | /* src = "generated/sv2v_out.v:17551.45-17551.82" */ illegal_csr_insn_i;
assign _0470_ = _0468_ | /* src = "generated/sv2v_out.v:17551.44-17551.103" */ illegal_dret_insn;
assign _0472_ = _0470_ | /* src = "generated/sv2v_out.v:17551.43-17551.125" */ illegal_umode_insn;
assign mem_resp_intg_err = lsu_load_resp_intg_err_i | /* src = "generated/sv2v_out.v:17552.29-17552.81" */ lsu_store_resp_intg_err_i;
assign multdiv_en_dec = mult_en_dec | /* src = "generated/sv2v_out.v:17624.26-17624.50" */ div_en_dec;
assign _0474_ = branch_set_raw | /* src = "generated/sv2v_out.v:17657.36-17657.65" */ jump_set_raw;
assign _0476_ = _0474_ | /* src = "generated/sv2v_out.v:17657.35-17657.91" */ branch_jump_set_done_q;
assign branch_taken = _0131_ | /* src = "generated/sv2v_out.v:17673.26-17673.61" */ \g_sec_branch_taken.branch_taken_q ;
assign _0478_ = branch_decision_i | /* src = "generated/sv2v_out.v:17722.27-17722.64" */ data_ind_timing_i;
assign _0480_ = stall_ld_hz | /* src = "generated/sv2v_out.v:17754.24-17754.47" */ stall_mem;
assign _0482_ = _0480_ | /* src = "generated/sv2v_out.v:17754.23-17754.64" */ stall_multdiv;
assign _0484_ = _0482_ | /* src = "generated/sv2v_out.v:17754.22-17754.78" */ stall_jump;
assign _0486_ = _0484_ | /* src = "generated/sv2v_out.v:17754.21-17754.94" */ stall_branch;
assign stall_id = _0486_ | /* src = "generated/sv2v_out.v:17754.20-17754.107" */ stall_alu;
assign _0488_ = outstanding_load_wb_i | /* src = "generated/sv2v_out.v:17767.40-17767.86" */ outstanding_store_wb_i;
assign _0490_ = instr_fetch_err_i | /* src = "generated/sv2v_out.v:17769.26-17769.58" */ wb_exception;
assign _0492_ = _0490_ | /* src = "generated/sv2v_out.v:17769.25-17769.74" */ id_exception;
assign \gen_stall_mem.instr_kill  = _0492_ | /* src = "generated/sv2v_out.v:17769.24-17769.93" */ _0461_;
assign _0494_ = \gen_stall_mem.outstanding_memory_access  | /* src = "generated/sv2v_out.v:17772.40-17772.99" */ _0069_;
assign _0496_ = \gen_stall_mem.rf_rd_a_hz  | /* src = "generated/sv2v_out.v:17781.50-17781.73" */ \gen_stall_mem.rf_rd_b_hz ;
assign _0498_ = \gen_stall_mem.outstanding_memory_access  | /* src = "generated/sv2v_out.v:17785.64-17785.103" */ stall_ld_hz;
/* src = "generated/sv2v_out.v:17668.4-17672.42" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$038d6e761af5e8bbfc2ed9b8473abfd849408d7b\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME \g_sec_branch_taken.branch_taken_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_sec_branch_taken.branch_taken_q  <= 1'h0;
else \g_sec_branch_taken.branch_taken_q  <= branch_decision_i;
/* src = "generated/sv2v_out.v:17649.4-17653.43" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$038d6e761af5e8bbfc2ed9b8473abfd849408d7b\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME branch_set_raw */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_set_raw <= 1'h0;
else branch_set_raw <= branch_set_raw_d;
/* src = "generated/sv2v_out.v:17658.2-17662.53" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$038d6e761af5e8bbfc2ed9b8473abfd849408d7b\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME branch_jump_set_done_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_jump_set_done_q <= 1'h0;
else branch_jump_set_done_q <= branch_jump_set_done_d;
assign _0500_ = imm_b_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17448.5-17457.12" */ 3'h5;
assign _0501_ = imm_b_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17448.5-17457.12" */ 3'h4;
assign _0502_ = imm_b_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17448.5-17457.12" */ 3'h3;
assign _0503_ = imm_b_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17448.5-17457.12" */ 3'h2;
assign _0504_ = imm_b_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17448.5-17457.12" */ 3'h1;
assign _0505_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17448.5-17457.12" */ imm_b_mux_sel;
assign _0046_ = _0061_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17742.10-17742.38|generated/sv2v_out.v:17742.6-17748.9" */ 1'h0 : 1'h1;
assign _0039_ = _0061_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17742.10-17742.38|generated/sv2v_out.v:17742.6-17748.9" */ 1'h0 : jump_in_dec;
assign _0037_ = _0061_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17742.10-17742.38|generated/sv2v_out.v:17742.6-17748.9" */ 1'h0 : branch_in_dec;
assign _0044_ = _0061_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17742.10-17742.38|generated/sv2v_out.v:17742.6-17748.9" */ 1'h0 : multdiv_en_dec;
assign _0042_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17740.10-17740.24|generated/sv2v_out.v:17740.6-17741.42" */ _0059_ : rf_we_dec;
assign _0035_ = ex_valid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17714.12-17714.23|generated/sv2v_out.v:17714.8-17718.11" */ rf_we_dec : 1'h0;
assign _0041_ = ex_valid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17714.12-17714.23|generated/sv2v_out.v:17714.8-17718.11" */ 1'h0 : 1'h1;
assign _0034_ = lsu_req_done_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17711.17-17711.32|generated/sv2v_out.v:17711.13-17712.25" */ 1'h0 : 1'h1;
assign _0507_ = jump_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h1 : _0506_;
assign _0508_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ _0546_ : _0507_;
assign _0509_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ _0041_ : _0508_;
assign _0023_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ _0034_ : _0509_;
assign _0506_ = alu_multicycle_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h1 : 1'h0;
assign _0510_ = jump_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0506_;
assign _0511_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0510_;
assign _0512_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0511_;
assign _0029_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0512_;
assign _0513_ = alu_multicycle_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : rf_we_dec;
assign _0515_ = jump_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ rf_we_dec : _0513_;
assign _0517_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ rf_we_dec : _0515_;
assign _0519_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ _0035_ : _0517_;
assign _0027_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ rf_we_dec : _0519_;
assign _0521_ = jump_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h1 : 1'h0;
assign _0522_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0521_;
assign _0523_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0522_;
assign _0030_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0523_;
assign _0524_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ _0478_ : 1'h0;
assign _0526_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0524_;
assign _0528_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ _0041_ : 1'h0;
assign _0031_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0528_;
assign _0529_ = jump_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ jump_set_dec : 1'h0;
assign _0531_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0529_;
assign _0533_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0531_;
assign _0024_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0533_;
assign _0535_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ _0032_ : 1'h0;
assign _0537_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0535_;
assign _0018_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0537_;
assign _0020_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0526_;
assign _0539_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h1 : 1'h0;
assign _0540_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0539_;
assign _0026_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17707.6-17738.13" */ 1'h0 : _0540_;
assign stall_alu = instr_executing_spec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17704.7-17704.27|generated/sv2v_out.v:17704.3-17751.11" */ _0011_ : 1'h0;
assign rf_we_raw = instr_executing_spec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17704.7-17704.27|generated/sv2v_out.v:17704.3-17751.11" */ _0009_ : rf_we_dec;
assign stall_jump = instr_executing_spec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17704.7-17704.27|generated/sv2v_out.v:17704.3-17751.11" */ _0014_ : 1'h0;
assign stall_branch = instr_executing_spec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17704.7-17704.27|generated/sv2v_out.v:17704.3-17751.11" */ _0012_ : 1'h0;
assign stall_multdiv = instr_executing_spec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17704.7-17704.27|generated/sv2v_out.v:17704.3-17751.11" */ _0016_ : 1'h0;
assign jump_set_raw = instr_executing_spec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17704.7-17704.27|generated/sv2v_out.v:17704.3-17751.11" */ _0006_ : 1'h0;
assign branch_not_set = instr_executing_spec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17704.7-17704.27|generated/sv2v_out.v:17704.3-17751.11" */ _0000_ : 1'h0;
assign branch_set_raw_d = instr_executing_spec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17704.7-17704.27|generated/sv2v_out.v:17704.3-17751.11" */ _0002_ : 1'h0;
assign perf_branch_o = instr_executing_spec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17704.7-17704.27|generated/sv2v_out.v:17704.3-17751.11" */ _0008_ : 1'h0;
assign _0033_ = _0451_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17546.8-17546.156|generated/sv2v_out.v:17546.4-17547.27" */ 1'h1 : 1'h0;
assign _0022_ = _0444_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17545.12-17545.55|generated/sv2v_out.v:17545.8-17547.27" */ _0033_ : 1'h0;
assign _0004_ = _0448_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17542.8-17542.154|generated/sv2v_out.v:17542.4-17543.27" */ 1'h1 : 1'h0;
assign csr_pipe_flush = _0443_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17541.7-17541.74|generated/sv2v_out.v:17541.3-17547.27" */ _0004_ : _0022_;
assign _0541_ = alu_op_a_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17399.3-17405.10" */ 2'h3;
assign _0542_ = alu_op_a_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17399.3-17405.10" */ 2'h2;
assign _0543_ = alu_op_a_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17399.3-17405.10" */ 2'h1;
assign _0544_ = | /* src = "generated/sv2v_out.v:17773.64-17773.77" */ rf_raddr_a_o;
assign _0545_ = | /* src = "generated/sv2v_out.v:17774.64-17774.77" */ rf_raddr_b_o;
assign alu_op_a_mux_sel = lsu_addr_incr_req_i ? /* src = "generated/sv2v_out.v:17394.29-17394.78" */ 2'h1 : alu_op_a_mux_sel_dec;
assign alu_op_b_mux_sel = lsu_addr_incr_req_i ? /* src = "generated/sv2v_out.v:17395.29-17395.78" */ 1'h1 : alu_op_b_mux_sel_dec;
assign imm_b_mux_sel = lsu_addr_incr_req_i ? /* src = "generated/sv2v_out.v:17396.26-17396.72" */ 3'h6 : imm_b_mux_sel_dec;
assign imm_a = imm_a_mux_sel ? /* src = "generated/sv2v_out.v:17397.18-17397.70" */ 32'd0 : zimm_rs1_type;
assign alu_operand_b_ex_o = alu_op_b_mux_sel ? /* src = "generated/sv2v_out.v:17461.26-17461.75" */ imm_b : lsu_wdata_o;
assign lsu_req_o = instr_executing ? /* src = "generated/sv2v_out.v:17625.20-17625.75" */ _0055_ : 1'h0;
assign mult_en_ex_o = instr_executing ? /* src = "generated/sv2v_out.v:17626.23-17626.59" */ mult_en_dec : 1'h0;
assign div_en_ex_o = instr_executing ? /* src = "generated/sv2v_out.v:17627.22-17627.57" */ div_en_dec : 1'h0;
assign _0145_ = instr_is_compressed_i ? /* src = "generated/sv2v_out.v:17679.41-17679.78" */ 32'd2 : 32'd4;
assign _0546_ = _0452_ ? /* src = "generated/sv2v_out.v:17720.20-17720.94" */ 1'h1 : 1'h0;
assign multicycle_done = lsu_req_dec ? /* src = "generated/sv2v_out.v:17766.30-17766.67" */ _0132_ : ex_valid_i;
assign multdiv_operand_a_ex_o = _0071_ ? /* src = "generated/sv2v_out.v:17779.29-17779.96" */ rf_wdata_fwd_wb_i : rf_rdata_a_i;
assign lsu_wdata_o = _0072_ ? /* src = "generated/sv2v_out.v:17780.29-17780.96" */ rf_wdata_fwd_wb_i : rf_rdata_b_i;
assign _0547_ = lsu_we_o ? /* src = "generated/sv2v_out.v:17782.53-17782.73" */ 2'h1 : 2'h0;
assign instr_type_wb_o = lsu_req_dec ? /* src = "generated/sv2v_out.v:17782.30-17782.74" */ _0547_ : 2'h2;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:17557.4-17623.3" */
\$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  controller_i (
.branch_not_set_i(branch_not_set),
.branch_not_set_i_t0(branch_not_set_t0),
.branch_set_i(branch_set),
.branch_set_i_t0(branch_set_t0),
.clk_i(clk_i),
.controller_run_o(controller_run),
.controller_run_o_t0(controller_run_t0),
.csr_mstatus_mie_i(csr_mstatus_mie_i),
.csr_mstatus_mie_i_t0(csr_mstatus_mie_i_t0),
.csr_mtval_o(csr_mtval_o),
.csr_mtval_o_t0(csr_mtval_o_t0),
.csr_pipe_flush_i(csr_pipe_flush),
.csr_pipe_flush_i_t0(1'h0),
.csr_restore_dret_id_o(csr_restore_dret_id_o),
.csr_restore_dret_id_o_t0(csr_restore_dret_id_o_t0),
.csr_restore_mret_id_o(csr_restore_mret_id_o),
.csr_restore_mret_id_o_t0(csr_restore_mret_id_o_t0),
.csr_save_cause_o(csr_save_cause_o),
.csr_save_cause_o_t0(csr_save_cause_o_t0),
.csr_save_id_o(csr_save_id_o),
.csr_save_id_o_t0(csr_save_id_o_t0),
.csr_save_if_o(csr_save_if_o),
.csr_save_if_o_t0(csr_save_if_o_t0),
.csr_save_wb_o(csr_save_wb_o),
.csr_save_wb_o_t0(csr_save_wb_o_t0),
.ctrl_busy_o(ctrl_busy_o),
.ctrl_busy_o_t0(ctrl_busy_o_t0),
.debug_cause_o(debug_cause_o),
.debug_cause_o_t0(debug_cause_o_t0),
.debug_csr_save_o(debug_csr_save_o),
.debug_csr_save_o_t0(debug_csr_save_o_t0),
.debug_ebreakm_i(debug_ebreakm_i),
.debug_ebreakm_i_t0(debug_ebreakm_i_t0),
.debug_ebreaku_i(debug_ebreaku_i),
.debug_ebreaku_i_t0(debug_ebreaku_i_t0),
.debug_mode_entering_o(debug_mode_entering_o),
.debug_mode_entering_o_t0(debug_mode_entering_o_t0),
.debug_mode_o(debug_mode_o),
.debug_mode_o_t0(debug_mode_o_t0),
.debug_req_i(debug_req_i),
.debug_req_i_t0(debug_req_i_t0),
.debug_single_step_i(debug_single_step_i),
.debug_single_step_i_t0(debug_single_step_i_t0),
.dret_insn_i(dret_insn_dec),
.dret_insn_i_t0(dret_insn_dec_t0),
.ebrk_insn_i(ebrk_insn),
.ebrk_insn_i_t0(ebrk_insn_t0),
.ecall_insn_i(ecall_insn_dec),
.ecall_insn_i_t0(ecall_insn_dec_t0),
.exc_cause_o(exc_cause_o),
.exc_cause_o_t0(exc_cause_o_t0),
.exc_pc_mux_o(exc_pc_mux_o),
.exc_pc_mux_o_t0(exc_pc_mux_o_t0),
.flush_id_o(flush_id),
.flush_id_o_t0(flush_id_t0),
.id_exception_o(id_exception),
.id_exception_o_t0(id_exception_t0),
.id_in_ready_o(id_in_ready_o),
.id_in_ready_o_t0(id_in_ready_o_t0),
.illegal_insn_i(illegal_insn_o),
.illegal_insn_i_t0(illegal_insn_o_t0),
.instr_bp_taken_i(instr_bp_taken_i),
.instr_bp_taken_i_t0(instr_bp_taken_i_t0),
.instr_compressed_i(instr_rdata_c_i),
.instr_compressed_i_t0(instr_rdata_c_i_t0),
.instr_exec_i(instr_exec_i),
.instr_exec_i_t0(instr_exec_i_t0),
.instr_fetch_err_i(instr_fetch_err_i),
.instr_fetch_err_i_t0(instr_fetch_err_i_t0),
.instr_fetch_err_plus2_i(instr_fetch_err_plus2_i),
.instr_fetch_err_plus2_i_t0(instr_fetch_err_plus2_i_t0),
.instr_i(instr_rdata_i),
.instr_i_t0(instr_rdata_i_t0),
.instr_is_compressed_i(instr_is_compressed_i),
.instr_is_compressed_i_t0(instr_is_compressed_i_t0),
.instr_req_o(instr_req_o),
.instr_req_o_t0(instr_req_o_t0),
.instr_valid_clear_o(instr_valid_clear_o),
.instr_valid_clear_o_t0(instr_valid_clear_o_t0),
.instr_valid_i(instr_valid_i),
.instr_valid_i_t0(instr_valid_i_t0),
.irq_nm_ext_i(irq_nm_i),
.irq_nm_ext_i_t0(irq_nm_i_t0),
.irq_pending_i(irq_pending_i),
.irq_pending_i_t0(irq_pending_i_t0),
.irqs_i(irqs_i),
.irqs_i_t0(irqs_i_t0),
.jump_set_i(jump_set),
.jump_set_i_t0(jump_set_t0),
.load_err_i(lsu_load_err_i),
.load_err_i_t0(lsu_load_err_i_t0),
.lsu_addr_last_i(lsu_addr_last_i),
.lsu_addr_last_i_t0(lsu_addr_last_i_t0),
.mem_resp_intg_err_i(mem_resp_intg_err),
.mem_resp_intg_err_i_t0(mem_resp_intg_err_t0),
.mret_insn_i(mret_insn_dec),
.mret_insn_i_t0(mret_insn_dec_t0),
.nmi_mode_o(nmi_mode_o),
.nmi_mode_o_t0(nmi_mode_o_t0),
.nt_branch_mispredict_o(nt_branch_mispredict_o),
.nt_branch_mispredict_o_t0(nt_branch_mispredict_o_t0),
.pc_id_i(pc_id_i),
.pc_id_i_t0(pc_id_i_t0),
.pc_mux_o(pc_mux_o),
.pc_mux_o_t0(pc_mux_o_t0),
.pc_set_o(pc_set_o),
.pc_set_o_t0(pc_set_o_t0),
.perf_jump_o(perf_jump_o),
.perf_jump_o_t0(perf_jump_o_t0),
.perf_tbranch_o(perf_tbranch_o),
.perf_tbranch_o_t0(perf_tbranch_o_t0),
.priv_mode_i(priv_mode_i),
.priv_mode_i_t0(priv_mode_i_t0),
.ready_wb_i(ready_wb_i),
.ready_wb_i_t0(ready_wb_i_t0),
.rst_ni(rst_ni),
.stall_id_i(stall_id),
.stall_id_i_t0(stall_id_t0),
.stall_wb_i(stall_wb),
.stall_wb_i_t0(stall_wb_t0),
.store_err_i(lsu_store_err_i),
.store_err_i_t0(lsu_store_err_i_t0),
.trigger_match_i(trigger_match_i),
.trigger_match_i_t0(trigger_match_i_t0),
.wb_exception_o(wb_exception),
.wb_exception_o_t0(wb_exception_t0),
.wfi_insn_i(wfi_insn_dec),
.wfi_insn_i_t0(wfi_insn_dec_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:17487.4-17538.3" */
\$paramod$5ffe4cc9ba21eb548f33468a0c4a93d38de3dae5\ibex_decoder  decoder_i (
.alu_multicycle_o(alu_multicycle_dec),
.alu_multicycle_o_t0(alu_multicycle_dec_t0),
.alu_op_a_mux_sel_o(alu_op_a_mux_sel_dec),
.alu_op_a_mux_sel_o_t0(alu_op_a_mux_sel_dec_t0),
.alu_op_b_mux_sel_o(alu_op_b_mux_sel_dec),
.alu_op_b_mux_sel_o_t0(alu_op_b_mux_sel_dec_t0),
.alu_operator_o(alu_operator_ex_o),
.alu_operator_o_t0(alu_operator_ex_o_t0),
.branch_in_dec_o(branch_in_dec),
.branch_in_dec_o_t0(branch_in_dec_t0),
.branch_taken_i(branch_taken),
.branch_taken_i_t0(branch_taken_t0),
.bt_a_mux_sel_o(bt_a_mux_sel),
.bt_a_mux_sel_o_t0(bt_a_mux_sel_t0),
.bt_b_mux_sel_o(bt_b_mux_sel),
.bt_b_mux_sel_o_t0(bt_b_mux_sel_t0),
.clk_i(clk_i),
.csr_access_o(csr_access_o),
.csr_access_o_t0(csr_access_o_t0),
.csr_op_o(csr_op_o),
.csr_op_o_t0(csr_op_o_t0),
.data_req_o(lsu_req_dec),
.data_req_o_t0(lsu_req_dec_t0),
.data_sign_extension_o(lsu_sign_ext_o),
.data_sign_extension_o_t0(lsu_sign_ext_o_t0),
.data_type_o(lsu_type_o),
.data_type_o_t0(lsu_type_o_t0),
.data_we_o(lsu_we_o),
.data_we_o_t0(lsu_we_o_t0),
.div_en_o(div_en_dec),
.div_en_o_t0(div_en_dec_t0),
.div_sel_o(div_sel_ex_o),
.div_sel_o_t0(div_sel_ex_o_t0),
.dret_insn_o(dret_insn_dec),
.dret_insn_o_t0(dret_insn_dec_t0),
.ebrk_insn_o(ebrk_insn),
.ebrk_insn_o_t0(ebrk_insn_t0),
.ecall_insn_o(ecall_insn_dec),
.ecall_insn_o_t0(ecall_insn_dec_t0),
.icache_inval_o(icache_inval_o),
.icache_inval_o_t0(icache_inval_o_t0),
.illegal_c_insn_i(illegal_c_insn_i),
.illegal_c_insn_i_t0(illegal_c_insn_i_t0),
.illegal_insn_o(illegal_insn_dec),
.illegal_insn_o_t0(illegal_insn_dec_t0),
.imm_a_mux_sel_o(imm_a_mux_sel),
.imm_a_mux_sel_o_t0(imm_a_mux_sel_t0),
.imm_b_mux_sel_o(imm_b_mux_sel_dec),
.imm_b_mux_sel_o_t0(imm_b_mux_sel_dec_t0),
.imm_b_type_o(imm_b_type),
.imm_b_type_o_t0(imm_b_type_t0),
.imm_i_type_o(imm_i_type),
.imm_i_type_o_t0(imm_i_type_t0),
.imm_j_type_o(imm_j_type),
.imm_j_type_o_t0(imm_j_type_t0),
.imm_s_type_o(imm_s_type),
.imm_s_type_o_t0(imm_s_type_t0),
.imm_u_type_o(imm_u_type),
.imm_u_type_o_t0(imm_u_type_t0),
.instr_first_cycle_i(instr_first_cycle_id_o),
.instr_first_cycle_i_t0(instr_first_cycle_id_o_t0),
.instr_rdata_alu_i(instr_rdata_alu_i),
.instr_rdata_alu_i_t0(instr_rdata_alu_i_t0),
.instr_rdata_i(instr_rdata_i),
.instr_rdata_i_t0(instr_rdata_i_t0),
.jump_in_dec_o(jump_in_dec),
.jump_in_dec_o_t0(jump_in_dec_t0),
.jump_set_o(jump_set_dec),
.jump_set_o_t0(jump_set_dec_t0),
.mret_insn_o(mret_insn_dec),
.mret_insn_o_t0(mret_insn_dec_t0),
.mult_en_o(mult_en_dec),
.mult_en_o_t0(mult_en_dec_t0),
.mult_sel_o(mult_sel_ex_o),
.mult_sel_o_t0(mult_sel_ex_o_t0),
.multdiv_operator_o(multdiv_operator_ex_o),
.multdiv_operator_o_t0(multdiv_operator_ex_o_t0),
.multdiv_signed_mode_o(multdiv_signed_mode_ex_o),
.multdiv_signed_mode_o_t0(multdiv_signed_mode_ex_o_t0),
.rf_raddr_a_o(rf_raddr_a_o),
.rf_raddr_a_o_t0(rf_raddr_a_o_t0),
.rf_raddr_b_o(rf_raddr_b_o),
.rf_raddr_b_o_t0(rf_raddr_b_o_t0),
.rf_ren_a_o(rf_ren_a_dec),
.rf_ren_a_o_t0(rf_ren_a_dec_t0),
.rf_ren_b_o(rf_ren_b_dec),
.rf_ren_b_o_t0(rf_ren_b_dec_t0),
.rf_waddr_o(rf_waddr_id_o),
.rf_waddr_o_t0(rf_waddr_id_o_t0),
.rf_wdata_sel_o(rf_wdata_sel),
.rf_wdata_sel_o_t0(rf_wdata_sel_t0),
.rf_we_o(rf_we_dec),
.rf_we_o_t0(rf_we_dec_t0),
.rst_ni(rst_ni),
.wfi_insn_o(wfi_insn_dec),
.wfi_insn_o_t0(wfi_insn_dec_t0),
.zimm_rs1_type_o(zimm_rs1_type),
.zimm_rs1_type_o_t0(zimm_rs1_type_t0)
);
assign bt_a_operand_o = 32'd0;
assign bt_a_operand_o_t0 = 32'd0;
assign bt_b_operand_o = 32'd0;
assign bt_b_operand_o_t0 = 32'd0;
assign instr_type_wb_o_t0 = 2'h0;
assign multdiv_operand_b_ex_o = lsu_wdata_o;
assign multdiv_operand_b_ex_o_t0 = lsu_wdata_o_t0;
assign multdiv_ready_id_o = ready_wb_i;
assign multdiv_ready_id_o_t0 = ready_wb_i_t0;
assign perf_branch_o_t0 = 1'h0;
assign rf_rd_a_wb_match_o_t0 = 1'h0;
assign rf_rd_b_wb_match_o_t0 = 1'h0;
endmodule

module \$paramod$34601000fe8707ce2501f5ed778e152043201712\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _0_;
wire [6:0] _1_;
wire [6:0] _2_;
wire [6:0] _3_;
/* src = "generated/sv2v_out.v:14936.13-14936.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14940.28-14940.37" */
output [6:0] rd_data_o;
reg [6:0] rd_data_o;
/* cellift = 32'd1 */
output [6:0] rd_data_o_t0;
reg [6:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14941.14-14941.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14937.13-14937.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14938.27-14938.36" */
input [6:0] wr_data_i;
wire [6:0] wr_data_i;
/* cellift = 32'd1 */
input [6:0] wr_data_i_t0;
wire [6:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14939.13-14939.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _0_ = ~ wr_en_i;
assign _1_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _2_ = { _0_, _0_, _0_, _0_, _0_, _0_, _0_ } & rd_data_o_t0;
assign _3_ = _1_ | _2_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$34601000fe8707ce2501f5ed778e152043201712\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 7'h00;
else rd_data_o_t0 <= _3_;
/* src = "generated/sv2v_out.v:14943.2-14947.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$34601000fe8707ce2501f5ed778e152043201712\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 7'h00;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$410b37fbfbfa994790f1902c150d2be939cadb3b\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _0_;
wire [2:0] _1_;
wire [2:0] _2_;
wire [2:0] _3_;
/* src = "generated/sv2v_out.v:14936.13-14936.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14940.28-14940.37" */
output [2:0] rd_data_o;
reg [2:0] rd_data_o;
/* cellift = 32'd1 */
output [2:0] rd_data_o_t0;
reg [2:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14941.14-14941.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14937.13-14937.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14938.27-14938.36" */
input [2:0] wr_data_i;
wire [2:0] wr_data_i;
/* cellift = 32'd1 */
input [2:0] wr_data_i_t0;
wire [2:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14939.13-14939.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _0_ = ~ wr_en_i;
assign _1_ = { wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _2_ = { _0_, _0_, _0_ } & rd_data_o_t0;
assign _3_ = _1_ | _2_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$410b37fbfbfa994790f1902c150d2be939cadb3b\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 3'h0;
else rd_data_o_t0 <= _3_;
/* src = "generated/sv2v_out.v:14943.2-14947.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$410b37fbfbfa994790f1902c150d2be939cadb3b\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 3'h4;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_flop (clk_i, rst_ni, d_i, q_o, d_i_t0, q_o_t0);
/* src = "generated/sv2v_out.v:24712.8-24712.13" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:24714.22-24714.25" */
input [3:0] d_i;
wire [3:0] d_i;
/* cellift = 32'd1 */
input [3:0] d_i_t0;
wire [3:0] d_i_t0;
/* src = "generated/sv2v_out.v:24715.28-24715.31" */
output [3:0] q_o;
wire [3:0] q_o;
/* cellift = 32'd1 */
output [3:0] q_o_t0;
wire [3:0] q_o_t0;
/* src = "generated/sv2v_out.v:24713.8-24713.14" */
input rst_ni;
wire rst_ni;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:24733.6-24738.5" */
\$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_generic_flop  \gen_generic.u_impl_generic  (
.clk_i(clk_i),
.d_i(d_i),
.d_i_t0(d_i_t0),
.q_o(q_o),
.q_o_t0(q_o_t0),
.rst_ni(rst_ni)
);
endmodule

module \$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_generic_flop (clk_i, rst_ni, d_i, q_o, d_i_t0, q_o_t0);
/* src = "generated/sv2v_out.v:24972.8-24972.13" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:24974.22-24974.25" */
input [3:0] d_i;
wire [3:0] d_i;
/* cellift = 32'd1 */
input [3:0] d_i_t0;
wire [3:0] d_i_t0;
/* src = "generated/sv2v_out.v:24975.27-24975.30" */
output [3:0] q_o;
reg [3:0] q_o;
/* cellift = 32'd1 */
output [3:0] q_o_t0;
reg [3:0] q_o_t0;
/* src = "generated/sv2v_out.v:24973.8-24973.14" */
input rst_ni;
wire rst_ni;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_generic_flop  */
/* PC_TAINT_INFO STATE_NAME q_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) q_o_t0 <= 4'h0;
else q_o_t0 <= d_i_t0;
/* src = "generated/sv2v_out.v:24976.2-24980.15" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_generic_flop  */
/* PC_TAINT_INFO STATE_NAME q_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) q_o <= 4'ha;
else q_o <= d_i;
endmodule

module \$paramod$4f46e25470a27719ee9ca03cee1a0827eff766f7\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _0_;
wire [31:0] _1_;
wire [31:0] _2_;
wire [31:0] _3_;
/* src = "generated/sv2v_out.v:14936.13-14936.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14940.28-14940.37" */
output [31:0] rd_data_o;
reg [31:0] rd_data_o;
/* cellift = 32'd1 */
output [31:0] rd_data_o_t0;
reg [31:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14941.14-14941.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14937.13-14937.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14938.27-14938.36" */
input [31:0] wr_data_i;
wire [31:0] wr_data_i;
/* cellift = 32'd1 */
input [31:0] wr_data_i_t0;
wire [31:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14939.13-14939.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _0_ = ~ wr_en_i;
assign _1_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _2_ = { _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_ } & rd_data_o_t0;
assign _3_ = _1_ | _2_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$4f46e25470a27719ee9ca03cee1a0827eff766f7\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 32'd0;
else rd_data_o_t0 <= _3_;
/* src = "generated/sv2v_out.v:14943.2-14947.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$4f46e25470a27719ee9ca03cee1a0827eff766f7\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 32'd1;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$501c60d7519704ee720c78ef16ad88cf05835059\ibex_dummy_instr (clk_i, rst_ni, dummy_instr_en_i, dummy_instr_mask_i, dummy_instr_seed_en_i, dummy_instr_seed_i, fetch_valid_i, id_in_ready_i, insert_dummy_instr_o, dummy_instr_data_o, insert_dummy_instr_o_t0, id_in_ready_i_t0, dummy_instr_seed_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_mask_i_t0, dummy_instr_en_i_t0, dummy_instr_data_o_t0, fetch_valid_i_t0);
/* src = "generated/sv2v_out.v:15916.25-15916.57" */
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire [31:0] _06_;
wire [31:0] _07_;
wire _08_;
wire [31:0] _09_;
wire [2:0] _10_;
/* src = "generated/sv2v_out.v:15922.50-15922.84" */
wire _11_;
/* src = "generated/sv2v_out.v:15916.62-15916.96" */
wire _12_;
wire _13_;
wire _14_;
wire _15_;
/* src = "generated/sv2v_out.v:15859.13-15859.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:15875.13-15875.24" */
wire [4:0] dummy_cnt_d;
/* src = "generated/sv2v_out.v:15877.7-15877.19" */
wire dummy_cnt_en;
/* src = "generated/sv2v_out.v:15873.13-15873.27" */
wire [4:0] dummy_cnt_incr;
/* src = "generated/sv2v_out.v:15876.12-15876.23" */
reg [4:0] dummy_cnt_q;
/* src = "generated/sv2v_out.v:15874.13-15874.32" */
wire [4:0] dummy_cnt_threshold;
/* src = "generated/sv2v_out.v:15868.21-15868.39" */
output [31:0] dummy_instr_data_o;
wire [31:0] dummy_instr_data_o;
/* cellift = 32'd1 */
output [31:0] dummy_instr_data_o_t0;
wire [31:0] dummy_instr_data_o_t0;
/* src = "generated/sv2v_out.v:15861.13-15861.29" */
input dummy_instr_en_i;
wire dummy_instr_en_i;
/* cellift = 32'd1 */
input dummy_instr_en_i_t0;
wire dummy_instr_en_i_t0;
/* src = "generated/sv2v_out.v:15862.19-15862.37" */
input [2:0] dummy_instr_mask_i;
wire [2:0] dummy_instr_mask_i;
/* cellift = 32'd1 */
input [2:0] dummy_instr_mask_i_t0;
wire [2:0] dummy_instr_mask_i_t0;
/* src = "generated/sv2v_out.v:15885.14-15885.32" */
wire [31:0] dummy_instr_seed_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15885.14-15885.32" */
wire [31:0] dummy_instr_seed_d_t0;
/* src = "generated/sv2v_out.v:15863.13-15863.34" */
input dummy_instr_seed_en_i;
wire dummy_instr_seed_en_i;
/* cellift = 32'd1 */
input dummy_instr_seed_en_i_t0;
wire dummy_instr_seed_en_i_t0;
/* src = "generated/sv2v_out.v:15864.20-15864.38" */
input [31:0] dummy_instr_seed_i;
wire [31:0] dummy_instr_seed_i;
/* cellift = 32'd1 */
input [31:0] dummy_instr_seed_i_t0;
wire [31:0] dummy_instr_seed_i_t0;
/* src = "generated/sv2v_out.v:15884.13-15884.31" */
reg [31:0] dummy_instr_seed_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15884.13-15884.31" */
reg [31:0] dummy_instr_seed_q_t0;
/* src = "generated/sv2v_out.v:15882.12-15882.24" */
wire [2:0] dummy_opcode;
/* src = "generated/sv2v_out.v:15881.12-15881.21" */
wire [6:0] dummy_set;
/* src = "generated/sv2v_out.v:15865.13-15865.26" */
input fetch_valid_i;
wire fetch_valid_i;
/* cellift = 32'd1 */
input fetch_valid_i_t0;
wire fetch_valid_i_t0;
/* src = "generated/sv2v_out.v:15866.13-15866.26" */
input id_in_ready_i;
wire id_in_ready_i;
/* cellift = 32'd1 */
input id_in_ready_i_t0;
wire id_in_ready_i_t0;
/* src = "generated/sv2v_out.v:15867.14-15867.34" */
output insert_dummy_instr_o;
wire insert_dummy_instr_o;
/* cellift = 32'd1 */
output insert_dummy_instr_o_t0;
wire insert_dummy_instr_o_t0;
/* src = "generated/sv2v_out.v:15872.14-15872.23" */
wire [16:0] lfsr_data;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15872.14-15872.23" */
/* unused_bits = "0 1 2 3 4 15 16" */
wire [16:0] lfsr_data_t0;
/* src = "generated/sv2v_out.v:15878.7-15878.14" */
wire lfsr_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15878.7-15878.14" */
wire lfsr_en_t0;
/* src = "generated/sv2v_out.v:15860.13-15860.19" */
input rst_ni;
wire rst_ni;
assign dummy_cnt_incr = dummy_cnt_q + /* src = "generated/sv2v_out.v:15914.26-15914.58" */ 5'h01;
assign lfsr_en = insert_dummy_instr_o & /* src = "generated/sv2v_out.v:15886.19-15886.53" */ id_in_ready_i;
assign dummy_cnt_threshold = lfsr_data[4:0] & /* src = "generated/sv2v_out.v:15913.31-15913.93" */ { dummy_instr_mask_i, 2'h3 };
assign _00_ = dummy_instr_en_i & /* src = "generated/sv2v_out.v:15916.25-15916.57" */ id_in_ready_i;
assign dummy_cnt_en = _00_ & /* src = "generated/sv2v_out.v:15916.24-15916.97" */ _12_;
assign insert_dummy_instr_o = dummy_instr_en_i & /* src = "generated/sv2v_out.v:15922.30-15922.85" */ _11_;
assign _01_ = ~ dummy_instr_seed_en_i;
assign _06_ = { dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i } & dummy_instr_seed_d_t0;
assign _07_ = { _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_, _01_ } & dummy_instr_seed_q_t0;
assign _09_ = _06_ | _07_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$501c60d7519704ee720c78ef16ad88cf05835059\ibex_dummy_instr  */
/* PC_TAINT_INFO STATE_NAME dummy_instr_seed_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_instr_seed_q_t0 <= 32'd0;
else dummy_instr_seed_q_t0 <= _09_;
assign _03_ = insert_dummy_instr_o_t0 & id_in_ready_i;
assign insert_dummy_instr_o_t0 = dummy_instr_en_i_t0 & _11_;
assign _04_ = id_in_ready_i_t0 & insert_dummy_instr_o;
assign _05_ = insert_dummy_instr_o_t0 & id_in_ready_i_t0;
assign _08_ = _03_ | _04_;
assign lfsr_en_t0 = _08_ | _05_;
/* src = "generated/sv2v_out.v:15917.2-15921.31" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$501c60d7519704ee720c78ef16ad88cf05835059\ibex_dummy_instr  */
/* PC_TAINT_INFO STATE_NAME dummy_cnt_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_cnt_q <= 5'h00;
else if (dummy_cnt_en) dummy_cnt_q <= dummy_cnt_d;
/* src = "generated/sv2v_out.v:15888.2-15892.45" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$501c60d7519704ee720c78ef16ad88cf05835059\ibex_dummy_instr  */
/* PC_TAINT_INFO STATE_NAME dummy_instr_seed_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_instr_seed_q <= 32'd0;
else if (dummy_instr_seed_en_i) dummy_instr_seed_q <= dummy_instr_seed_d;
assign _02_ = | { _15_, _13_ };
assign _10_ = _14_ ? 3'h4 : 3'h0;
assign dummy_opcode = _13_ ? 3'h7 : _10_;
assign dummy_set = _02_ ? 7'h00 : 7'h01;
assign dummy_instr_seed_d_t0 = dummy_instr_seed_q_t0 | dummy_instr_seed_i_t0;
assign _11_ = dummy_cnt_q == /* src = "generated/sv2v_out.v:15922.50-15922.84" */ dummy_cnt_threshold;
assign _12_ = fetch_valid_i | /* src = "generated/sv2v_out.v:15916.62-15916.96" */ insert_dummy_instr_o;
assign _13_ = lfsr_data[16:15] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15924.3-15945.10" */ 2'h3;
assign _14_ = lfsr_data[16:15] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15924.3-15945.10" */ 2'h2;
assign _15_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15924.3-15945.10" */ lfsr_data[16:15];
assign dummy_cnt_d = insert_dummy_instr_o ? /* src = "generated/sv2v_out.v:15915.24-15915.73" */ 5'h00 : dummy_cnt_incr;
assign dummy_instr_seed_d = dummy_instr_seed_q ^ /* src = "generated/sv2v_out.v:15887.30-15887.69" */ dummy_instr_seed_i;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:15899.4-15907.3" */
\$paramod$5fd3ce2f8a67228d339c5f62898ff83b3c2a14f0\prim_lfsr  lfsr_i (
.clk_i(clk_i),
.entropy_i(8'h00),
.entropy_i_t0(8'h00),
.lfsr_en_i(lfsr_en),
.lfsr_en_i_t0(lfsr_en_t0),
.rst_ni(rst_ni),
.seed_en_i(dummy_instr_seed_en_i),
.seed_en_i_t0(dummy_instr_seed_en_i_t0),
.seed_i(dummy_instr_seed_d),
.seed_i_t0(dummy_instr_seed_d_t0),
.state_o(lfsr_data),
.state_o_t0(lfsr_data_t0)
);
assign dummy_instr_data_o = { dummy_set, lfsr_data[14:5], dummy_opcode, 12'h033 };
assign dummy_instr_data_o_t0 = { 7'h00, lfsr_data_t0[14:5], 15'h0000 };
endmodule

module \$paramod$5714e31d82f2b8816750797f158ebea69a089104\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _0_;
wire [5:0] _1_;
wire [5:0] _2_;
wire [5:0] _3_;
/* src = "generated/sv2v_out.v:14936.13-14936.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14940.28-14940.37" */
output [5:0] rd_data_o;
reg [5:0] rd_data_o;
/* cellift = 32'd1 */
output [5:0] rd_data_o_t0;
reg [5:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14941.14-14941.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14937.13-14937.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14938.27-14938.36" */
input [5:0] wr_data_i;
wire [5:0] wr_data_i;
/* cellift = 32'd1 */
input [5:0] wr_data_i_t0;
wire [5:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14939.13-14939.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _0_ = ~ wr_en_i;
assign _1_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _2_ = { _0_, _0_, _0_, _0_, _0_, _0_ } & rd_data_o_t0;
assign _3_ = _1_ | _2_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$5714e31d82f2b8816750797f158ebea69a089104\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 6'h00;
else rd_data_o_t0 <= _3_;
/* src = "generated/sv2v_out.v:14943.2-14947.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$5714e31d82f2b8816750797f158ebea69a089104\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 6'h10;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$5fd3ce2f8a67228d339c5f62898ff83b3c2a14f0\prim_lfsr (clk_i, rst_ni, seed_en_i, seed_i, lfsr_en_i, entropy_i, state_o, state_o_t0, seed_i_t0, seed_en_i_t0, lfsr_en_i_t0, entropy_i_t0);
wire _00_;
wire [31:0] _01_;
wire [31:0] _02_;
wire _03_;
wire [31:0] _04_;
wire [31:0] _05_;
wire [31:0] _06_;
wire [31:0] _07_;
wire [31:0] _08_;
/* src = "generated/sv2v_out.v:25540.41-25540.60" */
wire _09_;
/* src = "generated/sv2v_out.v:25522.22-25522.29" */
wire _10_;
/* src = "generated/sv2v_out.v:25540.83-25540.119" */
wire [31:0] _11_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25540.83-25540.119" */
wire [31:0] _12_;
/* src = "generated/sv2v_out.v:25540.41-25540.120" */
wire [31:0] _13_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25540.41-25540.120" */
wire [31:0] _14_;
/* src = "generated/sv2v_out.v:25521.30-25521.90" */
wire [31:0] _15_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25521.30-25521.90" */
wire [31:0] _16_;
/* src = "generated/sv2v_out.v:25488.8-25488.13" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:25493.26-25493.35" */
input [7:0] entropy_i;
wire [7:0] entropy_i;
/* cellift = 32'd1 */
input [7:0] entropy_i_t0;
wire [7:0] entropy_i_t0;
/* src = "generated/sv2v_out.v:25500.22-25500.28" */
wire [31:0] lfsr_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25500.22-25500.28" */
wire [31:0] lfsr_d_t0;
/* src = "generated/sv2v_out.v:25492.8-25492.17" */
input lfsr_en_i;
wire lfsr_en_i;
/* cellift = 32'd1 */
input lfsr_en_i_t0;
wire lfsr_en_i_t0;
/* src = "generated/sv2v_out.v:25501.21-25501.27" */
reg [31:0] lfsr_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25501.21-25501.27" */
reg [31:0] lfsr_q_t0;
/* src = "generated/sv2v_out.v:25499.7-25499.13" */
wire lockup;
/* src = "generated/sv2v_out.v:25502.22-25502.37" */
wire [31:0] next_lfsr_state;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25502.22-25502.37" */
wire [31:0] next_lfsr_state_t0;
/* src = "generated/sv2v_out.v:25489.8-25489.14" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:25490.8-25490.17" */
input seed_en_i;
wire seed_en_i;
/* cellift = 32'd1 */
input seed_en_i_t0;
wire seed_en_i_t0;
/* src = "generated/sv2v_out.v:25491.23-25491.29" */
input [31:0] seed_i;
wire [31:0] seed_i;
/* cellift = 32'd1 */
input [31:0] seed_i_t0;
wire [31:0] seed_i_t0;
/* src = "generated/sv2v_out.v:25494.33-25494.40" */
output [16:0] state_o;
wire [16:0] state_o;
/* cellift = 32'd1 */
output [16:0] state_o_t0;
wire [16:0] state_o_t0;
assign _00_ = ~ _03_;
assign _04_ = { _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_ } & lfsr_d_t0;
assign _05_ = { _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_ } & lfsr_q_t0;
assign _08_ = _04_ | _05_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$5fd3ce2f8a67228d339c5f62898ff83b3c2a14f0\prim_lfsr  */
/* PC_TAINT_INFO STATE_NAME lfsr_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) lfsr_q_t0 <= 32'd0;
else lfsr_q_t0 <= _08_;
/* src = "generated/sv2v_out.v:25619.2-25624.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$5fd3ce2f8a67228d339c5f62898ff83b3c2a14f0\prim_lfsr  */
/* PC_TAINT_INFO STATE_NAME lfsr_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) lfsr_q <= 32'd2891135988;
else if (_03_) lfsr_q <= lfsr_d;
assign _01_ = ~ { _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_, _09_ };
assign _02_ = ~ { seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i };
assign _14_ = _01_ & _12_;
assign _06_ = _02_ & _14_;
assign _12_ = { lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i } & next_lfsr_state_t0;
assign _07_ = { seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i } & seed_i_t0;
assign lfsr_d_t0 = _06_ | _07_;
assign _03_ = | { lfsr_en_i, seed_en_i, _09_ };
assign _16_ = { 24'h000000, entropy_i_t0 } | { lfsr_q_t0[0], 24'h000000, lfsr_q_t0[0], 1'h0, lfsr_q_t0[0], 1'h0, lfsr_q_t0[0], lfsr_q_t0[0], lfsr_q_t0[0] };
assign next_lfsr_state_t0 = _16_ | { 1'h0, lfsr_q_t0[31:1] };
assign _09_ = lfsr_en_i && /* src = "generated/sv2v_out.v:25540.41-25540.60" */ lockup;
assign lockup = ~ /* src = "generated/sv2v_out.v:25522.20-25522.30" */ _10_;
assign _10_ = | /* src = "generated/sv2v_out.v:25522.22-25522.29" */ lfsr_q;
assign _11_ = lfsr_en_i ? /* src = "generated/sv2v_out.v:25540.83-25540.119" */ next_lfsr_state : 32'hxxxxxxxx;
assign _13_ = _09_ ? /* src = "generated/sv2v_out.v:25540.41-25540.120" */ 32'd2891135988 : _11_;
assign lfsr_d = seed_en_i ? /* src = "generated/sv2v_out.v:25540.19-25540.121" */ seed_i : _13_;
assign _15_ = { 24'h000000, entropy_i } ^ /* src = "generated/sv2v_out.v:25521.30-25521.90" */ { lfsr_q[0], 24'h000000, lfsr_q[0], 1'h0, lfsr_q[0], 1'h0, lfsr_q[0], lfsr_q[0], lfsr_q[0] };
assign next_lfsr_state = _15_ ^ /* src = "generated/sv2v_out.v:25521.29-25521.107" */ { 1'h0, lfsr_q[31:1] };
assign state_o = { lfsr_q[21], lfsr_q[16], lfsr_q[5], lfsr_q[9], lfsr_q[12], lfsr_q[0], lfsr_q[19], lfsr_q[29], lfsr_q[4], lfsr_q[7], lfsr_q[1], lfsr_q[28], lfsr_q[10], lfsr_q[17], lfsr_q[22], lfsr_q[23], lfsr_q[13] };
assign state_o_t0 = { lfsr_q_t0[21], lfsr_q_t0[16], lfsr_q_t0[5], lfsr_q_t0[9], lfsr_q_t0[12], lfsr_q_t0[0], lfsr_q_t0[19], lfsr_q_t0[29], lfsr_q_t0[4], lfsr_q_t0[7], lfsr_q_t0[1], lfsr_q_t0[28], lfsr_q_t0[10], lfsr_q_t0[17], lfsr_q_t0[22], lfsr_q_t0[23], lfsr_q_t0[13] };
endmodule

module \$paramod$5ffe4cc9ba21eb548f33468a0c4a93d38de3dae5\ibex_decoder (clk_i, rst_ni, illegal_insn_o, ebrk_insn_o, mret_insn_o, dret_insn_o, ecall_insn_o, wfi_insn_o, jump_set_o, branch_taken_i, icache_inval_o, instr_first_cycle_i, instr_rdata_i, instr_rdata_alu_i, illegal_c_insn_i, imm_a_mux_sel_o, imm_b_mux_sel_o, bt_a_mux_sel_o, bt_b_mux_sel_o, imm_i_type_o, imm_s_type_o
, imm_b_type_o, imm_u_type_o, imm_j_type_o, zimm_rs1_type_o, rf_wdata_sel_o, rf_we_o, rf_raddr_a_o, rf_raddr_b_o, rf_waddr_o, rf_ren_a_o, rf_ren_b_o, alu_operator_o, alu_op_a_mux_sel_o, alu_op_b_mux_sel_o, alu_multicycle_o, mult_en_o, div_en_o, mult_sel_o, div_sel_o, multdiv_operator_o, multdiv_signed_mode_o
, csr_access_o, csr_op_o, data_req_o, data_we_o, data_type_o, data_sign_extension_o, jump_in_dec_o, branch_in_dec_o, zimm_rs1_type_o_t0, wfi_insn_o_t0, rf_we_o_t0, rf_wdata_sel_o_t0, rf_waddr_o_t0, rf_ren_b_o_t0, rf_ren_a_o_t0, rf_raddr_b_o_t0, rf_raddr_a_o_t0, multdiv_signed_mode_o_t0, multdiv_operator_o_t0, mult_sel_o_t0, mult_en_o_t0
, mret_insn_o_t0, jump_set_o_t0, jump_in_dec_o_t0, instr_rdata_alu_i_t0, instr_first_cycle_i_t0, imm_u_type_o_t0, imm_s_type_o_t0, imm_j_type_o_t0, imm_i_type_o_t0, imm_b_type_o_t0, imm_b_mux_sel_o_t0, imm_a_mux_sel_o_t0, illegal_insn_o_t0, illegal_c_insn_i_t0, icache_inval_o_t0, ecall_insn_o_t0, ebrk_insn_o_t0, dret_insn_o_t0, div_sel_o_t0, div_en_o_t0, data_we_o_t0
, data_type_o_t0, data_sign_extension_o_t0, data_req_o_t0, csr_op_o_t0, csr_access_o_t0, bt_b_mux_sel_o_t0, bt_a_mux_sel_o_t0, branch_taken_i_t0, branch_in_dec_o_t0, alu_operator_o_t0, alu_op_b_mux_sel_o_t0, alu_op_a_mux_sel_o_t0, alu_multicycle_o_t0, instr_rdata_i_t0);
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [6:0] _000_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [6:0] _001_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [6:0] _002_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _003_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [6:0] _004_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _005_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [6:0] _006_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _007_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _008_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _009_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _010_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _011_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _012_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _013_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _014_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _015_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _016_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _017_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _018_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _019_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _020_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire [1:0] _021_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire [1:0] _022_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire _023_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _024_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _025_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _026_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _027_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _028_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire _029_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [2:0] _030_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _031_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _032_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _033_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire _034_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire [1:0] _035_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire [1:0] _036_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _037_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _038_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _039_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [1:0] _040_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _041_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire [1:0] _042_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire _043_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _044_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _045_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _046_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _047_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [2:0] _048_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _049_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire _050_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire [1:0] _051_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire [1:0] _052_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _053_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _054_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [6:0] _055_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _056_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [2:0] _057_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [6:0] _058_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _059_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [2:0] _060_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [1:0] _061_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire _062_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _063_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [2:0] _064_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [6:0] _065_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [2:0] _066_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [1:0] _067_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _068_;
/* src = "generated/sv2v_out.v:15384.2-15835.5" */
wire [1:0] _069_;
/* src = "generated/sv2v_out.v:15132.2-15383.5" */
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire [1:0] _114_;
wire [6:0] _115_;
wire [6:0] _116_;
wire [6:0] _117_;
wire [6:0] _118_;
wire [6:0] _119_;
wire [6:0] _120_;
wire [6:0] _121_;
wire [6:0] _122_;
wire [6:0] _123_;
wire [6:0] _124_;
wire [6:0] _125_;
wire [6:0] _126_;
wire [6:0] _127_;
wire [6:0] _128_;
wire [6:0] _129_;
wire [6:0] _130_;
wire [6:0] _131_;
wire [6:0] _132_;
wire [6:0] _133_;
wire _134_;
wire _135_;
wire [1:0] _136_;
wire [1:0] _137_;
wire [1:0] _138_;
wire [1:0] _139_;
wire [6:0] _140_;
wire [6:0] _141_;
wire [6:0] _142_;
wire [6:0] _143_;
wire [2:0] _144_;
wire [2:0] _145_;
wire [2:0] _146_;
wire [2:0] _147_;
wire [2:0] _148_;
wire [1:0] _149_;
wire [1:0] _150_;
wire [1:0] _151_;
wire [1:0] _152_;
wire [1:0] _153_;
wire _154_;
wire [1:0] _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
/* src = "generated/sv2v_out.v:15129.9-15129.23" */
wire _170_;
/* src = "generated/sv2v_out.v:15129.29-15129.43" */
wire _171_;
/* src = "generated/sv2v_out.v:15129.50-15129.74" */
wire _172_;
/* src = "generated/sv2v_out.v:15227.34-15227.55" */
wire _173_;
/* src = "generated/sv2v_out.v:15279.9-15279.44" */
wire _174_;
/* src = "generated/sv2v_out.v:15344.9-15344.31" */
wire _175_;
/* src = "generated/sv2v_out.v:15589.16-15589.44" */
wire _176_;
/* src = "generated/sv2v_out.v:15591.16-15591.44" */
wire _177_;
/* src = "generated/sv2v_out.v:15819.9-15819.35" */
wire _178_;
/* src = "generated/sv2v_out.v:15129.7-15129.75" */
wire _179_;
/* src = "generated/sv2v_out.v:15129.8-15129.44" */
wire _180_;
/* src = "generated/sv2v_out.v:15353.10-15353.59" */
wire _181_;
/* src = "generated/sv2v_out.v:15175.9-15175.31" */
wire _182_;
/* src = "generated/sv2v_out.v:15353.11-15353.32" */
wire _183_;
/* src = "generated/sv2v_out.v:15353.38-15353.58" */
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire [9:0] _239_;
wire _240_;
wire _241_;
wire _242_;
wire [1:0] _243_;
wire _244_;
/* unused_bits = "1 2" */
wire [5:0] _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
/* src = "generated/sv2v_out.v:15227.34-15227.69" */
wire _255_;
/* src = "generated/sv2v_out.v:15055.13-15055.29" */
output alu_multicycle_o;
wire alu_multicycle_o;
/* cellift = 32'd1 */
output alu_multicycle_o_t0;
wire alu_multicycle_o_t0;
/* src = "generated/sv2v_out.v:15053.19-15053.37" */
output [1:0] alu_op_a_mux_sel_o;
wire [1:0] alu_op_a_mux_sel_o;
/* cellift = 32'd1 */
output [1:0] alu_op_a_mux_sel_o_t0;
wire [1:0] alu_op_a_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:15054.13-15054.31" */
output alu_op_b_mux_sel_o;
wire alu_op_b_mux_sel_o;
/* cellift = 32'd1 */
output alu_op_b_mux_sel_o_t0;
wire alu_op_b_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:15052.19-15052.33" */
output [6:0] alu_operator_o;
wire [6:0] alu_operator_o;
/* cellift = 32'd1 */
output [6:0] alu_operator_o_t0;
wire [6:0] alu_operator_o_t0;
/* src = "generated/sv2v_out.v:15069.13-15069.28" */
output branch_in_dec_o;
wire branch_in_dec_o;
/* cellift = 32'd1 */
output branch_in_dec_o_t0;
wire branch_in_dec_o_t0;
/* src = "generated/sv2v_out.v:15029.13-15029.27" */
input branch_taken_i;
wire branch_taken_i;
/* cellift = 32'd1 */
input branch_taken_i_t0;
wire branch_taken_i_t0;
/* src = "generated/sv2v_out.v:15037.19-15037.33" */
output [1:0] bt_a_mux_sel_o;
wire [1:0] bt_a_mux_sel_o;
/* cellift = 32'd1 */
output [1:0] bt_a_mux_sel_o_t0;
wire [1:0] bt_a_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:15038.19-15038.33" */
output [2:0] bt_b_mux_sel_o;
wire [2:0] bt_b_mux_sel_o;
/* cellift = 32'd1 */
output [2:0] bt_b_mux_sel_o_t0;
wire [2:0] bt_b_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:15020.13-15020.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:15062.13-15062.25" */
output csr_access_o;
wire csr_access_o;
/* cellift = 32'd1 */
output csr_access_o_t0;
wire csr_access_o_t0;
/* src = "generated/sv2v_out.v:15083.12-15083.18" */
wire [1:0] csr_op;
/* src = "generated/sv2v_out.v:15063.19-15063.27" */
output [1:0] csr_op_o;
wire [1:0] csr_op_o;
/* cellift = 32'd1 */
output [1:0] csr_op_o_t0;
wire [1:0] csr_op_o_t0;
/* src = "generated/sv2v_out.v:15064.13-15064.23" */
output data_req_o;
wire data_req_o;
/* cellift = 32'd1 */
output data_req_o_t0;
wire data_req_o_t0;
/* src = "generated/sv2v_out.v:15067.13-15067.34" */
output data_sign_extension_o;
wire data_sign_extension_o;
/* cellift = 32'd1 */
output data_sign_extension_o_t0;
wire data_sign_extension_o_t0;
/* src = "generated/sv2v_out.v:15066.19-15066.30" */
output [1:0] data_type_o;
wire [1:0] data_type_o;
/* cellift = 32'd1 */
output [1:0] data_type_o_t0;
wire [1:0] data_type_o_t0;
/* src = "generated/sv2v_out.v:15065.13-15065.22" */
output data_we_o;
wire data_we_o;
/* cellift = 32'd1 */
output data_we_o_t0;
wire data_we_o_t0;
/* src = "generated/sv2v_out.v:15057.14-15057.22" */
output div_en_o;
wire div_en_o;
/* cellift = 32'd1 */
output div_en_o_t0;
wire div_en_o_t0;
/* src = "generated/sv2v_out.v:15059.13-15059.22" */
output div_sel_o;
wire div_sel_o;
/* cellift = 32'd1 */
output div_sel_o_t0;
wire div_sel_o_t0;
/* src = "generated/sv2v_out.v:15025.13-15025.24" */
output dret_insn_o;
wire dret_insn_o;
/* cellift = 32'd1 */
output dret_insn_o_t0;
wire dret_insn_o_t0;
/* src = "generated/sv2v_out.v:15023.13-15023.24" */
output ebrk_insn_o;
wire ebrk_insn_o;
/* cellift = 32'd1 */
output ebrk_insn_o_t0;
wire ebrk_insn_o_t0;
/* src = "generated/sv2v_out.v:15026.13-15026.25" */
output ecall_insn_o;
wire ecall_insn_o;
/* cellift = 32'd1 */
output ecall_insn_o_t0;
wire ecall_insn_o_t0;
/* src = "generated/sv2v_out.v:15030.13-15030.27" */
output icache_inval_o;
wire icache_inval_o;
/* cellift = 32'd1 */
output icache_inval_o_t0;
wire icache_inval_o_t0;
/* src = "generated/sv2v_out.v:15034.13-15034.29" */
input illegal_c_insn_i;
wire illegal_c_insn_i;
/* cellift = 32'd1 */
input illegal_c_insn_i_t0;
wire illegal_c_insn_i_t0;
/* src = "generated/sv2v_out.v:15022.14-15022.28" */
output illegal_insn_o;
wire illegal_insn_o;
/* cellift = 32'd1 */
output illegal_insn_o_t0;
wire illegal_insn_o_t0;
/* src = "generated/sv2v_out.v:15035.13-15035.28" */
output imm_a_mux_sel_o;
wire imm_a_mux_sel_o;
/* cellift = 32'd1 */
output imm_a_mux_sel_o_t0;
wire imm_a_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:15036.19-15036.34" */
output [2:0] imm_b_mux_sel_o;
wire [2:0] imm_b_mux_sel_o;
/* cellift = 32'd1 */
output [2:0] imm_b_mux_sel_o_t0;
wire [2:0] imm_b_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:15041.21-15041.33" */
output [31:0] imm_b_type_o;
wire [31:0] imm_b_type_o;
/* cellift = 32'd1 */
output [31:0] imm_b_type_o_t0;
wire [31:0] imm_b_type_o_t0;
/* src = "generated/sv2v_out.v:15039.21-15039.33" */
output [31:0] imm_i_type_o;
wire [31:0] imm_i_type_o;
/* cellift = 32'd1 */
output [31:0] imm_i_type_o_t0;
wire [31:0] imm_i_type_o_t0;
/* src = "generated/sv2v_out.v:15043.21-15043.33" */
output [31:0] imm_j_type_o;
wire [31:0] imm_j_type_o;
/* cellift = 32'd1 */
output [31:0] imm_j_type_o_t0;
wire [31:0] imm_j_type_o_t0;
/* src = "generated/sv2v_out.v:15040.21-15040.33" */
output [31:0] imm_s_type_o;
wire [31:0] imm_s_type_o;
/* cellift = 32'd1 */
output [31:0] imm_s_type_o_t0;
wire [31:0] imm_s_type_o_t0;
/* src = "generated/sv2v_out.v:15042.21-15042.33" */
output [31:0] imm_u_type_o;
wire [31:0] imm_u_type_o;
/* cellift = 32'd1 */
output [31:0] imm_u_type_o_t0;
wire [31:0] imm_u_type_o_t0;
/* src = "generated/sv2v_out.v:15031.13-15031.32" */
input instr_first_cycle_i;
wire instr_first_cycle_i;
/* cellift = 32'd1 */
input instr_first_cycle_i_t0;
wire instr_first_cycle_i_t0;
/* src = "generated/sv2v_out.v:15033.20-15033.37" */
input [31:0] instr_rdata_alu_i;
wire [31:0] instr_rdata_alu_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_alu_i_t0;
wire [31:0] instr_rdata_alu_i_t0;
/* src = "generated/sv2v_out.v:15032.20-15032.33" */
input [31:0] instr_rdata_i;
wire [31:0] instr_rdata_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_i_t0;
wire [31:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:15068.13-15068.26" */
output jump_in_dec_o;
wire jump_in_dec_o;
/* cellift = 32'd1 */
output jump_in_dec_o_t0;
wire jump_in_dec_o_t0;
/* src = "generated/sv2v_out.v:15028.13-15028.23" */
output jump_set_o;
wire jump_set_o;
/* cellift = 32'd1 */
output jump_set_o_t0;
wire jump_set_o_t0;
/* src = "generated/sv2v_out.v:15024.13-15024.24" */
output mret_insn_o;
wire mret_insn_o;
/* cellift = 32'd1 */
output mret_insn_o_t0;
wire mret_insn_o_t0;
/* src = "generated/sv2v_out.v:15056.14-15056.23" */
output mult_en_o;
wire mult_en_o;
/* cellift = 32'd1 */
output mult_en_o_t0;
wire mult_en_o_t0;
/* src = "generated/sv2v_out.v:15058.13-15058.23" */
output mult_sel_o;
wire mult_sel_o;
/* cellift = 32'd1 */
output mult_sel_o_t0;
wire mult_sel_o_t0;
/* src = "generated/sv2v_out.v:15060.19-15060.37" */
output [1:0] multdiv_operator_o;
wire [1:0] multdiv_operator_o;
/* cellift = 32'd1 */
output [1:0] multdiv_operator_o_t0;
wire [1:0] multdiv_operator_o_t0;
/* src = "generated/sv2v_out.v:15061.19-15061.40" */
output [1:0] multdiv_signed_mode_o;
wire [1:0] multdiv_signed_mode_o;
/* cellift = 32'd1 */
output [1:0] multdiv_signed_mode_o_t0;
wire [1:0] multdiv_signed_mode_o_t0;
/* src = "generated/sv2v_out.v:15047.20-15047.32" */
output [4:0] rf_raddr_a_o;
wire [4:0] rf_raddr_a_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_a_o_t0;
wire [4:0] rf_raddr_a_o_t0;
/* src = "generated/sv2v_out.v:15048.20-15048.32" */
output [4:0] rf_raddr_b_o;
wire [4:0] rf_raddr_b_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_b_o_t0;
wire [4:0] rf_raddr_b_o_t0;
/* src = "generated/sv2v_out.v:15050.13-15050.23" */
output rf_ren_a_o;
wire rf_ren_a_o;
/* cellift = 32'd1 */
output rf_ren_a_o_t0;
wire rf_ren_a_o_t0;
/* src = "generated/sv2v_out.v:15051.13-15051.23" */
output rf_ren_b_o;
wire rf_ren_b_o;
/* cellift = 32'd1 */
output rf_ren_b_o_t0;
wire rf_ren_b_o_t0;
/* src = "generated/sv2v_out.v:15049.20-15049.30" */
output [4:0] rf_waddr_o;
wire [4:0] rf_waddr_o;
/* cellift = 32'd1 */
output [4:0] rf_waddr_o_t0;
wire [4:0] rf_waddr_o_t0;
/* src = "generated/sv2v_out.v:15045.13-15045.27" */
output rf_wdata_sel_o;
wire rf_wdata_sel_o;
/* cellift = 32'd1 */
output rf_wdata_sel_o_t0;
wire rf_wdata_sel_o_t0;
/* src = "generated/sv2v_out.v:15046.14-15046.21" */
output rf_we_o;
wire rf_we_o;
/* cellift = 32'd1 */
output rf_we_o_t0;
wire rf_we_o_t0;
/* src = "generated/sv2v_out.v:15021.13-15021.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:15027.13-15027.23" */
output wfi_insn_o;
wire wfi_insn_o;
/* cellift = 32'd1 */
output wfi_insn_o_t0;
wire wfi_insn_o_t0;
/* src = "generated/sv2v_out.v:15044.21-15044.36" */
output [31:0] zimm_rs1_type_o;
wire [31:0] zimm_rs1_type_o;
/* cellift = 32'd1 */
output [31:0] zimm_rs1_type_o_t0;
wire [31:0] zimm_rs1_type_o_t0;
assign _071_ = ~ instr_rdata_i[14];
assign data_sign_extension_o_t0 = _246_ & instr_rdata_i_t0[14];
assign _083_ = | { _229_, _175_ };
assign _084_ = | { _217_, _216_ };
assign _085_ = | { _250_, _248_, _240_ };
assign _086_ = | { _228_, _227_, _226_, _225_, _224_ };
assign _087_ = | { _254_, _253_, _242_, _240_ };
assign _089_ = | { _251_, _250_, _248_, _246_, _242_, _240_ };
assign _090_ = | { _195_, _194_, _193_, _192_ };
assign _091_ = | { _191_, _190_, _189_, _188_ };
assign _092_ = | { _232_, _231_ };
assign _093_ = | { _234_, _233_ };
assign _094_ = | { _237_, _236_, _235_ };
assign _095_ = | { _204_, _195_, _194_, _193_, _192_, _191_, _190_, _189_, _188_ };
assign _096_ = | { _237_, _234_, _232_ };
assign _097_ = | { _219_, _217_ };
assign _098_ = | { _219_, _218_, _217_, _216_, _215_, _213_ };
assign _100_ = | { _239_, _238_, _237_, _236_, _235_, _234_, _233_, _232_, _231_ };
assign _101_ = | { _215_, _214_ };
assign _088_ = | { _252_, _251_ };
assign _099_ = | { _248_, _246_ };
assign _072_ = | { _186_, _178_ };
assign _073_ = | { _222_, _221_, _220_ };
assign _074_ = | { _247_, _222_ };
assign _075_ = | { _247_, _222_, _221_ };
assign _102_ = _196_ | _095_;
assign _103_ = _201_ | _200_;
assign _104_ = _186_ | _206_;
assign _105_ = _211_ | _210_;
assign _106_ = _186_ | _210_;
assign _107_ = _213_ | _205_;
assign _108_ = _215_ | _214_;
assign _109_ = _221_ | _220_;
assign _110_ = _093_ | _092_;
assign _111_ = _087_ | _223_;
assign _112_ = _230_ | _223_;
assign _113_ = _248_ | _246_;
assign _076_ = | { _102_, _199_, _198_, _197_ };
assign _077_ = | { _209_, _208_, _104_ };
assign _078_ = | { _209_, _208_, _206_ };
assign _079_ = | { _218_, _213_, _207_, _205_, _187_, _185_ };
assign _080_ = | { _207_, _205_, _187_ };
assign _081_ = | { _219_, _217_, _213_, _187_ };
assign _082_ = | { _112_, _254_, _253_, _252_, _242_, _240_ };
assign _114_ = _178_ ? 2'h0 : 2'h3;
assign _061_ = _186_ ? 2'h2 : _114_;
assign _115_ = _095_ ? 7'h00 : 7'h08;
assign _116_ = _198_ ? 7'h0a : 7'h04;
assign _117_ = _197_ ? 7'h09 : _116_;
assign _118_ = _102_ ? _115_ : _117_;
assign _119_ = _200_ ? 7'h03 : 7'h02;
assign _120_ = _203_ ? 7'h01 : 7'h2c;
assign _121_ = _202_ ? 7'h2b : _120_;
assign _122_ = _103_ ? _119_ : _121_;
assign _004_ = _076_ ? _118_ : _122_;
assign _123_ = _206_ ? _000_ : 7'h0a;
assign _124_ = _208_ ? 7'h04 : 7'h03;
assign _125_ = _104_ ? _123_ : _124_;
assign _126_ = _210_ ? 7'h02 : 7'h2c;
assign _127_ = _212_ ? 7'h2b : 7'h00;
assign _128_ = _105_ ? _126_ : _127_;
assign _065_ = _077_ ? _125_ : _128_;
assign _129_ = _209_ ? 7'h1a : 7'h1b;
assign _130_ = _208_ ? 7'h1c : _129_;
assign _131_ = _210_ ? 7'h19 : 7'h1e;
assign _132_ = _178_ ? 7'h1d : 7'h2c;
assign _133_ = _106_ ? _131_ : _132_;
assign _055_ = _078_ ? _130_ : _133_;
assign _134_ = _205_ ? 1'h0 : _062_;
assign _135_ = _214_ ? _038_ : 1'h1;
assign alu_op_b_mux_sel_o = _107_ ? _134_ : _135_;
assign _136_ = _187_ ? _061_ : 2'h0;
assign _137_ = _185_ ? _067_ : _136_;
assign _138_ = _101_ ? _040_ : 2'h3;
assign _139_ = _084_ ? 2'h2 : _138_;
assign alu_op_a_mux_sel_o = _079_ ? _137_ : _139_;
assign _140_ = _205_ ? _002_ : _065_;
assign _141_ = _187_ ? _006_ : _140_;
assign _142_ = _214_ ? _058_ : 7'h2c;
assign _143_ = _098_ ? 7'h00 : _142_;
assign alu_operator_o = _080_ ? _141_ : _143_;
assign _144_ = _097_ ? 3'h3 : _064_;
assign _145_ = _187_ ? _066_ : _144_;
assign _146_ = _214_ ? _057_ : _048_;
assign _147_ = _216_ ? _030_ : 3'h0;
assign _148_ = _108_ ? _146_ : _147_;
assign imm_b_mux_sel_o = _081_ ? _145_ : _148_;
assign _149_ = _220_ ? 2'h3 : 2'h2;
assign _150_ = _222_ ? 2'h1 : 2'h0;
assign _042_ = _109_ ? _149_ : _150_;
assign _151_ = _236_ ? 2'h1 : 2'h0;
assign _052_ = _096_ ? 2'h3 : _151_;
assign _152_ = _092_ ? 2'h3 : 2'h2;
assign _153_ = _094_ ? 2'h1 : 2'h0;
assign _051_ = _110_ ? _152_ : _153_;
assign _154_ = _229_ ? _070_ : 1'h0;
assign _068_ = _241_ ? _003_ : _154_;
assign _155_ = _247_ ? 2'h2 : 2'h0;
assign _022_ = _222_ ? 2'h1 : _155_;
assign _156_ = _074_ ? 1'h0 : 1'h1;
assign _063_ = _221_ ? _056_ : _156_;
assign _157_ = _223_ ? _020_ : 1'h1;
assign _158_ = _088_ ? _038_ : 1'h0;
assign _014_ = _111_ ? _157_ : _158_;
assign _159_ = _088_ ? _032_ : 1'h0;
assign _013_ = _230_ ? _027_ : _159_;
assign _160_ = _088_ ? 1'h1 : 1'h0;
assign _012_ = _230_ ? _031_ : _160_;
assign _161_ = _223_ ? _017_ : _016_;
assign _162_ = _242_ ? _068_ : 1'h0;
assign _163_ = _240_ ? _007_ : _162_;
assign _164_ = _112_ ? _161_ : _163_;
assign _165_ = _246_ ? _063_ : _059_;
assign _166_ = _251_ ? _028_ : 1'h1;
assign _167_ = _250_ ? _047_ : _166_;
assign _168_ = _113_ ? _165_ : _167_;
assign _011_ = _082_ ? _164_ : _168_;
assign _169_ = _089_ ? 1'h1 : 1'h0;
assign rf_ren_a_o = _223_ ? _037_ : _169_;
assign _170_ = csr_op == /* src = "generated/sv2v_out.v:15129.9-15129.23" */ 2'h2;
assign _171_ = csr_op == /* src = "generated/sv2v_out.v:15129.29-15129.43" */ 2'h3;
assign _172_ = ! /* src = "generated/sv2v_out.v:15129.50-15129.74" */ instr_rdata_i[19:15];
assign _174_ = { instr_rdata_i[26], instr_rdata_i[13:12] } == /* src = "generated/sv2v_out.v:15279.9-15279.44" */ 3'h5;
assign _176_ = ! /* src = "generated/sv2v_out.v:15589.16-15589.44" */ instr_rdata_alu_i[31:27];
assign _177_ = instr_rdata_alu_i[31:27] == /* src = "generated/sv2v_out.v:15591.16-15591.44" */ 5'h08;
assign _179_ = _180_ && /* src = "generated/sv2v_out.v:15129.7-15129.75" */ _172_;
assign _180_ = _170_ || /* src = "generated/sv2v_out.v:15129.8-15129.44" */ _171_;
assign _181_ = _183_ || /* src = "generated/sv2v_out.v:15353.10-15353.59" */ _184_;
assign _182_ = | /* src = "generated/sv2v_out.v:15175.9-15175.31" */ instr_rdata_i[14:12];
assign _183_ = | /* src = "generated/sv2v_out.v:15353.11-15353.32" */ instr_rdata_i[19:15];
assign _184_ = | /* src = "generated/sv2v_out.v:15353.38-15353.58" */ instr_rdata_i[11:7];
assign _069_ = instr_rdata_alu_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15827.10-15827.23|generated/sv2v_out.v:15827.6-15830.33" */ 2'h3 : 2'h0;
assign _067_ = _178_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15819.9-15819.35|generated/sv2v_out.v:15819.5-15831.8" */ 2'h0 : _069_;
assign _029_ = _178_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15819.9-15819.35|generated/sv2v_out.v:15819.5-15831.8" */ 1'h1 : 1'h0;
assign _006_ = _072_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15798.5-15817.12" */ 7'h00 : 7'h2c;
assign _066_ = _186_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15798.5-15817.12" */ 3'h5 : 3'h0;
assign _196_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 10'h105;
assign _197_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 10'h005;
assign _198_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 10'h001;
assign _199_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 10'h007;
assign _200_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 10'h006;
assign _201_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 10'h004;
assign _202_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 10'h002;
assign _203_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 10'h100;
assign _204_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] };
assign _043_ = _091_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 1'h1 : 1'h0;
assign _188_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 10'h00f;
assign _189_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 10'h00e;
assign _190_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 10'h00d;
assign _191_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 10'h00c;
assign _050_ = _090_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 1'h1 : 1'h0;
assign _192_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 10'h00b;
assign _193_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 10'h00a;
assign _194_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 10'h009;
assign _195_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15640.6-15795.13" */ 10'h008;
assign _023_ = instr_rdata_alu_i[26] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15600.9-15600.22|generated/sv2v_out.v:15600.5-15795.13" */ 1'h0 : _043_;
assign _034_ = instr_rdata_alu_i[26] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15600.9-15600.22|generated/sv2v_out.v:15600.5-15795.13" */ 1'h0 : _050_;
assign _002_ = instr_rdata_alu_i[26] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15600.9-15600.22|generated/sv2v_out.v:15600.5-15795.13" */ 7'h2c : _004_;
assign _001_ = _177_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15591.16-15591.44|generated/sv2v_out.v:15591.12-15592.30" */ 7'h08 : 7'h2c;
assign _000_ = _176_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15589.16-15589.44|generated/sv2v_out.v:15589.12-15592.30" */ 7'h09 : _001_;
assign _211_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15492.5-15595.12" */ 3'h3;
assign _212_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15492.5-15595.12" */ 3'h2;
assign _062_ = instr_rdata_alu_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15464.9-15464.23|generated/sv2v_out.v:15464.5-15467.8" */ 1'h0 : 1'h1;
assign _064_ = instr_rdata_alu_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15464.9-15464.23|generated/sv2v_out.v:15464.5-15467.8" */ 3'h0 : 3'h1;
assign _038_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15449.9-15449.28|generated/sv2v_out.v:15449.5-15458.8" */ 1'h0 : 1'h1;
assign _058_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15449.9-15449.28|generated/sv2v_out.v:15449.5-15458.8" */ _055_ : 7'h00;
assign _057_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15449.9-15449.28|generated/sv2v_out.v:15449.5-15458.8" */ 3'h0 : _060_;
assign _208_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15435.5-15444.12" */ 3'h7;
assign _209_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15435.5-15444.12" */ 3'h6;
assign _206_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15435.5-15444.12" */ 3'h5;
assign _210_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15435.5-15444.12" */ 3'h4;
assign _186_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15435.5-15444.12" */ 3'h1;
assign _178_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15435.5-15444.12" */ instr_rdata_alu_i[14:12];
assign _048_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15421.9-15421.48|generated/sv2v_out.v:15421.5-15432.8" */ 3'h0 : 3'h5;
assign _040_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15421.9-15421.48|generated/sv2v_out.v:15421.5-15432.8" */ 2'h0 : 2'h2;
assign _030_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15403.9-15403.48|generated/sv2v_out.v:15403.5-15414.8" */ 3'h4 : 3'h5;
assign _207_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15397.3-15834.10" */ 7'h13;
assign _218_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15397.3-15834.10" */ 7'h03;
assign _187_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15397.3-15834.10" */ 7'h0f;
assign _217_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15397.3-15834.10" */ 7'h17;
assign _219_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15397.3-15834.10" */ 7'h37;
assign _213_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15397.3-15834.10" */ 7'h23;
assign _214_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15397.3-15834.10" */ 7'h63;
assign _215_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15397.3-15834.10" */ 7'h67;
assign _216_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15397.3-15834.10" */ 7'h6f;
assign div_sel_o = _205_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15397.3-15834.10" */ _023_ : 1'h0;
assign mult_sel_o = _205_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15397.3-15834.10" */ _034_ : 1'h0;
assign _205_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15397.3-15834.10" */ 7'h33;
assign imm_a_mux_sel_o = _185_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15397.3-15834.10" */ _029_ : 1'h1;
assign _185_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15397.3-15834.10" */ 7'h73;
assign csr_access_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15374.7-15374.19|generated/sv2v_out.v:15374.3-15382.6" */ 1'h0 : rf_wdata_sel_o;
assign branch_in_dec_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15374.7-15374.19|generated/sv2v_out.v:15374.3-15382.6" */ 1'h0 : _008_;
assign jump_set_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15374.7-15374.19|generated/sv2v_out.v:15374.3-15382.6" */ 1'h0 : _013_;
assign jump_in_dec_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15374.7-15374.19|generated/sv2v_out.v:15374.3-15382.6" */ 1'h0 : _012_;
assign data_we_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15374.7-15374.19|generated/sv2v_out.v:15374.3-15382.6" */ 1'h0 : _010_;
assign data_req_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15374.7-15374.19|generated/sv2v_out.v:15374.3-15382.6" */ 1'h0 : _009_;
assign rf_we_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15374.7-15374.19|generated/sv2v_out.v:15374.3-15382.6" */ 1'h0 : _014_;
assign illegal_insn_o = illegal_c_insn_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15372.7-15372.23|generated/sv2v_out.v:15372.3-15373.24" */ 1'h1 : _011_;
assign _041_ = _073_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15362.6-15367.13" */ 1'h0 : 1'h1;
assign _220_ = instr_rdata_i[13:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15362.6-15367.13" */ 2'h3;
assign _053_ = instr_rdata_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15360.10-15360.20|generated/sv2v_out.v:15360.6-15361.25" */ 1'h0 : 1'h1;
assign _019_ = _181_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15353.10-15353.59|generated/sv2v_out.v:15353.6-15354.27" */ 1'h1 : _018_;
assign _046_ = _224_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15345.6-15352.13" */ 1'h1 : 1'h0;
assign _018_ = _086_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15345.6-15352.13" */ 1'h0 : 1'h1;
assign _224_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15345.6-15352.13" */ instr_rdata_i[31:20];
assign _054_ = _225_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15345.6-15352.13" */ 1'h1 : 1'h0;
assign _225_ = instr_rdata_i[31:20] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15345.6-15352.13" */ 12'h105;
assign _044_ = _226_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15345.6-15352.13" */ 1'h1 : 1'h0;
assign _226_ = instr_rdata_i[31:20] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15345.6-15352.13" */ 12'h7b2;
assign _049_ = _227_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15345.6-15352.13" */ 1'h1 : 1'h0;
assign _227_ = instr_rdata_i[31:20] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15345.6-15352.13" */ 12'h302;
assign _045_ = _228_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15345.6-15352.13" */ 1'h1 : 1'h0;
assign _228_ = instr_rdata_i[31:20] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15345.6-15352.13" */ 12'h001;
assign _017_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15344.9-15344.31|generated/sv2v_out.v:15344.5-15369.8" */ _019_ : _041_;
assign _039_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15344.9-15344.31|generated/sv2v_out.v:15344.5-15369.8" */ _054_ : 1'h0;
assign _026_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15344.9-15344.31|generated/sv2v_out.v:15344.5-15369.8" */ _046_ : 1'h0;
assign _024_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15344.9-15344.31|generated/sv2v_out.v:15344.5-15369.8" */ _044_ : 1'h0;
assign _033_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15344.9-15344.31|generated/sv2v_out.v:15344.5-15369.8" */ _049_ : 1'h0;
assign _025_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15344.9-15344.31|generated/sv2v_out.v:15344.5-15369.8" */ _045_ : 1'h0;
assign _037_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15344.9-15344.31|generated/sv2v_out.v:15344.5-15369.8" */ 1'h0 : _053_;
assign _020_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15344.9-15344.31|generated/sv2v_out.v:15344.5-15369.8" */ 1'h0 : 1'h1;
assign _021_ = _175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15344.9-15344.31|generated/sv2v_out.v:15344.5-15369.8" */ 2'h0 : _042_;
assign _016_ = _083_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15331.5-15342.12" */ 1'h0 : 1'h1;
assign _031_ = _229_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15331.5-15342.12" */ 1'h1 : 1'h0;
assign _027_ = _229_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15331.5-15342.12" */ _032_ : 1'h0;
assign _015_ = _100_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 1'h0 : 1'h1;
assign _238_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h008;
assign _239_[0] = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ { instr_rdata_i[31:25], instr_rdata_i[14:12] };
assign _239_[1] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h100;
assign _239_[2] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h002;
assign _239_[3] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h003;
assign _239_[4] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h004;
assign _239_[5] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h006;
assign _239_[6] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h007;
assign _239_[7] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h001;
assign _239_[8] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h005;
assign _239_[9] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h105;
assign _231_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h00f;
assign _232_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h00e;
assign _233_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h00d;
assign _234_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h00c;
assign _235_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h00b;
assign _236_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h00a;
assign _237_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15282.6-15328.13" */ 10'h009;
assign _007_ = _174_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15279.9-15279.44|generated/sv2v_out.v:15279.5-15328.13" */ 1'h1 : _015_;
assign _036_ = _174_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15279.9-15279.44|generated/sv2v_out.v:15279.5-15328.13" */ 2'h0 : _052_;
assign _035_ = _174_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15279.9-15279.44|generated/sv2v_out.v:15279.5-15328.13" */ 2'h0 : _051_;
assign _005_ = _244_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15247.8-15271.15" */ _255_ : 1'h1;
assign _244_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15247.8-15271.15" */ _243_;
assign _243_[1] = instr_rdata_i[31:27] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15247.8-15271.15" */ 5'h08;
assign _003_ = instr_rdata_i[26] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15244.11-15244.20|generated/sv2v_out.v:15244.7-15271.15" */ 1'h1 : _005_;
assign _173_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15236.9-15240.16" */ instr_rdata_i[26:25];
assign _070_ = _243_[0] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15226.7-15242.14" */ _255_ : 1'h1;
assign _243_[0] = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15226.7-15242.14" */ instr_rdata_i[31:27];
assign _056_ = instr_rdata_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15212.11-15212.20|generated/sv2v_out.v:15212.7-15213.28" */ 1'h1 : 1'h0;
assign _059_ = _075_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15195.5-15200.12" */ _056_ : 1'h1;
assign _221_ = instr_rdata_i[13:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15195.5-15200.12" */ 2'h2;
assign _222_ = instr_rdata_i[13:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15195.5-15200.12" */ 2'h1;
assign _247_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15195.5-15200.12" */ instr_rdata_i[13:12];
assign _047_ = _249_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15181.5-15184.12" */ 1'h0 : 1'h1;
assign _249_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15181.5-15184.12" */ { _245_[5:3], _241_, _229_, _175_ };
assign _175_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15181.5-15184.12" */ instr_rdata_i[14:12];
assign _229_ = instr_rdata_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15181.5-15184.12" */ 3'h1;
assign _245_[3] = instr_rdata_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15181.5-15184.12" */ 3'h4;
assign _241_ = instr_rdata_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15181.5-15184.12" */ 3'h5;
assign _245_[4] = instr_rdata_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15181.5-15184.12" */ 3'h6;
assign _245_[5] = instr_rdata_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15181.5-15184.12" */ 3'h7;
assign _028_ = _182_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15175.9-15175.31|generated/sv2v_out.v:15175.5-15176.26" */ 1'h1 : 1'h0;
assign _032_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15169.9-15169.28|generated/sv2v_out.v:15169.5-15174.19" */ 1'h1 : 1'h0;
assign _253_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ 7'h17;
assign _254_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ 7'h37;
assign _252_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ 7'h6f;
assign _008_ = _250_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ 1'h1 : 1'h0;
assign data_sign_extension_o = _246_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ _071_ : 1'h0;
assign data_type_o = _099_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ _022_ : 2'h0;
assign multdiv_signed_mode_o = _240_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ _036_ : 2'h0;
assign multdiv_operator_o = _240_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ _035_ : 2'h0;
assign rf_wdata_sel_o = _223_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ _020_ : 1'h0;
assign wfi_insn_o = _223_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ _039_ : 1'h0;
assign ecall_insn_o = _223_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ _026_ : 1'h0;
assign dret_insn_o = _223_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ _024_ : 1'h0;
assign mret_insn_o = _223_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ _033_ : 1'h0;
assign ebrk_insn_o = _223_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ _025_ : 1'h0;
assign rf_ren_b_o = _085_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ 1'h1 : 1'h0;
assign _240_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ 7'h33;
assign _242_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ 7'h13;
assign _246_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ 7'h03;
assign _248_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ 7'h23;
assign _250_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ 7'h63;
assign _251_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ 7'h67;
assign icache_inval_o = _230_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ _027_ : 1'h0;
assign _230_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ 7'h0f;
assign csr_op = _223_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ _021_ : 2'h0;
assign _223_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ 7'h73;
assign _010_ = _248_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ 1'h1 : 1'h0;
assign _009_ = _099_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15157.3-15371.10" */ 1'h1 : 1'h0;
assign csr_op_o = _179_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15129.7-15129.75|generated/sv2v_out.v:15129.3-15130.20" */ 2'h0 : csr_op;
assign _255_ = _173_ ? /* src = "generated/sv2v_out.v:15248.45-15248.80" */ 1'h0 : 1'h1;
assign _060_ = branch_taken_i ? /* src = "generated/sv2v_out.v:15456.25-15456.53" */ 3'h2 : 3'h5;
assign mult_en_o = illegal_insn_o ? /* src = "generated/sv2v_out.v:15836.22-15836.54" */ 1'h0 : mult_sel_o;
assign div_en_o = illegal_insn_o ? /* src = "generated/sv2v_out.v:15837.21-15837.52" */ 1'h0 : div_sel_o;
assign _245_[0] = _175_;
assign alu_multicycle_o = 1'h0;
assign alu_multicycle_o_t0 = 1'h0;
assign alu_op_a_mux_sel_o_t0 = 2'h0;
assign alu_op_b_mux_sel_o_t0 = 1'h0;
assign alu_operator_o_t0 = 7'h00;
assign branch_in_dec_o_t0 = 1'h0;
assign bt_a_mux_sel_o = 2'h2;
assign bt_a_mux_sel_o_t0 = 2'h0;
assign bt_b_mux_sel_o = 3'h0;
assign bt_b_mux_sel_o_t0 = 3'h0;
assign csr_access_o_t0 = 1'h0;
assign csr_op_o_t0 = 2'h0;
assign data_req_o_t0 = 1'h0;
assign data_type_o_t0 = 2'h0;
assign data_we_o_t0 = 1'h0;
assign div_en_o_t0 = 1'h0;
assign div_sel_o_t0 = 1'h0;
assign dret_insn_o_t0 = 1'h0;
assign ebrk_insn_o_t0 = 1'h0;
assign ecall_insn_o_t0 = 1'h0;
assign icache_inval_o_t0 = 1'h0;
assign illegal_insn_o_t0 = 1'h0;
assign imm_a_mux_sel_o_t0 = 1'h0;
assign imm_b_mux_sel_o_t0 = 3'h0;
assign imm_b_type_o = { instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[7], instr_rdata_i[30:25], instr_rdata_i[11:8], 1'h0 };
assign imm_b_type_o_t0 = { instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[7], instr_rdata_i_t0[30:25], instr_rdata_i_t0[11:8], 1'h0 };
assign imm_i_type_o = { instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31:20] };
assign imm_i_type_o_t0 = { instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31:20] };
assign imm_j_type_o = { instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[19:12], instr_rdata_i[20], instr_rdata_i[30:21], 1'h0 };
assign imm_j_type_o_t0 = { instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[19:12], instr_rdata_i_t0[20], instr_rdata_i_t0[30:21], 1'h0 };
assign imm_s_type_o = { instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31:25], instr_rdata_i[11:7] };
assign imm_s_type_o_t0 = { instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31:25], instr_rdata_i_t0[11:7] };
assign imm_u_type_o = { instr_rdata_i[31:12], 12'h000 };
assign imm_u_type_o_t0 = { instr_rdata_i_t0[31:12], 12'h000 };
assign jump_in_dec_o_t0 = 1'h0;
assign jump_set_o_t0 = 1'h0;
assign mret_insn_o_t0 = 1'h0;
assign mult_en_o_t0 = 1'h0;
assign mult_sel_o_t0 = 1'h0;
assign multdiv_operator_o_t0 = 2'h0;
assign multdiv_signed_mode_o_t0 = 2'h0;
assign rf_raddr_a_o = instr_rdata_i[19:15];
assign rf_raddr_a_o_t0 = instr_rdata_i_t0[19:15];
assign rf_raddr_b_o = instr_rdata_i[24:20];
assign rf_raddr_b_o_t0 = instr_rdata_i_t0[24:20];
assign rf_ren_a_o_t0 = 1'h0;
assign rf_ren_b_o_t0 = 1'h0;
assign rf_waddr_o = instr_rdata_i[11:7];
assign rf_waddr_o_t0 = instr_rdata_i_t0[11:7];
assign rf_wdata_sel_o_t0 = 1'h0;
assign rf_we_o_t0 = 1'h0;
assign wfi_insn_o_t0 = 1'h0;
assign zimm_rs1_type_o = { 27'h0000000, instr_rdata_i[19:15] };
assign zimm_rs1_type_o_t0 = { 27'h0000000, instr_rdata_i_t0[19:15] };
endmodule

module \$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _0_;
wire [31:0] _1_;
wire [31:0] _2_;
wire [31:0] _3_;
/* src = "generated/sv2v_out.v:14936.13-14936.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14940.28-14940.37" */
output [31:0] rd_data_o;
reg [31:0] rd_data_o;
/* cellift = 32'd1 */
output [31:0] rd_data_o_t0;
reg [31:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14941.14-14941.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14937.13-14937.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14938.27-14938.36" */
input [31:0] wr_data_i;
wire [31:0] wr_data_i;
/* cellift = 32'd1 */
input [31:0] wr_data_i_t0;
wire [31:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14939.13-14939.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _0_ = ~ wr_en_i;
assign _1_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _2_ = { _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_ } & rd_data_o_t0;
assign _3_ = _1_ | _2_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 32'd0;
else rd_data_o_t0 <= _3_;
/* src = "generated/sv2v_out.v:14943.2-14947.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 32'd0;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$8d906854a94bfc59042b9faf57c7a7f19e3f03e7\ibex_core (clk_i, rst_ni, hart_id_i, boot_addr_i, instr_req_o, instr_gnt_i, instr_rvalid_i, instr_addr_o, instr_rdata_i, instr_err_i, data_req_o, data_gnt_i, data_rvalid_i, data_we_o, data_be_o, data_addr_o, data_wdata_o, data_rdata_i, data_err_i, dummy_instr_id_o, dummy_instr_wb_o
, rf_raddr_a_o, rf_raddr_b_o, rf_waddr_wb_o, rf_we_wb_o, rf_wdata_wb_ecc_o, rf_rdata_a_ecc_i, rf_rdata_b_ecc_i, ic_tag_req_o, ic_tag_write_o, ic_tag_addr_o, ic_tag_wdata_o, ic_tag_rdata_i, ic_data_req_o, ic_data_write_o, ic_data_addr_o, ic_data_wdata_o, ic_data_rdata_i, ic_scr_key_valid_i, ic_scr_key_req_o, irq_software_i, irq_timer_i
, irq_external_i, irq_fast_i, irq_nm_i, irq_pending_o, debug_req_i, crash_dump_o, double_fault_seen_o, fetch_enable_i, alert_minor_o, alert_major_internal_o, alert_major_bus_o, core_busy_o, debug_req_i_t0, ic_tag_write_o_t0, ic_tag_wdata_o_t0, ic_tag_req_o_t0, ic_tag_rdata_i_t0, ic_tag_addr_o_t0, ic_scr_key_valid_i_t0, ic_scr_key_req_o_t0, ic_data_write_o_t0
, ic_data_wdata_o_t0, ic_data_req_o_t0, ic_data_rdata_i_t0, ic_data_addr_o_t0, dummy_instr_id_o_t0, boot_addr_i_t0, irq_nm_i_t0, rf_raddr_b_o_t0, rf_raddr_a_o_t0, data_we_o_t0, data_req_o_t0, instr_rvalid_i_t0, instr_req_o_t0, instr_rdata_i_t0, instr_gnt_i_t0, instr_err_i_t0, instr_addr_o_t0, data_addr_o_t0, data_be_o_t0, data_gnt_i_t0, data_rdata_i_t0
, data_rvalid_i_t0, data_wdata_o_t0, dummy_instr_wb_o_t0, rf_waddr_wb_o_t0, rf_we_wb_o_t0, double_fault_seen_o_t0, hart_id_i_t0, irq_external_i_t0, irq_fast_i_t0, irq_pending_o_t0, irq_software_i_t0, irq_timer_i_t0, alert_major_bus_o_t0, alert_major_internal_o_t0, alert_minor_o_t0, core_busy_o_t0, crash_dump_o_t0, data_err_i_t0, fetch_enable_i_t0, rf_rdata_a_ecc_i_t0, rf_rdata_b_ecc_i_t0
, rf_wdata_wb_ecc_o_t0);
/* src = "generated/sv2v_out.v:13479.30-13479.54" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13479.30-13479.54" */
wire _001_;
/* src = "generated/sv2v_out.v:13480.30-13480.54" */
wire _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13480.30-13480.54" */
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
/* src = "generated/sv2v_out.v:13206.41-13206.56" */
wire _056_;
/* src = "generated/sv2v_out.v:13479.58-13479.75" */
wire _057_;
/* src = "generated/sv2v_out.v:13480.58-13480.75" */
wire _058_;
/* src = "generated/sv2v_out.v:13481.47-13481.80" */
wire _059_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13481.47-13481.80" */
wire _060_;
/* src = "generated/sv2v_out.v:13505.35-13505.70" */
wire _061_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13505.35-13505.70" */
wire _062_;
/* src = "generated/sv2v_out.v:13506.30-13506.78" */
wire _063_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13506.30-13506.78" */
wire _064_;
/* src = "generated/sv2v_out.v:13118.30-13118.81" */
wire _065_;
/* src = "generated/sv2v_out.v:13118.30-13118.81" */
wire _066_;
/* src = "generated/sv2v_out.v:13479.30-13479.43" */
wire _067_;
/* src = "generated/sv2v_out.v:13480.30-13480.43" */
wire _068_;
/* src = "generated/sv2v_out.v:12939.14-12939.31" */
output alert_major_bus_o;
wire alert_major_bus_o;
/* cellift = 32'd1 */
output alert_major_bus_o_t0;
wire alert_major_bus_o_t0;
/* src = "generated/sv2v_out.v:12938.14-12938.36" */
output alert_major_internal_o;
wire alert_major_internal_o;
/* cellift = 32'd1 */
output alert_major_internal_o_t0;
wire alert_major_internal_o_t0;
/* src = "generated/sv2v_out.v:12937.14-12937.27" */
output alert_minor_o;
wire alert_minor_o;
/* cellift = 32'd1 */
output alert_minor_o_t0;
wire alert_minor_o_t0;
/* src = "generated/sv2v_out.v:13016.14-13016.33" */
wire [31:0] alu_adder_result_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13016.14-13016.33" */
wire [31:0] alu_adder_result_ex_t0;
/* src = "generated/sv2v_out.v:13012.14-13012.30" */
wire [31:0] alu_operand_a_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13012.14-13012.30" */
wire [31:0] alu_operand_a_ex_t0;
/* src = "generated/sv2v_out.v:13013.14-13013.30" */
wire [31:0] alu_operand_b_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13013.14-13013.30" */
wire [31:0] alu_operand_b_ex_t0;
/* src = "generated/sv2v_out.v:13011.13-13011.28" */
wire [6:0] alu_operator_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13011.13-13011.28" */
wire [6:0] alu_operator_ex_t0;
/* src = "generated/sv2v_out.v:12890.20-12890.31" */
input [31:0] boot_addr_i;
wire [31:0] boot_addr_i;
/* cellift = 32'd1 */
input [31:0] boot_addr_i_t0;
wire [31:0] boot_addr_i_t0;
/* src = "generated/sv2v_out.v:12989.7-12989.22" */
wire branch_decision;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12989.7-12989.22" */
wire branch_decision_t0;
/* src = "generated/sv2v_out.v:12988.14-12988.30" */
wire [31:0] branch_target_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12988.14-12988.30" */
wire [31:0] branch_target_ex_t0;
/* src = "generated/sv2v_out.v:13014.14-13014.26" */
wire [31:0] bt_a_operand;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13014.14-13014.26" */
wire [31:0] bt_a_operand_t0;
/* src = "generated/sv2v_out.v:13015.14-13015.26" */
wire [31:0] bt_b_operand;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13015.14-13015.26" */
wire [31:0] bt_b_operand_t0;
/* src = "generated/sv2v_out.v:12887.13-12887.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:12940.20-12940.31" */
output [3:0] core_busy_o;
wire [3:0] core_busy_o;
/* cellift = 32'd1 */
output [3:0] core_busy_o_t0;
wire [3:0] core_busy_o_t0;
/* src = "generated/sv2v_out.v:13498.14-13498.30" */
wire [31:0] crash_dump_mtval;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13498.14-13498.30" */
wire [31:0] crash_dump_mtval_t0;
/* src = "generated/sv2v_out.v:12934.22-12934.34" */
output [159:0] crash_dump_o;
wire [159:0] crash_dump_o;
/* cellift = 32'd1 */
output [159:0] crash_dump_o_t0;
wire [159:0] crash_dump_o_t0;
/* src = "generated/sv2v_out.v:13027.7-13027.17" */
wire csr_access;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13027.7-13027.17" */
wire csr_access_t0;
/* src = "generated/sv2v_out.v:13030.14-13030.22" */
wire [11:0] csr_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13030.14-13030.22" */
wire [11:0] csr_addr_t0;
/* src = "generated/sv2v_out.v:13058.14-13058.22" */
wire [31:0] csr_depc;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13058.14-13058.22" */
wire [31:0] csr_depc_t0;
/* src = "generated/sv2v_out.v:13057.14-13057.22" */
wire [31:0] csr_mepc;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13057.14-13057.22" */
wire [31:0] csr_mepc_t0;
/* src = "generated/sv2v_out.v:13056.7-13056.22" */
wire csr_mstatus_mie;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13056.7-13056.22" */
wire csr_mstatus_mie_t0;
/* src = "generated/sv2v_out.v:13073.7-13073.21" */
wire csr_mstatus_tw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13073.7-13073.21" */
wire csr_mstatus_tw_t0;
/* src = "generated/sv2v_out.v:13072.14-13072.23" */
wire [31:0] csr_mtval;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13072.14-13072.23" */
wire [31:0] csr_mtval_t0;
/* src = "generated/sv2v_out.v:13071.14-13071.23" */
wire [31:0] csr_mtvec;
/* src = "generated/sv2v_out.v:13070.7-13070.21" */
wire csr_mtvec_init;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13070.7-13070.21" */
wire csr_mtvec_init_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13071.14-13071.23" */
wire [31:0] csr_mtvec_t0;
/* src = "generated/sv2v_out.v:13028.13-13028.19" */
wire [1:0] csr_op;
/* src = "generated/sv2v_out.v:13029.7-13029.16" */
wire csr_op_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13029.7-13029.16" */
wire csr_op_en_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13028.13-13028.19" */
wire [1:0] csr_op_t0;
/* src = "generated/sv2v_out.v:13059.36-13059.48" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135" */
wire [135:0] csr_pmp_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13059.36-13059.48" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135" */
wire [135:0] csr_pmp_addr_t0;
/* src = "generated/sv2v_out.v:13060.35-13060.46" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23" */
wire [23:0] csr_pmp_cfg;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13060.35-13060.46" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23" */
wire [23:0] csr_pmp_cfg_t0;
/* src = "generated/sv2v_out.v:13061.13-13061.28" */
/* unused_bits = "0 1 2" */
wire [2:0] csr_pmp_mseccfg;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13061.13-13061.28" */
/* unused_bits = "0 1 2" */
wire [2:0] csr_pmp_mseccfg_t0;
/* src = "generated/sv2v_out.v:13031.14-13031.23" */
wire [31:0] csr_rdata;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13031.14-13031.23" */
wire [31:0] csr_rdata_t0;
/* src = "generated/sv2v_out.v:13068.7-13068.26" */
wire csr_restore_dret_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13068.7-13068.26" */
wire csr_restore_dret_id_t0;
/* src = "generated/sv2v_out.v:13067.7-13067.26" */
wire csr_restore_mret_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13067.7-13067.26" */
wire csr_restore_mret_id_t0;
/* src = "generated/sv2v_out.v:13069.7-13069.21" */
wire csr_save_cause;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13069.7-13069.21" */
wire csr_save_cause_t0;
/* src = "generated/sv2v_out.v:13065.7-13065.18" */
wire csr_save_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13065.7-13065.18" */
wire csr_save_id_t0;
/* src = "generated/sv2v_out.v:13064.7-13064.18" */
wire csr_save_if;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13064.7-13064.18" */
wire csr_save_if_t0;
/* src = "generated/sv2v_out.v:13066.7-13066.18" */
wire csr_save_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13066.7-13066.18" */
wire csr_save_wb_t0;
/* src = "generated/sv2v_out.v:12972.7-12972.21" */
wire csr_shadow_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12972.7-12972.21" */
wire csr_shadow_err_t0;
/* src = "generated/sv2v_out.v:12990.7-12990.16" */
wire ctrl_busy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12990.7-12990.16" */
wire ctrl_busy_t0;
/* src = "generated/sv2v_out.v:12902.21-12902.32" */
output [31:0] data_addr_o;
wire [31:0] data_addr_o;
/* cellift = 32'd1 */
output [31:0] data_addr_o_t0;
wire [31:0] data_addr_o_t0;
/* src = "generated/sv2v_out.v:12901.20-12901.29" */
output [3:0] data_be_o;
wire [3:0] data_be_o;
/* cellift = 32'd1 */
output [3:0] data_be_o_t0;
wire [3:0] data_be_o_t0;
/* src = "generated/sv2v_out.v:12905.13-12905.23" */
input data_err_i;
wire data_err_i;
/* cellift = 32'd1 */
input data_err_i_t0;
wire data_err_i_t0;
/* src = "generated/sv2v_out.v:12898.13-12898.23" */
input data_gnt_i;
wire data_gnt_i;
/* cellift = 32'd1 */
input data_gnt_i_t0;
wire data_gnt_i_t0;
/* src = "generated/sv2v_out.v:12963.7-12963.22" */
wire data_ind_timing;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12963.7-12963.22" */
wire data_ind_timing_t0;
/* src = "generated/sv2v_out.v:12904.34-12904.46" */
input [38:0] data_rdata_i;
wire [38:0] data_rdata_i;
/* cellift = 32'd1 */
input [38:0] data_rdata_i_t0;
wire [38:0] data_rdata_i_t0;
/* src = "generated/sv2v_out.v:12897.14-12897.24" */
output data_req_o;
wire data_req_o;
/* cellift = 32'd1 */
output data_req_o_t0;
wire data_req_o_t0;
/* src = "generated/sv2v_out.v:12899.13-12899.26" */
input data_rvalid_i;
wire data_rvalid_i;
/* cellift = 32'd1 */
input data_rvalid_i_t0;
wire data_rvalid_i_t0;
/* src = "generated/sv2v_out.v:12903.35-12903.47" */
output [38:0] data_wdata_o;
wire [38:0] data_wdata_o;
/* cellift = 32'd1 */
output [38:0] data_wdata_o_t0;
wire [38:0] data_wdata_o_t0;
/* src = "generated/sv2v_out.v:12900.14-12900.23" */
output data_we_o;
wire data_we_o;
/* cellift = 32'd1 */
output data_we_o_t0;
wire data_we_o_t0;
/* src = "generated/sv2v_out.v:13078.13-13078.24" */
wire [2:0] debug_cause;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13078.13-13078.24" */
wire [2:0] debug_cause_t0;
/* src = "generated/sv2v_out.v:13079.7-13079.21" */
wire debug_csr_save;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13079.7-13079.21" */
wire debug_csr_save_t0;
/* src = "generated/sv2v_out.v:13081.7-13081.20" */
wire debug_ebreakm;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13081.7-13081.20" */
wire debug_ebreakm_t0;
/* src = "generated/sv2v_out.v:13082.7-13082.20" */
wire debug_ebreaku;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13082.7-13082.20" */
wire debug_ebreaku_t0;
/* src = "generated/sv2v_out.v:13076.7-13076.17" */
wire debug_mode;
/* src = "generated/sv2v_out.v:13077.7-13077.26" */
wire debug_mode_entering;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13077.7-13077.26" */
wire debug_mode_entering_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13076.7-13076.17" */
wire debug_mode_t0;
/* src = "generated/sv2v_out.v:12933.13-12933.24" */
input debug_req_i;
wire debug_req_i;
/* cellift = 32'd1 */
input debug_req_i_t0;
wire debug_req_i_t0;
/* src = "generated/sv2v_out.v:13080.7-13080.24" */
wire debug_single_step;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13080.7-13080.24" */
wire debug_single_step_t0;
/* src = "generated/sv2v_out.v:13019.7-13019.16" */
wire div_en_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13019.7-13019.16" */
wire div_en_ex_t0;
/* src = "generated/sv2v_out.v:13021.7-13021.17" */
wire div_sel_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13021.7-13021.17" */
wire div_sel_ex_t0;
/* src = "generated/sv2v_out.v:12935.14-12935.33" */
output double_fault_seen_o;
wire double_fault_seen_o;
/* cellift = 32'd1 */
output double_fault_seen_o_t0;
wire double_fault_seen_o_t0;
/* src = "generated/sv2v_out.v:12964.7-12964.21" */
wire dummy_instr_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12964.7-12964.21" */
wire dummy_instr_en_t0;
/* src = "generated/sv2v_out.v:12906.14-12906.30" */
output dummy_instr_id_o;
wire dummy_instr_id_o;
/* cellift = 32'd1 */
output dummy_instr_id_o_t0;
wire dummy_instr_id_o_t0;
/* src = "generated/sv2v_out.v:12965.13-12965.29" */
wire [2:0] dummy_instr_mask;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12965.13-12965.29" */
wire [2:0] dummy_instr_mask_t0;
/* src = "generated/sv2v_out.v:12967.14-12967.30" */
wire [31:0] dummy_instr_seed;
/* src = "generated/sv2v_out.v:12966.7-12966.26" */
wire dummy_instr_seed_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12966.7-12966.26" */
wire dummy_instr_seed_en_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12967.14-12967.30" */
wire [31:0] dummy_instr_seed_t0;
/* src = "generated/sv2v_out.v:12907.14-12907.30" */
output dummy_instr_wb_o;
wire dummy_instr_wb_o;
/* cellift = 32'd1 */
output dummy_instr_wb_o_t0;
wire dummy_instr_wb_o_t0;
/* src = "generated/sv2v_out.v:13047.7-13047.12" */
wire en_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13047.7-13047.12" */
wire en_wb_t0;
/* src = "generated/sv2v_out.v:13041.7-13041.15" */
wire ex_valid;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13041.7-13041.15" */
wire ex_valid_t0;
/* src = "generated/sv2v_out.v:12980.13-12980.22" */
wire [6:0] exc_cause;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12980.13-12980.22" */
wire [6:0] exc_cause_t0;
/* src = "generated/sv2v_out.v:12979.13-12979.26" */
wire [1:0] exc_pc_mux_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12979.13-12979.26" */
wire [1:0] exc_pc_mux_id_t0;
/* src = "generated/sv2v_out.v:12936.19-12936.33" */
input [3:0] fetch_enable_i;
wire [3:0] fetch_enable_i;
/* cellift = 32'd1 */
input [3:0] fetch_enable_i_t0;
wire [3:0] fetch_enable_i_t0;
/* src = "generated/sv2v_out.v:13107.16-13107.29" */
wire [11:0] \g_core_busy_secure.busy_bits_buf ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13107.16-13107.29" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11" */
wire [11:0] \g_core_busy_secure.busy_bits_buf_t0 ;
/* src = "generated/sv2v_out.v:13632.15-13632.33" */
/* unused_bits = "0 1" */
wire [1:0] \g_no_pmp.unused_priv_lvl_ls ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13632.15-13632.33" */
/* unused_bits = "0 1" */
wire [1:0] \g_no_pmp.unused_priv_lvl_ls_t0 ;
/* src = "generated/sv2v_out.v:13461.15-13461.27" */
wire [1:0] \gen_regfile_ecc.rf_ecc_err_a ;
/* src = "generated/sv2v_out.v:13463.9-13463.24" */
wire \gen_regfile_ecc.rf_ecc_err_a_id ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13463.9-13463.24" */
wire \gen_regfile_ecc.rf_ecc_err_a_id_t0 ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13461.15-13461.27" */
/* unused_bits = "0 1" */
wire [1:0] \gen_regfile_ecc.rf_ecc_err_a_t0 ;
/* src = "generated/sv2v_out.v:13462.15-13462.27" */
wire [1:0] \gen_regfile_ecc.rf_ecc_err_b ;
/* src = "generated/sv2v_out.v:13464.9-13464.24" */
wire \gen_regfile_ecc.rf_ecc_err_b_id ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13464.9-13464.24" */
wire \gen_regfile_ecc.rf_ecc_err_b_id_t0 ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13462.15-13462.27" */
/* unused_bits = "0 1" */
wire [1:0] \gen_regfile_ecc.rf_ecc_err_b_t0 ;
/* src = "generated/sv2v_out.v:12889.20-12889.29" */
input [31:0] hart_id_i;
wire [31:0] hart_id_i;
/* cellift = 32'd1 */
input [31:0] hart_id_i_t0;
wire [31:0] hart_id_i_t0;
/* src = "generated/sv2v_out.v:12922.42-12922.56" */
output [7:0] ic_data_addr_o;
wire [7:0] ic_data_addr_o;
/* cellift = 32'd1 */
output [7:0] ic_data_addr_o_t0;
wire [7:0] ic_data_addr_o_t0;
/* src = "generated/sv2v_out.v:12924.58-12924.73" */
input [127:0] ic_data_rdata_i;
wire [127:0] ic_data_rdata_i;
/* cellift = 32'd1 */
input [127:0] ic_data_rdata_i_t0;
wire [127:0] ic_data_rdata_i_t0;
/* src = "generated/sv2v_out.v:12920.20-12920.33" */
output [1:0] ic_data_req_o;
wire [1:0] ic_data_req_o;
/* cellift = 32'd1 */
output [1:0] ic_data_req_o_t0;
wire [1:0] ic_data_req_o_t0;
/* src = "generated/sv2v_out.v:12923.34-12923.49" */
output [63:0] ic_data_wdata_o;
wire [63:0] ic_data_wdata_o;
/* cellift = 32'd1 */
output [63:0] ic_data_wdata_o_t0;
wire [63:0] ic_data_wdata_o_t0;
/* src = "generated/sv2v_out.v:12921.14-12921.29" */
output ic_data_write_o;
wire ic_data_write_o;
/* cellift = 32'd1 */
output ic_data_write_o_t0;
wire ic_data_write_o_t0;
/* src = "generated/sv2v_out.v:12926.14-12926.30" */
output ic_scr_key_req_o;
wire ic_scr_key_req_o;
/* cellift = 32'd1 */
output ic_scr_key_req_o_t0;
wire ic_scr_key_req_o_t0;
/* src = "generated/sv2v_out.v:12925.13-12925.31" */
input ic_scr_key_valid_i;
wire ic_scr_key_valid_i;
/* cellift = 32'd1 */
input ic_scr_key_valid_i_t0;
wire ic_scr_key_valid_i_t0;
/* src = "generated/sv2v_out.v:12917.42-12917.55" */
output [7:0] ic_tag_addr_o;
wire [7:0] ic_tag_addr_o;
/* cellift = 32'd1 */
output [7:0] ic_tag_addr_o_t0;
wire [7:0] ic_tag_addr_o_t0;
/* src = "generated/sv2v_out.v:12919.57-12919.71" */
input [43:0] ic_tag_rdata_i;
wire [43:0] ic_tag_rdata_i;
/* cellift = 32'd1 */
input [43:0] ic_tag_rdata_i_t0;
wire [43:0] ic_tag_rdata_i_t0;
/* src = "generated/sv2v_out.v:12915.20-12915.32" */
output [1:0] ic_tag_req_o;
wire [1:0] ic_tag_req_o;
/* cellift = 32'd1 */
output [1:0] ic_tag_req_o_t0;
wire [1:0] ic_tag_req_o_t0;
/* src = "generated/sv2v_out.v:12918.33-12918.47" */
output [21:0] ic_tag_wdata_o;
wire [21:0] ic_tag_wdata_o;
/* cellift = 32'd1 */
output [21:0] ic_tag_wdata_o_t0;
wire [21:0] ic_tag_wdata_o_t0;
/* src = "generated/sv2v_out.v:12916.14-12916.28" */
output ic_tag_write_o;
wire ic_tag_write_o;
/* cellift = 32'd1 */
output ic_tag_write_o_t0;
wire ic_tag_write_o_t0;
/* src = "generated/sv2v_out.v:12968.7-12968.20" */
wire icache_enable;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12968.7-12968.20" */
wire icache_enable_t0;
/* src = "generated/sv2v_out.v:12969.7-12969.19" */
wire icache_inval;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12969.7-12969.19" */
wire icache_inval_t0;
/* src = "generated/sv2v_out.v:13040.7-13040.18" */
wire id_in_ready;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13040.7-13040.18" */
wire id_in_ready_t0;
/* src = "generated/sv2v_out.v:12991.7-12991.14" */
wire if_busy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12991.7-12991.14" */
wire if_busy_t0;
/* src = "generated/sv2v_out.v:12956.7-12956.24" */
wire illegal_c_insn_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12956.7-12956.24" */
wire illegal_c_insn_id_t0;
/* src = "generated/sv2v_out.v:13033.7-13033.26" */
wire illegal_csr_insn_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13033.7-13033.26" */
wire illegal_csr_insn_id_t0;
/* src = "generated/sv2v_out.v:13099.7-13099.22" */
/* unused_bits = "0" */
wire illegal_insn_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13099.7-13099.22" */
/* unused_bits = "0" */
wire illegal_insn_id_t0;
/* src = "generated/sv2v_out.v:12960.14-12960.26" */
wire [67:0] imd_val_d_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12960.14-12960.26" */
wire [67:0] imd_val_d_ex_t0;
/* src = "generated/sv2v_out.v:12961.14-12961.26" */
wire [67:0] imd_val_q_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12961.14-12961.26" */
wire [67:0] imd_val_q_ex_t0;
/* src = "generated/sv2v_out.v:12962.13-12962.26" */
wire [1:0] imd_val_we_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12962.13-12962.26" */
wire [1:0] imd_val_we_ex_t0;
/* src = "generated/sv2v_out.v:12894.21-12894.33" */
output [31:0] instr_addr_o;
wire [31:0] instr_addr_o;
/* cellift = 32'd1 */
output [31:0] instr_addr_o_t0;
wire [31:0] instr_addr_o_t0;
/* src = "generated/sv2v_out.v:12953.7-12953.24" */
wire instr_bp_taken_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12953.7-12953.24" */
wire instr_bp_taken_id_t0;
/* src = "generated/sv2v_out.v:13085.7-13085.20" */
/* unused_bits = "0" */
wire instr_done_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13085.7-13085.20" */
/* unused_bits = "0" */
wire instr_done_wb_t0;
/* src = "generated/sv2v_out.v:12896.13-12896.24" */
input instr_err_i;
wire instr_err_i;
/* cellift = 32'd1 */
input instr_err_i_t0;
wire instr_err_i_t0;
/* src = "generated/sv2v_out.v:13046.7-13046.17" */
wire instr_exec;
/* src = "generated/sv2v_out.v:12954.7-12954.22" */
wire instr_fetch_err;
/* src = "generated/sv2v_out.v:12955.7-12955.28" */
wire instr_fetch_err_plus2;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12955.7-12955.28" */
wire instr_fetch_err_plus2_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12954.7-12954.22" */
wire instr_fetch_err_t0;
/* src = "generated/sv2v_out.v:12973.7-12973.27" */
wire instr_first_cycle_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12973.7-12973.27" */
wire instr_first_cycle_id_t0;
/* src = "generated/sv2v_out.v:12892.13-12892.24" */
input instr_gnt_i;
wire instr_gnt_i;
/* cellift = 32'd1 */
input instr_gnt_i_t0;
wire instr_gnt_i_t0;
/* src = "generated/sv2v_out.v:13084.7-13084.20" */
/* unused_bits = "0" */
wire instr_id_done;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13084.7-13084.20" */
/* unused_bits = "0" */
wire instr_id_done_t0;
/* src = "generated/sv2v_out.v:12981.7-12981.21" */
wire instr_intg_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12981.7-12981.21" */
wire instr_intg_err_t0;
/* src = "generated/sv2v_out.v:12951.7-12951.29" */
wire instr_is_compressed_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12951.7-12951.29" */
wire instr_is_compressed_id_t0;
/* src = "generated/sv2v_out.v:12947.7-12947.19" */
/* unused_bits = "0" */
wire instr_new_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12947.7-12947.19" */
/* unused_bits = "0" */
wire instr_new_id_t0;
/* src = "generated/sv2v_out.v:12952.7-12952.26" */
wire instr_perf_count_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12952.7-12952.26" */
wire instr_perf_count_id_t0;
/* src = "generated/sv2v_out.v:12949.14-12949.32" */
wire [31:0] instr_rdata_alu_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12949.14-12949.32" */
wire [31:0] instr_rdata_alu_id_t0;
/* src = "generated/sv2v_out.v:12950.14-12950.30" */
wire [15:0] instr_rdata_c_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12950.14-12950.30" */
wire [15:0] instr_rdata_c_id_t0;
/* src = "generated/sv2v_out.v:12895.34-12895.47" */
input [38:0] instr_rdata_i;
wire [38:0] instr_rdata_i;
/* cellift = 32'd1 */
input [38:0] instr_rdata_i_t0;
wire [38:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:12948.14-12948.28" */
wire [31:0] instr_rdata_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12948.14-12948.28" */
wire [31:0] instr_rdata_id_t0;
/* src = "generated/sv2v_out.v:13045.7-13045.22" */
wire instr_req_gated;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13045.7-13045.22" */
wire instr_req_gated_t0;
/* src = "generated/sv2v_out.v:13044.7-13044.20" */
wire instr_req_int;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13044.7-13044.20" */
wire instr_req_int_t0;
/* src = "generated/sv2v_out.v:12891.14-12891.25" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:12893.13-12893.27" */
input instr_rvalid_i;
wire instr_rvalid_i;
/* cellift = 32'd1 */
input instr_rvalid_i_t0;
wire instr_rvalid_i_t0;
/* src = "generated/sv2v_out.v:13048.13-13048.26" */
wire [1:0] instr_type_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13048.13-13048.26" */
wire [1:0] instr_type_wb_t0;
/* src = "generated/sv2v_out.v:12974.7-12974.24" */
wire instr_valid_clear;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12974.7-12974.24" */
wire instr_valid_clear_t0;
/* src = "generated/sv2v_out.v:12946.7-12946.21" */
wire instr_valid_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12946.7-12946.21" */
wire instr_valid_id_t0;
/* src = "generated/sv2v_out.v:12929.13-12929.27" */
input irq_external_i;
wire irq_external_i;
/* cellift = 32'd1 */
input irq_external_i_t0;
wire irq_external_i_t0;
/* src = "generated/sv2v_out.v:12930.20-12930.30" */
input [14:0] irq_fast_i;
wire [14:0] irq_fast_i;
/* cellift = 32'd1 */
input [14:0] irq_fast_i_t0;
wire [14:0] irq_fast_i_t0;
/* src = "generated/sv2v_out.v:12931.13-12931.21" */
input irq_nm_i;
wire irq_nm_i;
/* cellift = 32'd1 */
input irq_nm_i_t0;
wire irq_nm_i_t0;
/* src = "generated/sv2v_out.v:12932.14-12932.27" */
output irq_pending_o;
wire irq_pending_o;
/* cellift = 32'd1 */
output irq_pending_o_t0;
wire irq_pending_o_t0;
/* src = "generated/sv2v_out.v:12927.13-12927.27" */
input irq_software_i;
wire irq_software_i;
/* cellift = 32'd1 */
input irq_software_i_t0;
wire irq_software_i_t0;
/* src = "generated/sv2v_out.v:12928.13-12928.24" */
input irq_timer_i;
wire irq_timer_i;
/* cellift = 32'd1 */
input irq_timer_i_t0;
wire irq_timer_i_t0;
/* src = "generated/sv2v_out.v:13055.14-13055.18" */
wire [17:0] irqs;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13055.14-13055.18" */
wire [17:0] irqs_t0;
/* src = "generated/sv2v_out.v:12986.7-12986.24" */
wire lsu_addr_incr_req;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12986.7-12986.24" */
wire lsu_addr_incr_req_t0;
/* src = "generated/sv2v_out.v:12987.14-12987.27" */
wire [31:0] lsu_addr_last;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12987.14-12987.27" */
wire [31:0] lsu_addr_last_t0;
/* src = "generated/sv2v_out.v:12992.7-12992.15" */
wire lsu_busy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12992.7-12992.15" */
wire lsu_busy_t0;
/* src = "generated/sv2v_out.v:12982.7-12982.19" */
wire lsu_load_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12982.7-12982.19" */
wire lsu_load_err_t0;
/* src = "generated/sv2v_out.v:12984.7-12984.29" */
wire lsu_load_resp_intg_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12984.7-12984.29" */
wire lsu_load_resp_intg_err_t0;
/* src = "generated/sv2v_out.v:13037.7-13037.14" */
wire lsu_req;
/* src = "generated/sv2v_out.v:13039.7-13039.19" */
wire lsu_req_done;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13039.7-13039.19" */
wire lsu_req_done_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13037.7-13037.14" */
wire lsu_req_t0;
/* src = "generated/sv2v_out.v:13043.7-13043.19" */
wire lsu_resp_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13043.7-13043.19" */
wire lsu_resp_err_t0;
/* src = "generated/sv2v_out.v:13042.7-13042.21" */
wire lsu_resp_valid;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13042.7-13042.21" */
wire lsu_resp_valid_t0;
/* src = "generated/sv2v_out.v:13036.7-13036.19" */
wire lsu_sign_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13036.7-13036.19" */
wire lsu_sign_ext_t0;
/* src = "generated/sv2v_out.v:12983.7-12983.20" */
wire lsu_store_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12983.7-12983.20" */
wire lsu_store_err_t0;
/* src = "generated/sv2v_out.v:12985.7-12985.30" */
wire lsu_store_resp_intg_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12985.7-12985.30" */
wire lsu_store_resp_intg_err_t0;
/* src = "generated/sv2v_out.v:13035.13-13035.21" */
wire [1:0] lsu_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13035.13-13035.21" */
wire [1:0] lsu_type_t0;
/* src = "generated/sv2v_out.v:13038.14-13038.23" */
wire [31:0] lsu_wdata;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13038.14-13038.23" */
wire [31:0] lsu_wdata_t0;
/* src = "generated/sv2v_out.v:13034.7-13034.13" */
wire lsu_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13034.7-13034.13" */
wire lsu_we_t0;
/* src = "generated/sv2v_out.v:13018.7-13018.17" */
wire mult_en_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13018.7-13018.17" */
wire mult_en_ex_t0;
/* src = "generated/sv2v_out.v:13020.7-13020.18" */
wire mult_sel_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13020.7-13020.18" */
wire mult_sel_ex_t0;
/* src = "generated/sv2v_out.v:13024.14-13024.34" */
wire [31:0] multdiv_operand_a_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13024.14-13024.34" */
wire [31:0] multdiv_operand_a_ex_t0;
/* src = "generated/sv2v_out.v:13025.14-13025.34" */
wire [31:0] multdiv_operand_b_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13025.14-13025.34" */
wire [31:0] multdiv_operand_b_ex_t0;
/* src = "generated/sv2v_out.v:13022.13-13022.32" */
wire [1:0] multdiv_operator_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13022.13-13022.32" */
wire [1:0] multdiv_operator_ex_t0;
/* src = "generated/sv2v_out.v:13026.7-13026.23" */
wire multdiv_ready_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13026.7-13026.23" */
wire multdiv_ready_id_t0;
/* src = "generated/sv2v_out.v:13023.13-13023.35" */
wire [1:0] multdiv_signed_mode_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13023.13-13023.35" */
wire [1:0] multdiv_signed_mode_ex_t0;
/* src = "generated/sv2v_out.v:13054.7-13054.15" */
wire nmi_mode;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13054.7-13054.15" */
wire nmi_mode_t0;
/* src = "generated/sv2v_out.v:12977.14-12977.28" */
wire [31:0] nt_branch_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12977.14-12977.28" */
wire [31:0] nt_branch_addr_t0;
/* src = "generated/sv2v_out.v:12976.7-12976.27" */
wire nt_branch_mispredict;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12976.7-12976.27" */
wire nt_branch_mispredict_t0;
/* src = "generated/sv2v_out.v:13051.7-13051.26" */
wire outstanding_load_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13051.7-13051.26" */
wire outstanding_load_wb_t0;
/* src = "generated/sv2v_out.v:13052.7-13052.27" */
wire outstanding_store_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13052.7-13052.27" */
wire outstanding_store_wb_t0;
/* src = "generated/sv2v_out.v:12958.14-12958.19" */
wire [31:0] pc_id /* verilator public */;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12958.14-12958.19" */
wire [31:0] pc_id_t0 /* verilator public */;
/* src = "generated/sv2v_out.v:12957.14-12957.19" */
wire [31:0] pc_if;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12957.14-12957.19" */
wire [31:0] pc_if_t0;
/* src = "generated/sv2v_out.v:12971.7-12971.24" */
wire pc_mismatch_alert;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12971.7-12971.24" */
wire pc_mismatch_alert_t0;
/* src = "generated/sv2v_out.v:12978.13-12978.22" */
wire [2:0] pc_mux_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12978.13-12978.22" */
wire [2:0] pc_mux_id_t0;
/* src = "generated/sv2v_out.v:12975.7-12975.13" */
wire pc_set;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12975.7-12975.13" */
wire pc_set_t0;
/* src = "generated/sv2v_out.v:12959.14-12959.19" */
wire [31:0] pc_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12959.14-12959.19" */
wire [31:0] pc_wb_t0;
/* src = "generated/sv2v_out.v:13095.7-13095.18" */
wire perf_branch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13095.7-13095.18" */
wire perf_branch_t0;
/* src = "generated/sv2v_out.v:13093.7-13093.20" */
wire perf_div_wait;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13093.7-13093.20" */
wire perf_div_wait_t0;
/* src = "generated/sv2v_out.v:13091.7-13091.22" */
wire perf_dside_wait;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13091.7-13091.22" */
wire perf_dside_wait_t0;
/* src = "generated/sv2v_out.v:13087.7-13087.35" */
wire perf_instr_ret_compressed_wb;
/* src = "generated/sv2v_out.v:13089.7-13089.40" */
wire perf_instr_ret_compressed_wb_spec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13089.7-13089.40" */
wire perf_instr_ret_compressed_wb_spec_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13087.7-13087.35" */
wire perf_instr_ret_compressed_wb_t0;
/* src = "generated/sv2v_out.v:13086.7-13086.24" */
wire perf_instr_ret_wb;
/* src = "generated/sv2v_out.v:13088.7-13088.29" */
wire perf_instr_ret_wb_spec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13088.7-13088.29" */
wire perf_instr_ret_wb_spec_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13086.7-13086.24" */
wire perf_instr_ret_wb_t0;
/* src = "generated/sv2v_out.v:13090.7-13090.22" */
wire perf_iside_wait;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13090.7-13090.22" */
wire perf_iside_wait_t0;
/* src = "generated/sv2v_out.v:13094.7-13094.16" */
wire perf_jump;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13094.7-13094.16" */
wire perf_jump_t0;
/* src = "generated/sv2v_out.v:13097.7-13097.16" */
wire perf_load;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13097.7-13097.16" */
wire perf_load_t0;
/* src = "generated/sv2v_out.v:13092.7-13092.20" */
wire perf_mul_wait;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13092.7-13092.20" */
wire perf_mul_wait_t0;
/* src = "generated/sv2v_out.v:13098.7-13098.17" */
wire perf_store;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13098.7-13098.17" */
wire perf_store_t0;
/* src = "generated/sv2v_out.v:13096.7-13096.19" */
wire perf_tbranch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13096.7-13096.19" */
wire perf_tbranch_t0;
/* src = "generated/sv2v_out.v:13074.13-13074.25" */
wire [1:0] priv_mode_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13074.13-13074.25" */
wire [1:0] priv_mode_id_t0;
/* src = "generated/sv2v_out.v:13049.7-13049.15" */
wire ready_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13049.7-13049.15" */
wire ready_wb_t0;
/* src = "generated/sv2v_out.v:13017.14-13017.23" */
wire [31:0] result_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13017.14-13017.23" */
wire [31:0] result_ex_t0;
/* src = "generated/sv2v_out.v:13005.7-13005.22" */
wire rf_ecc_err_comb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13005.7-13005.22" */
wire rf_ecc_err_comb_t0;
/* src = "generated/sv2v_out.v:12908.20-12908.32" */
output [4:0] rf_raddr_a_o;
wire [4:0] rf_raddr_a_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_a_o_t0;
wire [4:0] rf_raddr_a_o_t0;
/* src = "generated/sv2v_out.v:12909.20-12909.32" */
output [4:0] rf_raddr_b_o;
wire [4:0] rf_raddr_b_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_b_o_t0;
wire [4:0] rf_raddr_b_o_t0;
/* src = "generated/sv2v_out.v:13009.7-13009.23" */
wire rf_rd_a_wb_match;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13009.7-13009.23" */
wire rf_rd_a_wb_match_t0;
/* src = "generated/sv2v_out.v:13010.7-13010.23" */
wire rf_rd_b_wb_match;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13010.7-13010.23" */
wire rf_rd_b_wb_match_t0;
/* src = "generated/sv2v_out.v:12913.38-12913.54" */
input [38:0] rf_rdata_a_ecc_i;
wire [38:0] rf_rdata_a_ecc_i;
/* cellift = 32'd1 */
input [38:0] rf_rdata_a_ecc_i_t0;
wire [38:0] rf_rdata_a_ecc_i_t0;
/* src = "generated/sv2v_out.v:12914.38-12914.54" */
input [38:0] rf_rdata_b_ecc_i;
wire [38:0] rf_rdata_b_ecc_i;
/* cellift = 32'd1 */
input [38:0] rf_rdata_b_ecc_i_t0;
wire [38:0] rf_rdata_b_ecc_i_t0;
/* src = "generated/sv2v_out.v:12997.7-12997.15" */
wire rf_ren_a;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12997.7-12997.15" */
wire rf_ren_a_t0;
/* src = "generated/sv2v_out.v:12998.7-12998.15" */
wire rf_ren_b;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12998.7-12998.15" */
wire rf_ren_b_t0;
/* src = "generated/sv2v_out.v:13006.13-13006.24" */
wire [4:0] rf_waddr_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13006.13-13006.24" */
wire [4:0] rf_waddr_id_t0;
/* src = "generated/sv2v_out.v:12910.20-12910.33" */
output [4:0] rf_waddr_wb_o;
wire [4:0] rf_waddr_wb_o;
/* cellift = 32'd1 */
output [4:0] rf_waddr_wb_o_t0;
wire [4:0] rf_waddr_wb_o_t0;
/* src = "generated/sv2v_out.v:13001.14-13001.29" */
wire [31:0] rf_wdata_fwd_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13001.14-13001.29" */
wire [31:0] rf_wdata_fwd_wb_t0;
/* src = "generated/sv2v_out.v:13007.14-13007.25" */
wire [31:0] rf_wdata_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13007.14-13007.25" */
wire [31:0] rf_wdata_id_t0;
/* src = "generated/sv2v_out.v:13002.14-13002.26" */
wire [31:0] rf_wdata_lsu;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13002.14-13002.26" */
wire [31:0] rf_wdata_lsu_t0;
/* src = "generated/sv2v_out.v:13000.14-13000.25" */
wire [31:0] rf_wdata_wb;
/* src = "generated/sv2v_out.v:12912.39-12912.56" */
output [38:0] rf_wdata_wb_ecc_o;
wire [38:0] rf_wdata_wb_ecc_o;
/* cellift = 32'd1 */
output [38:0] rf_wdata_wb_ecc_o_t0;
wire [38:0] rf_wdata_wb_ecc_o_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13000.14-13000.25" */
wire [31:0] rf_wdata_wb_t0;
/* src = "generated/sv2v_out.v:13008.7-13008.15" */
wire rf_we_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13008.7-13008.15" */
wire rf_we_id_t0;
/* src = "generated/sv2v_out.v:13004.7-13004.16" */
wire rf_we_lsu;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13004.7-13004.16" */
wire rf_we_lsu_t0;
/* src = "generated/sv2v_out.v:12911.14-12911.24" */
output rf_we_wb_o;
wire rf_we_wb_o;
/* cellift = 32'd1 */
output rf_we_wb_o_t0;
wire rf_we_wb_o_t0;
/* src = "generated/sv2v_out.v:13050.7-13050.18" */
wire rf_write_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13050.7-13050.18" */
wire rf_write_wb_t0;
/* src = "generated/sv2v_out.v:12888.13-12888.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:13083.7-13083.20" */
wire trigger_match;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13083.7-13083.20" */
wire trigger_match_t0;
assign perf_iside_wait = id_in_ready & /* src = "generated/sv2v_out.v:13206.27-13206.56" */ _056_;
assign instr_req_gated = instr_req_int & /* src = "generated/sv2v_out.v:13209.29-13209.84" */ instr_exec;
assign _000_ = _067_ & /* src = "generated/sv2v_out.v:13479.30-13479.54" */ rf_ren_a;
assign \gen_regfile_ecc.rf_ecc_err_a_id  = _000_ & /* src = "generated/sv2v_out.v:13479.29-13479.75" */ _057_;
assign _002_ = _068_ & /* src = "generated/sv2v_out.v:13480.30-13480.54" */ rf_ren_b;
assign \gen_regfile_ecc.rf_ecc_err_b_id  = _002_ & /* src = "generated/sv2v_out.v:13480.29-13480.75" */ _058_;
assign rf_ecc_err_comb = instr_valid_id & /* src = "generated/sv2v_out.v:13481.29-13481.81" */ _059_;
assign _016_ = id_in_ready_t0 & _056_;
assign instr_req_gated_t0 = instr_req_int_t0 & instr_exec;
assign _019_ = _001_ & _057_;
assign _022_ = _003_ & _058_;
assign _025_ = instr_valid_id_t0 & _059_;
assign _017_ = instr_valid_id_t0 & id_in_ready;
assign _001_ = rf_ren_a_t0 & _067_;
assign _020_ = rf_rd_a_wb_match_t0 & _000_;
assign _003_ = rf_ren_b_t0 & _068_;
assign _023_ = rf_rd_b_wb_match_t0 & _002_;
assign _026_ = _060_ & instr_valid_id;
assign _018_ = id_in_ready_t0 & instr_valid_id_t0;
assign _021_ = _001_ & rf_rd_a_wb_match_t0;
assign _024_ = _003_ & rf_rd_b_wb_match_t0;
assign _027_ = instr_valid_id_t0 & _060_;
assign _046_ = _016_ | _017_;
assign _047_ = _019_ | _020_;
assign _048_ = _022_ | _023_;
assign _049_ = _025_ | _026_;
assign perf_iside_wait_t0 = _046_ | _018_;
assign \gen_regfile_ecc.rf_ecc_err_a_id_t0  = _047_ | _021_;
assign \gen_regfile_ecc.rf_ecc_err_b_id_t0  = _048_ | _024_;
assign rf_ecc_err_comb_t0 = _049_ | _027_;
assign csr_addr_t0 = { csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access } & alu_operand_b_ex_t0[11:0];
assign _004_ = ~ lsu_load_err;
assign _005_ = ~ \gen_regfile_ecc.rf_ecc_err_a_id ;
assign _006_ = ~ rf_ecc_err_comb;
assign _007_ = ~ _061_;
assign _008_ = ~ lsu_load_resp_intg_err;
assign _009_ = ~ _063_;
assign _010_ = ~ lsu_store_err;
assign _011_ = ~ \gen_regfile_ecc.rf_ecc_err_b_id ;
assign _012_ = ~ pc_mismatch_alert;
assign _013_ = ~ csr_shadow_err;
assign _014_ = ~ lsu_store_resp_intg_err;
assign _015_ = ~ instr_intg_err;
assign _028_ = lsu_load_err_t0 & _010_;
assign _031_ = \gen_regfile_ecc.rf_ecc_err_a_id_t0  & _011_;
assign _034_ = rf_ecc_err_comb_t0 & _012_;
assign _037_ = _062_ & _013_;
assign _040_ = lsu_load_resp_intg_err_t0 & _014_;
assign _043_ = _064_ & _015_;
assign _029_ = lsu_store_err_t0 & _004_;
assign _032_ = \gen_regfile_ecc.rf_ecc_err_b_id_t0  & _005_;
assign _035_ = pc_mismatch_alert_t0 & _006_;
assign _038_ = csr_shadow_err_t0 & _007_;
assign _041_ = lsu_store_resp_intg_err_t0 & _008_;
assign _044_ = instr_intg_err_t0 & _009_;
assign _030_ = lsu_load_err_t0 & lsu_store_err_t0;
assign _033_ = \gen_regfile_ecc.rf_ecc_err_a_id_t0  & \gen_regfile_ecc.rf_ecc_err_b_id_t0 ;
assign _036_ = rf_ecc_err_comb_t0 & pc_mismatch_alert_t0;
assign _039_ = _062_ & csr_shadow_err_t0;
assign _042_ = lsu_load_resp_intg_err_t0 & lsu_store_resp_intg_err_t0;
assign _045_ = _064_ & instr_intg_err_t0;
assign _050_ = _028_ | _029_;
assign _051_ = _031_ | _032_;
assign _052_ = _034_ | _035_;
assign _053_ = _037_ | _038_;
assign _054_ = _040_ | _041_;
assign _055_ = _043_ | _044_;
assign lsu_resp_err_t0 = _050_ | _030_;
assign _060_ = _051_ | _033_;
assign _062_ = _052_ | _036_;
assign alert_major_internal_o_t0 = _053_ | _039_;
assign _064_ = _054_ | _042_;
assign alert_major_bus_o_t0 = _055_ | _045_;
assign instr_exec = fetch_enable_i == /* src = "generated/sv2v_out.v:13210.24-13210.61" */ 4'h5;
assign core_busy_o[1] = ! /* src = "generated/sv2v_out.v:13118.30-13118.81" */ _065_;
assign core_busy_o[3] = ! /* src = "generated/sv2v_out.v:13118.30-13118.81" */ _066_;
assign _056_ = ~ /* src = "generated/sv2v_out.v:13206.41-13206.56" */ instr_valid_id;
assign _057_ = ~ /* src = "generated/sv2v_out.v:13479.58-13479.75" */ rf_rd_a_wb_match;
assign _058_ = ~ /* src = "generated/sv2v_out.v:13480.58-13480.75" */ rf_rd_b_wb_match;
assign lsu_resp_err = lsu_load_err | /* src = "generated/sv2v_out.v:13380.24-13380.52" */ lsu_store_err;
assign _059_ = \gen_regfile_ecc.rf_ecc_err_a_id  | /* src = "generated/sv2v_out.v:13481.47-13481.80" */ \gen_regfile_ecc.rf_ecc_err_b_id ;
assign _061_ = rf_ecc_err_comb | /* src = "generated/sv2v_out.v:13505.35-13505.70" */ pc_mismatch_alert;
assign alert_major_internal_o = _061_ | /* src = "generated/sv2v_out.v:13505.34-13505.88" */ csr_shadow_err;
assign _063_ = lsu_load_resp_intg_err | /* src = "generated/sv2v_out.v:13506.30-13506.78" */ lsu_store_resp_intg_err;
assign alert_major_bus_o = _063_ | /* src = "generated/sv2v_out.v:13506.29-13506.96" */ instr_intg_err;
assign core_busy_o[0] = | /* src = "generated/sv2v_out.v:13115.30-13115.80" */ \g_core_busy_secure.busy_bits_buf [2:0];
assign core_busy_o[2] = | /* src = "generated/sv2v_out.v:13115.30-13115.80" */ \g_core_busy_secure.busy_bits_buf [8:6];
assign _065_ = | /* src = "generated/sv2v_out.v:13118.30-13118.81" */ \g_core_busy_secure.busy_bits_buf [5:3];
assign _066_ = | /* src = "generated/sv2v_out.v:13118.30-13118.81" */ \g_core_busy_secure.busy_bits_buf [11:9];
assign _067_ = | /* src = "generated/sv2v_out.v:13479.30-13479.43" */ \gen_regfile_ecc.rf_ecc_err_a ;
assign _068_ = | /* src = "generated/sv2v_out.v:13480.30-13480.43" */ \gen_regfile_ecc.rf_ecc_err_b ;
assign csr_addr = csr_access ? /* src = "generated/sv2v_out.v:13512.34-13512.88" */ alu_operand_b_ex[11:0] : 12'h000;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13528.4-13600.3" */
\$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers  cs_registers_i (
.boot_addr_i(boot_addr_i),
.boot_addr_i_t0(boot_addr_i_t0),
.branch_i(perf_branch),
.branch_i_t0(perf_branch_t0),
.branch_taken_i(perf_tbranch),
.branch_taken_i_t0(perf_tbranch_t0),
.clk_i(clk_i),
.csr_access_i(csr_access),
.csr_access_i_t0(csr_access_t0),
.csr_addr_i(csr_addr),
.csr_addr_i_t0(csr_addr_t0),
.csr_depc_o(csr_depc),
.csr_depc_o_t0(csr_depc_t0),
.csr_mcause_i(exc_cause),
.csr_mcause_i_t0(exc_cause_t0),
.csr_mepc_o(csr_mepc),
.csr_mepc_o_t0(csr_mepc_t0),
.csr_mstatus_mie_o(csr_mstatus_mie),
.csr_mstatus_mie_o_t0(csr_mstatus_mie_t0),
.csr_mstatus_tw_o(csr_mstatus_tw),
.csr_mstatus_tw_o_t0(csr_mstatus_tw_t0),
.csr_mtval_i(csr_mtval),
.csr_mtval_i_t0(csr_mtval_t0),
.csr_mtval_o(crash_dump_mtval),
.csr_mtval_o_t0(crash_dump_mtval_t0),
.csr_mtvec_init_i(csr_mtvec_init),
.csr_mtvec_init_i_t0(csr_mtvec_init_t0),
.csr_mtvec_o(csr_mtvec),
.csr_mtvec_o_t0(csr_mtvec_t0),
.csr_op_en_i(csr_op_en),
.csr_op_en_i_t0(csr_op_en_t0),
.csr_op_i(csr_op),
.csr_op_i_t0(csr_op_t0),
.csr_pmp_addr_o(csr_pmp_addr),
.csr_pmp_addr_o_t0(csr_pmp_addr_t0),
.csr_pmp_cfg_o(csr_pmp_cfg),
.csr_pmp_cfg_o_t0(csr_pmp_cfg_t0),
.csr_pmp_mseccfg_o(csr_pmp_mseccfg),
.csr_pmp_mseccfg_o_t0(csr_pmp_mseccfg_t0),
.csr_rdata_o(csr_rdata),
.csr_rdata_o_t0(csr_rdata_t0),
.csr_restore_dret_i(csr_restore_dret_id),
.csr_restore_dret_i_t0(csr_restore_dret_id_t0),
.csr_restore_mret_i(csr_restore_mret_id),
.csr_restore_mret_i_t0(csr_restore_mret_id_t0),
.csr_save_cause_i(csr_save_cause),
.csr_save_cause_i_t0(csr_save_cause_t0),
.csr_save_id_i(csr_save_id),
.csr_save_id_i_t0(csr_save_id_t0),
.csr_save_if_i(csr_save_if),
.csr_save_if_i_t0(csr_save_if_t0),
.csr_save_wb_i(csr_save_wb),
.csr_save_wb_i_t0(csr_save_wb_t0),
.csr_shadow_err_o(csr_shadow_err),
.csr_shadow_err_o_t0(csr_shadow_err_t0),
.csr_wdata_i(alu_operand_a_ex),
.csr_wdata_i_t0(alu_operand_a_ex_t0),
.data_ind_timing_o(data_ind_timing),
.data_ind_timing_o_t0(data_ind_timing_t0),
.debug_cause_i(debug_cause),
.debug_cause_i_t0(debug_cause_t0),
.debug_csr_save_i(debug_csr_save),
.debug_csr_save_i_t0(debug_csr_save_t0),
.debug_ebreakm_o(debug_ebreakm),
.debug_ebreakm_o_t0(debug_ebreakm_t0),
.debug_ebreaku_o(debug_ebreaku),
.debug_ebreaku_o_t0(debug_ebreaku_t0),
.debug_mode_entering_i(debug_mode_entering),
.debug_mode_entering_i_t0(debug_mode_entering_t0),
.debug_mode_i(debug_mode),
.debug_mode_i_t0(debug_mode_t0),
.debug_single_step_o(debug_single_step),
.debug_single_step_o_t0(debug_single_step_t0),
.div_wait_i(perf_div_wait),
.div_wait_i_t0(perf_div_wait_t0),
.double_fault_seen_o(double_fault_seen_o),
.double_fault_seen_o_t0(double_fault_seen_o_t0),
.dside_wait_i(perf_dside_wait),
.dside_wait_i_t0(perf_dside_wait_t0),
.dummy_instr_en_o(dummy_instr_en),
.dummy_instr_en_o_t0(dummy_instr_en_t0),
.dummy_instr_mask_o(dummy_instr_mask),
.dummy_instr_mask_o_t0(dummy_instr_mask_t0),
.dummy_instr_seed_en_o(dummy_instr_seed_en),
.dummy_instr_seed_en_o_t0(dummy_instr_seed_en_t0),
.dummy_instr_seed_o(dummy_instr_seed),
.dummy_instr_seed_o_t0(dummy_instr_seed_t0),
.hart_id_i(hart_id_i),
.hart_id_i_t0(hart_id_i_t0),
.ic_scr_key_valid_i(ic_scr_key_valid_i),
.ic_scr_key_valid_i_t0(ic_scr_key_valid_i_t0),
.icache_enable_o(icache_enable),
.icache_enable_o_t0(icache_enable_t0),
.illegal_csr_insn_o(illegal_csr_insn_id),
.illegal_csr_insn_o_t0(illegal_csr_insn_id_t0),
.instr_ret_compressed_i(perf_instr_ret_compressed_wb),
.instr_ret_compressed_i_t0(perf_instr_ret_compressed_wb_t0),
.instr_ret_compressed_spec_i(perf_instr_ret_compressed_wb_spec),
.instr_ret_compressed_spec_i_t0(perf_instr_ret_compressed_wb_spec_t0),
.instr_ret_i(perf_instr_ret_wb),
.instr_ret_i_t0(perf_instr_ret_wb_t0),
.instr_ret_spec_i(perf_instr_ret_wb_spec),
.instr_ret_spec_i_t0(perf_instr_ret_wb_spec_t0),
.irq_external_i(irq_external_i),
.irq_external_i_t0(irq_external_i_t0),
.irq_fast_i(irq_fast_i),
.irq_fast_i_t0(irq_fast_i_t0),
.irq_pending_o(irq_pending_o),
.irq_pending_o_t0(irq_pending_o_t0),
.irq_software_i(irq_software_i),
.irq_software_i_t0(irq_software_i_t0),
.irq_timer_i(irq_timer_i),
.irq_timer_i_t0(irq_timer_i_t0),
.irqs_o(irqs),
.irqs_o_t0(irqs_t0),
.iside_wait_i(perf_iside_wait),
.iside_wait_i_t0(perf_iside_wait_t0),
.jump_i(perf_jump),
.jump_i_t0(perf_jump_t0),
.mem_load_i(perf_load),
.mem_load_i_t0(perf_load_t0),
.mem_store_i(perf_store),
.mem_store_i_t0(perf_store_t0),
.mul_wait_i(perf_mul_wait),
.mul_wait_i_t0(perf_mul_wait_t0),
.nmi_mode_i(nmi_mode),
.nmi_mode_i_t0(nmi_mode_t0),
.pc_id_i(pc_id),
.pc_id_i_t0(pc_id_t0),
.pc_if_i(pc_if),
.pc_if_i_t0(pc_if_t0),
.pc_wb_i(pc_wb),
.pc_wb_i_t0(pc_wb_t0),
.priv_mode_id_o(priv_mode_id),
.priv_mode_id_o_t0(priv_mode_id_t0),
.priv_mode_lsu_o(\g_no_pmp.unused_priv_lvl_ls ),
.priv_mode_lsu_o_t0(\g_no_pmp.unused_priv_lvl_ls_t0 ),
.rst_ni(rst_ni),
.trigger_match_o(trigger_match),
.trigger_match_o_t0(trigger_match_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13350.4-13377.3" */
\$paramod$a308247794889ee6093207090edbf289adef8be1\ibex_ex_block  ex_block_i (
.alu_adder_result_ex_o(alu_adder_result_ex),
.alu_adder_result_ex_o_t0(alu_adder_result_ex_t0),
.alu_instr_first_cycle_i(instr_first_cycle_id),
.alu_instr_first_cycle_i_t0(instr_first_cycle_id_t0),
.alu_operand_a_i(alu_operand_a_ex),
.alu_operand_a_i_t0(alu_operand_a_ex_t0),
.alu_operand_b_i(alu_operand_b_ex),
.alu_operand_b_i_t0(alu_operand_b_ex_t0),
.alu_operator_i(alu_operator_ex),
.alu_operator_i_t0(alu_operator_ex_t0),
.branch_decision_o(branch_decision),
.branch_decision_o_t0(branch_decision_t0),
.branch_target_o(branch_target_ex),
.branch_target_o_t0(branch_target_ex_t0),
.bt_a_operand_i(bt_a_operand),
.bt_a_operand_i_t0(bt_a_operand_t0),
.bt_b_operand_i(bt_b_operand),
.bt_b_operand_i_t0(bt_b_operand_t0),
.clk_i(clk_i),
.data_ind_timing_i(data_ind_timing),
.data_ind_timing_i_t0(data_ind_timing_t0),
.div_en_i(div_en_ex),
.div_en_i_t0(div_en_ex_t0),
.div_sel_i(div_sel_ex),
.div_sel_i_t0(div_sel_ex_t0),
.ex_valid_o(ex_valid),
.ex_valid_o_t0(ex_valid_t0),
.imd_val_d_o(imd_val_d_ex),
.imd_val_d_o_t0(imd_val_d_ex_t0),
.imd_val_q_i(imd_val_q_ex),
.imd_val_q_i_t0(imd_val_q_ex_t0),
.imd_val_we_o(imd_val_we_ex),
.imd_val_we_o_t0(imd_val_we_ex_t0),
.mult_en_i(mult_en_ex),
.mult_en_i_t0(mult_en_ex_t0),
.mult_sel_i(mult_sel_ex),
.mult_sel_i_t0(mult_sel_ex_t0),
.multdiv_operand_a_i(multdiv_operand_a_ex),
.multdiv_operand_a_i_t0(multdiv_operand_a_ex_t0),
.multdiv_operand_b_i(multdiv_operand_b_ex),
.multdiv_operand_b_i_t0(multdiv_operand_b_ex_t0),
.multdiv_operator_i(multdiv_operator_ex),
.multdiv_operator_i_t0(multdiv_operator_ex_t0),
.multdiv_ready_id_i(multdiv_ready_id),
.multdiv_ready_id_i_t0(multdiv_ready_id_t0),
.multdiv_signed_mode_i(multdiv_signed_mode_ex),
.multdiv_signed_mode_i_t0(multdiv_signed_mode_ex_t0),
.result_ex_o(result_ex),
.result_ex_o_t0(result_ex_t0),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13108.36-13111.5" */
\$paramod\prim_buf\Width=32'00000000000000000000000000001100  \g_core_busy_secure.u_fetch_enable_buf  (
.in_i({ ctrl_busy, if_busy, lsu_busy, ctrl_busy, if_busy, lsu_busy, ctrl_busy, if_busy, lsu_busy, ctrl_busy, if_busy, lsu_busy }),
.in_i_t0({ ctrl_busy_t0, if_busy_t0, lsu_busy_t0, ctrl_busy_t0, if_busy_t0, lsu_busy_t0, ctrl_busy_t0, if_busy_t0, lsu_busy_t0, ctrl_busy_t0, if_busy_t0, lsu_busy_t0 }),
.out_o(\g_core_busy_secure.busy_bits_buf ),
.out_o_t0(\g_core_busy_secure.busy_bits_buf_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13469.30-13472.5" */
prim_secded_inv_39_32_dec \gen_regfile_ecc.regfile_ecc_dec_a  (
.data_i(rf_rdata_a_ecc_i),
.data_i_t0(rf_rdata_a_ecc_i_t0),
.err_o(\gen_regfile_ecc.rf_ecc_err_a ),
.err_o_t0(\gen_regfile_ecc.rf_ecc_err_a_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13473.30-13476.5" */
prim_secded_inv_39_32_dec \gen_regfile_ecc.regfile_ecc_dec_b  (
.data_i(rf_rdata_b_ecc_i),
.data_i_t0(rf_rdata_b_ecc_i_t0),
.err_o(\gen_regfile_ecc.rf_ecc_err_b ),
.err_o_t0(\gen_regfile_ecc.rf_ecc_err_b_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13465.30-13468.5" */
prim_secded_inv_39_32_enc \gen_regfile_ecc.regfile_ecc_enc  (
.data_i(rf_wdata_wb),
.data_i_t0(rf_wdata_wb_t0),
.data_o(rf_wdata_wb_ecc_o),
.data_o_t0(rf_wdata_wb_ecc_o_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13228.4-13344.3" */
\$paramod$038d6e761af5e8bbfc2ed9b8473abfd849408d7b\ibex_id_stage  id_stage_i (
.alu_operand_a_ex_o(alu_operand_a_ex),
.alu_operand_a_ex_o_t0(alu_operand_a_ex_t0),
.alu_operand_b_ex_o(alu_operand_b_ex),
.alu_operand_b_ex_o_t0(alu_operand_b_ex_t0),
.alu_operator_ex_o(alu_operator_ex),
.alu_operator_ex_o_t0(alu_operator_ex_t0),
.branch_decision_i(branch_decision),
.branch_decision_i_t0(branch_decision_t0),
.bt_a_operand_o(bt_a_operand),
.bt_a_operand_o_t0(bt_a_operand_t0),
.bt_b_operand_o(bt_b_operand),
.bt_b_operand_o_t0(bt_b_operand_t0),
.clk_i(clk_i),
.csr_access_o(csr_access),
.csr_access_o_t0(csr_access_t0),
.csr_mstatus_mie_i(csr_mstatus_mie),
.csr_mstatus_mie_i_t0(csr_mstatus_mie_t0),
.csr_mstatus_tw_i(csr_mstatus_tw),
.csr_mstatus_tw_i_t0(csr_mstatus_tw_t0),
.csr_mtval_o(csr_mtval),
.csr_mtval_o_t0(csr_mtval_t0),
.csr_op_en_o(csr_op_en),
.csr_op_en_o_t0(csr_op_en_t0),
.csr_op_o(csr_op),
.csr_op_o_t0(csr_op_t0),
.csr_rdata_i(csr_rdata),
.csr_rdata_i_t0(csr_rdata_t0),
.csr_restore_dret_id_o(csr_restore_dret_id),
.csr_restore_dret_id_o_t0(csr_restore_dret_id_t0),
.csr_restore_mret_id_o(csr_restore_mret_id),
.csr_restore_mret_id_o_t0(csr_restore_mret_id_t0),
.csr_save_cause_o(csr_save_cause),
.csr_save_cause_o_t0(csr_save_cause_t0),
.csr_save_id_o(csr_save_id),
.csr_save_id_o_t0(csr_save_id_t0),
.csr_save_if_o(csr_save_if),
.csr_save_if_o_t0(csr_save_if_t0),
.csr_save_wb_o(csr_save_wb),
.csr_save_wb_o_t0(csr_save_wb_t0),
.ctrl_busy_o(ctrl_busy),
.ctrl_busy_o_t0(ctrl_busy_t0),
.data_ind_timing_i(data_ind_timing),
.data_ind_timing_i_t0(data_ind_timing_t0),
.debug_cause_o(debug_cause),
.debug_cause_o_t0(debug_cause_t0),
.debug_csr_save_o(debug_csr_save),
.debug_csr_save_o_t0(debug_csr_save_t0),
.debug_ebreakm_i(debug_ebreakm),
.debug_ebreakm_i_t0(debug_ebreakm_t0),
.debug_ebreaku_i(debug_ebreaku),
.debug_ebreaku_i_t0(debug_ebreaku_t0),
.debug_mode_entering_o(debug_mode_entering),
.debug_mode_entering_o_t0(debug_mode_entering_t0),
.debug_mode_o(debug_mode),
.debug_mode_o_t0(debug_mode_t0),
.debug_req_i(debug_req_i),
.debug_req_i_t0(debug_req_i_t0),
.debug_single_step_i(debug_single_step),
.debug_single_step_i_t0(debug_single_step_t0),
.div_en_ex_o(div_en_ex),
.div_en_ex_o_t0(div_en_ex_t0),
.div_sel_ex_o(div_sel_ex),
.div_sel_ex_o_t0(div_sel_ex_t0),
.en_wb_o(en_wb),
.en_wb_o_t0(en_wb_t0),
.ex_valid_i(ex_valid),
.ex_valid_i_t0(ex_valid_t0),
.exc_cause_o(exc_cause),
.exc_cause_o_t0(exc_cause_t0),
.exc_pc_mux_o(exc_pc_mux_id),
.exc_pc_mux_o_t0(exc_pc_mux_id_t0),
.icache_inval_o(icache_inval),
.icache_inval_o_t0(icache_inval_t0),
.id_in_ready_o(id_in_ready),
.id_in_ready_o_t0(id_in_ready_t0),
.illegal_c_insn_i(illegal_c_insn_id),
.illegal_c_insn_i_t0(illegal_c_insn_id_t0),
.illegal_csr_insn_i(illegal_csr_insn_id),
.illegal_csr_insn_i_t0(illegal_csr_insn_id_t0),
.illegal_insn_o(illegal_insn_id),
.illegal_insn_o_t0(illegal_insn_id_t0),
.imd_val_d_ex_i(imd_val_d_ex),
.imd_val_d_ex_i_t0(imd_val_d_ex_t0),
.imd_val_q_ex_o(imd_val_q_ex),
.imd_val_q_ex_o_t0(imd_val_q_ex_t0),
.imd_val_we_ex_i(imd_val_we_ex),
.imd_val_we_ex_i_t0(imd_val_we_ex_t0),
.instr_bp_taken_i(instr_bp_taken_id),
.instr_bp_taken_i_t0(instr_bp_taken_id_t0),
.instr_exec_i(instr_exec),
.instr_exec_i_t0(1'h0),
.instr_fetch_err_i(instr_fetch_err),
.instr_fetch_err_i_t0(instr_fetch_err_t0),
.instr_fetch_err_plus2_i(instr_fetch_err_plus2),
.instr_fetch_err_plus2_i_t0(instr_fetch_err_plus2_t0),
.instr_first_cycle_id_o(instr_first_cycle_id),
.instr_first_cycle_id_o_t0(instr_first_cycle_id_t0),
.instr_id_done_o(instr_id_done),
.instr_id_done_o_t0(instr_id_done_t0),
.instr_is_compressed_i(instr_is_compressed_id),
.instr_is_compressed_i_t0(instr_is_compressed_id_t0),
.instr_perf_count_id_o(instr_perf_count_id),
.instr_perf_count_id_o_t0(instr_perf_count_id_t0),
.instr_rdata_alu_i(instr_rdata_alu_id),
.instr_rdata_alu_i_t0(instr_rdata_alu_id_t0),
.instr_rdata_c_i(instr_rdata_c_id),
.instr_rdata_c_i_t0(instr_rdata_c_id_t0),
.instr_rdata_i(instr_rdata_id),
.instr_rdata_i_t0(instr_rdata_id_t0),
.instr_req_o(instr_req_int),
.instr_req_o_t0(instr_req_int_t0),
.instr_type_wb_o(instr_type_wb),
.instr_type_wb_o_t0(instr_type_wb_t0),
.instr_valid_clear_o(instr_valid_clear),
.instr_valid_clear_o_t0(instr_valid_clear_t0),
.instr_valid_i(instr_valid_id),
.instr_valid_i_t0(instr_valid_id_t0),
.irq_nm_i(irq_nm_i),
.irq_nm_i_t0(irq_nm_i_t0),
.irq_pending_i(irq_pending_o),
.irq_pending_i_t0(irq_pending_o_t0),
.irqs_i(irqs),
.irqs_i_t0(irqs_t0),
.lsu_addr_incr_req_i(lsu_addr_incr_req),
.lsu_addr_incr_req_i_t0(lsu_addr_incr_req_t0),
.lsu_addr_last_i(lsu_addr_last),
.lsu_addr_last_i_t0(lsu_addr_last_t0),
.lsu_load_err_i(lsu_load_err),
.lsu_load_err_i_t0(lsu_load_err_t0),
.lsu_load_resp_intg_err_i(lsu_load_resp_intg_err),
.lsu_load_resp_intg_err_i_t0(lsu_load_resp_intg_err_t0),
.lsu_req_done_i(lsu_req_done),
.lsu_req_done_i_t0(lsu_req_done_t0),
.lsu_req_o(lsu_req),
.lsu_req_o_t0(lsu_req_t0),
.lsu_resp_valid_i(lsu_resp_valid),
.lsu_resp_valid_i_t0(lsu_resp_valid_t0),
.lsu_sign_ext_o(lsu_sign_ext),
.lsu_sign_ext_o_t0(lsu_sign_ext_t0),
.lsu_store_err_i(lsu_store_err),
.lsu_store_err_i_t0(lsu_store_err_t0),
.lsu_store_resp_intg_err_i(lsu_store_resp_intg_err),
.lsu_store_resp_intg_err_i_t0(lsu_store_resp_intg_err_t0),
.lsu_type_o(lsu_type),
.lsu_type_o_t0(lsu_type_t0),
.lsu_wdata_o(lsu_wdata),
.lsu_wdata_o_t0(lsu_wdata_t0),
.lsu_we_o(lsu_we),
.lsu_we_o_t0(lsu_we_t0),
.mult_en_ex_o(mult_en_ex),
.mult_en_ex_o_t0(mult_en_ex_t0),
.mult_sel_ex_o(mult_sel_ex),
.mult_sel_ex_o_t0(mult_sel_ex_t0),
.multdiv_operand_a_ex_o(multdiv_operand_a_ex),
.multdiv_operand_a_ex_o_t0(multdiv_operand_a_ex_t0),
.multdiv_operand_b_ex_o(multdiv_operand_b_ex),
.multdiv_operand_b_ex_o_t0(multdiv_operand_b_ex_t0),
.multdiv_operator_ex_o(multdiv_operator_ex),
.multdiv_operator_ex_o_t0(multdiv_operator_ex_t0),
.multdiv_ready_id_o(multdiv_ready_id),
.multdiv_ready_id_o_t0(multdiv_ready_id_t0),
.multdiv_signed_mode_ex_o(multdiv_signed_mode_ex),
.multdiv_signed_mode_ex_o_t0(multdiv_signed_mode_ex_t0),
.nmi_mode_o(nmi_mode),
.nmi_mode_o_t0(nmi_mode_t0),
.nt_branch_addr_o(nt_branch_addr),
.nt_branch_addr_o_t0(nt_branch_addr_t0),
.nt_branch_mispredict_o(nt_branch_mispredict),
.nt_branch_mispredict_o_t0(nt_branch_mispredict_t0),
.outstanding_load_wb_i(outstanding_load_wb),
.outstanding_load_wb_i_t0(outstanding_load_wb_t0),
.outstanding_store_wb_i(outstanding_store_wb),
.outstanding_store_wb_i_t0(outstanding_store_wb_t0),
.pc_id_i(pc_id),
.pc_id_i_t0(pc_id_t0),
.pc_mux_o(pc_mux_id),
.pc_mux_o_t0(pc_mux_id_t0),
.pc_set_o(pc_set),
.pc_set_o_t0(pc_set_t0),
.perf_branch_o(perf_branch),
.perf_branch_o_t0(perf_branch_t0),
.perf_div_wait_o(perf_div_wait),
.perf_div_wait_o_t0(perf_div_wait_t0),
.perf_dside_wait_o(perf_dside_wait),
.perf_dside_wait_o_t0(perf_dside_wait_t0),
.perf_jump_o(perf_jump),
.perf_jump_o_t0(perf_jump_t0),
.perf_mul_wait_o(perf_mul_wait),
.perf_mul_wait_o_t0(perf_mul_wait_t0),
.perf_tbranch_o(perf_tbranch),
.perf_tbranch_o_t0(perf_tbranch_t0),
.priv_mode_i(priv_mode_id),
.priv_mode_i_t0(priv_mode_id_t0),
.ready_wb_i(ready_wb),
.ready_wb_i_t0(ready_wb_t0),
.result_ex_i(result_ex),
.result_ex_i_t0(result_ex_t0),
.rf_raddr_a_o(rf_raddr_a_o),
.rf_raddr_a_o_t0(rf_raddr_a_o_t0),
.rf_raddr_b_o(rf_raddr_b_o),
.rf_raddr_b_o_t0(rf_raddr_b_o_t0),
.rf_rd_a_wb_match_o(rf_rd_a_wb_match),
.rf_rd_a_wb_match_o_t0(rf_rd_a_wb_match_t0),
.rf_rd_b_wb_match_o(rf_rd_b_wb_match),
.rf_rd_b_wb_match_o_t0(rf_rd_b_wb_match_t0),
.rf_rdata_a_i(rf_rdata_a_ecc_i[31:0]),
.rf_rdata_a_i_t0(rf_rdata_a_ecc_i_t0[31:0]),
.rf_rdata_b_i(rf_rdata_b_ecc_i[31:0]),
.rf_rdata_b_i_t0(rf_rdata_b_ecc_i_t0[31:0]),
.rf_ren_a_o(rf_ren_a),
.rf_ren_a_o_t0(rf_ren_a_t0),
.rf_ren_b_o(rf_ren_b),
.rf_ren_b_o_t0(rf_ren_b_t0),
.rf_waddr_id_o(rf_waddr_id),
.rf_waddr_id_o_t0(rf_waddr_id_t0),
.rf_waddr_wb_i(rf_waddr_wb_o),
.rf_waddr_wb_i_t0(rf_waddr_wb_o_t0),
.rf_wdata_fwd_wb_i(rf_wdata_fwd_wb),
.rf_wdata_fwd_wb_i_t0(rf_wdata_fwd_wb_t0),
.rf_wdata_id_o(rf_wdata_id),
.rf_wdata_id_o_t0(rf_wdata_id_t0),
.rf_we_id_o(rf_we_id),
.rf_we_id_o_t0(rf_we_id_t0),
.rf_write_wb_i(rf_write_wb),
.rf_write_wb_i_t0(rf_write_wb_t0),
.rst_ni(rst_ni),
.trigger_match_i(trigger_match),
.trigger_match_i_t0(trigger_match_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13144.4-13205.3" */
\$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  if_stage_i (
.boot_addr_i(boot_addr_i),
.boot_addr_i_t0(boot_addr_i_t0),
.branch_target_ex_i(branch_target_ex),
.branch_target_ex_i_t0(branch_target_ex_t0),
.clk_i(clk_i),
.csr_depc_i(csr_depc),
.csr_depc_i_t0(csr_depc_t0),
.csr_mepc_i(csr_mepc),
.csr_mepc_i_t0(csr_mepc_t0),
.csr_mtvec_i(csr_mtvec),
.csr_mtvec_i_t0(csr_mtvec_t0),
.csr_mtvec_init_o(csr_mtvec_init),
.csr_mtvec_init_o_t0(csr_mtvec_init_t0),
.dummy_instr_en_i(dummy_instr_en),
.dummy_instr_en_i_t0(dummy_instr_en_t0),
.dummy_instr_id_o(dummy_instr_id_o),
.dummy_instr_id_o_t0(dummy_instr_id_o_t0),
.dummy_instr_mask_i(dummy_instr_mask),
.dummy_instr_mask_i_t0(dummy_instr_mask_t0),
.dummy_instr_seed_en_i(dummy_instr_seed_en),
.dummy_instr_seed_en_i_t0(dummy_instr_seed_en_t0),
.dummy_instr_seed_i(dummy_instr_seed),
.dummy_instr_seed_i_t0(dummy_instr_seed_t0),
.exc_cause(exc_cause),
.exc_cause_t0(exc_cause_t0),
.exc_pc_mux_i(exc_pc_mux_id),
.exc_pc_mux_i_t0(exc_pc_mux_id_t0),
.ic_data_addr_o(ic_data_addr_o),
.ic_data_addr_o_t0(ic_data_addr_o_t0),
.ic_data_rdata_i(ic_data_rdata_i),
.ic_data_rdata_i_t0(ic_data_rdata_i_t0),
.ic_data_req_o(ic_data_req_o),
.ic_data_req_o_t0(ic_data_req_o_t0),
.ic_data_wdata_o(ic_data_wdata_o),
.ic_data_wdata_o_t0(ic_data_wdata_o_t0),
.ic_data_write_o(ic_data_write_o),
.ic_data_write_o_t0(ic_data_write_o_t0),
.ic_scr_key_req_o(ic_scr_key_req_o),
.ic_scr_key_req_o_t0(ic_scr_key_req_o_t0),
.ic_scr_key_valid_i(ic_scr_key_valid_i),
.ic_scr_key_valid_i_t0(ic_scr_key_valid_i_t0),
.ic_tag_addr_o(ic_tag_addr_o),
.ic_tag_addr_o_t0(ic_tag_addr_o_t0),
.ic_tag_rdata_i(ic_tag_rdata_i),
.ic_tag_rdata_i_t0(ic_tag_rdata_i_t0),
.ic_tag_req_o(ic_tag_req_o),
.ic_tag_req_o_t0(ic_tag_req_o_t0),
.ic_tag_wdata_o(ic_tag_wdata_o),
.ic_tag_wdata_o_t0(ic_tag_wdata_o_t0),
.ic_tag_write_o(ic_tag_write_o),
.ic_tag_write_o_t0(ic_tag_write_o_t0),
.icache_ecc_error_o(alert_minor_o),
.icache_ecc_error_o_t0(alert_minor_o_t0),
.icache_enable_i(icache_enable),
.icache_enable_i_t0(icache_enable_t0),
.icache_inval_i(icache_inval),
.icache_inval_i_t0(icache_inval_t0),
.id_in_ready_i(id_in_ready),
.id_in_ready_i_t0(id_in_ready_t0),
.if_busy_o(if_busy),
.if_busy_o_t0(if_busy_t0),
.illegal_c_insn_id_o(illegal_c_insn_id),
.illegal_c_insn_id_o_t0(illegal_c_insn_id_t0),
.instr_addr_o(instr_addr_o),
.instr_addr_o_t0(instr_addr_o_t0),
.instr_bp_taken_o(instr_bp_taken_id),
.instr_bp_taken_o_t0(instr_bp_taken_id_t0),
.instr_bus_err_i(instr_err_i),
.instr_bus_err_i_t0(instr_err_i_t0),
.instr_fetch_err_o(instr_fetch_err),
.instr_fetch_err_o_t0(instr_fetch_err_t0),
.instr_fetch_err_plus2_o(instr_fetch_err_plus2),
.instr_fetch_err_plus2_o_t0(instr_fetch_err_plus2_t0),
.instr_gnt_i(instr_gnt_i),
.instr_gnt_i_t0(instr_gnt_i_t0),
.instr_intg_err_o(instr_intg_err),
.instr_intg_err_o_t0(instr_intg_err_t0),
.instr_is_compressed_id_o(instr_is_compressed_id),
.instr_is_compressed_id_o_t0(instr_is_compressed_id_t0),
.instr_new_id_o(instr_new_id),
.instr_new_id_o_t0(instr_new_id_t0),
.instr_rdata_alu_id_o(instr_rdata_alu_id),
.instr_rdata_alu_id_o_t0(instr_rdata_alu_id_t0),
.instr_rdata_c_id_o(instr_rdata_c_id),
.instr_rdata_c_id_o_t0(instr_rdata_c_id_t0),
.instr_rdata_i(instr_rdata_i),
.instr_rdata_i_t0(instr_rdata_i_t0),
.instr_rdata_id_o(instr_rdata_id),
.instr_rdata_id_o_t0(instr_rdata_id_t0),
.instr_req_o(instr_req_o),
.instr_req_o_t0(instr_req_o_t0),
.instr_rvalid_i(instr_rvalid_i),
.instr_rvalid_i_t0(instr_rvalid_i_t0),
.instr_valid_clear_i(instr_valid_clear),
.instr_valid_clear_i_t0(instr_valid_clear_t0),
.instr_valid_id_o(instr_valid_id),
.instr_valid_id_o_t0(instr_valid_id_t0),
.nt_branch_addr_i(nt_branch_addr),
.nt_branch_addr_i_t0(nt_branch_addr_t0),
.nt_branch_mispredict_i(nt_branch_mispredict),
.nt_branch_mispredict_i_t0(nt_branch_mispredict_t0),
.pc_id_o(pc_id),
.pc_id_o_t0(pc_id_t0),
.pc_if_o(pc_if),
.pc_if_o_t0(pc_if_t0),
.pc_mismatch_alert_o(pc_mismatch_alert),
.pc_mismatch_alert_o_t0(pc_mismatch_alert_t0),
.pc_mux_i(pc_mux_id),
.pc_mux_i_t0(pc_mux_id_t0),
.pc_set_i(pc_set),
.pc_set_i_t0(pc_set_t0),
.pmp_err_if_i(1'h0),
.pmp_err_if_i_t0(1'h0),
.pmp_err_if_plus2_i(1'h0),
.pmp_err_if_plus2_i_t0(1'h0),
.req_i(instr_req_gated),
.req_i_t0(instr_req_gated_t0),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13384.4-13416.3" */
\$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  load_store_unit_i (
.adder_result_ex_i(alu_adder_result_ex),
.adder_result_ex_i_t0(alu_adder_result_ex_t0),
.addr_incr_req_o(lsu_addr_incr_req),
.addr_incr_req_o_t0(lsu_addr_incr_req_t0),
.addr_last_o(lsu_addr_last),
.addr_last_o_t0(lsu_addr_last_t0),
.busy_o(lsu_busy),
.busy_o_t0(lsu_busy_t0),
.clk_i(clk_i),
.data_addr_o(data_addr_o),
.data_addr_o_t0(data_addr_o_t0),
.data_be_o(data_be_o),
.data_be_o_t0(data_be_o_t0),
.data_bus_err_i(data_err_i),
.data_bus_err_i_t0(data_err_i_t0),
.data_gnt_i(data_gnt_i),
.data_gnt_i_t0(data_gnt_i_t0),
.data_pmp_err_i(1'h0),
.data_pmp_err_i_t0(1'h0),
.data_rdata_i(data_rdata_i),
.data_rdata_i_t0(data_rdata_i_t0),
.data_req_o(data_req_o),
.data_req_o_t0(data_req_o_t0),
.data_rvalid_i(data_rvalid_i),
.data_rvalid_i_t0(data_rvalid_i_t0),
.data_wdata_o(data_wdata_o),
.data_wdata_o_t0(data_wdata_o_t0),
.data_we_o(data_we_o),
.data_we_o_t0(data_we_o_t0),
.load_err_o(lsu_load_err),
.load_err_o_t0(lsu_load_err_t0),
.load_resp_intg_err_o(lsu_load_resp_intg_err),
.load_resp_intg_err_o_t0(lsu_load_resp_intg_err_t0),
.lsu_rdata_o(rf_wdata_lsu),
.lsu_rdata_o_t0(rf_wdata_lsu_t0),
.lsu_rdata_valid_o(rf_we_lsu),
.lsu_rdata_valid_o_t0(rf_we_lsu_t0),
.lsu_req_done_o(lsu_req_done),
.lsu_req_done_o_t0(lsu_req_done_t0),
.lsu_req_i(lsu_req),
.lsu_req_i_t0(lsu_req_t0),
.lsu_resp_valid_o(lsu_resp_valid),
.lsu_resp_valid_o_t0(lsu_resp_valid_t0),
.lsu_sign_ext_i(lsu_sign_ext),
.lsu_sign_ext_i_t0(lsu_sign_ext_t0),
.lsu_type_i(lsu_type),
.lsu_type_i_t0(lsu_type_t0),
.lsu_wdata_i(lsu_wdata),
.lsu_wdata_i_t0(lsu_wdata_t0),
.lsu_we_i(lsu_we),
.lsu_we_i_t0(lsu_we_t0),
.perf_load_o(perf_load),
.perf_load_o_t0(perf_load_t0),
.perf_store_o(perf_store),
.perf_store_o_t0(perf_store_t0),
.rst_ni(rst_ni),
.store_err_o(lsu_store_err),
.store_err_o_t0(lsu_store_err_t0),
.store_resp_intg_err_o(lsu_store_resp_intg_err),
.store_resp_intg_err_o_t0(lsu_store_resp_intg_err_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13421.4-13452.3" */
\$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  wb_stage_i (
.clk_i(clk_i),
.dummy_instr_id_i(dummy_instr_id_o),
.dummy_instr_id_i_t0(dummy_instr_id_o_t0),
.dummy_instr_wb_o(dummy_instr_wb_o),
.dummy_instr_wb_o_t0(dummy_instr_wb_o_t0),
.en_wb_i(en_wb),
.en_wb_i_t0(en_wb_t0),
.instr_done_wb_o(instr_done_wb),
.instr_done_wb_o_t0(instr_done_wb_t0),
.instr_is_compressed_id_i(instr_is_compressed_id),
.instr_is_compressed_id_i_t0(instr_is_compressed_id_t0),
.instr_perf_count_id_i(instr_perf_count_id),
.instr_perf_count_id_i_t0(instr_perf_count_id_t0),
.instr_type_wb_i(instr_type_wb),
.instr_type_wb_i_t0(instr_type_wb_t0),
.lsu_resp_err_i(lsu_resp_err),
.lsu_resp_err_i_t0(lsu_resp_err_t0),
.lsu_resp_valid_i(lsu_resp_valid),
.lsu_resp_valid_i_t0(lsu_resp_valid_t0),
.outstanding_load_wb_o(outstanding_load_wb),
.outstanding_load_wb_o_t0(outstanding_load_wb_t0),
.outstanding_store_wb_o(outstanding_store_wb),
.outstanding_store_wb_o_t0(outstanding_store_wb_t0),
.pc_id_i(pc_id),
.pc_id_i_t0(pc_id_t0),
.pc_wb_o(pc_wb),
.pc_wb_o_t0(pc_wb_t0),
.perf_instr_ret_compressed_wb_o(perf_instr_ret_compressed_wb),
.perf_instr_ret_compressed_wb_o_t0(perf_instr_ret_compressed_wb_t0),
.perf_instr_ret_compressed_wb_spec_o(perf_instr_ret_compressed_wb_spec),
.perf_instr_ret_compressed_wb_spec_o_t0(perf_instr_ret_compressed_wb_spec_t0),
.perf_instr_ret_wb_o(perf_instr_ret_wb),
.perf_instr_ret_wb_o_t0(perf_instr_ret_wb_t0),
.perf_instr_ret_wb_spec_o(perf_instr_ret_wb_spec),
.perf_instr_ret_wb_spec_o_t0(perf_instr_ret_wb_spec_t0),
.ready_wb_o(ready_wb),
.ready_wb_o_t0(ready_wb_t0),
.rf_waddr_id_i(rf_waddr_id),
.rf_waddr_id_i_t0(rf_waddr_id_t0),
.rf_waddr_wb_o(rf_waddr_wb_o),
.rf_waddr_wb_o_t0(rf_waddr_wb_o_t0),
.rf_wdata_fwd_wb_o(rf_wdata_fwd_wb),
.rf_wdata_fwd_wb_o_t0(rf_wdata_fwd_wb_t0),
.rf_wdata_id_i(rf_wdata_id),
.rf_wdata_id_i_t0(rf_wdata_id_t0),
.rf_wdata_lsu_i(rf_wdata_lsu),
.rf_wdata_lsu_i_t0(rf_wdata_lsu_t0),
.rf_wdata_wb_o(rf_wdata_wb),
.rf_wdata_wb_o_t0(rf_wdata_wb_t0),
.rf_we_id_i(rf_we_id),
.rf_we_id_i_t0(rf_we_id_t0),
.rf_we_lsu_i(rf_we_lsu),
.rf_we_lsu_i_t0(rf_we_lsu_t0),
.rf_we_wb_o(rf_we_wb_o),
.rf_we_wb_o_t0(rf_we_wb_o_t0),
.rf_write_wb_o(rf_write_wb),
.rf_write_wb_o_t0(rf_write_wb_t0),
.rst_ni(rst_ni)
);
assign core_busy_o_t0 = 4'h0;
assign crash_dump_o = { pc_id, pc_if, lsu_addr_last, csr_mepc, crash_dump_mtval };
assign crash_dump_o_t0 = { pc_id_t0, pc_if_t0, lsu_addr_last_t0, csr_mepc_t0, crash_dump_mtval_t0 };
endmodule

module \$paramod$916c47de983e2a42946808797a4a11650abb788f\prim_onehot_check (clk_i, rst_ni, oh_i, addr_i, en_i, err_o, addr_i_t0, en_i_t0, err_o_t0, oh_i_t0);
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _000_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _001_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _002_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _003_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _004_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _005_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _006_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _007_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _008_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _009_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _010_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _011_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _012_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _013_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _014_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _015_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _016_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _017_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _018_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _019_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _020_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _021_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _022_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _023_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _024_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _025_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _026_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _027_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _028_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _029_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _030_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _031_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _032_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _033_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _034_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _035_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _036_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _037_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _038_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _039_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _040_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _041_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _042_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _043_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _044_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _045_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _046_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _047_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _048_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _049_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _050_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _051_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _052_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _053_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _054_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _055_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _056_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _057_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _058_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _059_;
/* src = "generated/sv2v_out.v:26549.29-26549.77" */
wire _060_;
/* src = "generated/sv2v_out.v:26549.83-26549.130" */
wire _061_;
/* src = "generated/sv2v_out.v:26550.30-26550.56" */
wire _062_;
/* src = "generated/sv2v_out.v:26550.30-26550.56" */
wire _063_;
/* src = "generated/sv2v_out.v:26550.30-26550.56" */
wire _064_;
/* src = "generated/sv2v_out.v:26550.30-26550.56" */
wire _065_;
/* src = "generated/sv2v_out.v:26550.30-26550.56" */
wire _066_;
/* src = "generated/sv2v_out.v:26550.30-26550.56" */
wire _067_;
/* src = "generated/sv2v_out.v:26550.30-26550.56" */
wire _068_;
/* src = "generated/sv2v_out.v:26550.30-26550.56" */
wire _069_;
/* src = "generated/sv2v_out.v:26550.30-26550.56" */
wire _070_;
/* src = "generated/sv2v_out.v:26550.30-26550.56" */
wire _071_;
/* src = "generated/sv2v_out.v:26550.30-26550.56" */
wire _072_;
/* src = "generated/sv2v_out.v:26550.30-26550.56" */
wire _073_;
/* src = "generated/sv2v_out.v:26550.30-26550.56" */
wire _074_;
/* src = "generated/sv2v_out.v:26550.30-26550.56" */
wire _075_;
/* src = "generated/sv2v_out.v:26550.30-26550.56" */
wire _076_;
/* src = "generated/sv2v_out.v:26549.29-26549.61" */
wire _077_;
/* src = "generated/sv2v_out.v:26549.29-26549.61" */
wire _078_;
/* src = "generated/sv2v_out.v:26549.29-26549.61" */
wire _079_;
/* src = "generated/sv2v_out.v:26549.29-26549.61" */
wire _080_;
/* src = "generated/sv2v_out.v:26549.29-26549.61" */
wire _081_;
/* src = "generated/sv2v_out.v:26550.29-26550.73" */
wire _082_;
/* src = "generated/sv2v_out.v:26550.29-26550.73" */
wire _083_;
/* src = "generated/sv2v_out.v:26550.29-26550.73" */
wire _084_;
/* src = "generated/sv2v_out.v:26550.29-26550.73" */
wire _085_;
/* src = "generated/sv2v_out.v:26550.29-26550.73" */
wire _086_;
/* src = "generated/sv2v_out.v:26550.29-26550.73" */
wire _087_;
/* src = "generated/sv2v_out.v:26550.29-26550.73" */
wire _088_;
/* src = "generated/sv2v_out.v:26550.29-26550.73" */
wire _089_;
/* src = "generated/sv2v_out.v:26550.29-26550.73" */
wire _090_;
/* src = "generated/sv2v_out.v:26550.29-26550.73" */
wire _091_;
/* src = "generated/sv2v_out.v:26550.29-26550.73" */
wire _092_;
/* src = "generated/sv2v_out.v:26550.29-26550.73" */
wire _093_;
/* src = "generated/sv2v_out.v:26550.29-26550.73" */
wire _094_;
/* src = "generated/sv2v_out.v:26550.29-26550.73" */
wire _095_;
/* src = "generated/sv2v_out.v:26550.29-26550.73" */
wire _096_;
/* src = "generated/sv2v_out.v:26558.18-26558.39" */
wire _097_;
/* src = "generated/sv2v_out.v:26556.7-26556.15" */
wire addr_err;
/* src = "generated/sv2v_out.v:26519.31-26519.37" */
input [4:0] addr_i;
wire [4:0] addr_i;
/* cellift = 32'd1 */
input [4:0] addr_i_t0;
wire [4:0] addr_i_t0;
/* src = "generated/sv2v_out.v:26524.38-26524.46" */
wire [62:0] and_tree;
/* src = "generated/sv2v_out.v:26516.8-26516.13" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:26520.13-26520.17" */
input en_i;
wire en_i;
/* cellift = 32'd1 */
input en_i_t0;
wire en_i_t0;
/* src = "generated/sv2v_out.v:26555.7-26555.17" */
wire enable_err;
/* src = "generated/sv2v_out.v:26521.14-26521.19" */
output err_o;
wire err_o;
/* cellift = 32'd1 */
output err_o_t0;
wire err_o_t0;
/* src = "generated/sv2v_out.v:26525.38-26525.46" */
wire [62:0] err_tree;
/* src = "generated/sv2v_out.v:26557.7-26557.14" */
wire oh0_err;
/* src = "generated/sv2v_out.v:26518.33-26518.37" */
input [31:0] oh_i;
wire [31:0] oh_i;
/* cellift = 32'd1 */
input [31:0] oh_i_t0;
wire [31:0] oh_i_t0;
/* src = "generated/sv2v_out.v:26523.38-26523.45" */
wire [62:0] or_tree;
/* src = "generated/sv2v_out.v:26517.8-26517.14" */
input rst_ni;
wire rst_ni;
assign _000_ = _077_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ and_tree[1];
assign _001_ = addr_i[4] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ and_tree[2];
assign _002_ = _078_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ and_tree[3];
assign _003_ = addr_i[3] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ and_tree[4];
assign _004_ = _078_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ and_tree[5];
assign _005_ = addr_i[3] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ and_tree[6];
assign _006_ = _079_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ and_tree[7];
assign _007_ = addr_i[2] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ and_tree[8];
assign _008_ = _079_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ and_tree[9];
assign _009_ = addr_i[2] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ and_tree[10];
assign _010_ = _079_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ and_tree[11];
assign _011_ = addr_i[2] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ and_tree[12];
assign _012_ = _079_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ and_tree[13];
assign _013_ = addr_i[2] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ and_tree[14];
assign _014_ = _080_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ and_tree[15];
assign _015_ = addr_i[1] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ and_tree[16];
assign _016_ = _080_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ and_tree[17];
assign _017_ = addr_i[1] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ and_tree[18];
assign _018_ = _080_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ and_tree[19];
assign _019_ = addr_i[1] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ and_tree[20];
assign _020_ = _080_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ and_tree[21];
assign _021_ = addr_i[1] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ and_tree[22];
assign _022_ = _080_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ and_tree[23];
assign _023_ = addr_i[1] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ and_tree[24];
assign _024_ = _080_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ and_tree[25];
assign _025_ = addr_i[1] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ and_tree[26];
assign _026_ = _080_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ and_tree[27];
assign _027_ = addr_i[1] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ and_tree[28];
assign _028_ = _080_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ and_tree[29];
assign _029_ = addr_i[1] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ and_tree[30];
assign _030_ = _081_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ oh_i[0];
assign _031_ = addr_i[0] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ oh_i[1];
assign _032_ = _081_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ oh_i[2];
assign _033_ = addr_i[0] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ oh_i[3];
assign _034_ = _081_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ oh_i[4];
assign _035_ = addr_i[0] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ oh_i[5];
assign _036_ = _081_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ oh_i[6];
assign _037_ = addr_i[0] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ oh_i[7];
assign _038_ = _081_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ oh_i[8];
assign _039_ = addr_i[0] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ oh_i[9];
assign _040_ = _081_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ oh_i[10];
assign _041_ = addr_i[0] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ oh_i[11];
assign _042_ = _081_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ oh_i[12];
assign _043_ = addr_i[0] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ oh_i[13];
assign _044_ = _081_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ oh_i[14];
assign _045_ = addr_i[0] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ oh_i[15];
assign _046_ = _081_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ oh_i[16];
assign _047_ = addr_i[0] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ oh_i[17];
assign _048_ = _081_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ oh_i[18];
assign _049_ = addr_i[0] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ oh_i[19];
assign _050_ = _081_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ oh_i[20];
assign _051_ = addr_i[0] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ oh_i[21];
assign _052_ = _081_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ oh_i[22];
assign _053_ = addr_i[0] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ oh_i[23];
assign _054_ = _081_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ oh_i[24];
assign _055_ = addr_i[0] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ oh_i[25];
assign _056_ = _081_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ oh_i[26];
assign _057_ = addr_i[0] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ oh_i[27];
assign _058_ = _081_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ oh_i[28];
assign _059_ = addr_i[0] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ oh_i[29];
assign _060_ = _081_ && /* src = "generated/sv2v_out.v:26549.29-26549.77" */ oh_i[30];
assign _061_ = addr_i[0] && /* src = "generated/sv2v_out.v:26549.83-26549.130" */ oh_i[31];
assign _062_ = or_tree[1] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ or_tree[2];
assign _063_ = or_tree[3] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ or_tree[4];
assign _064_ = or_tree[5] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ or_tree[6];
assign _065_ = or_tree[7] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ or_tree[8];
assign _066_ = or_tree[9] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ or_tree[10];
assign _067_ = or_tree[11] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ or_tree[12];
assign _068_ = or_tree[13] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ or_tree[14];
assign _069_ = or_tree[15] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ or_tree[16];
assign _070_ = or_tree[17] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ or_tree[18];
assign _071_ = or_tree[19] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ or_tree[20];
assign _072_ = or_tree[21] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ or_tree[22];
assign _073_ = or_tree[23] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ or_tree[24];
assign _074_ = or_tree[25] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ or_tree[26];
assign _075_ = or_tree[27] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ or_tree[28];
assign _076_ = or_tree[29] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ or_tree[30];
assign err_tree[15] = oh_i[0] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ oh_i[1];
assign err_tree[16] = oh_i[2] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ oh_i[3];
assign err_tree[17] = oh_i[4] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ oh_i[5];
assign err_tree[18] = oh_i[6] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ oh_i[7];
assign err_tree[19] = oh_i[8] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ oh_i[9];
assign err_tree[20] = oh_i[10] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ oh_i[11];
assign err_tree[21] = oh_i[12] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ oh_i[13];
assign err_tree[22] = oh_i[14] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ oh_i[15];
assign err_tree[23] = oh_i[16] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ oh_i[17];
assign err_tree[24] = oh_i[18] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ oh_i[19];
assign err_tree[25] = oh_i[20] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ oh_i[21];
assign err_tree[26] = oh_i[22] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ oh_i[23];
assign err_tree[27] = oh_i[24] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ oh_i[25];
assign err_tree[28] = oh_i[26] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ oh_i[27];
assign err_tree[29] = oh_i[28] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ oh_i[29];
assign err_tree[30] = oh_i[30] && /* src = "generated/sv2v_out.v:26550.30-26550.56" */ oh_i[31];
assign _077_ = ! /* src = "generated/sv2v_out.v:26549.29-26549.61" */ addr_i[4];
assign _078_ = ! /* src = "generated/sv2v_out.v:26549.29-26549.61" */ addr_i[3];
assign _079_ = ! /* src = "generated/sv2v_out.v:26549.29-26549.61" */ addr_i[2];
assign _080_ = ! /* src = "generated/sv2v_out.v:26549.29-26549.61" */ addr_i[1];
assign _081_ = ! /* src = "generated/sv2v_out.v:26549.29-26549.61" */ addr_i[0];
assign or_tree[0] = or_tree[1] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ or_tree[2];
assign or_tree[1] = or_tree[3] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ or_tree[4];
assign or_tree[2] = or_tree[5] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ or_tree[6];
assign or_tree[3] = or_tree[7] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ or_tree[8];
assign or_tree[4] = or_tree[9] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ or_tree[10];
assign or_tree[5] = or_tree[11] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ or_tree[12];
assign or_tree[6] = or_tree[13] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ or_tree[14];
assign or_tree[7] = or_tree[15] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ or_tree[16];
assign or_tree[8] = or_tree[17] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ or_tree[18];
assign or_tree[9] = or_tree[19] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ or_tree[20];
assign or_tree[10] = or_tree[21] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ or_tree[22];
assign or_tree[11] = or_tree[23] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ or_tree[24];
assign or_tree[12] = or_tree[25] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ or_tree[26];
assign or_tree[13] = or_tree[27] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ or_tree[28];
assign or_tree[14] = or_tree[29] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ or_tree[30];
assign or_tree[15] = oh_i[0] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ oh_i[1];
assign or_tree[16] = oh_i[2] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ oh_i[3];
assign or_tree[17] = oh_i[4] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ oh_i[5];
assign or_tree[18] = oh_i[6] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ oh_i[7];
assign or_tree[19] = oh_i[8] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ oh_i[9];
assign or_tree[20] = oh_i[10] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ oh_i[11];
assign or_tree[21] = oh_i[12] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ oh_i[13];
assign or_tree[22] = oh_i[14] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ oh_i[15];
assign or_tree[23] = oh_i[16] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ oh_i[17];
assign or_tree[24] = oh_i[18] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ oh_i[19];
assign or_tree[25] = oh_i[20] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ oh_i[21];
assign or_tree[26] = oh_i[22] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ oh_i[23];
assign or_tree[27] = oh_i[24] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ oh_i[25];
assign or_tree[28] = oh_i[26] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ oh_i[27];
assign or_tree[29] = oh_i[28] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ oh_i[29];
assign or_tree[30] = oh_i[30] || /* src = "generated/sv2v_out.v:26548.27-26548.53" */ oh_i[31];
assign and_tree[0] = _000_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _001_;
assign and_tree[1] = _002_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _003_;
assign and_tree[2] = _004_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _005_;
assign and_tree[3] = _006_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _007_;
assign and_tree[4] = _008_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _009_;
assign and_tree[5] = _010_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _011_;
assign and_tree[6] = _012_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _013_;
assign and_tree[7] = _014_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _015_;
assign and_tree[8] = _016_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _017_;
assign and_tree[9] = _018_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _019_;
assign and_tree[10] = _020_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _021_;
assign and_tree[11] = _022_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _023_;
assign and_tree[12] = _024_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _025_;
assign and_tree[13] = _026_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _027_;
assign and_tree[14] = _028_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _029_;
assign and_tree[15] = _030_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _031_;
assign and_tree[16] = _032_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _033_;
assign and_tree[17] = _034_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _035_;
assign and_tree[18] = _036_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _037_;
assign and_tree[19] = _038_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _039_;
assign and_tree[20] = _040_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _041_;
assign and_tree[21] = _042_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _043_;
assign and_tree[22] = _044_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _045_;
assign and_tree[23] = _046_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _047_;
assign and_tree[24] = _048_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _049_;
assign and_tree[25] = _050_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _051_;
assign and_tree[26] = _052_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _053_;
assign and_tree[27] = _054_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _055_;
assign and_tree[28] = _056_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _057_;
assign and_tree[29] = _058_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _059_;
assign and_tree[30] = _060_ || /* src = "generated/sv2v_out.v:26549.28-26549.131" */ _061_;
assign _082_ = _062_ || /* src = "generated/sv2v_out.v:26550.29-26550.73" */ err_tree[1];
assign oh0_err = _082_ || /* src = "generated/sv2v_out.v:26550.28-26550.90" */ err_tree[2];
assign _083_ = _063_ || /* src = "generated/sv2v_out.v:26550.29-26550.73" */ err_tree[3];
assign err_tree[1] = _083_ || /* src = "generated/sv2v_out.v:26550.28-26550.90" */ err_tree[4];
assign _084_ = _064_ || /* src = "generated/sv2v_out.v:26550.29-26550.73" */ err_tree[5];
assign err_tree[2] = _084_ || /* src = "generated/sv2v_out.v:26550.28-26550.90" */ err_tree[6];
assign _085_ = _065_ || /* src = "generated/sv2v_out.v:26550.29-26550.73" */ err_tree[7];
assign err_tree[3] = _085_ || /* src = "generated/sv2v_out.v:26550.28-26550.90" */ err_tree[8];
assign _086_ = _066_ || /* src = "generated/sv2v_out.v:26550.29-26550.73" */ err_tree[9];
assign err_tree[4] = _086_ || /* src = "generated/sv2v_out.v:26550.28-26550.90" */ err_tree[10];
assign _087_ = _067_ || /* src = "generated/sv2v_out.v:26550.29-26550.73" */ err_tree[11];
assign err_tree[5] = _087_ || /* src = "generated/sv2v_out.v:26550.28-26550.90" */ err_tree[12];
assign _088_ = _068_ || /* src = "generated/sv2v_out.v:26550.29-26550.73" */ err_tree[13];
assign err_tree[6] = _088_ || /* src = "generated/sv2v_out.v:26550.28-26550.90" */ err_tree[14];
assign _089_ = _069_ || /* src = "generated/sv2v_out.v:26550.29-26550.73" */ err_tree[15];
assign err_tree[7] = _089_ || /* src = "generated/sv2v_out.v:26550.28-26550.90" */ err_tree[16];
assign _090_ = _070_ || /* src = "generated/sv2v_out.v:26550.29-26550.73" */ err_tree[17];
assign err_tree[8] = _090_ || /* src = "generated/sv2v_out.v:26550.28-26550.90" */ err_tree[18];
assign _091_ = _071_ || /* src = "generated/sv2v_out.v:26550.29-26550.73" */ err_tree[19];
assign err_tree[9] = _091_ || /* src = "generated/sv2v_out.v:26550.28-26550.90" */ err_tree[20];
assign _092_ = _072_ || /* src = "generated/sv2v_out.v:26550.29-26550.73" */ err_tree[21];
assign err_tree[10] = _092_ || /* src = "generated/sv2v_out.v:26550.28-26550.90" */ err_tree[22];
assign _093_ = _073_ || /* src = "generated/sv2v_out.v:26550.29-26550.73" */ err_tree[23];
assign err_tree[11] = _093_ || /* src = "generated/sv2v_out.v:26550.28-26550.90" */ err_tree[24];
assign _094_ = _074_ || /* src = "generated/sv2v_out.v:26550.29-26550.73" */ err_tree[25];
assign err_tree[12] = _094_ || /* src = "generated/sv2v_out.v:26550.28-26550.90" */ err_tree[26];
assign _095_ = _075_ || /* src = "generated/sv2v_out.v:26550.29-26550.73" */ err_tree[27];
assign err_tree[13] = _095_ || /* src = "generated/sv2v_out.v:26550.28-26550.90" */ err_tree[28];
assign _096_ = _076_ || /* src = "generated/sv2v_out.v:26550.29-26550.73" */ err_tree[29];
assign err_tree[14] = _096_ || /* src = "generated/sv2v_out.v:26550.28-26550.90" */ err_tree[30];
assign _097_ = oh0_err || /* src = "generated/sv2v_out.v:26558.18-26558.39" */ enable_err;
assign err_o = _097_ || /* src = "generated/sv2v_out.v:26558.17-26558.52" */ addr_err;
assign enable_err = or_tree[0] ^ /* src = "generated/sv2v_out.v:26563.25-26563.42" */ en_i;
assign addr_err = or_tree[0] ^ /* src = "generated/sv2v_out.v:26575.22-26575.46" */ and_tree[0];
assign and_tree[62:31] = oh_i;
assign err_o_t0 = 1'h0;
assign { err_tree[62:31], err_tree[0] } = { 32'h00000000, oh0_err };
assign or_tree[62:31] = oh_i;
endmodule

module \$paramod$9a435d8f6db004a67362aa9a56f32ea481a74dbe\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _0_;
wire [31:0] _1_;
wire [31:0] _2_;
wire [31:0] _3_;
/* src = "generated/sv2v_out.v:14936.13-14936.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14940.28-14940.37" */
output [31:0] rd_data_o;
reg [31:0] rd_data_o;
/* cellift = 32'd1 */
output [31:0] rd_data_o_t0;
reg [31:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14941.14-14941.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14937.13-14937.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14938.27-14938.36" */
input [31:0] wr_data_i;
wire [31:0] wr_data_i;
/* cellift = 32'd1 */
input [31:0] wr_data_i_t0;
wire [31:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14939.13-14939.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _0_ = ~ wr_en_i;
assign _1_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _2_ = { _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_ } & rd_data_o_t0;
assign _3_ = _1_ | _2_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$9a435d8f6db004a67362aa9a56f32ea481a74dbe\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 32'd0;
else rd_data_o_t0 <= _3_;
/* src = "generated/sv2v_out.v:14943.2-14947.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$9a435d8f6db004a67362aa9a56f32ea481a74dbe\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 32'd1073741827;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$a088b13b9337f1e1fba58a671f47d7c7701ffa49\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _0_;
wire [7:0] _1_;
wire [7:0] _2_;
wire [7:0] _3_;
/* src = "generated/sv2v_out.v:14936.13-14936.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14940.28-14940.37" */
output [7:0] rd_data_o;
reg [7:0] rd_data_o;
/* cellift = 32'd1 */
output [7:0] rd_data_o_t0;
reg [7:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14941.14-14941.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14937.13-14937.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14938.27-14938.36" */
input [7:0] wr_data_i;
wire [7:0] wr_data_i;
/* cellift = 32'd1 */
input [7:0] wr_data_i_t0;
wire [7:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14939.13-14939.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _0_ = ~ wr_en_i;
assign _1_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _2_ = { _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_ } & rd_data_o_t0;
assign _3_ = _1_ | _2_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a088b13b9337f1e1fba58a671f47d7c7701ffa49\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 8'h00;
else rd_data_o_t0 <= _3_;
/* src = "generated/sv2v_out.v:14943.2-14947.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a088b13b9337f1e1fba58a671f47d7c7701ffa49\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 8'h00;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$a308247794889ee6093207090edbf289adef8be1\ibex_ex_block (clk_i, rst_ni, alu_operator_i, alu_operand_a_i, alu_operand_b_i, alu_instr_first_cycle_i, bt_a_operand_i, bt_b_operand_i, multdiv_operator_i, mult_en_i, div_en_i, mult_sel_i, div_sel_i, multdiv_signed_mode_i, multdiv_operand_a_i, multdiv_operand_b_i, multdiv_ready_id_i, data_ind_timing_i, imd_val_we_o, imd_val_d_o, imd_val_q_i
, alu_adder_result_ex_o, result_ex_o, branch_target_o, branch_decision_o, ex_valid_o, multdiv_operand_a_i_t0, multdiv_operand_b_i_t0, data_ind_timing_i_t0, div_en_i_t0, div_sel_i_t0, imd_val_d_o_t0, imd_val_q_i_t0, imd_val_we_o_t0, mult_en_i_t0, mult_sel_i_t0, multdiv_ready_id_i_t0, alu_adder_result_ex_o_t0, alu_instr_first_cycle_i_t0, alu_operand_a_i_t0, alu_operand_b_i_t0, alu_operator_i_t0
, branch_decision_o_t0, branch_target_o_t0, bt_a_operand_i_t0, bt_b_operand_i_t0, ex_valid_o_t0, multdiv_operator_i_t0, multdiv_signed_mode_i_t0, result_ex_o_t0);
wire [33:0] _00_;
wire [1:0] _01_;
wire [31:0] _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire [33:0] _08_;
wire [33:0] _09_;
wire [33:0] _10_;
wire [33:0] _11_;
wire [1:0] _12_;
wire [1:0] _13_;
wire [31:0] _14_;
wire [31:0] _15_;
wire _16_;
/* src = "generated/sv2v_out.v:16122.53-16122.71" */
wire _17_;
/* src = "generated/sv2v_out.v:16122.55-16122.70" */
wire _18_;
/* src = "generated/sv2v_out.v:16002.21-16002.42" */
output [31:0] alu_adder_result_ex_o;
wire [31:0] alu_adder_result_ex_o;
/* cellift = 32'd1 */
output [31:0] alu_adder_result_ex_o_t0;
wire [31:0] alu_adder_result_ex_o_t0;
/* src = "generated/sv2v_out.v:16011.14-16011.34" */
wire [33:0] alu_adder_result_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16011.14-16011.34" */
wire [33:0] alu_adder_result_ext_t0;
/* src = "generated/sv2v_out.v:16017.14-16017.27" */
wire [63:0] alu_imd_val_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16017.14-16017.27" */
wire [63:0] alu_imd_val_d_t0;
/* src = "generated/sv2v_out.v:16018.13-16018.27" */
wire [1:0] alu_imd_val_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16018.13-16018.27" */
wire [1:0] alu_imd_val_we_t0;
/* src = "generated/sv2v_out.v:15986.13-15986.36" */
input alu_instr_first_cycle_i;
wire alu_instr_first_cycle_i;
/* cellift = 32'd1 */
input alu_instr_first_cycle_i_t0;
wire alu_instr_first_cycle_i_t0;
/* src = "generated/sv2v_out.v:16013.7-16013.26" */
wire alu_is_equal_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16013.7-16013.26" */
wire alu_is_equal_result_t0;
/* src = "generated/sv2v_out.v:15984.20-15984.35" */
input [31:0] alu_operand_a_i;
wire [31:0] alu_operand_a_i;
/* cellift = 32'd1 */
input [31:0] alu_operand_a_i_t0;
wire [31:0] alu_operand_a_i_t0;
/* src = "generated/sv2v_out.v:15985.20-15985.35" */
input [31:0] alu_operand_b_i;
wire [31:0] alu_operand_b_i;
/* cellift = 32'd1 */
input [31:0] alu_operand_b_i_t0;
wire [31:0] alu_operand_b_i_t0;
/* src = "generated/sv2v_out.v:15983.19-15983.33" */
input [6:0] alu_operator_i;
wire [6:0] alu_operator_i;
/* cellift = 32'd1 */
input [6:0] alu_operator_i_t0;
wire [6:0] alu_operator_i_t0;
/* src = "generated/sv2v_out.v:16007.14-16007.24" */
wire [31:0] alu_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16007.14-16007.24" */
wire [31:0] alu_result_t0;
/* src = "generated/sv2v_out.v:16005.14-16005.31" */
output branch_decision_o;
wire branch_decision_o;
/* cellift = 32'd1 */
output branch_decision_o_t0;
wire branch_decision_o_t0;
/* src = "generated/sv2v_out.v:16004.21-16004.36" */
output [31:0] branch_target_o;
wire [31:0] branch_target_o;
/* cellift = 32'd1 */
output [31:0] branch_target_o_t0;
wire [31:0] branch_target_o_t0;
/* src = "generated/sv2v_out.v:15987.20-15987.34" */
input [31:0] bt_a_operand_i;
wire [31:0] bt_a_operand_i;
/* cellift = 32'd1 */
input [31:0] bt_a_operand_i_t0;
wire [31:0] bt_a_operand_i_t0;
/* src = "generated/sv2v_out.v:15988.20-15988.34" */
input [31:0] bt_b_operand_i;
wire [31:0] bt_b_operand_i;
/* cellift = 32'd1 */
input [31:0] bt_b_operand_i_t0;
wire [31:0] bt_b_operand_i_t0;
/* src = "generated/sv2v_out.v:15981.13-15981.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:15998.13-15998.30" */
input data_ind_timing_i;
wire data_ind_timing_i;
/* cellift = 32'd1 */
input data_ind_timing_i_t0;
wire data_ind_timing_i_t0;
/* src = "generated/sv2v_out.v:15991.13-15991.21" */
input div_en_i;
wire div_en_i;
/* cellift = 32'd1 */
input div_en_i_t0;
wire div_en_i_t0;
/* src = "generated/sv2v_out.v:15993.13-15993.22" */
input div_sel_i;
wire div_sel_i;
/* cellift = 32'd1 */
input div_sel_i_t0;
wire div_sel_i_t0;
/* src = "generated/sv2v_out.v:16006.14-16006.24" */
output ex_valid_o;
wire ex_valid_o;
/* cellift = 32'd1 */
output ex_valid_o_t0;
wire ex_valid_o_t0;
/* src = "generated/sv2v_out.v:16000.21-16000.32" */
output [67:0] imd_val_d_o;
wire [67:0] imd_val_d_o;
/* cellift = 32'd1 */
output [67:0] imd_val_d_o_t0;
wire [67:0] imd_val_d_o_t0;
/* src = "generated/sv2v_out.v:16001.20-16001.31" */
input [67:0] imd_val_q_i;
wire [67:0] imd_val_q_i;
/* cellift = 32'd1 */
input [67:0] imd_val_q_i_t0;
wire [67:0] imd_val_q_i_t0;
/* src = "generated/sv2v_out.v:15999.20-15999.32" */
output [1:0] imd_val_we_o;
wire [1:0] imd_val_we_o;
/* cellift = 32'd1 */
output [1:0] imd_val_we_o_t0;
wire [1:0] imd_val_we_o_t0;
/* src = "generated/sv2v_out.v:15990.13-15990.22" */
input mult_en_i;
wire mult_en_i;
/* cellift = 32'd1 */
input mult_en_i_t0;
wire mult_en_i_t0;
/* src = "generated/sv2v_out.v:15992.13-15992.23" */
input mult_sel_i;
wire mult_sel_i;
/* cellift = 32'd1 */
input mult_sel_i_t0;
wire mult_sel_i_t0;
/* src = "generated/sv2v_out.v:16010.14-16010.35" */
wire [32:0] multdiv_alu_operand_a;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16010.14-16010.35" */
wire [32:0] multdiv_alu_operand_a_t0;
/* src = "generated/sv2v_out.v:16009.14-16009.35" */
wire [32:0] multdiv_alu_operand_b;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16009.14-16009.35" */
wire [32:0] multdiv_alu_operand_b_t0;
/* src = "generated/sv2v_out.v:16019.14-16019.31" */
wire [67:0] multdiv_imd_val_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16019.14-16019.31" */
wire [67:0] multdiv_imd_val_d_t0;
/* src = "generated/sv2v_out.v:16020.13-16020.31" */
wire [1:0] multdiv_imd_val_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16020.13-16020.31" */
wire [1:0] multdiv_imd_val_we_t0;
/* src = "generated/sv2v_out.v:15995.20-15995.39" */
input [31:0] multdiv_operand_a_i;
wire [31:0] multdiv_operand_a_i;
/* cellift = 32'd1 */
input [31:0] multdiv_operand_a_i_t0;
wire [31:0] multdiv_operand_a_i_t0;
/* src = "generated/sv2v_out.v:15996.20-15996.39" */
input [31:0] multdiv_operand_b_i;
wire [31:0] multdiv_operand_b_i;
/* cellift = 32'd1 */
input [31:0] multdiv_operand_b_i_t0;
wire [31:0] multdiv_operand_b_i_t0;
/* src = "generated/sv2v_out.v:15989.19-15989.37" */
input [1:0] multdiv_operator_i;
wire [1:0] multdiv_operator_i;
/* cellift = 32'd1 */
input [1:0] multdiv_operator_i_t0;
wire [1:0] multdiv_operator_i_t0;
/* src = "generated/sv2v_out.v:15997.13-15997.31" */
input multdiv_ready_id_i;
wire multdiv_ready_id_i;
/* cellift = 32'd1 */
input multdiv_ready_id_i_t0;
wire multdiv_ready_id_i_t0;
/* src = "generated/sv2v_out.v:16008.14-16008.28" */
wire [31:0] multdiv_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16008.14-16008.28" */
wire [31:0] multdiv_result_t0;
/* src = "generated/sv2v_out.v:16015.7-16015.18" */
wire multdiv_sel;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16015.7-16015.18" */
wire multdiv_sel_t0;
/* src = "generated/sv2v_out.v:15994.19-15994.40" */
input [1:0] multdiv_signed_mode_i;
wire [1:0] multdiv_signed_mode_i;
/* cellift = 32'd1 */
input [1:0] multdiv_signed_mode_i_t0;
wire [1:0] multdiv_signed_mode_i_t0;
/* src = "generated/sv2v_out.v:16014.7-16014.20" */
wire multdiv_valid;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16014.7-16014.20" */
wire multdiv_valid_t0;
/* src = "generated/sv2v_out.v:16003.21-16003.32" */
output [31:0] result_ex_o;
wire [31:0] result_ex_o;
/* cellift = 32'd1 */
output [31:0] result_ex_o_t0;
wire [31:0] result_ex_o_t0;
/* src = "generated/sv2v_out.v:15982.13-15982.19" */
input rst_ni;
wire rst_ni;
assign _00_ = ~ { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel };
assign _01_ = ~ { multdiv_sel, multdiv_sel };
assign _02_ = ~ { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel };
assign _08_ = _00_ & { 2'h0, alu_imd_val_d_t0[63:32] };
assign _10_ = _00_ & { 2'h0, alu_imd_val_d_t0[31:0] };
assign _12_ = _01_ & alu_imd_val_we_t0;
assign _14_ = _02_ & alu_result_t0;
assign _09_ = { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel } & multdiv_imd_val_d_t0[67:34];
assign _11_ = { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel } & multdiv_imd_val_d_t0[33:0];
assign _13_ = { multdiv_sel, multdiv_sel } & multdiv_imd_val_we_t0;
assign _15_ = { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel } & multdiv_result_t0;
assign ex_valid_o_t0 = multdiv_sel & multdiv_valid_t0;
assign imd_val_d_o_t0[67:34] = _08_ | _09_;
assign imd_val_d_o_t0[33:0] = _10_ | _11_;
assign imd_val_we_o_t0 = _12_ | _13_;
assign result_ex_o_t0 = _14_ | _15_;
assign _03_ = ~ mult_sel_i;
assign _04_ = ~ div_sel_i;
assign _05_ = mult_sel_i_t0 & _04_;
assign _06_ = div_sel_i_t0 & _03_;
assign _07_ = mult_sel_i_t0 & div_sel_i_t0;
assign _16_ = _05_ | _06_;
assign multdiv_sel_t0 = _16_ | _07_;
assign _17_ = ~ /* src = "generated/sv2v_out.v:16122.53-16122.71" */ _18_;
assign multdiv_sel = mult_sel_i | /* src = "generated/sv2v_out.v:16023.25-16023.47" */ div_sel_i;
assign _18_ = | /* src = "generated/sv2v_out.v:16122.55-16122.70" */ alu_imd_val_we;
assign imd_val_d_o[67:34] = multdiv_sel ? /* src = "generated/sv2v_out.v:16029.32-16029.104" */ multdiv_imd_val_d[67:34] : { 2'h0, alu_imd_val_d[63:32] };
assign imd_val_d_o[33:0] = multdiv_sel ? /* src = "generated/sv2v_out.v:16030.31-16030.101" */ multdiv_imd_val_d[33:0] : { 2'h0, alu_imd_val_d[31:0] };
assign imd_val_we_o = multdiv_sel ? /* src = "generated/sv2v_out.v:16031.25-16031.74" */ multdiv_imd_val_we : alu_imd_val_we;
assign result_ex_o = multdiv_sel ? /* src = "generated/sv2v_out.v:16033.24-16033.65" */ multdiv_result : alu_result;
assign ex_valid_o = multdiv_sel ? /* src = "generated/sv2v_out.v:16122.23-16122.71" */ multdiv_valid : _17_;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:16051.28-16067.3" */
\$paramod\ibex_alu\RV32B=s32'00000000000000000000000000000000  alu_i (
.adder_result_ext_o(alu_adder_result_ext),
.adder_result_ext_o_t0(alu_adder_result_ext_t0),
.adder_result_o(alu_adder_result_ex_o),
.adder_result_o_t0(alu_adder_result_ex_o_t0),
.comparison_result_o(branch_decision_o),
.comparison_result_o_t0(branch_decision_o_t0),
.imd_val_d_o(alu_imd_val_d),
.imd_val_d_o_t0(alu_imd_val_d_t0),
.imd_val_q_i({ imd_val_q_i[65:34], imd_val_q_i[31:0] }),
.imd_val_q_i_t0({ imd_val_q_i_t0[65:34], imd_val_q_i_t0[31:0] }),
.imd_val_we_o(alu_imd_val_we),
.imd_val_we_o_t0(alu_imd_val_we_t0),
.instr_first_cycle_i(alu_instr_first_cycle_i),
.instr_first_cycle_i_t0(alu_instr_first_cycle_i_t0),
.is_equal_result_o(alu_is_equal_result),
.is_equal_result_o_t0(alu_is_equal_result_t0),
.multdiv_operand_a_i(multdiv_alu_operand_a),
.multdiv_operand_a_i_t0(multdiv_alu_operand_a_t0),
.multdiv_operand_b_i(multdiv_alu_operand_b),
.multdiv_operand_b_i_t0(multdiv_alu_operand_b_t0),
.multdiv_sel_i(multdiv_sel),
.multdiv_sel_i_t0(multdiv_sel_t0),
.operand_a_i(alu_operand_a_i),
.operand_a_i_t0(alu_operand_a_i_t0),
.operand_b_i(alu_operand_b_i),
.operand_b_i_t0(alu_operand_b_i_t0),
.operator_i(alu_operator_i),
.operator_i_t0(alu_operator_i_t0),
.result_o(alu_result),
.result_o_t0(alu_result_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:16070.22-16093.5" */
ibex_multdiv_slow \gen_multdiv_slow.multdiv_i  (
.alu_adder_ext_i(alu_adder_result_ext),
.alu_adder_ext_i_t0(alu_adder_result_ext_t0),
.alu_adder_i(alu_adder_result_ex_o),
.alu_adder_i_t0(alu_adder_result_ex_o_t0),
.alu_operand_a_o(multdiv_alu_operand_a),
.alu_operand_a_o_t0(multdiv_alu_operand_a_t0),
.alu_operand_b_o(multdiv_alu_operand_b),
.alu_operand_b_o_t0(multdiv_alu_operand_b_t0),
.clk_i(clk_i),
.data_ind_timing_i(data_ind_timing_i),
.data_ind_timing_i_t0(data_ind_timing_i_t0),
.div_en_i(div_en_i),
.div_en_i_t0(div_en_i_t0),
.div_sel_i(div_sel_i),
.div_sel_i_t0(div_sel_i_t0),
.equal_to_zero_i(alu_is_equal_result),
.equal_to_zero_i_t0(alu_is_equal_result_t0),
.imd_val_d_o(multdiv_imd_val_d),
.imd_val_d_o_t0(multdiv_imd_val_d_t0),
.imd_val_q_i(imd_val_q_i),
.imd_val_q_i_t0(imd_val_q_i_t0),
.imd_val_we_o(multdiv_imd_val_we),
.imd_val_we_o_t0(multdiv_imd_val_we_t0),
.mult_en_i(mult_en_i),
.mult_en_i_t0(mult_en_i_t0),
.mult_sel_i(mult_sel_i),
.mult_sel_i_t0(mult_sel_i_t0),
.multdiv_ready_id_i(multdiv_ready_id_i),
.multdiv_ready_id_i_t0(multdiv_ready_id_i_t0),
.multdiv_result_o(multdiv_result),
.multdiv_result_o_t0(multdiv_result_t0),
.op_a_i(multdiv_operand_a_i),
.op_a_i_t0(multdiv_operand_a_i_t0),
.op_b_i(multdiv_operand_b_i),
.op_b_i_t0(multdiv_operand_b_i_t0),
.operator_i(multdiv_operator_i),
.operator_i_t0(multdiv_operator_i_t0),
.rst_ni(rst_ni),
.signed_mode_i(multdiv_signed_mode_i),
.signed_mode_i_t0(multdiv_signed_mode_i_t0),
.valid_o(multdiv_valid),
.valid_o_t0(multdiv_valid_t0)
);
assign branch_target_o = alu_adder_result_ex_o;
assign branch_target_o_t0 = alu_adder_result_ex_o_t0;
endmodule

module \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff (clk_i, rst_ni, test_en_i, dummy_instr_id_i, dummy_instr_wb_i, raddr_a_i, rdata_a_o, raddr_b_i, rdata_b_o, waddr_a_i, wdata_a_i, we_a_i, err_o, test_en_i_t0, err_o_t0, dummy_instr_id_i_t0, dummy_instr_wb_i_t0, raddr_a_i_t0, raddr_b_i_t0, rdata_a_o_t0, rdata_b_o_t0
, waddr_a_i_t0, wdata_a_i_t0, we_a_i_t0);
wire _0000_;
wire _0001_;
wire _0002_;
wire _0003_;
wire _0004_;
wire _0005_;
wire _0006_;
wire _0007_;
wire _0008_;
wire _0009_;
wire _0010_;
wire _0011_;
wire _0012_;
wire _0013_;
wire _0014_;
wire _0015_;
wire _0016_;
wire _0017_;
wire _0018_;
wire _0019_;
wire _0020_;
wire _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire _0026_;
wire _0027_;
wire _0028_;
wire _0029_;
wire _0030_;
wire _0031_;
wire [38:0] _0032_;
wire [38:0] _0033_;
wire [38:0] _0034_;
wire [38:0] _0035_;
wire [38:0] _0036_;
wire [38:0] _0037_;
wire [38:0] _0038_;
wire [38:0] _0039_;
wire [38:0] _0040_;
wire [38:0] _0041_;
wire [38:0] _0042_;
wire [38:0] _0043_;
wire [38:0] _0044_;
wire [38:0] _0045_;
wire [38:0] _0046_;
wire [38:0] _0047_;
wire [38:0] _0048_;
wire [38:0] _0049_;
wire [38:0] _0050_;
wire [38:0] _0051_;
wire [38:0] _0052_;
wire [38:0] _0053_;
wire [38:0] _0054_;
wire [38:0] _0055_;
wire [38:0] _0056_;
wire [38:0] _0057_;
wire [38:0] _0058_;
wire [38:0] _0059_;
wire [38:0] _0060_;
wire [38:0] _0061_;
wire [38:0] _0062_;
wire [38:0] _0063_;
wire [38:0] _0064_;
wire [38:0] _0065_;
wire [38:0] _0066_;
wire [38:0] _0067_;
wire [38:0] _0068_;
wire [38:0] _0069_;
wire [38:0] _0070_;
wire [38:0] _0071_;
wire [38:0] _0072_;
wire [38:0] _0073_;
wire [38:0] _0074_;
wire [38:0] _0075_;
wire [38:0] _0076_;
wire [38:0] _0077_;
wire [38:0] _0078_;
wire [38:0] _0079_;
wire [38:0] _0080_;
wire [38:0] _0081_;
wire [38:0] _0082_;
wire [38:0] _0083_;
wire [38:0] _0084_;
wire [38:0] _0085_;
wire [38:0] _0086_;
wire [38:0] _0087_;
wire [38:0] _0088_;
wire [38:0] _0089_;
wire [38:0] _0090_;
wire [38:0] _0091_;
wire [38:0] _0092_;
wire [38:0] _0093_;
wire _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire [38:0] _0108_;
wire [38:0] _0109_;
wire [38:0] _0110_;
wire [38:0] _0111_;
wire [38:0] _0112_;
wire [38:0] _0113_;
wire [38:0] _0114_;
wire [38:0] _0115_;
wire [38:0] _0116_;
wire [38:0] _0117_;
wire [38:0] _0118_;
wire [38:0] _0119_;
wire [38:0] _0120_;
wire [38:0] _0121_;
wire [38:0] _0122_;
wire [38:0] _0123_;
wire [38:0] _0124_;
wire [38:0] _0125_;
wire [38:0] _0126_;
wire [38:0] _0127_;
wire [38:0] _0128_;
wire [38:0] _0129_;
wire [38:0] _0130_;
wire [38:0] _0131_;
wire [38:0] _0132_;
wire [38:0] _0133_;
wire [38:0] _0134_;
wire [38:0] _0135_;
wire [38:0] _0136_;
wire [38:0] _0137_;
wire [38:0] _0138_;
wire [38:0] _0139_;
wire [38:0] _0140_;
wire [38:0] _0141_;
wire [38:0] _0142_;
wire [38:0] _0143_;
wire [38:0] _0144_;
wire [38:0] _0145_;
wire [38:0] _0146_;
wire [38:0] _0147_;
wire [38:0] _0148_;
wire [38:0] _0149_;
wire [38:0] _0150_;
wire [38:0] _0151_;
wire [38:0] _0152_;
wire [38:0] _0153_;
wire [38:0] _0154_;
wire [38:0] _0155_;
wire [38:0] _0156_;
wire [38:0] _0157_;
wire [38:0] _0158_;
wire [38:0] _0159_;
wire [38:0] _0160_;
wire [38:0] _0161_;
wire [38:0] _0162_;
wire [38:0] _0163_;
wire [38:0] _0164_;
wire [38:0] _0165_;
wire [38:0] _0166_;
wire [38:0] _0167_;
wire [38:0] _0168_;
wire [38:0] _0169_;
wire [38:0] _0170_;
wire [38:0] _0171_;
wire [38:0] _0172_;
wire [38:0] _0173_;
wire [38:0] _0174_;
wire [38:0] _0175_;
wire [38:0] _0176_;
wire [38:0] _0177_;
wire [38:0] _0178_;
wire [38:0] _0179_;
wire [38:0] _0180_;
wire [38:0] _0181_;
wire [38:0] _0182_;
wire [38:0] _0183_;
wire [38:0] _0184_;
wire [38:0] _0185_;
wire [38:0] _0186_;
wire [38:0] _0187_;
wire [38:0] _0188_;
wire [38:0] _0189_;
wire [38:0] _0190_;
wire [38:0] _0191_;
wire [38:0] _0192_;
wire [38:0] _0193_;
wire [38:0] _0194_;
wire [38:0] _0195_;
wire [38:0] _0196_;
wire [38:0] _0197_;
wire [38:0] _0198_;
wire [38:0] _0199_;
wire [38:0] _0200_;
wire [38:0] _0201_;
wire [38:0] _0202_;
wire [38:0] _0203_;
wire [38:0] _0204_;
wire [38:0] _0205_;
wire [38:0] _0206_;
wire [38:0] _0207_;
wire [38:0] _0208_;
wire [38:0] _0209_;
wire [38:0] _0210_;
wire [38:0] _0211_;
wire [38:0] _0212_;
wire [38:0] _0213_;
wire [38:0] _0214_;
wire [38:0] _0215_;
wire [38:0] _0216_;
wire [38:0] _0217_;
wire [38:0] _0218_;
wire [38:0] _0219_;
wire [38:0] _0220_;
wire [38:0] _0221_;
wire [38:0] _0222_;
wire [38:0] _0223_;
wire [38:0] _0224_;
wire [38:0] _0225_;
wire [38:0] _0226_;
wire [38:0] _0227_;
wire [38:0] _0228_;
wire [38:0] _0229_;
wire [38:0] _0230_;
wire [38:0] _0231_;
wire [38:0] _0232_;
wire [38:0] _0233_;
wire [38:0] _0234_;
wire [38:0] _0235_;
wire [38:0] _0236_;
wire [38:0] _0237_;
wire [38:0] _0238_;
wire [38:0] _0239_;
wire [38:0] _0240_;
wire [38:0] _0241_;
wire [38:0] _0242_;
wire [38:0] _0243_;
wire [38:0] _0244_;
wire [38:0] _0245_;
wire [38:0] _0246_;
wire [38:0] _0247_;
wire [38:0] _0248_;
wire [38:0] _0249_;
wire [38:0] _0250_;
wire [38:0] _0251_;
wire [38:0] _0252_;
wire [38:0] _0253_;
wire [38:0] _0254_;
wire [38:0] _0255_;
wire [38:0] _0256_;
wire [38:0] _0257_;
wire [38:0] _0258_;
wire [38:0] _0259_;
wire [38:0] _0260_;
wire [38:0] _0261_;
wire [38:0] _0262_;
wire [38:0] _0263_;
wire [38:0] _0264_;
wire [38:0] _0265_;
wire [38:0] _0266_;
wire [38:0] _0267_;
wire [38:0] _0268_;
wire [38:0] _0269_;
wire [38:0] _0270_;
wire [38:0] _0271_;
wire [38:0] _0272_;
wire [38:0] _0273_;
wire [38:0] _0274_;
wire [38:0] _0275_;
wire [38:0] _0276_;
wire [38:0] _0277_;
wire [38:0] _0278_;
wire [38:0] _0279_;
wire [38:0] _0280_;
wire [38:0] _0281_;
wire [38:0] _0282_;
wire [38:0] _0283_;
wire [38:0] _0284_;
wire [38:0] _0285_;
wire [38:0] _0286_;
wire [38:0] _0287_;
wire [38:0] _0288_;
wire [38:0] _0289_;
wire [38:0] _0290_;
wire [38:0] _0291_;
wire [38:0] _0292_;
wire [38:0] _0293_;
wire [38:0] _0294_;
wire [38:0] _0295_;
wire _0296_;
wire _0297_;
wire _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire [38:0] _0310_;
wire [38:0] _0311_;
wire [38:0] _0312_;
wire [38:0] _0313_;
wire [38:0] _0314_;
wire [38:0] _0315_;
wire [38:0] _0316_;
wire [38:0] _0317_;
wire [38:0] _0318_;
wire [38:0] _0319_;
wire [38:0] _0320_;
wire [38:0] _0321_;
wire [38:0] _0322_;
wire [38:0] _0323_;
wire [38:0] _0324_;
wire [38:0] _0325_;
wire [38:0] _0326_;
wire [38:0] _0327_;
wire [38:0] _0328_;
wire [38:0] _0329_;
wire [38:0] _0330_;
wire [38:0] _0331_;
wire [38:0] _0332_;
wire [38:0] _0333_;
wire [38:0] _0334_;
wire [38:0] _0335_;
wire [38:0] _0336_;
wire [38:0] _0337_;
wire [38:0] _0338_;
wire [38:0] _0339_;
wire [38:0] _0340_;
wire [38:0] _0341_;
wire _0342_;
wire _0343_;
wire [38:0] _0344_;
/* cellift = 32'd1 */
wire [38:0] _0345_;
wire [38:0] _0346_;
/* cellift = 32'd1 */
wire [38:0] _0347_;
wire [38:0] _0348_;
/* cellift = 32'd1 */
wire [38:0] _0349_;
wire [38:0] _0350_;
/* cellift = 32'd1 */
wire [38:0] _0351_;
wire [38:0] _0352_;
/* cellift = 32'd1 */
wire [38:0] _0353_;
wire [38:0] _0354_;
/* cellift = 32'd1 */
wire [38:0] _0355_;
wire [38:0] _0356_;
/* cellift = 32'd1 */
wire [38:0] _0357_;
wire [38:0] _0358_;
/* cellift = 32'd1 */
wire [38:0] _0359_;
wire [38:0] _0360_;
/* cellift = 32'd1 */
wire [38:0] _0361_;
wire [38:0] _0362_;
/* cellift = 32'd1 */
wire [38:0] _0363_;
wire [38:0] _0364_;
/* cellift = 32'd1 */
wire [38:0] _0365_;
wire [38:0] _0366_;
/* cellift = 32'd1 */
wire [38:0] _0367_;
wire [38:0] _0368_;
/* cellift = 32'd1 */
wire [38:0] _0369_;
wire [38:0] _0370_;
/* cellift = 32'd1 */
wire [38:0] _0371_;
wire [38:0] _0372_;
/* cellift = 32'd1 */
wire [38:0] _0373_;
wire [38:0] _0374_;
/* cellift = 32'd1 */
wire [38:0] _0375_;
wire [38:0] _0376_;
/* cellift = 32'd1 */
wire [38:0] _0377_;
wire [38:0] _0378_;
/* cellift = 32'd1 */
wire [38:0] _0379_;
wire [38:0] _0380_;
/* cellift = 32'd1 */
wire [38:0] _0381_;
wire [38:0] _0382_;
/* cellift = 32'd1 */
wire [38:0] _0383_;
wire [38:0] _0384_;
/* cellift = 32'd1 */
wire [38:0] _0385_;
wire [38:0] _0386_;
/* cellift = 32'd1 */
wire [38:0] _0387_;
wire [38:0] _0388_;
/* cellift = 32'd1 */
wire [38:0] _0389_;
wire [38:0] _0390_;
/* cellift = 32'd1 */
wire [38:0] _0391_;
wire [38:0] _0392_;
/* cellift = 32'd1 */
wire [38:0] _0393_;
wire [38:0] _0394_;
/* cellift = 32'd1 */
wire [38:0] _0395_;
wire [38:0] _0396_;
/* cellift = 32'd1 */
wire [38:0] _0397_;
wire [38:0] _0398_;
/* cellift = 32'd1 */
wire [38:0] _0399_;
wire [38:0] _0400_;
/* cellift = 32'd1 */
wire [38:0] _0401_;
wire [38:0] _0402_;
/* cellift = 32'd1 */
wire [38:0] _0403_;
wire [38:0] _0404_;
/* cellift = 32'd1 */
wire [38:0] _0405_;
wire [38:0] _0406_;
/* cellift = 32'd1 */
wire [38:0] _0407_;
wire [38:0] _0408_;
/* cellift = 32'd1 */
wire [38:0] _0409_;
wire [38:0] _0410_;
/* cellift = 32'd1 */
wire [38:0] _0411_;
wire [38:0] _0412_;
/* cellift = 32'd1 */
wire [38:0] _0413_;
wire [38:0] _0414_;
/* cellift = 32'd1 */
wire [38:0] _0415_;
wire [38:0] _0416_;
/* cellift = 32'd1 */
wire [38:0] _0417_;
wire [38:0] _0418_;
/* cellift = 32'd1 */
wire [38:0] _0419_;
wire [38:0] _0420_;
/* cellift = 32'd1 */
wire [38:0] _0421_;
wire [38:0] _0422_;
/* cellift = 32'd1 */
wire [38:0] _0423_;
wire [38:0] _0424_;
/* cellift = 32'd1 */
wire [38:0] _0425_;
wire [38:0] _0426_;
/* cellift = 32'd1 */
wire [38:0] _0427_;
wire [38:0] _0428_;
/* cellift = 32'd1 */
wire [38:0] _0429_;
wire [38:0] _0430_;
/* cellift = 32'd1 */
wire [38:0] _0431_;
wire [38:0] _0432_;
/* cellift = 32'd1 */
wire [38:0] _0433_;
wire [38:0] _0434_;
/* cellift = 32'd1 */
wire [38:0] _0435_;
wire [38:0] _0436_;
/* cellift = 32'd1 */
wire [38:0] _0437_;
wire [38:0] _0438_;
/* cellift = 32'd1 */
wire [38:0] _0439_;
wire [38:0] _0440_;
/* cellift = 32'd1 */
wire [38:0] _0441_;
wire [38:0] _0442_;
/* cellift = 32'd1 */
wire [38:0] _0443_;
wire [38:0] _0444_;
/* cellift = 32'd1 */
wire [38:0] _0445_;
wire [38:0] _0446_;
/* cellift = 32'd1 */
wire [38:0] _0447_;
wire [38:0] _0448_;
/* cellift = 32'd1 */
wire [38:0] _0449_;
wire [38:0] _0450_;
/* cellift = 32'd1 */
wire [38:0] _0451_;
wire [38:0] _0452_;
/* cellift = 32'd1 */
wire [38:0] _0453_;
wire [38:0] _0454_;
/* cellift = 32'd1 */
wire [38:0] _0455_;
wire [38:0] _0456_;
/* cellift = 32'd1 */
wire [38:0] _0457_;
wire [38:0] _0458_;
/* cellift = 32'd1 */
wire [38:0] _0459_;
wire [38:0] _0460_;
/* cellift = 32'd1 */
wire [38:0] _0461_;
wire [38:0] _0462_;
/* cellift = 32'd1 */
wire [38:0] _0463_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0464_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0465_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0466_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0467_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0468_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0469_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0470_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0471_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0472_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0473_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0474_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0475_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0476_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0477_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0478_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0479_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0480_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0481_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0482_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0483_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0484_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0485_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0486_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0487_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0488_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0489_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0490_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0491_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0492_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0493_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0494_;
/* src = "generated/sv2v_out.v:20139.20-20139.47" */
wire _0495_;
wire _0496_;
wire _0497_;
wire _0498_;
wire _0499_;
wire _0500_;
wire _0501_;
wire _0502_;
wire _0503_;
wire _0504_;
wire _0505_;
wire _0506_;
wire _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0517_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
wire _0525_;
wire _0526_;
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire _0534_;
wire _0535_;
wire _0536_;
wire _0537_;
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0542_;
wire _0543_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
/* src = "generated/sv2v_out.v:20114.13-20114.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:20117.13-20117.29" */
input dummy_instr_id_i;
wire dummy_instr_id_i;
/* cellift = 32'd1 */
input dummy_instr_id_i_t0;
wire dummy_instr_id_i_t0;
/* src = "generated/sv2v_out.v:20118.13-20118.29" */
input dummy_instr_wb_i;
wire dummy_instr_wb_i;
/* cellift = 32'd1 */
input dummy_instr_wb_i_t0;
wire dummy_instr_wb_i_t0;
/* src = "generated/sv2v_out.v:20126.14-20126.19" */
output err_o;
wire err_o;
/* cellift = 32'd1 */
output err_o_t0;
wire err_o_t0;
/* src = "generated/sv2v_out.v:20181.26-20181.33" */
reg [38:0] \g_dummy_r0.rf_r0_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20181.26-20181.33" */
reg [38:0] \g_dummy_r0.rf_r0_q_t0 ;
/* src = "generated/sv2v_out.v:20180.9-20180.20" */
wire \g_dummy_r0.we_r0_dummy ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[10].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[10].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[11].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[11].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[12].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[12].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[13].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[13].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[14].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[14].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[15].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[15].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[16].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[16].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[17].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[17].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[18].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[18].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[19].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[19].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[1].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[1].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[20].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[20].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[21].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[21].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[22].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[22].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[23].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[23].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[24].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[24].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[25].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[25].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[26].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[26].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[27].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[27].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[28].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[28].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[29].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[29].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[2].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[2].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[30].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[30].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[31].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[31].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[3].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[3].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[4].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[4].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[5].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[5].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[6].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[6].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[7].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[7].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[8].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[8].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[9].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20171.26-20171.34" */
reg [38:0] \g_rf_flops[9].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20144.27-20144.39" */
wire [31:0] \gen_wren_check.we_a_dec_buf ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20144.27-20144.39" */
wire [31:0] \gen_wren_check.we_a_dec_buf_t0 ;
/* src = "generated/sv2v_out.v:20119.19-20119.28" */
input [4:0] raddr_a_i;
wire [4:0] raddr_a_i;
/* cellift = 32'd1 */
input [4:0] raddr_a_i_t0;
wire [4:0] raddr_a_i_t0;
/* src = "generated/sv2v_out.v:20121.19-20121.28" */
input [4:0] raddr_b_i;
wire [4:0] raddr_b_i;
/* cellift = 32'd1 */
input [4:0] raddr_b_i_t0;
wire [4:0] raddr_b_i_t0;
/* src = "generated/sv2v_out.v:20120.32-20120.41" */
output [38:0] rdata_a_o;
wire [38:0] rdata_a_o;
/* cellift = 32'd1 */
output [38:0] rdata_a_o_t0;
wire [38:0] rdata_a_o_t0;
/* src = "generated/sv2v_out.v:20122.32-20122.41" */
output [38:0] rdata_b_o;
wire [38:0] rdata_b_o;
/* cellift = 32'd1 */
output [38:0] rdata_b_o_t0;
wire [38:0] rdata_b_o_t0;
/* src = "generated/sv2v_out.v:20129.25-20129.31" */
wire [38:0] \rf_reg[0] ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20129.25-20129.31" */
wire [38:0] \rf_reg[0]_t0 ;
/* src = "generated/sv2v_out.v:20115.13-20115.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:20116.13-20116.22" */
input test_en_i;
wire test_en_i;
/* cellift = 32'd1 */
input test_en_i_t0;
wire test_en_i_t0;
/* src = "generated/sv2v_out.v:20123.19-20123.28" */
input [4:0] waddr_a_i;
wire [4:0] waddr_a_i;
/* cellift = 32'd1 */
input [4:0] waddr_a_i_t0;
wire [4:0] waddr_a_i_t0;
/* src = "generated/sv2v_out.v:20124.31-20124.40" */
input [38:0] wdata_a_i;
wire [38:0] wdata_a_i;
/* cellift = 32'd1 */
input [38:0] wdata_a_i_t0;
wire [38:0] wdata_a_i_t0;
/* src = "generated/sv2v_out.v:20130.24-20130.32" */
wire [31:0] we_a_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20130.24-20130.32" */
wire [31:0] we_a_dec_t0;
/* src = "generated/sv2v_out.v:20125.13-20125.19" */
input we_a_i;
wire we_a_i;
/* cellift = 32'd1 */
input we_a_i_t0;
wire we_a_i_t0;
assign \g_dummy_r0.we_r0_dummy  = we_a_i & /* src = "generated/sv2v_out.v:20182.25-20182.50" */ dummy_instr_wb_i;
assign _0000_ = ~ we_a_dec[31];
assign _0001_ = ~ we_a_dec[30];
assign _0002_ = ~ we_a_dec[29];
assign _0003_ = ~ we_a_dec[28];
assign _0004_ = ~ we_a_dec[27];
assign _0005_ = ~ we_a_dec[26];
assign _0006_ = ~ we_a_dec[25];
assign _0007_ = ~ we_a_dec[24];
assign _0008_ = ~ we_a_dec[23];
assign _0009_ = ~ we_a_dec[22];
assign _0010_ = ~ we_a_dec[21];
assign _0011_ = ~ we_a_dec[20];
assign _0012_ = ~ we_a_dec[19];
assign _0013_ = ~ we_a_dec[18];
assign _0014_ = ~ we_a_dec[17];
assign _0015_ = ~ we_a_dec[16];
assign _0016_ = ~ we_a_dec[15];
assign _0017_ = ~ we_a_dec[14];
assign _0018_ = ~ we_a_dec[13];
assign _0019_ = ~ we_a_dec[12];
assign _0020_ = ~ we_a_dec[11];
assign _0021_ = ~ we_a_dec[10];
assign _0022_ = ~ we_a_dec[9];
assign _0023_ = ~ we_a_dec[8];
assign _0024_ = ~ we_a_dec[7];
assign _0025_ = ~ we_a_dec[6];
assign _0026_ = ~ we_a_dec[5];
assign _0027_ = ~ we_a_dec[4];
assign _0028_ = ~ we_a_dec[3];
assign _0029_ = ~ we_a_dec[2];
assign _0030_ = ~ we_a_dec[1];
assign _0031_ = ~ \g_dummy_r0.we_r0_dummy ;
assign _0108_ = { we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31] } & wdata_a_i_t0;
assign _0110_ = { we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30] } & wdata_a_i_t0;
assign _0112_ = { we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29] } & wdata_a_i_t0;
assign _0114_ = { we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28] } & wdata_a_i_t0;
assign _0116_ = { we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27] } & wdata_a_i_t0;
assign _0118_ = { we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26] } & wdata_a_i_t0;
assign _0120_ = { we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25] } & wdata_a_i_t0;
assign _0122_ = { we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24] } & wdata_a_i_t0;
assign _0124_ = { we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23] } & wdata_a_i_t0;
assign _0126_ = { we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22] } & wdata_a_i_t0;
assign _0128_ = { we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21] } & wdata_a_i_t0;
assign _0130_ = { we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20] } & wdata_a_i_t0;
assign _0132_ = { we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19] } & wdata_a_i_t0;
assign _0134_ = { we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18] } & wdata_a_i_t0;
assign _0136_ = { we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17] } & wdata_a_i_t0;
assign _0138_ = { we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16] } & wdata_a_i_t0;
assign _0140_ = { we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15] } & wdata_a_i_t0;
assign _0142_ = { we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14] } & wdata_a_i_t0;
assign _0144_ = { we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13] } & wdata_a_i_t0;
assign _0146_ = { we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12] } & wdata_a_i_t0;
assign _0148_ = { we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11] } & wdata_a_i_t0;
assign _0150_ = { we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10] } & wdata_a_i_t0;
assign _0152_ = { we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9] } & wdata_a_i_t0;
assign _0154_ = { we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8] } & wdata_a_i_t0;
assign _0156_ = { we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7] } & wdata_a_i_t0;
assign _0158_ = { we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6] } & wdata_a_i_t0;
assign _0160_ = { we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5] } & wdata_a_i_t0;
assign _0162_ = { we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4] } & wdata_a_i_t0;
assign _0164_ = { we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3] } & wdata_a_i_t0;
assign _0166_ = { we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2] } & wdata_a_i_t0;
assign _0168_ = { we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1] } & wdata_a_i_t0;
assign _0170_ = { \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy  } & wdata_a_i_t0;
assign _0109_ = { _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_ } & \g_rf_flops[31].rf_reg_q_t0 ;
assign _0111_ = { _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_ } & \g_rf_flops[30].rf_reg_q_t0 ;
assign _0113_ = { _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_ } & \g_rf_flops[29].rf_reg_q_t0 ;
assign _0115_ = { _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_ } & \g_rf_flops[28].rf_reg_q_t0 ;
assign _0117_ = { _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_ } & \g_rf_flops[27].rf_reg_q_t0 ;
assign _0119_ = { _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_ } & \g_rf_flops[26].rf_reg_q_t0 ;
assign _0121_ = { _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_ } & \g_rf_flops[25].rf_reg_q_t0 ;
assign _0123_ = { _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_ } & \g_rf_flops[24].rf_reg_q_t0 ;
assign _0125_ = { _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_ } & \g_rf_flops[23].rf_reg_q_t0 ;
assign _0127_ = { _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_ } & \g_rf_flops[22].rf_reg_q_t0 ;
assign _0129_ = { _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_ } & \g_rf_flops[21].rf_reg_q_t0 ;
assign _0131_ = { _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_ } & \g_rf_flops[20].rf_reg_q_t0 ;
assign _0133_ = { _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_ } & \g_rf_flops[19].rf_reg_q_t0 ;
assign _0135_ = { _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_ } & \g_rf_flops[18].rf_reg_q_t0 ;
assign _0137_ = { _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_ } & \g_rf_flops[17].rf_reg_q_t0 ;
assign _0139_ = { _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_ } & \g_rf_flops[16].rf_reg_q_t0 ;
assign _0141_ = { _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_ } & \g_rf_flops[15].rf_reg_q_t0 ;
assign _0143_ = { _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_ } & \g_rf_flops[14].rf_reg_q_t0 ;
assign _0145_ = { _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_ } & \g_rf_flops[13].rf_reg_q_t0 ;
assign _0147_ = { _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_ } & \g_rf_flops[12].rf_reg_q_t0 ;
assign _0149_ = { _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_ } & \g_rf_flops[11].rf_reg_q_t0 ;
assign _0151_ = { _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_ } & \g_rf_flops[10].rf_reg_q_t0 ;
assign _0153_ = { _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_ } & \g_rf_flops[9].rf_reg_q_t0 ;
assign _0155_ = { _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_ } & \g_rf_flops[8].rf_reg_q_t0 ;
assign _0157_ = { _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_ } & \g_rf_flops[7].rf_reg_q_t0 ;
assign _0159_ = { _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_ } & \g_rf_flops[6].rf_reg_q_t0 ;
assign _0161_ = { _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_ } & \g_rf_flops[5].rf_reg_q_t0 ;
assign _0163_ = { _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_ } & \g_rf_flops[4].rf_reg_q_t0 ;
assign _0165_ = { _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_ } & \g_rf_flops[3].rf_reg_q_t0 ;
assign _0167_ = { _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_ } & \g_rf_flops[2].rf_reg_q_t0 ;
assign _0169_ = { _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_ } & \g_rf_flops[1].rf_reg_q_t0 ;
assign _0171_ = { _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_ } & \g_dummy_r0.rf_r0_q_t0 ;
assign _0310_ = _0108_ | _0109_;
assign _0311_ = _0110_ | _0111_;
assign _0312_ = _0112_ | _0113_;
assign _0313_ = _0114_ | _0115_;
assign _0314_ = _0116_ | _0117_;
assign _0315_ = _0118_ | _0119_;
assign _0316_ = _0120_ | _0121_;
assign _0317_ = _0122_ | _0123_;
assign _0318_ = _0124_ | _0125_;
assign _0319_ = _0126_ | _0127_;
assign _0320_ = _0128_ | _0129_;
assign _0321_ = _0130_ | _0131_;
assign _0322_ = _0132_ | _0133_;
assign _0323_ = _0134_ | _0135_;
assign _0324_ = _0136_ | _0137_;
assign _0325_ = _0138_ | _0139_;
assign _0326_ = _0140_ | _0141_;
assign _0327_ = _0142_ | _0143_;
assign _0328_ = _0144_ | _0145_;
assign _0329_ = _0146_ | _0147_;
assign _0330_ = _0148_ | _0149_;
assign _0331_ = _0150_ | _0151_;
assign _0332_ = _0152_ | _0153_;
assign _0333_ = _0154_ | _0155_;
assign _0334_ = _0156_ | _0157_;
assign _0335_ = _0158_ | _0159_;
assign _0336_ = _0160_ | _0161_;
assign _0337_ = _0162_ | _0163_;
assign _0338_ = _0164_ | _0165_;
assign _0339_ = _0166_ | _0167_;
assign _0340_ = _0168_ | _0169_;
assign _0341_ = _0170_ | _0171_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[31].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[31].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[31].rf_reg_q_t0  <= _0310_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[30].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[30].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[30].rf_reg_q_t0  <= _0311_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[29].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[29].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[29].rf_reg_q_t0  <= _0312_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[28].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[28].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[28].rf_reg_q_t0  <= _0313_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[27].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[27].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[27].rf_reg_q_t0  <= _0314_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[26].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[26].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[26].rf_reg_q_t0  <= _0315_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[25].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[25].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[25].rf_reg_q_t0  <= _0316_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[24].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[24].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[24].rf_reg_q_t0  <= _0317_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[23].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[23].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[23].rf_reg_q_t0  <= _0318_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[22].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[22].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[22].rf_reg_q_t0  <= _0319_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[21].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[21].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[21].rf_reg_q_t0  <= _0320_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[20].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[20].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[20].rf_reg_q_t0  <= _0321_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[19].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[19].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[19].rf_reg_q_t0  <= _0322_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[18].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[18].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[18].rf_reg_q_t0  <= _0323_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[17].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[17].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[17].rf_reg_q_t0  <= _0324_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[16].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[16].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[16].rf_reg_q_t0  <= _0325_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[15].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[15].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[15].rf_reg_q_t0  <= _0326_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[14].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[14].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[14].rf_reg_q_t0  <= _0327_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[13].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[13].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[13].rf_reg_q_t0  <= _0328_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[12].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[12].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[12].rf_reg_q_t0  <= _0329_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[11].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[11].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[11].rf_reg_q_t0  <= _0330_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[10].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[10].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[10].rf_reg_q_t0  <= _0331_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[9].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[9].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[9].rf_reg_q_t0  <= _0332_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[8].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[8].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[8].rf_reg_q_t0  <= _0333_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[7].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[7].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[7].rf_reg_q_t0  <= _0334_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[6].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[6].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[6].rf_reg_q_t0  <= _0335_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[5].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[5].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[5].rf_reg_q_t0  <= _0336_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[4].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[4].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[4].rf_reg_q_t0  <= _0337_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[3].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[3].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[3].rf_reg_q_t0  <= _0338_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[2].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[2].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[2].rf_reg_q_t0  <= _0339_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[1].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[1].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[1].rf_reg_q_t0  <= _0340_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_dummy_r0.rf_r0_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_dummy_r0.rf_r0_q_t0  <= 39'h0000000000;
else \g_dummy_r0.rf_r0_q_t0  <= _0341_;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[31].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[31].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[31]) \g_rf_flops[31].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[30].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[30].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[30]) \g_rf_flops[30].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[29].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[29].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[29]) \g_rf_flops[29].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[28].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[28].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[28]) \g_rf_flops[28].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[27].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[27].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[27]) \g_rf_flops[27].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[26].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[26].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[26]) \g_rf_flops[26].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[25].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[25].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[25]) \g_rf_flops[25].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[24].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[24].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[24]) \g_rf_flops[24].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[23].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[23].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[23]) \g_rf_flops[23].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[22].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[22].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[22]) \g_rf_flops[22].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[21].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[21].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[21]) \g_rf_flops[21].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[20].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[20].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[20]) \g_rf_flops[20].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[19].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[19].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[19]) \g_rf_flops[19].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[18].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[18].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[18]) \g_rf_flops[18].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[17].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[17].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[17]) \g_rf_flops[17].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[16].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[16].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[16]) \g_rf_flops[16].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[15].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[15].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[15]) \g_rf_flops[15].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[14].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[14].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[14]) \g_rf_flops[14].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[13].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[13].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[13]) \g_rf_flops[13].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[12].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[12].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[12]) \g_rf_flops[12].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[11].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[11].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[11]) \g_rf_flops[11].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[10].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[10].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[10]) \g_rf_flops[10].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[9].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[9].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[9]) \g_rf_flops[9].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[8].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[8].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[8]) \g_rf_flops[8].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[7].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[7].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[7]) \g_rf_flops[7].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[6].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[6].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[6]) \g_rf_flops[6].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[5].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[5].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[5]) \g_rf_flops[5].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[4].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[4].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[4]) \g_rf_flops[4].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[3].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[3].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[3]) \g_rf_flops[3].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[2].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[2].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[2]) \g_rf_flops[2].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20172.4-20176.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[1].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[1].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[1]) \g_rf_flops[1].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20183.4-20187.27" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_dummy_r0.rf_r0_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_dummy_r0.rf_r0_q  <= 39'h2a00000000;
else if (\g_dummy_r0.we_r0_dummy ) \g_dummy_r0.rf_r0_q  <= wdata_a_i;
assign _0032_ = ~ { _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_ };
assign _0033_ = ~ { _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_ };
assign _0034_ = ~ { _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_ };
assign _0035_ = ~ { _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_ };
assign _0036_ = ~ { _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_ };
assign _0037_ = ~ { _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_ };
assign _0038_ = ~ { _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_ };
assign _0039_ = ~ { _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_ };
assign _0040_ = ~ { _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_ };
assign _0041_ = ~ { _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_ };
assign _0042_ = ~ { _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_ };
assign _0043_ = ~ { _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_ };
assign _0044_ = ~ { _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_ };
assign _0045_ = ~ { _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_ };
assign _0046_ = ~ { _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_ };
assign _0047_ = ~ { _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_ };
assign _0048_ = ~ { _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_ };
assign _0049_ = ~ { _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_ };
assign _0050_ = ~ { _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_ };
assign _0051_ = ~ { _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_ };
assign _0052_ = ~ { _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_ };
assign _0053_ = ~ { _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_ };
assign _0054_ = ~ { _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_ };
assign _0055_ = ~ { _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_ };
assign _0056_ = ~ { _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_ };
assign _0057_ = ~ { _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_ };
assign _0058_ = ~ { _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_ };
assign _0059_ = ~ { _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_ };
assign _0060_ = ~ { _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_ };
assign _0061_ = ~ { _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_ };
assign _0062_ = ~ { _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_ };
assign _0063_ = ~ { _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_ };
assign _0064_ = ~ { _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_ };
assign _0065_ = ~ { _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_ };
assign _0066_ = ~ { _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_ };
assign _0067_ = ~ { _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_ };
assign _0068_ = ~ { _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_ };
assign _0069_ = ~ { _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_ };
assign _0070_ = ~ { _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_ };
assign _0071_ = ~ { _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_ };
assign _0072_ = ~ { _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_ };
assign _0073_ = ~ { _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_ };
assign _0074_ = ~ { _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_ };
assign _0075_ = ~ { _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_ };
assign _0076_ = ~ { _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_ };
assign _0077_ = ~ { _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_ };
assign _0078_ = ~ { _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_ };
assign _0079_ = ~ { _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_ };
assign _0080_ = ~ { _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_ };
assign _0081_ = ~ { _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_ };
assign _0082_ = ~ { _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_ };
assign _0083_ = ~ { _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_ };
assign _0084_ = ~ { _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_ };
assign _0085_ = ~ { _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_ };
assign _0086_ = ~ { _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_ };
assign _0087_ = ~ { _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_ };
assign _0088_ = ~ { _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_ };
assign _0089_ = ~ { _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_ };
assign _0090_ = ~ { _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_ };
assign _0091_ = ~ { _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_ };
assign _0092_ = ~ { _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_ };
assign _0093_ = ~ { _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_ };
assign _0172_ = _0032_ & _0463_;
assign _0174_ = _0033_ & \g_rf_flops[22].rf_reg_q_t0 ;
assign _0176_ = _0034_ & \g_rf_flops[20].rf_reg_q_t0 ;
assign _0178_ = _0035_ & _0349_;
assign _0180_ = _0036_ & \g_rf_flops[18].rf_reg_q_t0 ;
assign _0182_ = _0037_ & \g_rf_flops[16].rf_reg_q_t0 ;
assign _0184_ = _0038_ & _0355_;
assign _0186_ = _0039_ & _0357_;
assign _0188_ = _0040_ & _0359_;
assign _0190_ = _0041_ & \g_rf_flops[14].rf_reg_q_t0 ;
assign _0192_ = _0042_ & \g_rf_flops[12].rf_reg_q_t0 ;
assign _0194_ = _0043_ & _0365_;
assign _0196_ = _0044_ & \g_rf_flops[10].rf_reg_q_t0 ;
assign _0198_ = _0045_ & \g_rf_flops[8].rf_reg_q_t0 ;
assign _0200_ = _0046_ & _0371_;
assign _0202_ = _0047_ & _0373_;
assign _0204_ = _0048_ & \g_rf_flops[6].rf_reg_q_t0 ;
assign _0206_ = _0049_ & \g_rf_flops[4].rf_reg_q_t0 ;
assign _0208_ = _0050_ & _0379_;
assign _0210_ = _0051_ & \g_rf_flops[2].rf_reg_q_t0 ;
assign _0212_ = _0052_ & \rf_reg[0]_t0 ;
assign _0214_ = _0053_ & _0385_;
assign _0216_ = _0054_ & _0387_;
assign _0218_ = _0055_ & _0389_;
assign _0220_ = _0056_ & _0391_;
assign _0222_ = _0057_ & \g_rf_flops[30].rf_reg_q_t0 ;
assign _0224_ = _0058_ & \g_rf_flops[28].rf_reg_q_t0 ;
assign _0226_ = _0059_ & _0395_;
assign _0228_ = _0060_ & \g_rf_flops[26].rf_reg_q_t0 ;
assign _0230_ = _0061_ & \g_rf_flops[24].rf_reg_q_t0 ;
assign _0232_ = _0062_ & _0401_;
assign _0234_ = _0063_ & _0403_;
assign _0236_ = _0064_ & \g_rf_flops[22].rf_reg_q_t0 ;
assign _0238_ = _0065_ & \g_rf_flops[20].rf_reg_q_t0 ;
assign _0240_ = _0066_ & _0409_;
assign _0242_ = _0067_ & \g_rf_flops[18].rf_reg_q_t0 ;
assign _0244_ = _0068_ & \g_rf_flops[16].rf_reg_q_t0 ;
assign _0246_ = _0069_ & _0415_;
assign _0248_ = _0070_ & _0417_;
assign _0250_ = _0071_ & _0419_;
assign _0252_ = _0072_ & \g_rf_flops[14].rf_reg_q_t0 ;
assign _0254_ = _0073_ & \g_rf_flops[12].rf_reg_q_t0 ;
assign _0256_ = _0074_ & _0425_;
assign _0258_ = _0075_ & \g_rf_flops[10].rf_reg_q_t0 ;
assign _0260_ = _0076_ & \g_rf_flops[8].rf_reg_q_t0 ;
assign _0262_ = _0077_ & _0431_;
assign _0264_ = _0078_ & _0433_;
assign _0266_ = _0079_ & \g_rf_flops[6].rf_reg_q_t0 ;
assign _0268_ = _0080_ & \g_rf_flops[4].rf_reg_q_t0 ;
assign _0270_ = _0081_ & _0439_;
assign _0272_ = _0082_ & \g_rf_flops[2].rf_reg_q_t0 ;
assign _0274_ = _0083_ & \rf_reg[0]_t0 ;
assign _0276_ = _0084_ & _0445_;
assign _0278_ = _0085_ & _0447_;
assign _0280_ = _0086_ & _0449_;
assign _0282_ = _0087_ & _0451_;
assign _0284_ = _0088_ & \g_rf_flops[30].rf_reg_q_t0 ;
assign _0286_ = _0089_ & \g_rf_flops[28].rf_reg_q_t0 ;
assign _0288_ = _0090_ & _0455_;
assign _0290_ = _0091_ & \g_rf_flops[26].rf_reg_q_t0 ;
assign _0292_ = _0092_ & \g_rf_flops[24].rf_reg_q_t0 ;
assign _0294_ = _0093_ & _0461_;
assign _0173_ = { _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_, _0094_ } & _0457_;
assign _0175_ = { _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_ } & \g_rf_flops[23].rf_reg_q_t0 ;
assign _0177_ = { _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_ } & \g_rf_flops[21].rf_reg_q_t0 ;
assign _0179_ = { _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_, _0296_ } & _0347_;
assign _0181_ = { _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_ } & \g_rf_flops[19].rf_reg_q_t0 ;
assign _0183_ = { _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_ } & \g_rf_flops[17].rf_reg_q_t0 ;
assign _0185_ = { _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_, _0297_ } & _0353_;
assign _0187_ = { _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_, _0095_ } & _0351_;
assign _0189_ = { _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_, _0096_ } & _0345_;
assign _0191_ = { _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_ } & \g_rf_flops[15].rf_reg_q_t0 ;
assign _0193_ = { _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_ } & \g_rf_flops[13].rf_reg_q_t0 ;
assign _0195_ = { _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_, _0298_ } & _0363_;
assign _0197_ = { _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_ } & \g_rf_flops[11].rf_reg_q_t0 ;
assign _0199_ = { _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_ } & \g_rf_flops[9].rf_reg_q_t0 ;
assign _0201_ = { _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_, _0299_ } & _0369_;
assign _0203_ = { _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_, _0097_ } & _0367_;
assign _0205_ = { _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_, _0520_ } & \g_rf_flops[7].rf_reg_q_t0 ;
assign _0207_ = { _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_, _0522_ } & \g_rf_flops[5].rf_reg_q_t0 ;
assign _0209_ = { _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_, _0300_ } & _0377_;
assign _0211_ = { _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_ } & \g_rf_flops[3].rf_reg_q_t0 ;
assign _0213_ = { _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_ } & \g_rf_flops[1].rf_reg_q_t0 ;
assign _0215_ = { _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_, _0301_ } & _0383_;
assign _0217_ = { _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_, _0098_ } & _0381_;
assign _0219_ = { _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_, _0099_ } & _0375_;
assign _0221_ = { _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_ } & _0361_;
assign _0223_ = { _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_ } & \g_rf_flops[31].rf_reg_q_t0 ;
assign _0225_ = { _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_, _0529_ } & \g_rf_flops[29].rf_reg_q_t0 ;
assign _0227_ = { _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_, _0302_ } & _0393_;
assign _0229_ = { _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_, _0531_ } & \g_rf_flops[27].rf_reg_q_t0 ;
assign _0231_ = { _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_, _0533_ } & \g_rf_flops[25].rf_reg_q_t0 ;
assign _0233_ = { _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_, _0303_ } & _0399_;
assign _0235_ = { _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_ } & _0397_;
assign _0237_ = { _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_, _0535_ } & \g_rf_flops[23].rf_reg_q_t0 ;
assign _0239_ = { _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_, _0537_ } & \g_rf_flops[21].rf_reg_q_t0 ;
assign _0241_ = { _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_, _0304_ } & _0407_;
assign _0243_ = { _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_, _0539_ } & \g_rf_flops[19].rf_reg_q_t0 ;
assign _0245_ = { _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_, _0541_ } & \g_rf_flops[17].rf_reg_q_t0 ;
assign _0247_ = { _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_, _0305_ } & _0413_;
assign _0249_ = { _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_, _0102_ } & _0411_;
assign _0251_ = { _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_, _0103_ } & _0405_;
assign _0253_ = { _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_, _0543_ } & \g_rf_flops[15].rf_reg_q_t0 ;
assign _0255_ = { _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_, _0545_ } & \g_rf_flops[13].rf_reg_q_t0 ;
assign _0257_ = { _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_, _0306_ } & _0423_;
assign _0259_ = { _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_, _0547_ } & \g_rf_flops[11].rf_reg_q_t0 ;
assign _0261_ = { _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_, _0549_ } & \g_rf_flops[9].rf_reg_q_t0 ;
assign _0263_ = { _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_, _0307_ } & _0429_;
assign _0265_ = { _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_, _0104_ } & _0427_;
assign _0267_ = { _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_, _0551_ } & \g_rf_flops[7].rf_reg_q_t0 ;
assign _0269_ = { _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_, _0553_ } & \g_rf_flops[5].rf_reg_q_t0 ;
assign _0271_ = { _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_, _0308_ } & _0437_;
assign _0273_ = { _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_, _0555_ } & \g_rf_flops[3].rf_reg_q_t0 ;
assign _0275_ = { _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_, _0557_ } & \g_rf_flops[1].rf_reg_q_t0 ;
assign _0277_ = { _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_, _0309_ } & _0443_;
assign _0279_ = { _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_, _0105_ } & _0441_;
assign _0281_ = { _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_, _0106_ } & _0435_;
assign _0283_ = { _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_, _0107_ } & _0421_;
assign _0285_ = { _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_, _0496_ } & \g_rf_flops[31].rf_reg_q_t0 ;
assign _0287_ = { _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_, _0498_ } & \g_rf_flops[29].rf_reg_q_t0 ;
assign _0289_ = { _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_, _0342_ } & _0453_;
assign _0291_ = { _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_ } & \g_rf_flops[27].rf_reg_q_t0 ;
assign _0293_ = { _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_, _0502_ } & \g_rf_flops[25].rf_reg_q_t0 ;
assign _0295_ = { _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_, _0343_ } & _0459_;
assign we_a_dec_t0[0] = _0464_ & we_a_i_t0;
assign we_a_dec_t0[1] = _0465_ & we_a_i_t0;
assign we_a_dec_t0[2] = _0466_ & we_a_i_t0;
assign we_a_dec_t0[3] = _0467_ & we_a_i_t0;
assign we_a_dec_t0[4] = _0468_ & we_a_i_t0;
assign we_a_dec_t0[5] = _0469_ & we_a_i_t0;
assign we_a_dec_t0[6] = _0470_ & we_a_i_t0;
assign we_a_dec_t0[7] = _0471_ & we_a_i_t0;
assign we_a_dec_t0[8] = _0472_ & we_a_i_t0;
assign we_a_dec_t0[9] = _0473_ & we_a_i_t0;
assign we_a_dec_t0[10] = _0474_ & we_a_i_t0;
assign we_a_dec_t0[11] = _0475_ & we_a_i_t0;
assign we_a_dec_t0[12] = _0476_ & we_a_i_t0;
assign we_a_dec_t0[13] = _0477_ & we_a_i_t0;
assign we_a_dec_t0[14] = _0478_ & we_a_i_t0;
assign we_a_dec_t0[15] = _0479_ & we_a_i_t0;
assign we_a_dec_t0[16] = _0480_ & we_a_i_t0;
assign we_a_dec_t0[17] = _0481_ & we_a_i_t0;
assign we_a_dec_t0[18] = _0482_ & we_a_i_t0;
assign we_a_dec_t0[19] = _0483_ & we_a_i_t0;
assign we_a_dec_t0[20] = _0484_ & we_a_i_t0;
assign we_a_dec_t0[21] = _0485_ & we_a_i_t0;
assign we_a_dec_t0[22] = _0486_ & we_a_i_t0;
assign we_a_dec_t0[23] = _0487_ & we_a_i_t0;
assign we_a_dec_t0[24] = _0488_ & we_a_i_t0;
assign we_a_dec_t0[25] = _0489_ & we_a_i_t0;
assign we_a_dec_t0[26] = _0490_ & we_a_i_t0;
assign we_a_dec_t0[27] = _0491_ & we_a_i_t0;
assign we_a_dec_t0[28] = _0492_ & we_a_i_t0;
assign we_a_dec_t0[29] = _0493_ & we_a_i_t0;
assign we_a_dec_t0[30] = _0494_ & we_a_i_t0;
assign we_a_dec_t0[31] = _0495_ & we_a_i_t0;
assign \rf_reg[0]_t0  = { dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i } & \g_dummy_r0.rf_r0_q_t0 ;
assign _0345_ = _0172_ | _0173_;
assign _0347_ = _0174_ | _0175_;
assign _0349_ = _0176_ | _0177_;
assign _0351_ = _0178_ | _0179_;
assign _0353_ = _0180_ | _0181_;
assign _0355_ = _0182_ | _0183_;
assign _0357_ = _0184_ | _0185_;
assign _0359_ = _0186_ | _0187_;
assign _0361_ = _0188_ | _0189_;
assign _0363_ = _0190_ | _0191_;
assign _0365_ = _0192_ | _0193_;
assign _0367_ = _0194_ | _0195_;
assign _0369_ = _0196_ | _0197_;
assign _0371_ = _0198_ | _0199_;
assign _0373_ = _0200_ | _0201_;
assign _0375_ = _0202_ | _0203_;
assign _0377_ = _0204_ | _0205_;
assign _0379_ = _0206_ | _0207_;
assign _0381_ = _0208_ | _0209_;
assign _0383_ = _0210_ | _0211_;
assign _0385_ = _0212_ | _0213_;
assign _0387_ = _0214_ | _0215_;
assign _0389_ = _0216_ | _0217_;
assign _0391_ = _0218_ | _0219_;
assign rdata_b_o_t0 = _0220_ | _0221_;
assign _0393_ = _0222_ | _0223_;
assign _0395_ = _0224_ | _0225_;
assign _0397_ = _0226_ | _0227_;
assign _0399_ = _0228_ | _0229_;
assign _0401_ = _0230_ | _0231_;
assign _0403_ = _0232_ | _0233_;
assign _0405_ = _0234_ | _0235_;
assign _0407_ = _0236_ | _0237_;
assign _0409_ = _0238_ | _0239_;
assign _0411_ = _0240_ | _0241_;
assign _0413_ = _0242_ | _0243_;
assign _0415_ = _0244_ | _0245_;
assign _0417_ = _0246_ | _0247_;
assign _0419_ = _0248_ | _0249_;
assign _0421_ = _0250_ | _0251_;
assign _0423_ = _0252_ | _0253_;
assign _0425_ = _0254_ | _0255_;
assign _0427_ = _0256_ | _0257_;
assign _0429_ = _0258_ | _0259_;
assign _0431_ = _0260_ | _0261_;
assign _0433_ = _0262_ | _0263_;
assign _0435_ = _0264_ | _0265_;
assign _0437_ = _0266_ | _0267_;
assign _0439_ = _0268_ | _0269_;
assign _0441_ = _0270_ | _0271_;
assign _0443_ = _0272_ | _0273_;
assign _0445_ = _0274_ | _0275_;
assign _0447_ = _0276_ | _0277_;
assign _0449_ = _0278_ | _0279_;
assign _0451_ = _0280_ | _0281_;
assign rdata_a_o_t0 = _0282_ | _0283_;
assign _0453_ = _0284_ | _0285_;
assign _0455_ = _0286_ | _0287_;
assign _0457_ = _0288_ | _0289_;
assign _0459_ = _0290_ | _0291_;
assign _0461_ = _0292_ | _0293_;
assign _0463_ = _0294_ | _0295_;
assign _0296_ = _0505_ | _0504_;
assign _0297_ = _0509_ | _0508_;
assign _0298_ = _0513_ | _0512_;
assign _0299_ = _0517_ | _0516_;
assign _0300_ = _0521_ | _0520_;
assign _0301_ = _0525_ | _0524_;
assign _0302_ = _0528_ | _0527_;
assign _0303_ = _0532_ | _0531_;
assign _0304_ = _0536_ | _0535_;
assign _0305_ = _0540_ | _0539_;
assign _0306_ = _0544_ | _0543_;
assign _0307_ = _0548_ | _0547_;
assign _0308_ = _0552_ | _0551_;
assign _0309_ = _0556_ | _0555_;
assign _0342_ = _0497_ | _0496_;
assign _0343_ = _0501_ | _0500_;
assign _0094_ = | { _0342_, _0499_, _0498_ };
assign _0095_ = | { _0296_, _0507_, _0506_ };
assign _0096_ = | { _0342_, _0343_, _0503_, _0502_, _0499_, _0498_ };
assign _0097_ = | { _0298_, _0514_, _0515_ };
assign _0098_ = | { _0300_, _0523_, _0522_ };
assign _0099_ = | { _0298_, _0299_, _0519_, _0518_, _0514_, _0515_ };
assign _0100_ = | { _0342_, _0343_, _0296_, _0297_, _0511_, _0510_, _0507_, _0506_, _0503_, _0502_, _0499_, _0498_ };
assign _0101_ = | { _0302_, _0530_, _0529_ };
assign _0102_ = | { _0304_, _0538_, _0537_ };
assign _0103_ = | { _0302_, _0303_, _0534_, _0533_, _0530_, _0529_ };
assign _0104_ = | { _0306_, _0546_, _0545_ };
assign _0105_ = | { _0308_, _0554_, _0553_ };
assign _0106_ = | { _0306_, _0307_, _0550_, _0549_, _0546_, _0545_ };
assign _0107_ = | { _0302_, _0303_, _0304_, _0305_, _0542_, _0541_, _0538_, _0537_, _0534_, _0533_, _0530_, _0529_ };
assign _0344_ = _0094_ ? _0456_ : _0462_;
assign _0346_ = _0504_ ? \g_rf_flops[23].rf_reg_q  : \g_rf_flops[22].rf_reg_q ;
assign _0348_ = _0506_ ? \g_rf_flops[21].rf_reg_q  : \g_rf_flops[20].rf_reg_q ;
assign _0350_ = _0296_ ? _0346_ : _0348_;
assign _0352_ = _0508_ ? \g_rf_flops[19].rf_reg_q  : \g_rf_flops[18].rf_reg_q ;
assign _0354_ = _0510_ ? \g_rf_flops[17].rf_reg_q  : \g_rf_flops[16].rf_reg_q ;
assign _0356_ = _0297_ ? _0352_ : _0354_;
assign _0358_ = _0095_ ? _0350_ : _0356_;
assign _0360_ = _0096_ ? _0344_ : _0358_;
assign _0362_ = _0512_ ? \g_rf_flops[15].rf_reg_q  : \g_rf_flops[14].rf_reg_q ;
assign _0364_ = _0514_ ? \g_rf_flops[13].rf_reg_q  : \g_rf_flops[12].rf_reg_q ;
assign _0366_ = _0298_ ? _0362_ : _0364_;
assign _0368_ = _0516_ ? \g_rf_flops[11].rf_reg_q  : \g_rf_flops[10].rf_reg_q ;
assign _0370_ = _0518_ ? \g_rf_flops[9].rf_reg_q  : \g_rf_flops[8].rf_reg_q ;
assign _0372_ = _0299_ ? _0368_ : _0370_;
assign _0374_ = _0097_ ? _0366_ : _0372_;
assign _0376_ = _0520_ ? \g_rf_flops[7].rf_reg_q  : \g_rf_flops[6].rf_reg_q ;
assign _0378_ = _0522_ ? \g_rf_flops[5].rf_reg_q  : \g_rf_flops[4].rf_reg_q ;
assign _0380_ = _0300_ ? _0376_ : _0378_;
assign _0382_ = _0524_ ? \g_rf_flops[3].rf_reg_q  : \g_rf_flops[2].rf_reg_q ;
assign _0384_ = _0526_ ? \g_rf_flops[1].rf_reg_q  : \rf_reg[0] ;
assign _0386_ = _0301_ ? _0382_ : _0384_;
assign _0388_ = _0098_ ? _0380_ : _0386_;
assign _0390_ = _0099_ ? _0374_ : _0388_;
assign rdata_b_o = _0100_ ? _0360_ : _0390_;
assign _0392_ = _0527_ ? \g_rf_flops[31].rf_reg_q  : \g_rf_flops[30].rf_reg_q ;
assign _0394_ = _0529_ ? \g_rf_flops[29].rf_reg_q  : \g_rf_flops[28].rf_reg_q ;
assign _0396_ = _0302_ ? _0392_ : _0394_;
assign _0398_ = _0531_ ? \g_rf_flops[27].rf_reg_q  : \g_rf_flops[26].rf_reg_q ;
assign _0400_ = _0533_ ? \g_rf_flops[25].rf_reg_q  : \g_rf_flops[24].rf_reg_q ;
assign _0402_ = _0303_ ? _0398_ : _0400_;
assign _0404_ = _0101_ ? _0396_ : _0402_;
assign _0406_ = _0535_ ? \g_rf_flops[23].rf_reg_q  : \g_rf_flops[22].rf_reg_q ;
assign _0408_ = _0537_ ? \g_rf_flops[21].rf_reg_q  : \g_rf_flops[20].rf_reg_q ;
assign _0410_ = _0304_ ? _0406_ : _0408_;
assign _0412_ = _0539_ ? \g_rf_flops[19].rf_reg_q  : \g_rf_flops[18].rf_reg_q ;
assign _0414_ = _0541_ ? \g_rf_flops[17].rf_reg_q  : \g_rf_flops[16].rf_reg_q ;
assign _0416_ = _0305_ ? _0412_ : _0414_;
assign _0418_ = _0102_ ? _0410_ : _0416_;
assign _0420_ = _0103_ ? _0404_ : _0418_;
assign _0422_ = _0543_ ? \g_rf_flops[15].rf_reg_q  : \g_rf_flops[14].rf_reg_q ;
assign _0424_ = _0545_ ? \g_rf_flops[13].rf_reg_q  : \g_rf_flops[12].rf_reg_q ;
assign _0426_ = _0306_ ? _0422_ : _0424_;
assign _0428_ = _0547_ ? \g_rf_flops[11].rf_reg_q  : \g_rf_flops[10].rf_reg_q ;
assign _0430_ = _0549_ ? \g_rf_flops[9].rf_reg_q  : \g_rf_flops[8].rf_reg_q ;
assign _0432_ = _0307_ ? _0428_ : _0430_;
assign _0434_ = _0104_ ? _0426_ : _0432_;
assign _0436_ = _0551_ ? \g_rf_flops[7].rf_reg_q  : \g_rf_flops[6].rf_reg_q ;
assign _0438_ = _0553_ ? \g_rf_flops[5].rf_reg_q  : \g_rf_flops[4].rf_reg_q ;
assign _0440_ = _0308_ ? _0436_ : _0438_;
assign _0442_ = _0555_ ? \g_rf_flops[3].rf_reg_q  : \g_rf_flops[2].rf_reg_q ;
assign _0444_ = _0557_ ? \g_rf_flops[1].rf_reg_q  : \rf_reg[0] ;
assign _0446_ = _0309_ ? _0442_ : _0444_;
assign _0448_ = _0105_ ? _0440_ : _0446_;
assign _0450_ = _0106_ ? _0434_ : _0448_;
assign rdata_a_o = _0107_ ? _0420_ : _0450_;
assign _0452_ = _0496_ ? \g_rf_flops[31].rf_reg_q  : \g_rf_flops[30].rf_reg_q ;
assign _0454_ = _0498_ ? \g_rf_flops[29].rf_reg_q  : \g_rf_flops[28].rf_reg_q ;
assign _0456_ = _0342_ ? _0452_ : _0454_;
assign _0458_ = _0500_ ? \g_rf_flops[27].rf_reg_q  : \g_rf_flops[26].rf_reg_q ;
assign _0460_ = _0502_ ? \g_rf_flops[25].rf_reg_q  : \g_rf_flops[24].rf_reg_q ;
assign _0462_ = _0343_ ? _0458_ : _0460_;
assign _0464_ = ! /* src = "generated/sv2v_out.v:20139.20-20139.47" */ waddr_a_i;
assign _0465_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h01;
assign _0466_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h02;
assign _0467_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h03;
assign _0468_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h04;
assign _0469_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h05;
assign _0470_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h06;
assign _0471_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h07;
assign _0472_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h08;
assign _0473_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h09;
assign _0474_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h0a;
assign _0475_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h0b;
assign _0476_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h0c;
assign _0477_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h0d;
assign _0478_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h0e;
assign _0479_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h0f;
assign _0480_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h10;
assign _0481_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h11;
assign _0482_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h12;
assign _0483_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h13;
assign _0484_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h14;
assign _0485_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h15;
assign _0486_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h16;
assign _0487_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h17;
assign _0488_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h18;
assign _0489_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h19;
assign _0490_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h1a;
assign _0491_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h1b;
assign _0492_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h1c;
assign _0493_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h1d;
assign _0494_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h1e;
assign _0495_ = waddr_a_i == /* src = "generated/sv2v_out.v:20139.20-20139.47" */ 5'h1f;
assign _0496_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1f;
assign _0497_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1e;
assign _0498_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1d;
assign _0499_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1c;
assign _0500_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1b;
assign _0501_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1a;
assign _0502_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h19;
assign _0503_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h18;
assign _0504_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h17;
assign _0505_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h16;
assign _0506_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h15;
assign _0507_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h14;
assign _0508_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h13;
assign _0509_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h12;
assign _0510_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h11;
assign _0511_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h10;
assign _0512_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0f;
assign _0513_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0e;
assign _0514_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0d;
assign _0515_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0c;
assign _0516_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0b;
assign _0517_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0a;
assign _0518_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h09;
assign _0519_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h08;
assign _0520_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h07;
assign _0521_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h06;
assign _0522_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h05;
assign _0523_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h04;
assign _0524_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h03;
assign _0525_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h02;
assign _0526_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h01;
assign _0527_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1f;
assign _0528_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1e;
assign _0529_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1d;
assign _0530_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1c;
assign _0531_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1b;
assign _0532_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1a;
assign _0533_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h19;
assign _0534_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h18;
assign _0535_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h17;
assign _0536_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h16;
assign _0537_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h15;
assign _0538_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h14;
assign _0539_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h13;
assign _0540_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h12;
assign _0541_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h11;
assign _0542_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h10;
assign _0543_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0f;
assign _0544_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0e;
assign _0545_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0d;
assign _0546_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0c;
assign _0547_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0b;
assign _0548_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0a;
assign _0549_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h09;
assign _0550_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h08;
assign _0551_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h07;
assign _0552_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h06;
assign _0553_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h05;
assign _0554_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h04;
assign _0555_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h03;
assign _0556_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h02;
assign _0557_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h01;
assign we_a_dec[0] = _0464_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[1] = _0465_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[2] = _0466_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[3] = _0467_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[4] = _0468_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[5] = _0469_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[6] = _0470_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[7] = _0471_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[8] = _0472_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[9] = _0473_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[10] = _0474_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[11] = _0475_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[12] = _0476_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[13] = _0477_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[14] = _0478_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[15] = _0479_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[16] = _0480_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[17] = _0481_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[18] = _0482_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[19] = _0483_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[20] = _0484_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[21] = _0485_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[22] = _0486_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[23] = _0487_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[24] = _0488_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[25] = _0489_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[26] = _0490_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[27] = _0491_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[28] = _0492_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[29] = _0493_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[30] = _0494_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign we_a_dec[31] = _0495_ ? /* src = "generated/sv2v_out.v:20139.20-20139.63" */ we_a_i : 1'h0;
assign \rf_reg[0]  = dummy_instr_id_i ? /* src = "generated/sv2v_out.v:20188.24-20188.64" */ \g_dummy_r0.rf_r0_q  : 39'h2a00000000;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20145.34-20148.5" */
\$paramod\prim_buf\Width=32'00000000000000000000000000100000  \gen_wren_check.u_prim_buf  (
.in_i(we_a_dec),
.in_i_t0(we_a_dec_t0),
.out_o(\gen_wren_check.we_a_dec_buf ),
.out_o_t0(\gen_wren_check.we_a_dec_buf_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20153.6-20160.5" */
\$paramod$916c47de983e2a42946808797a4a11650abb788f\prim_onehot_check  \gen_wren_check.u_prim_onehot_check  (
.addr_i(waddr_a_i),
.addr_i_t0(waddr_a_i_t0),
.clk_i(clk_i),
.en_i(we_a_i),
.en_i_t0(we_a_i_t0),
.err_o(err_o),
.err_o_t0(err_o_t0),
.oh_i(\gen_wren_check.we_a_dec_buf ),
.oh_i_t0(\gen_wren_check.we_a_dec_buf_t0 ),
.rst_ni(rst_ni)
);
endmodule

module \$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers (clk_i, rst_ni, hart_id_i, priv_mode_id_o, priv_mode_lsu_o, csr_mstatus_tw_o, csr_mtvec_o, csr_mtvec_init_i, boot_addr_i, csr_access_i, csr_addr_i, csr_wdata_i, csr_op_i, csr_op_en_i, csr_rdata_o, irq_software_i, irq_timer_i, irq_external_i, irq_fast_i, nmi_mode_i, irq_pending_o
, irqs_o, csr_mstatus_mie_o, csr_mepc_o, csr_mtval_o, csr_pmp_cfg_o, csr_pmp_addr_o, csr_pmp_mseccfg_o, debug_mode_i, debug_mode_entering_i, debug_cause_i, debug_csr_save_i, csr_depc_o, debug_single_step_o, debug_ebreakm_o, debug_ebreaku_o, trigger_match_o, pc_if_i, pc_id_i, pc_wb_i, data_ind_timing_o, dummy_instr_en_o
, dummy_instr_mask_o, dummy_instr_seed_en_o, dummy_instr_seed_o, icache_enable_o, csr_shadow_err_o, ic_scr_key_valid_i, csr_save_if_i, csr_save_id_i, csr_save_wb_i, csr_restore_mret_i, csr_restore_dret_i, csr_save_cause_i, csr_mcause_i, csr_mtval_i, illegal_csr_insn_o, double_fault_seen_o, instr_ret_i, instr_ret_compressed_i, instr_ret_spec_i, instr_ret_compressed_spec_i, iside_wait_i
, jump_i, branch_i, branch_taken_i, mem_load_i, mem_store_i, dside_wait_i, mul_wait_i, div_wait_i, pc_id_i_t0, csr_mtval_o_t0, ic_scr_key_valid_i_t0, boot_addr_i_t0, branch_taken_i_t0, branch_i_t0, csr_access_i_t0, csr_addr_i_t0, csr_depc_o_t0, csr_mcause_i_t0, csr_mepc_o_t0, csr_mstatus_mie_o_t0, csr_mstatus_tw_o_t0
, csr_mtval_i_t0, csr_mtvec_init_i_t0, csr_mtvec_o_t0, csr_op_en_i_t0, csr_op_i_t0, csr_pmp_addr_o_t0, csr_pmp_cfg_o_t0, csr_pmp_mseccfg_o_t0, csr_rdata_o_t0, csr_restore_dret_i_t0, csr_restore_mret_i_t0, csr_save_cause_i_t0, csr_save_id_i_t0, csr_save_if_i_t0, csr_save_wb_i_t0, csr_shadow_err_o_t0, csr_wdata_i_t0, data_ind_timing_o_t0, debug_cause_i_t0, debug_csr_save_i_t0, debug_ebreakm_o_t0
, debug_ebreaku_o_t0, debug_mode_entering_i_t0, debug_mode_i_t0, debug_single_step_o_t0, div_wait_i_t0, double_fault_seen_o_t0, dside_wait_i_t0, dummy_instr_en_o_t0, dummy_instr_mask_o_t0, dummy_instr_seed_en_o_t0, dummy_instr_seed_o_t0, hart_id_i_t0, icache_enable_o_t0, illegal_csr_insn_o_t0, instr_ret_compressed_i_t0, instr_ret_compressed_spec_i_t0, instr_ret_i_t0, instr_ret_spec_i_t0, irq_external_i_t0, irq_fast_i_t0, irq_pending_o_t0
, irq_software_i_t0, irq_timer_i_t0, irqs_o_t0, iside_wait_i_t0, jump_i_t0, mem_load_i_t0, mem_store_i_t0, mul_wait_i_t0, nmi_mode_i_t0, pc_if_i_t0, pc_wb_i_t0, priv_mode_id_o_t0, priv_mode_lsu_o_t0, trigger_match_o_t0);
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [7:0] _0000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [7:0] _0001_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0002_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0003_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0004_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0005_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0006_;
/* src = "generated/sv2v_out.v:14024.2-14154.5" */
wire _0007_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0008_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0009_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [5:0] _0010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [5:0] _0011_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0012_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0013_;
/* src = "generated/sv2v_out.v:14024.2-14154.5" */
wire [63:0] _0014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14024.2-14154.5" */
wire [63:0] _0015_;
/* src = "generated/sv2v_out.v:14024.2-14154.5" */
wire [31:0] _0016_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [7:0] _0017_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [7:0] _0018_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0019_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0021_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0022_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0023_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0024_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0025_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0026_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0027_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0028_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0029_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0030_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [6:0] _0031_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [6:0] _0032_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0033_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0034_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0035_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0036_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0037_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0038_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0039_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0040_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0041_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0042_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0043_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0044_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [5:0] _0045_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [5:0] _0046_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0047_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0048_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0049_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0050_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0051_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0052_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [1:0] _0053_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [1:0] _0054_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0055_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [6:0] _0056_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [6:0] _0057_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0058_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0059_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0060_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [1:0] _0061_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [1:0] _0062_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0063_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0064_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [1:0] _0065_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [1:0] _0066_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0067_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0068_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0069_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0070_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [6:0] _0071_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [6:0] _0072_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0073_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0074_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [31:0] _0075_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0076_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0077_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0078_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [1:0] _0079_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [1:0] _0080_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0081_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0082_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0083_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0084_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [3:0] _0085_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [3:0] _0086_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0087_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0088_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [1:0] _0089_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [1:0] _0090_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0091_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [1:0] _0092_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [1:0] _0093_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0094_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0095_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [3:0] _0096_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [3:0] _0097_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0098_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0099_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [2:0] _0100_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [2:0] _0101_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0102_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire _0103_;
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [2:0] _0104_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14159.2-14298.5" */
wire [2:0] _0105_;
/* src = "generated/sv2v_out.v:14310.26-14310.52" */
wire [31:0] _0106_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14310.26-14310.52" */
wire [31:0] _0107_;
/* src = "generated/sv2v_out.v:14315.23-14315.43" */
wire _0108_;
/* src = "generated/sv2v_out.v:14687.18-14687.57" */
wire _0109_;
/* src = "generated/sv2v_out.v:14699.18-14699.57" */
wire _0110_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14699.18-14699.57" */
wire _0111_;
/* src = "generated/sv2v_out.v:14706.27-14706.63" */
wire _0112_;
wire _0113_;
wire _0114_;
wire [31:0] _0115_;
wire [31:0] _0116_;
wire _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire [2:0] _0139_;
wire [2:0] _0140_;
wire [2:0] _0141_;
wire [2:0] _0142_;
wire [2:0] _0143_;
wire [2:0] _0144_;
wire [2:0] _0145_;
wire [2:0] _0146_;
wire [2:0] _0147_;
wire [2:0] _0148_;
wire [2:0] _0149_;
wire [2:0] _0150_;
wire [2:0] _0151_;
wire [2:0] _0152_;
wire [2:0] _0153_;
wire [2:0] _0154_;
wire [2:0] _0155_;
wire [2:0] _0156_;
wire [2:0] _0157_;
wire [2:0] _0158_;
wire [2:0] _0159_;
wire [2:0] _0160_;
wire [2:0] _0161_;
wire [2:0] _0162_;
wire [2:0] _0163_;
wire [2:0] _0164_;
wire [2:0] _0165_;
wire [2:0] _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire [2:0] _0178_;
wire [2:0] _0179_;
wire [2:0] _0180_;
wire [2:0] _0181_;
wire [8:0] _0182_;
wire [8:0] _0183_;
wire [8:0] _0184_;
wire [8:0] _0185_;
wire [8:0] _0186_;
wire [8:0] _0187_;
wire [8:0] _0188_;
wire [8:0] _0189_;
wire [8:0] _0190_;
wire [8:0] _0191_;
wire [8:0] _0192_;
wire [8:0] _0193_;
wire [8:0] _0194_;
wire [8:0] _0195_;
wire [63:0] _0196_;
wire [63:0] _0197_;
wire _0198_;
wire [31:0] _0199_;
wire _0200_;
wire [2:0] _0201_;
wire [2:0] _0202_;
wire [2:0] _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire [1:0] _0209_;
wire [6:0] _0210_;
wire [31:0] _0211_;
wire [31:0] _0212_;
wire [2:0] _0213_;
wire [1:0] _0214_;
wire [6:0] _0215_;
wire [3:0] _0216_;
wire [31:0] _0217_;
wire [31:0] _0218_;
wire [31:0] _0219_;
wire [31:0] _0220_;
wire [1:0] _0221_;
wire [6:0] _0222_;
wire [6:0] _0223_;
wire [6:0] _0224_;
wire [31:0] _0225_;
wire [31:0] _0226_;
wire [6:0] _0227_;
wire [1:0] _0228_;
wire [3:0] _0229_;
wire [1:0] _0230_;
wire [11:0] _0231_;
wire [1:0] _0232_;
wire [1:0] _0233_;
wire [1:0] _0234_;
wire [7:0] _0235_;
wire _0236_;
wire [7:0] _0237_;
wire [31:0] _0238_;
wire [5:0] _0239_;
wire [31:0] _0240_;
wire [1:0] _0241_;
wire [63:0] _0242_;
wire _0243_;
wire _0244_;
wire [31:0] _0245_;
wire _0246_;
wire _0247_;
wire _0248_;
wire [31:0] _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire _0271_;
wire _0272_;
wire _0273_;
wire [31:0] _0274_;
wire [31:0] _0275_;
wire [31:0] _0276_;
wire [17:0] _0277_;
wire [17:0] _0278_;
wire [17:0] _0279_;
wire _0280_;
wire _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire _0285_;
wire [1:0] _0286_;
wire [1:0] _0287_;
wire [1:0] _0288_;
wire [1:0] _0289_;
wire [31:0] _0290_;
wire [31:0] _0291_;
wire [31:0] _0292_;
wire [31:0] _0293_;
wire _0294_;
wire _0295_;
wire _0296_;
wire _0297_;
wire _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire _0324_;
wire _0325_;
wire _0326_;
wire _0327_;
wire _0328_;
wire _0329_;
wire _0330_;
wire _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire _0335_;
wire _0336_;
wire _0337_;
wire _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire [2:0] _0344_;
wire [2:0] _0345_;
wire [2:0] _0346_;
wire [2:0] _0347_;
wire [2:0] _0348_;
wire [2:0] _0349_;
wire [2:0] _0350_;
wire [2:0] _0351_;
wire [2:0] _0352_;
wire [2:0] _0353_;
wire [2:0] _0354_;
wire [2:0] _0355_;
wire [2:0] _0356_;
wire [2:0] _0357_;
wire [2:0] _0358_;
wire [2:0] _0359_;
wire [2:0] _0360_;
wire [2:0] _0361_;
wire [2:0] _0362_;
wire [2:0] _0363_;
wire [2:0] _0364_;
wire [2:0] _0365_;
wire [2:0] _0366_;
wire [2:0] _0367_;
wire _0368_;
wire _0369_;
wire _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire _0376_;
wire _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire _0382_;
wire _0383_;
wire _0384_;
wire _0385_;
wire _0386_;
wire _0387_;
wire _0388_;
wire _0389_;
wire _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire [2:0] _0398_;
wire [2:0] _0399_;
wire [2:0] _0400_;
wire [2:0] _0401_;
wire [2:0] _0402_;
wire [2:0] _0403_;
wire [2:0] _0404_;
wire [2:0] _0405_;
wire [2:0] _0406_;
wire [2:0] _0407_;
wire [2:0] _0408_;
wire [2:0] _0409_;
wire [2:0] _0410_;
wire [2:0] _0411_;
wire [2:0] _0412_;
wire [2:0] _0413_;
wire [2:0] _0414_;
wire [2:0] _0415_;
wire [2:0] _0416_;
wire [2:0] _0417_;
wire [2:0] _0418_;
wire [2:0] _0419_;
wire [2:0] _0420_;
wire [2:0] _0421_;
wire [2:0] _0422_;
wire [2:0] _0423_;
wire [2:0] _0424_;
wire [2:0] _0425_;
wire [2:0] _0426_;
wire [2:0] _0427_;
wire [2:0] _0428_;
wire [2:0] _0429_;
wire [2:0] _0430_;
wire [2:0] _0431_;
wire [2:0] _0432_;
wire [2:0] _0433_;
wire [2:0] _0434_;
wire [2:0] _0435_;
wire [2:0] _0436_;
wire [2:0] _0437_;
wire [2:0] _0438_;
wire [2:0] _0439_;
wire [2:0] _0440_;
wire [2:0] _0441_;
wire [2:0] _0442_;
wire [2:0] _0443_;
wire [2:0] _0444_;
wire [2:0] _0445_;
wire [2:0] _0446_;
wire [2:0] _0447_;
wire [2:0] _0448_;
wire [2:0] _0449_;
wire [2:0] _0450_;
wire [2:0] _0451_;
wire [2:0] _0452_;
wire [2:0] _0453_;
wire [2:0] _0454_;
wire [2:0] _0455_;
wire [2:0] _0456_;
wire [2:0] _0457_;
wire [2:0] _0458_;
wire [2:0] _0459_;
wire [2:0] _0460_;
wire [2:0] _0461_;
wire [2:0] _0462_;
wire [2:0] _0463_;
wire [2:0] _0464_;
wire [2:0] _0465_;
wire [2:0] _0466_;
wire [2:0] _0467_;
wire _0468_;
wire _0469_;
wire _0470_;
wire _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire _0477_;
wire _0478_;
wire _0479_;
wire _0480_;
wire _0481_;
wire _0482_;
wire _0483_;
wire _0484_;
wire _0485_;
wire _0486_;
wire _0487_;
wire _0488_;
wire _0489_;
wire _0490_;
wire _0491_;
wire _0492_;
wire _0493_;
wire _0494_;
wire _0495_;
wire _0496_;
wire _0497_;
wire _0498_;
wire _0499_;
wire _0500_;
wire _0501_;
wire _0502_;
wire _0503_;
wire _0504_;
wire _0505_;
wire _0506_;
wire _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire [2:0] _0516_;
wire [2:0] _0517_;
wire [2:0] _0518_;
wire [2:0] _0519_;
wire [2:0] _0520_;
wire [2:0] _0521_;
wire [2:0] _0522_;
wire [2:0] _0523_;
wire [2:0] _0524_;
wire [2:0] _0525_;
wire [2:0] _0526_;
wire [2:0] _0527_;
wire [2:0] _0528_;
wire [2:0] _0529_;
wire [2:0] _0530_;
wire [2:0] _0531_;
wire [2:0] _0532_;
wire [2:0] _0533_;
wire [2:0] _0534_;
wire [2:0] _0535_;
wire _0536_;
wire _0537_;
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0542_;
wire _0543_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire [8:0] _0560_;
wire [8:0] _0561_;
wire [8:0] _0562_;
wire [8:0] _0563_;
wire [8:0] _0564_;
wire [8:0] _0565_;
wire [8:0] _0566_;
wire [8:0] _0567_;
wire [8:0] _0568_;
wire [8:0] _0569_;
wire [8:0] _0570_;
wire [8:0] _0571_;
wire [8:0] _0572_;
wire [8:0] _0573_;
wire [8:0] _0574_;
wire [8:0] _0575_;
wire [8:0] _0576_;
wire [8:0] _0577_;
wire [8:0] _0578_;
wire [8:0] _0579_;
wire [8:0] _0580_;
wire [8:0] _0581_;
wire [8:0] _0582_;
wire [8:0] _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire _0596_;
wire _0597_;
wire _0598_;
wire _0599_;
wire _0600_;
wire _0601_;
wire _0602_;
wire _0603_;
wire _0604_;
wire _0605_;
wire _0606_;
wire _0607_;
wire _0608_;
wire _0609_;
wire [63:0] _0610_;
wire [63:0] _0611_;
wire _0612_;
wire _0613_;
wire _0614_;
wire _0615_;
wire _0616_;
wire _0617_;
wire _0618_;
wire _0619_;
wire _0620_;
wire _0621_;
wire _0622_;
wire _0623_;
wire _0624_;
wire _0625_;
wire _0626_;
wire _0627_;
wire _0628_;
wire _0629_;
wire _0630_;
wire _0631_;
wire _0632_;
wire _0633_;
wire _0634_;
wire _0635_;
wire _0636_;
wire _0637_;
wire _0638_;
wire _0639_;
wire _0640_;
wire [31:0] _0641_;
wire _0642_;
wire _0643_;
wire _0644_;
wire _0645_;
wire _0646_;
wire _0647_;
wire _0648_;
wire _0649_;
wire _0650_;
wire _0651_;
wire _0652_;
wire [31:0] _0653_;
wire [31:0] _0654_;
wire [2:0] _0655_;
wire [2:0] _0656_;
wire [2:0] _0657_;
wire [2:0] _0658_;
wire [2:0] _0659_;
wire [2:0] _0660_;
wire _0661_;
wire _0662_;
wire _0663_;
wire _0664_;
wire _0665_;
wire _0666_;
wire _0667_;
wire _0668_;
wire _0669_;
wire _0670_;
wire _0671_;
wire _0672_;
wire [1:0] _0673_;
wire [1:0] _0674_;
wire [6:0] _0675_;
wire [6:0] _0676_;
wire [31:0] _0677_;
wire [31:0] _0678_;
wire _0679_;
wire _0680_;
wire [1:0] _0681_;
wire [1:0] _0682_;
wire _0683_;
wire _0684_;
wire [31:0] _0685_;
wire [31:0] _0686_;
wire [31:0] _0687_;
wire [31:0] _0688_;
wire [2:0] _0689_;
wire [2:0] _0690_;
wire [1:0] _0691_;
wire [1:0] _0692_;
wire [1:0] _0693_;
wire [1:0] _0694_;
wire [31:0] _0695_;
wire [31:0] _0696_;
wire [6:0] _0697_;
wire [6:0] _0698_;
wire [31:0] _0699_;
wire [31:0] _0700_;
wire [3:0] _0701_;
wire [3:0] _0702_;
wire [31:0] _0703_;
wire [31:0] _0704_;
wire [31:0] _0705_;
wire [31:0] _0706_;
wire [31:0] _0707_;
wire [31:0] _0708_;
wire _0709_;
wire _0710_;
wire _0711_;
wire _0712_;
wire [31:0] _0713_;
wire [31:0] _0714_;
wire [2:0] _0715_;
wire [2:0] _0716_;
wire [1:0] _0717_;
wire [1:0] _0718_;
wire [31:0] _0719_;
wire [31:0] _0720_;
wire [6:0] _0721_;
wire [6:0] _0722_;
wire [6:0] _0723_;
wire [6:0] _0724_;
wire [6:0] _0725_;
wire [6:0] _0726_;
wire [31:0] _0727_;
wire [31:0] _0728_;
wire [31:0] _0729_;
wire [31:0] _0730_;
wire [31:0] _0731_;
wire [31:0] _0732_;
wire [6:0] _0733_;
wire [6:0] _0734_;
wire [1:0] _0735_;
wire [1:0] _0736_;
wire [1:0] _0737_;
wire [1:0] _0738_;
wire [1:0] _0739_;
wire [1:0] _0740_;
wire _0741_;
wire _0742_;
wire [1:0] _0743_;
wire [1:0] _0744_;
wire [1:0] _0745_;
wire [1:0] _0746_;
wire _0747_;
wire _0748_;
wire [1:0] _0749_;
wire [1:0] _0750_;
wire [7:0] _0751_;
wire [7:0] _0752_;
wire [7:0] _0753_;
wire [7:0] _0754_;
wire [31:0] _0755_;
wire [31:0] _0756_;
wire _0757_;
wire _0758_;
wire [5:0] _0759_;
wire [5:0] _0760_;
wire [31:0] _0761_;
wire [31:0] _0762_;
wire [1:0] _0763_;
wire [1:0] _0764_;
wire [63:0] _0765_;
wire [63:0] _0766_;
wire _0767_;
wire _0768_;
wire _0769_;
wire _0770_;
wire _0771_;
wire _0772_;
wire _0773_;
wire _0774_;
wire _0775_;
wire _0776_;
wire _0777_;
wire _0778_;
wire _0779_;
wire [31:0] _0780_;
wire [17:0] _0781_;
wire _0782_;
wire _0783_;
wire [1:0] _0784_;
wire [1:0] _0785_;
wire _0786_;
wire [31:0] _0787_;
wire _0788_;
wire _0789_;
wire _0790_;
wire [31:0] _0791_;
/* cellift = 32'd1 */
wire [31:0] _0792_;
wire _0793_;
/* cellift = 32'd1 */
wire _0794_;
wire _0795_;
/* cellift = 32'd1 */
wire _0796_;
wire _0797_;
/* cellift = 32'd1 */
wire _0798_;
wire _0799_;
/* cellift = 32'd1 */
wire _0800_;
wire _0801_;
/* cellift = 32'd1 */
wire _0802_;
wire _0803_;
/* cellift = 32'd1 */
wire _0804_;
wire _0805_;
/* cellift = 32'd1 */
wire _0806_;
wire _0807_;
/* cellift = 32'd1 */
wire _0808_;
wire _0809_;
/* cellift = 32'd1 */
wire _0810_;
wire _0811_;
/* cellift = 32'd1 */
wire _0812_;
wire _0813_;
/* cellift = 32'd1 */
wire _0814_;
wire _0815_;
/* cellift = 32'd1 */
wire _0816_;
wire _0817_;
/* cellift = 32'd1 */
wire _0818_;
wire _0819_;
/* cellift = 32'd1 */
wire _0820_;
wire _0821_;
/* cellift = 32'd1 */
wire _0822_;
wire _0823_;
/* cellift = 32'd1 */
wire _0824_;
wire _0825_;
/* cellift = 32'd1 */
wire _0826_;
wire _0827_;
/* cellift = 32'd1 */
wire _0828_;
wire _0829_;
/* cellift = 32'd1 */
wire _0830_;
wire _0831_;
/* cellift = 32'd1 */
wire _0832_;
wire _0833_;
/* cellift = 32'd1 */
wire _0834_;
wire _0835_;
/* cellift = 32'd1 */
wire _0836_;
wire _0837_;
/* cellift = 32'd1 */
wire _0838_;
wire _0839_;
/* cellift = 32'd1 */
wire _0840_;
wire _0841_;
/* cellift = 32'd1 */
wire _0842_;
wire _0843_;
/* cellift = 32'd1 */
wire _0844_;
wire _0845_;
/* cellift = 32'd1 */
wire _0846_;
wire _0847_;
/* cellift = 32'd1 */
wire _0848_;
wire [2:0] _0849_;
/* cellift = 32'd1 */
wire [2:0] _0850_;
wire [2:0] _0851_;
/* cellift = 32'd1 */
wire [2:0] _0852_;
wire [2:0] _0853_;
/* cellift = 32'd1 */
wire [2:0] _0854_;
wire [2:0] _0855_;
/* cellift = 32'd1 */
wire [2:0] _0856_;
wire [2:0] _0857_;
/* cellift = 32'd1 */
wire [2:0] _0858_;
wire [2:0] _0859_;
/* cellift = 32'd1 */
wire [2:0] _0860_;
wire [2:0] _0861_;
/* cellift = 32'd1 */
wire [2:0] _0862_;
wire [2:0] _0863_;
/* cellift = 32'd1 */
wire [2:0] _0864_;
wire [2:0] _0865_;
/* cellift = 32'd1 */
wire [2:0] _0866_;
wire [2:0] _0867_;
/* cellift = 32'd1 */
wire [2:0] _0868_;
wire [2:0] _0869_;
/* cellift = 32'd1 */
wire [2:0] _0870_;
wire [2:0] _0871_;
wire [2:0] _0872_;
/* cellift = 32'd1 */
wire [2:0] _0873_;
wire [2:0] _0874_;
/* cellift = 32'd1 */
wire [2:0] _0875_;
wire _0876_;
/* cellift = 32'd1 */
wire _0877_;
wire _0878_;
/* cellift = 32'd1 */
wire _0879_;
wire _0880_;
/* cellift = 32'd1 */
wire _0881_;
wire _0882_;
/* cellift = 32'd1 */
wire _0883_;
wire _0884_;
/* cellift = 32'd1 */
wire _0885_;
wire _0886_;
/* cellift = 32'd1 */
wire _0887_;
wire _0888_;
/* cellift = 32'd1 */
wire _0889_;
wire _0890_;
/* cellift = 32'd1 */
wire _0891_;
wire _0892_;
/* cellift = 32'd1 */
wire _0893_;
wire _0894_;
/* cellift = 32'd1 */
wire _0895_;
wire _0896_;
/* cellift = 32'd1 */
wire _0897_;
wire _0898_;
/* cellift = 32'd1 */
wire _0899_;
wire _0900_;
/* cellift = 32'd1 */
wire _0901_;
wire _0902_;
/* cellift = 32'd1 */
wire _0903_;
wire _0904_;
/* cellift = 32'd1 */
wire _0905_;
wire _0906_;
/* cellift = 32'd1 */
wire _0907_;
wire [2:0] _0908_;
/* cellift = 32'd1 */
wire [2:0] _0909_;
wire [2:0] _0910_;
/* cellift = 32'd1 */
wire [2:0] _0911_;
wire [2:0] _0912_;
/* cellift = 32'd1 */
wire [2:0] _0913_;
wire [2:0] _0914_;
/* cellift = 32'd1 */
wire [2:0] _0915_;
wire [2:0] _0916_;
/* cellift = 32'd1 */
wire [2:0] _0917_;
wire [2:0] _0918_;
/* cellift = 32'd1 */
wire [2:0] _0919_;
wire [2:0] _0920_;
/* cellift = 32'd1 */
wire [2:0] _0921_;
wire [2:0] _0922_;
/* cellift = 32'd1 */
wire [2:0] _0923_;
wire [2:0] _0924_;
/* cellift = 32'd1 */
wire [2:0] _0925_;
wire [2:0] _0926_;
/* cellift = 32'd1 */
wire [2:0] _0927_;
wire [2:0] _0928_;
/* cellift = 32'd1 */
wire [2:0] _0929_;
wire [2:0] _0930_;
/* cellift = 32'd1 */
wire [2:0] _0931_;
wire [2:0] _0932_;
wire [2:0] _0933_;
/* cellift = 32'd1 */
wire [2:0] _0934_;
wire [2:0] _0935_;
/* cellift = 32'd1 */
wire [2:0] _0936_;
wire [2:0] _0937_;
/* cellift = 32'd1 */
wire [2:0] _0938_;
wire [2:0] _0939_;
/* cellift = 32'd1 */
wire [2:0] _0940_;
wire [2:0] _0941_;
/* cellift = 32'd1 */
wire [2:0] _0942_;
wire [2:0] _0943_;
/* cellift = 32'd1 */
wire [2:0] _0944_;
wire [2:0] _0945_;
/* cellift = 32'd1 */
wire [2:0] _0946_;
wire [2:0] _0947_;
/* cellift = 32'd1 */
wire [2:0] _0948_;
wire [2:0] _0949_;
/* cellift = 32'd1 */
wire [2:0] _0950_;
wire [2:0] _0951_;
/* cellift = 32'd1 */
wire [2:0] _0952_;
wire [2:0] _0953_;
/* cellift = 32'd1 */
wire [2:0] _0954_;
wire [2:0] _0955_;
/* cellift = 32'd1 */
wire [2:0] _0956_;
wire [2:0] _0957_;
/* cellift = 32'd1 */
wire [2:0] _0958_;
wire [2:0] _0959_;
/* cellift = 32'd1 */
wire [2:0] _0960_;
wire [2:0] _0961_;
/* cellift = 32'd1 */
wire [2:0] _0962_;
wire [2:0] _0963_;
/* cellift = 32'd1 */
wire [2:0] _0964_;
wire [2:0] _0965_;
/* cellift = 32'd1 */
wire [2:0] _0966_;
wire [2:0] _0967_;
/* cellift = 32'd1 */
wire [2:0] _0968_;
wire [2:0] _0969_;
/* cellift = 32'd1 */
wire [2:0] _0970_;
wire [2:0] _0971_;
/* cellift = 32'd1 */
wire [2:0] _0972_;
wire [2:0] _0973_;
/* cellift = 32'd1 */
wire [2:0] _0974_;
wire [2:0] _0975_;
/* cellift = 32'd1 */
wire [2:0] _0976_;
wire [2:0] _0977_;
/* cellift = 32'd1 */
wire [2:0] _0978_;
wire [2:0] _0979_;
/* cellift = 32'd1 */
wire [2:0] _0980_;
wire [2:0] _0981_;
/* cellift = 32'd1 */
wire [2:0] _0982_;
wire [2:0] _0983_;
/* cellift = 32'd1 */
wire [2:0] _0984_;
wire [2:0] _0985_;
/* cellift = 32'd1 */
wire [2:0] _0986_;
wire [2:0] _0987_;
/* cellift = 32'd1 */
wire [2:0] _0988_;
wire [2:0] _0989_;
/* cellift = 32'd1 */
wire [2:0] _0990_;
wire [2:0] _0991_;
/* cellift = 32'd1 */
wire [2:0] _0992_;
wire [2:0] _0993_;
/* cellift = 32'd1 */
wire [2:0] _0994_;
wire _0995_;
/* cellift = 32'd1 */
wire _0996_;
wire _0997_;
/* cellift = 32'd1 */
wire _0998_;
wire _0999_;
/* cellift = 32'd1 */
wire _1000_;
wire _1001_;
/* cellift = 32'd1 */
wire _1002_;
wire _1003_;
/* cellift = 32'd1 */
wire _1004_;
wire _1005_;
/* cellift = 32'd1 */
wire _1006_;
wire _1007_;
/* cellift = 32'd1 */
wire _1008_;
wire _1009_;
/* cellift = 32'd1 */
wire _1010_;
wire _1011_;
/* cellift = 32'd1 */
wire _1012_;
wire _1013_;
/* cellift = 32'd1 */
wire _1014_;
wire _1015_;
/* cellift = 32'd1 */
wire _1016_;
wire _1017_;
/* cellift = 32'd1 */
wire _1018_;
wire _1019_;
/* cellift = 32'd1 */
wire _1020_;
wire _1021_;
/* cellift = 32'd1 */
wire _1022_;
wire _1023_;
/* cellift = 32'd1 */
wire _1024_;
wire _1025_;
/* cellift = 32'd1 */
wire _1026_;
wire _1027_;
/* cellift = 32'd1 */
wire _1028_;
wire _1029_;
/* cellift = 32'd1 */
wire _1030_;
wire _1031_;
/* cellift = 32'd1 */
wire _1032_;
wire _1033_;
/* cellift = 32'd1 */
wire _1034_;
wire _1035_;
/* cellift = 32'd1 */
wire _1036_;
wire _1037_;
/* cellift = 32'd1 */
wire _1038_;
wire _1039_;
/* cellift = 32'd1 */
wire _1040_;
wire _1041_;
/* cellift = 32'd1 */
wire _1042_;
wire _1043_;
/* cellift = 32'd1 */
wire _1044_;
wire _1045_;
/* cellift = 32'd1 */
wire _1046_;
wire _1047_;
/* cellift = 32'd1 */
wire _1048_;
wire _1049_;
/* cellift = 32'd1 */
wire _1050_;
wire _1051_;
/* cellift = 32'd1 */
wire _1052_;
wire [2:0] _1053_;
/* cellift = 32'd1 */
wire [2:0] _1054_;
wire [2:0] _1055_;
/* cellift = 32'd1 */
wire [2:0] _1056_;
wire [2:0] _1057_;
/* cellift = 32'd1 */
wire [2:0] _1058_;
wire [2:0] _1059_;
/* cellift = 32'd1 */
wire [2:0] _1060_;
wire [2:0] _1061_;
/* cellift = 32'd1 */
wire [2:0] _1062_;
wire [2:0] _1063_;
/* cellift = 32'd1 */
wire [2:0] _1064_;
wire [2:0] _1065_;
/* cellift = 32'd1 */
wire [2:0] _1066_;
wire [2:0] _1067_;
/* cellift = 32'd1 */
wire [2:0] _1068_;
wire [2:0] _1069_;
/* cellift = 32'd1 */
wire [2:0] _1070_;
wire [2:0] _1071_;
/* cellift = 32'd1 */
wire [2:0] _1072_;
wire [2:0] _1073_;
/* cellift = 32'd1 */
wire [2:0] _1074_;
wire [2:0] _1075_;
/* cellift = 32'd1 */
wire [2:0] _1076_;
wire _1077_;
/* cellift = 32'd1 */
wire _1078_;
wire _1079_;
/* cellift = 32'd1 */
wire _1080_;
wire _1081_;
/* cellift = 32'd1 */
wire _1082_;
wire _1083_;
/* cellift = 32'd1 */
wire _1084_;
wire _1085_;
/* cellift = 32'd1 */
wire _1086_;
wire _1087_;
/* cellift = 32'd1 */
wire _1088_;
wire _1089_;
/* cellift = 32'd1 */
wire _1090_;
wire _1091_;
/* cellift = 32'd1 */
wire _1092_;
wire _1093_;
/* cellift = 32'd1 */
wire _1094_;
wire _1095_;
/* cellift = 32'd1 */
wire _1096_;
wire _1097_;
/* cellift = 32'd1 */
wire _1098_;
wire _1099_;
/* cellift = 32'd1 */
wire _1100_;
wire _1101_;
/* cellift = 32'd1 */
wire _1102_;
wire _1103_;
/* cellift = 32'd1 */
wire _1104_;
wire [8:0] _1105_;
/* cellift = 32'd1 */
wire [8:0] _1106_;
wire [8:0] _1107_;
/* cellift = 32'd1 */
wire [8:0] _1108_;
wire [8:0] _1109_;
/* cellift = 32'd1 */
wire [8:0] _1110_;
wire [8:0] _1111_;
/* cellift = 32'd1 */
wire [8:0] _1112_;
wire [8:0] _1113_;
/* cellift = 32'd1 */
wire [8:0] _1114_;
wire [8:0] _1115_;
/* cellift = 32'd1 */
wire [8:0] _1116_;
wire [8:0] _1117_;
/* cellift = 32'd1 */
wire [8:0] _1118_;
wire [8:0] _1119_;
/* cellift = 32'd1 */
wire [8:0] _1120_;
wire [8:0] _1121_;
/* cellift = 32'd1 */
wire [8:0] _1122_;
wire [8:0] _1123_;
/* cellift = 32'd1 */
wire [8:0] _1124_;
wire [8:0] _1125_;
/* cellift = 32'd1 */
wire [8:0] _1126_;
wire [8:0] _1127_;
/* cellift = 32'd1 */
wire [8:0] _1128_;
wire [8:0] _1129_;
/* cellift = 32'd1 */
wire [8:0] _1130_;
wire [8:0] _1131_;
/* cellift = 32'd1 */
wire [8:0] _1132_;
wire [8:0] _1133_;
/* cellift = 32'd1 */
wire [8:0] _1134_;
wire _1135_;
/* cellift = 32'd1 */
wire _1136_;
wire _1137_;
/* cellift = 32'd1 */
wire _1138_;
wire _1139_;
/* cellift = 32'd1 */
wire _1140_;
wire _1141_;
/* cellift = 32'd1 */
wire _1142_;
wire _1143_;
/* cellift = 32'd1 */
wire _1144_;
wire _1145_;
/* cellift = 32'd1 */
wire _1146_;
wire _1147_;
/* cellift = 32'd1 */
wire _1148_;
wire _1149_;
/* cellift = 32'd1 */
wire _1150_;
wire _1151_;
/* cellift = 32'd1 */
wire _1152_;
wire _1153_;
/* cellift = 32'd1 */
wire _1154_;
wire _1155_;
/* cellift = 32'd1 */
wire _1156_;
wire _1157_;
/* cellift = 32'd1 */
wire _1158_;
wire _1159_;
/* cellift = 32'd1 */
wire _1160_;
wire _1161_;
/* cellift = 32'd1 */
wire _1162_;
wire _1163_;
/* cellift = 32'd1 */
wire _1164_;
wire [63:0] _1165_;
/* cellift = 32'd1 */
wire [63:0] _1166_;
wire _1167_;
/* cellift = 32'd1 */
wire _1168_;
wire _1169_;
/* cellift = 32'd1 */
wire _1170_;
wire _1171_;
/* cellift = 32'd1 */
wire _1172_;
wire _1173_;
/* cellift = 32'd1 */
wire _1174_;
wire _1175_;
/* cellift = 32'd1 */
wire _1176_;
wire _1177_;
/* cellift = 32'd1 */
wire _1178_;
wire _1179_;
/* cellift = 32'd1 */
wire _1180_;
wire _1181_;
/* cellift = 32'd1 */
wire _1182_;
wire _1183_;
/* cellift = 32'd1 */
wire _1184_;
wire _1185_;
/* cellift = 32'd1 */
wire _1186_;
wire _1187_;
/* cellift = 32'd1 */
wire _1188_;
wire _1189_;
/* cellift = 32'd1 */
wire _1190_;
wire _1191_;
/* cellift = 32'd1 */
wire _1192_;
wire _1193_;
/* cellift = 32'd1 */
wire _1194_;
wire _1195_;
/* cellift = 32'd1 */
wire _1196_;
/* src = "generated/sv2v_out.v:14000.30-14000.54" */
wire _1197_;
/* src = "generated/sv2v_out.v:14152.409-14152.428" */
wire _1198_;
/* src = "generated/sv2v_out.v:14152.388-14152.407" */
wire _1199_;
/* src = "generated/sv2v_out.v:14152.367-14152.386" */
wire _1200_;
/* src = "generated/sv2v_out.v:14152.346-14152.365" */
wire _1201_;
/* src = "generated/sv2v_out.v:14152.325-14152.344" */
wire _1202_;
/* src = "generated/sv2v_out.v:14152.304-14152.323" */
wire _1203_;
/* src = "generated/sv2v_out.v:14152.283-14152.302" */
wire _1204_;
/* src = "generated/sv2v_out.v:14152.262-14152.281" */
wire _1205_;
/* src = "generated/sv2v_out.v:14152.241-14152.260" */
wire _1206_;
/* src = "generated/sv2v_out.v:14152.220-14152.239" */
wire _1207_;
/* src = "generated/sv2v_out.v:14152.199-14152.218" */
wire _1208_;
/* src = "generated/sv2v_out.v:14152.178-14152.197" */
wire _1209_;
/* src = "generated/sv2v_out.v:14152.157-14152.176" */
wire _1210_;
/* src = "generated/sv2v_out.v:14152.136-14152.155" */
wire _1211_;
/* src = "generated/sv2v_out.v:14152.115-14152.134" */
wire _1212_;
/* src = "generated/sv2v_out.v:14152.94-14152.113" */
wire _1213_;
/* src = "generated/sv2v_out.v:14152.73-14152.92" */
wire _1214_;
/* src = "generated/sv2v_out.v:14152.52-14152.71" */
wire _1215_;
/* src = "generated/sv2v_out.v:14152.31-14152.50" */
wire _1216_;
/* src = "generated/sv2v_out.v:14152.10-14152.29" */
wire _1217_;
/* src = "generated/sv2v_out.v:14169.46-14169.75" */
wire _1218_;
/* src = "generated/sv2v_out.v:14169.15-14169.44" */
wire _1219_;
/* src = "generated/sv2v_out.v:14314.56-14314.72" */
wire _1220_;
/* src = "generated/sv2v_out.v:14314.38-14314.54" */
wire _1221_;
/* src = "generated/sv2v_out.v:14314.20-14314.36" */
wire _1222_;
/* src = "generated/sv2v_out.v:14866.50-14866.69" */
wire _1223_;
/* src = "generated/sv2v_out.v:14196.10-14196.66" */
wire _1224_;
/* src = "generated/sv2v_out.v:14208.10-14208.60" */
wire _1225_;
/* src = "generated/sv2v_out.v:14263.12-14263.38" */
wire _1226_;
/* src = "generated/sv2v_out.v:14196.11-14196.35" */
wire _1227_;
/* src = "generated/sv2v_out.v:14196.41-14196.65" */
wire _1228_;
/* src = "generated/sv2v_out.v:14208.11-14208.32" */
wire _1229_;
/* src = "generated/sv2v_out.v:14208.38-14208.59" */
wire _1230_;
/* src = "generated/sv2v_out.v:14278.9-14278.33" */
wire _1231_;
/* src = "generated/sv2v_out.v:0.0-0.0" */
wire [31:0] _1232_;
/* src = "generated/sv2v_out.v:14315.47-14315.66" */
wire _1233_;
/* src = "generated/sv2v_out.v:14699.40-14699.57" */
wire _1234_;
/* src = "generated/sv2v_out.v:14910.50-14910.89" */
wire _1235_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14910.50-14910.89" */
wire _1236_;
/* src = "generated/sv2v_out.v:0.0-0.0" */
wire [31:0] _1237_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:0.0-0.0" */
wire [31:0] _1238_;
/* src = "generated/sv2v_out.v:14001.48-14001.79" */
wire _1239_;
/* src = "generated/sv2v_out.v:14001.47-14001.99" */
wire _1240_;
/* src = "generated/sv2v_out.v:14001.46-14001.118" */
wire _1241_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14001.46-14001.118" */
wire _1242_;
/* src = "generated/sv2v_out.v:14056.30-14056.55" */
wire _1243_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14056.30-14056.55" */
wire _1244_;
/* src = "generated/sv2v_out.v:14309.26-14309.51" */
wire [31:0] _1245_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14309.26-14309.51" */
wire [31:0] _1246_;
/* src = "generated/sv2v_out.v:14910.52-14910.88" */
wire _1247_;
/* src = "generated/sv2v_out.v:14923.31-14923.54" */
wire _1248_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14923.31-14923.54" */
wire _1249_;
wire _1250_;
wire [2:0] _1251_;
/* cellift = 32'd1 */
wire [2:0] _1252_;
wire [2:0] _1253_;
/* cellift = 32'd1 */
wire [2:0] _1254_;
wire _1255_;
/* cellift = 32'd1 */
wire _1256_;
wire _1257_;
/* cellift = 32'd1 */
wire _1258_;
wire _1259_;
/* cellift = 32'd1 */
wire _1260_;
wire _1261_;
/* cellift = 32'd1 */
wire _1262_;
wire [31:0] _1263_;
/* cellift = 32'd1 */
wire [31:0] _1264_;
wire [31:0] _1265_;
/* cellift = 32'd1 */
wire [31:0] _1266_;
wire _1267_;
wire _1268_;
wire _1269_;
/* cellift = 32'd1 */
wire _1270_;
wire _1271_;
/* cellift = 32'd1 */
wire _1272_;
wire _1273_;
wire _1274_;
wire [6:0] _1275_;
/* cellift = 32'd1 */
wire [6:0] _1276_;
wire [6:0] _1277_;
/* cellift = 32'd1 */
wire [6:0] _1278_;
wire _1279_;
wire _1280_;
wire [31:0] _1281_;
/* cellift = 32'd1 */
wire [31:0] _1282_;
wire [31:0] _1283_;
/* cellift = 32'd1 */
wire [31:0] _1284_;
wire _1285_;
wire _1286_;
wire [1:0] _1287_;
/* cellift = 32'd1 */
wire [1:0] _1288_;
wire [1:0] _1289_;
/* cellift = 32'd1 */
wire [1:0] _1290_;
wire _1291_;
wire _1292_;
wire [30:0] _1293_;
wire _1294_;
wire [30:0] _1295_;
wire _1296_;
wire _1297_;
wire _1298_;
wire _1299_;
wire _1300_;
wire _1301_;
wire _1302_;
wire _1303_;
wire _1304_;
wire _1305_;
wire _1306_;
wire _1307_;
wire _1308_;
wire [28:0] _1309_;
wire _1310_;
wire _1311_;
wire _1312_;
wire _1313_;
wire _1314_;
wire _1315_;
wire _1316_;
wire _1317_;
wire _1318_;
wire _1319_;
wire _1320_;
wire _1321_;
wire _1322_;
wire _1323_;
wire _1324_;
wire _1325_;
wire _1326_;
wire _1327_;
wire _1328_;
wire _1329_;
wire _1330_;
wire _1331_;
wire _1332_;
wire _1333_;
wire _1334_;
wire _1335_;
wire _1336_;
wire _1337_;
wire _1338_;
wire _1339_;
wire _1340_;
wire _1341_;
wire _1342_;
wire _1343_;
wire _1344_;
wire _1345_;
wire _1346_;
wire _1347_;
wire [1:0] _1348_;
wire _1349_;
wire _1350_;
wire _1351_;
wire _1352_;
/* src = "generated/sv2v_out.v:14056.58-14056.116" */
wire [25:0] _1353_;
/* src = "generated/sv2v_out.v:13820.20-13820.31" */
input [31:0] boot_addr_i;
wire [31:0] boot_addr_i;
/* cellift = 32'd1 */
input [31:0] boot_addr_i_t0;
wire [31:0] boot_addr_i_t0;
/* src = "generated/sv2v_out.v:13876.13-13876.21" */
input branch_i;
wire branch_i;
/* cellift = 32'd1 */
input branch_i_t0;
wire branch_i_t0;
/* src = "generated/sv2v_out.v:13877.13-13877.27" */
input branch_taken_i;
wire branch_taken_i;
/* cellift = 32'd1 */
input branch_taken_i_t0;
wire branch_taken_i_t0;
/* src = "generated/sv2v_out.v:13812.13-13812.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:13975.12-13975.29" */
wire [7:0] cpuctrlsts_part_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13975.12-13975.29" */
wire [7:0] cpuctrlsts_part_d_t0;
/* src = "generated/sv2v_out.v:13979.7-13979.26" */
wire cpuctrlsts_part_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13979.7-13979.26" */
wire cpuctrlsts_part_err_t0;
/* src = "generated/sv2v_out.v:13974.13-13974.30" */
wire [7:0] cpuctrlsts_part_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13974.13-13974.30" */
wire [7:0] cpuctrlsts_part_q_t0;
/* src = "generated/sv2v_out.v:13978.6-13978.24" */
wire cpuctrlsts_part_we;
/* src = "generated/sv2v_out.v:13821.13-13821.25" */
input csr_access_i;
wire csr_access_i;
/* cellift = 32'd1 */
input csr_access_i_t0;
wire csr_access_i_t0;
/* src = "generated/sv2v_out.v:13822.20-13822.30" */
input [11:0] csr_addr_i;
wire [11:0] csr_addr_i;
/* cellift = 32'd1 */
input [11:0] csr_addr_i_t0;
wire [11:0] csr_addr_i_t0;
/* src = "generated/sv2v_out.v:13844.21-13844.31" */
output [31:0] csr_depc_o;
wire [31:0] csr_depc_o;
/* cellift = 32'd1 */
output [31:0] csr_depc_o_t0;
wire [31:0] csr_depc_o_t0;
/* src = "generated/sv2v_out.v:13866.19-13866.31" */
input [6:0] csr_mcause_i;
wire [6:0] csr_mcause_i;
/* cellift = 32'd1 */
input [6:0] csr_mcause_i_t0;
wire [6:0] csr_mcause_i_t0;
/* src = "generated/sv2v_out.v:13835.21-13835.31" */
output [31:0] csr_mepc_o;
wire [31:0] csr_mepc_o;
/* cellift = 32'd1 */
output [31:0] csr_mepc_o_t0;
wire [31:0] csr_mepc_o_t0;
/* src = "generated/sv2v_out.v:13834.14-13834.31" */
output csr_mstatus_mie_o;
wire csr_mstatus_mie_o;
/* cellift = 32'd1 */
output csr_mstatus_mie_o_t0;
wire csr_mstatus_mie_o_t0;
/* src = "generated/sv2v_out.v:13817.14-13817.30" */
output csr_mstatus_tw_o;
wire csr_mstatus_tw_o;
/* cellift = 32'd1 */
output csr_mstatus_tw_o_t0;
wire csr_mstatus_tw_o_t0;
/* src = "generated/sv2v_out.v:13867.20-13867.31" */
input [31:0] csr_mtval_i;
wire [31:0] csr_mtval_i;
/* cellift = 32'd1 */
input [31:0] csr_mtval_i_t0;
wire [31:0] csr_mtval_i_t0;
/* src = "generated/sv2v_out.v:13836.21-13836.32" */
output [31:0] csr_mtval_o;
wire [31:0] csr_mtval_o;
/* cellift = 32'd1 */
output [31:0] csr_mtval_o_t0;
wire [31:0] csr_mtval_o_t0;
/* src = "generated/sv2v_out.v:13819.13-13819.29" */
input csr_mtvec_init_i;
wire csr_mtvec_init_i;
/* cellift = 32'd1 */
input csr_mtvec_init_i_t0;
wire csr_mtvec_init_i_t0;
/* src = "generated/sv2v_out.v:13818.21-13818.32" */
output [31:0] csr_mtvec_o;
wire [31:0] csr_mtvec_o;
/* cellift = 32'd1 */
output [31:0] csr_mtvec_o_t0;
wire [31:0] csr_mtvec_o_t0;
/* src = "generated/sv2v_out.v:13825.8-13825.19" */
input csr_op_en_i;
wire csr_op_en_i;
/* cellift = 32'd1 */
input csr_op_en_i_t0;
wire csr_op_en_i_t0;
/* src = "generated/sv2v_out.v:13824.19-13824.27" */
input [1:0] csr_op_i;
wire [1:0] csr_op_i;
/* cellift = 32'd1 */
input [1:0] csr_op_i_t0;
wire [1:0] csr_op_i_t0;
/* src = "generated/sv2v_out.v:13838.43-13838.57" */
output [135:0] csr_pmp_addr_o;
wire [135:0] csr_pmp_addr_o;
/* cellift = 32'd1 */
output [135:0] csr_pmp_addr_o_t0;
wire [135:0] csr_pmp_addr_o_t0;
/* src = "generated/sv2v_out.v:13837.42-13837.55" */
output [23:0] csr_pmp_cfg_o;
wire [23:0] csr_pmp_cfg_o;
/* cellift = 32'd1 */
output [23:0] csr_pmp_cfg_o_t0;
wire [23:0] csr_pmp_cfg_o_t0;
/* src = "generated/sv2v_out.v:13839.20-13839.37" */
output [2:0] csr_pmp_mseccfg_o;
wire [2:0] csr_pmp_mseccfg_o;
/* cellift = 32'd1 */
output [2:0] csr_pmp_mseccfg_o_t0;
wire [2:0] csr_pmp_mseccfg_o_t0;
/* src = "generated/sv2v_out.v:13826.21-13826.32" */
output [31:0] csr_rdata_o;
wire [31:0] csr_rdata_o;
/* cellift = 32'd1 */
output [31:0] csr_rdata_o_t0;
wire [31:0] csr_rdata_o_t0;
/* src = "generated/sv2v_out.v:13864.13-13864.31" */
input csr_restore_dret_i;
wire csr_restore_dret_i;
/* cellift = 32'd1 */
input csr_restore_dret_i_t0;
wire csr_restore_dret_i_t0;
/* src = "generated/sv2v_out.v:13863.13-13863.31" */
input csr_restore_mret_i;
wire csr_restore_mret_i;
/* cellift = 32'd1 */
input csr_restore_mret_i_t0;
wire csr_restore_mret_i_t0;
/* src = "generated/sv2v_out.v:13865.13-13865.29" */
input csr_save_cause_i;
wire csr_save_cause_i;
/* cellift = 32'd1 */
input csr_save_cause_i_t0;
wire csr_save_cause_i_t0;
/* src = "generated/sv2v_out.v:13861.13-13861.26" */
input csr_save_id_i;
wire csr_save_id_i;
/* cellift = 32'd1 */
input csr_save_id_i_t0;
wire csr_save_id_i_t0;
/* src = "generated/sv2v_out.v:13860.13-13860.26" */
input csr_save_if_i;
wire csr_save_if_i;
/* cellift = 32'd1 */
input csr_save_if_i_t0;
wire csr_save_if_i_t0;
/* src = "generated/sv2v_out.v:13862.13-13862.26" */
input csr_save_wb_i;
wire csr_save_wb_i;
/* cellift = 32'd1 */
input csr_save_wb_i_t0;
wire csr_save_wb_i_t0;
/* src = "generated/sv2v_out.v:13858.14-13858.30" */
output csr_shadow_err_o;
wire csr_shadow_err_o;
/* cellift = 32'd1 */
output csr_shadow_err_o_t0;
wire csr_shadow_err_o_t0;
/* src = "generated/sv2v_out.v:13823.20-13823.31" */
input [31:0] csr_wdata_i;
wire [31:0] csr_wdata_i;
/* cellift = 32'd1 */
input [31:0] csr_wdata_i_t0;
wire [31:0] csr_wdata_i_t0;
/* src = "generated/sv2v_out.v:13984.7-13984.17" */
wire csr_we_int;
/* src = "generated/sv2v_out.v:13985.7-13985.13" */
wire csr_wr;
/* src = "generated/sv2v_out.v:13852.14-13852.31" */
output data_ind_timing_o;
wire data_ind_timing_o;
/* cellift = 32'd1 */
output data_ind_timing_o_t0;
wire data_ind_timing_o_t0;
/* src = "generated/sv2v_out.v:13986.6-13986.13" */
wire dbg_csr;
/* src = "generated/sv2v_out.v:13934.13-13934.19" */
wire [31:0] dcsr_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13934.13-13934.19" */
wire [31:0] dcsr_d_t0;
/* src = "generated/sv2v_out.v:13935.6-13935.13" */
wire dcsr_en;
/* src = "generated/sv2v_out.v:13933.14-13933.20" */
wire [31:0] dcsr_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13933.14-13933.20" */
wire [31:0] dcsr_q_t0;
/* src = "generated/sv2v_out.v:13842.19-13842.32" */
input [2:0] debug_cause_i;
wire [2:0] debug_cause_i;
/* cellift = 32'd1 */
input [2:0] debug_cause_i_t0;
wire [2:0] debug_cause_i_t0;
/* src = "generated/sv2v_out.v:13843.13-13843.29" */
input debug_csr_save_i;
wire debug_csr_save_i;
/* cellift = 32'd1 */
input debug_csr_save_i_t0;
wire debug_csr_save_i_t0;
/* src = "generated/sv2v_out.v:13846.14-13846.29" */
output debug_ebreakm_o;
wire debug_ebreakm_o;
/* cellift = 32'd1 */
output debug_ebreakm_o_t0;
wire debug_ebreakm_o_t0;
/* src = "generated/sv2v_out.v:13847.14-13847.29" */
output debug_ebreaku_o;
wire debug_ebreaku_o;
/* cellift = 32'd1 */
output debug_ebreaku_o_t0;
wire debug_ebreaku_o_t0;
/* src = "generated/sv2v_out.v:13841.13-13841.34" */
input debug_mode_entering_i;
wire debug_mode_entering_i;
/* cellift = 32'd1 */
input debug_mode_entering_i_t0;
wire debug_mode_entering_i_t0;
/* src = "generated/sv2v_out.v:13840.13-13840.25" */
input debug_mode_i;
wire debug_mode_i;
/* cellift = 32'd1 */
input debug_mode_i_t0;
wire debug_mode_i_t0;
/* src = "generated/sv2v_out.v:13845.14-13845.33" */
output debug_single_step_o;
wire debug_single_step_o;
/* cellift = 32'd1 */
output debug_single_step_o_t0;
wire debug_single_step_o_t0;
/* src = "generated/sv2v_out.v:13937.13-13937.19" */
wire [31:0] depc_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13937.13-13937.19" */
wire [31:0] depc_d_t0;
/* src = "generated/sv2v_out.v:13938.6-13938.13" */
wire depc_en;
/* src = "generated/sv2v_out.v:13882.13-13882.23" */
input div_wait_i;
wire div_wait_i;
/* cellift = 32'd1 */
input div_wait_i_t0;
wire div_wait_i_t0;
/* src = "generated/sv2v_out.v:13869.13-13869.32" */
output double_fault_seen_o;
wire double_fault_seen_o;
/* cellift = 32'd1 */
output double_fault_seen_o_t0;
wire double_fault_seen_o_t0;
/* src = "generated/sv2v_out.v:13941.6-13941.18" */
wire dscratch0_en;
/* src = "generated/sv2v_out.v:13939.14-13939.25" */
wire [31:0] dscratch0_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13939.14-13939.25" */
wire [31:0] dscratch0_q_t0;
/* src = "generated/sv2v_out.v:13942.6-13942.18" */
wire dscratch1_en;
/* src = "generated/sv2v_out.v:13940.14-13940.25" */
wire [31:0] dscratch1_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13940.14-13940.25" */
wire [31:0] dscratch1_q_t0;
/* src = "generated/sv2v_out.v:13880.13-13880.25" */
input dside_wait_i;
wire dside_wait_i;
/* cellift = 32'd1 */
input dside_wait_i_t0;
wire dside_wait_i_t0;
/* src = "generated/sv2v_out.v:13853.14-13853.30" */
output dummy_instr_en_o;
wire dummy_instr_en_o;
/* cellift = 32'd1 */
output dummy_instr_en_o_t0;
wire dummy_instr_en_o_t0;
/* src = "generated/sv2v_out.v:13854.20-13854.38" */
output [2:0] dummy_instr_mask_o;
wire [2:0] dummy_instr_mask_o;
/* cellift = 32'd1 */
output [2:0] dummy_instr_mask_o_t0;
wire [2:0] dummy_instr_mask_o_t0;
/* src = "generated/sv2v_out.v:13855.14-13855.35" */
output dummy_instr_seed_en_o;
wire dummy_instr_seed_en_o;
/* cellift = 32'd1 */
output dummy_instr_seed_en_o_t0;
wire dummy_instr_seed_en_o_t0;
/* src = "generated/sv2v_out.v:13856.21-13856.39" */
output [31:0] dummy_instr_seed_o;
wire [31:0] dummy_instr_seed_o;
/* cellift = 32'd1 */
output [31:0] dummy_instr_seed_o_t0;
wire [31:0] dummy_instr_seed_o_t0;
/* src = "generated/sv2v_out.v:13814.20-13814.29" */
input [31:0] hart_id_i;
wire [31:0] hart_id_i;
/* cellift = 32'd1 */
input [31:0] hart_id_i_t0;
wire [31:0] hart_id_i_t0;
/* src = "generated/sv2v_out.v:13859.13-13859.31" */
input ic_scr_key_valid_i;
wire ic_scr_key_valid_i;
/* cellift = 32'd1 */
input ic_scr_key_valid_i_t0;
wire ic_scr_key_valid_i_t0;
/* src = "generated/sv2v_out.v:13857.14-13857.29" */
output icache_enable_o;
wire icache_enable_o;
/* cellift = 32'd1 */
output icache_enable_o_t0;
wire icache_enable_o_t0;
/* src = "generated/sv2v_out.v:13987.6-13987.17" */
wire illegal_csr;
/* src = "generated/sv2v_out.v:13989.7-13989.22" */
wire illegal_csr_dbg;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13989.7-13989.22" */
wire illegal_csr_dbg_t0;
/* src = "generated/sv2v_out.v:13868.14-13868.32" */
output illegal_csr_insn_o;
wire illegal_csr_insn_o;
/* cellift = 32'd1 */
output illegal_csr_insn_o_t0;
wire illegal_csr_insn_o_t0;
/* src = "generated/sv2v_out.v:13988.7-13988.23" */
wire illegal_csr_priv;
/* src = "generated/sv2v_out.v:13990.7-13990.24" */
wire illegal_csr_write;
/* src = "generated/sv2v_out.v:13871.13-13871.35" */
input instr_ret_compressed_i;
wire instr_ret_compressed_i;
/* cellift = 32'd1 */
input instr_ret_compressed_i_t0;
wire instr_ret_compressed_i_t0;
/* src = "generated/sv2v_out.v:13873.13-13873.40" */
input instr_ret_compressed_spec_i;
wire instr_ret_compressed_spec_i;
/* cellift = 32'd1 */
input instr_ret_compressed_spec_i_t0;
wire instr_ret_compressed_spec_i_t0;
/* src = "generated/sv2v_out.v:13870.13-13870.24" */
input instr_ret_i;
wire instr_ret_i;
/* cellift = 32'd1 */
input instr_ret_i_t0;
wire instr_ret_i_t0;
/* src = "generated/sv2v_out.v:13872.13-13872.29" */
input instr_ret_spec_i;
wire instr_ret_spec_i;
/* cellift = 32'd1 */
input instr_ret_spec_i_t0;
wire instr_ret_spec_i_t0;
/* src = "generated/sv2v_out.v:13829.13-13829.27" */
input irq_external_i;
wire irq_external_i;
/* cellift = 32'd1 */
input irq_external_i_t0;
wire irq_external_i_t0;
/* src = "generated/sv2v_out.v:13830.20-13830.30" */
input [14:0] irq_fast_i;
wire [14:0] irq_fast_i;
/* cellift = 32'd1 */
input [14:0] irq_fast_i_t0;
wire [14:0] irq_fast_i_t0;
/* src = "generated/sv2v_out.v:13832.14-13832.27" */
output irq_pending_o;
wire irq_pending_o;
/* cellift = 32'd1 */
output irq_pending_o_t0;
wire irq_pending_o_t0;
/* src = "generated/sv2v_out.v:13827.13-13827.27" */
input irq_software_i;
wire irq_software_i;
/* cellift = 32'd1 */
input irq_software_i_t0;
wire irq_software_i_t0;
/* src = "generated/sv2v_out.v:13828.13-13828.24" */
input irq_timer_i;
wire irq_timer_i;
/* cellift = 32'd1 */
input irq_timer_i_t0;
wire irq_timer_i_t0;
/* src = "generated/sv2v_out.v:13833.21-13833.27" */
output [17:0] irqs_o;
wire [17:0] irqs_o;
/* cellift = 32'd1 */
output [17:0] irqs_o_t0;
wire [17:0] irqs_o_t0;
/* src = "generated/sv2v_out.v:13874.13-13874.25" */
input iside_wait_i;
wire iside_wait_i;
/* cellift = 32'd1 */
input iside_wait_i_t0;
wire iside_wait_i_t0;
/* src = "generated/sv2v_out.v:13875.13-13875.19" */
input jump_i;
wire jump_i;
/* cellift = 32'd1 */
input jump_i_t0;
wire jump_i_t0;
/* src = "generated/sv2v_out.v:13923.12-13923.20" */
wire [6:0] mcause_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13923.12-13923.20" */
wire [6:0] mcause_d_t0;
/* src = "generated/sv2v_out.v:13924.6-13924.15" */
wire mcause_en;
/* src = "generated/sv2v_out.v:13922.13-13922.21" */
wire [6:0] mcause_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13922.13-13922.21" */
wire [6:0] mcause_q_t0;
/* src = "generated/sv2v_out.v:13956.14-13956.27" */
wire [31:0] mcountinhibit;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13956.14-13956.27" */
wire [31:0] mcountinhibit_t0;
/* src = "generated/sv2v_out.v:13959.6-13959.22" */
wire mcountinhibit_we;
/* src = "generated/sv2v_out.v:13878.13-13878.23" */
input mem_load_i;
wire mem_load_i;
/* cellift = 32'd1 */
input mem_load_i_t0;
wire mem_load_i_t0;
/* src = "generated/sv2v_out.v:13879.13-13879.24" */
input mem_store_i;
wire mem_store_i;
/* cellift = 32'd1 */
input mem_store_i_t0;
wire mem_store_i_t0;
/* src = "generated/sv2v_out.v:13920.13-13920.19" */
wire [31:0] mepc_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13920.13-13920.19" */
wire [31:0] mepc_d_t0;
/* src = "generated/sv2v_out.v:13921.6-13921.13" */
wire mepc_en;
/* src = "generated/sv2v_out.v:13960.14-13960.25" */
wire [63:0] \mhpmcounter[0] ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13960.14-13960.25" */
wire [63:0] \mhpmcounter[0]_t0 ;
/* src = "generated/sv2v_out.v:13960.14-13960.25" */
wire [63:0] \mhpmcounter[2] ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13960.14-13960.25" */
wire [63:0] \mhpmcounter[2]_t0 ;
/* src = "generated/sv2v_out.v:13961.13-13961.27" */
/* unused_bits = "1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] mhpmcounter_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13961.13-13961.27" */
/* unused_bits = "1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] mhpmcounter_we_t0;
/* src = "generated/sv2v_out.v:13962.13-13962.28" */
/* unused_bits = "1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] mhpmcounterh_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13962.13-13962.28" */
/* unused_bits = "1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] mhpmcounterh_we_t0;
/* src = "generated/sv2v_out.v:13916.6-13916.12" */
wire mie_en;
/* src = "generated/sv2v_out.v:13914.14-13914.19" */
wire [17:0] mie_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13914.14-13914.19" */
wire [17:0] mie_q_t0;
/* src = "generated/sv2v_out.v:13969.14-13969.27" */
wire [63:0] minstret_next;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13969.14-13969.27" */
wire [63:0] minstret_next_t0;
/* src = "generated/sv2v_out.v:13970.14-13970.26" */
wire [63:0] minstret_raw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13970.14-13970.26" */
wire [63:0] minstret_raw_t0;
/* src = "generated/sv2v_out.v:13918.6-13918.17" */
wire mscratch_en;
/* src = "generated/sv2v_out.v:13917.14-13917.24" */
wire [31:0] mscratch_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13917.14-13917.24" */
wire [31:0] mscratch_q_t0;
/* src = "generated/sv2v_out.v:13948.13-13948.27" */
wire [6:0] mstack_cause_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13948.13-13948.27" */
wire [6:0] mstack_cause_q_t0;
/* src = "generated/sv2v_out.v:13945.6-13945.15" */
wire mstack_en;
/* src = "generated/sv2v_out.v:13946.14-13946.26" */
wire [31:0] mstack_epc_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13946.14-13946.26" */
wire [31:0] mstack_epc_q_t0;
/* src = "generated/sv2v_out.v:13943.13-13943.21" */
wire [2:0] mstack_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13943.13-13943.21" */
wire [2:0] mstack_q_t0;
/* src = "generated/sv2v_out.v:13911.12-13911.21" */
wire [5:0] mstatus_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13911.12-13911.21" */
wire [5:0] mstatus_d_t0;
/* src = "generated/sv2v_out.v:13913.6-13913.16" */
wire mstatus_en;
/* src = "generated/sv2v_out.v:13912.7-13912.18" */
wire mstatus_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13912.7-13912.18" */
wire mstatus_err_t0;
/* src = "generated/sv2v_out.v:13910.13-13910.22" */
wire [5:0] mstatus_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13910.13-13910.22" */
wire [5:0] mstatus_q_t0;
/* src = "generated/sv2v_out.v:13926.13-13926.20" */
wire [31:0] mtval_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13926.13-13926.20" */
wire [31:0] mtval_d_t0;
/* src = "generated/sv2v_out.v:13927.6-13927.14" */
wire mtval_en;
/* src = "generated/sv2v_out.v:13929.13-13929.20" */
wire [31:0] mtvec_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13929.13-13929.20" */
wire [31:0] mtvec_d_t0;
/* src = "generated/sv2v_out.v:13931.6-13931.14" */
wire mtvec_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13931.6-13931.14" */
wire mtvec_en_t0;
/* src = "generated/sv2v_out.v:13930.7-13930.16" */
wire mtvec_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13930.7-13930.16" */
wire mtvec_err_t0;
/* src = "generated/sv2v_out.v:13881.13-13881.23" */
input mul_wait_i;
wire mul_wait_i;
/* cellift = 32'd1 */
input mul_wait_i_t0;
wire mul_wait_i_t0;
/* src = "generated/sv2v_out.v:13831.13-13831.23" */
input nmi_mode_i;
wire nmi_mode_i;
/* cellift = 32'd1 */
input nmi_mode_i_t0;
wire nmi_mode_i_t0;
/* src = "generated/sv2v_out.v:13850.20-13850.27" */
input [31:0] pc_id_i;
wire [31:0] pc_id_i;
/* cellift = 32'd1 */
input [31:0] pc_id_i_t0;
wire [31:0] pc_id_i_t0;
/* src = "generated/sv2v_out.v:13849.20-13849.27" */
input [31:0] pc_if_i;
wire [31:0] pc_if_i;
/* cellift = 32'd1 */
input [31:0] pc_if_i_t0;
wire [31:0] pc_if_i_t0;
/* src = "generated/sv2v_out.v:13851.20-13851.27" */
input [31:0] pc_wb_i;
wire [31:0] pc_wb_i;
/* cellift = 32'd1 */
input [31:0] pc_wb_i_t0;
wire [31:0] pc_wb_i_t0;
/* src = "generated/sv2v_out.v:13909.12-13909.22" */
wire [1:0] priv_lvl_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13909.12-13909.22" */
wire [1:0] priv_lvl_d_t0;
/* src = "generated/sv2v_out.v:13815.20-13815.34" */
output [1:0] priv_mode_id_o;
reg [1:0] priv_mode_id_o;
/* cellift = 32'd1 */
output [1:0] priv_mode_id_o_t0;
reg [1:0] priv_mode_id_o_t0;
/* src = "generated/sv2v_out.v:13816.20-13816.35" */
output [1:0] priv_mode_lsu_o;
wire [1:0] priv_mode_lsu_o;
/* cellift = 32'd1 */
output [1:0] priv_mode_lsu_o_t0;
wire [1:0] priv_mode_lsu_o_t0;
/* src = "generated/sv2v_out.v:13813.13-13813.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:13848.14-13848.29" */
output trigger_match_o;
wire trigger_match_o;
/* cellift = 32'd1 */
output trigger_match_o_t0;
wire trigger_match_o_t0;
assign illegal_csr_dbg = dbg_csr & /* src = "generated/sv2v_out.v:13998.27-13998.50" */ _0208_;
assign illegal_csr_insn_o = csr_access_i & /* src = "generated/sv2v_out.v:14001.30-14001.119" */ _1241_;
assign _0106_ = _0245_ & /* src = "generated/sv2v_out.v:14310.26-14310.52" */ csr_rdata_o;
assign _0108_ = csr_wr & /* src = "generated/sv2v_out.v:14315.23-14315.43" */ csr_op_en_i;
assign csr_we_int = _0108_ & /* src = "generated/sv2v_out.v:14315.22-14315.66" */ _1233_;
assign irqs_o = { irq_software_i, irq_timer_i, irq_external_i, irq_fast_i } & /* src = "generated/sv2v_out.v:14326.18-14326.29" */ mie_q;
assign _0110_ = instr_ret_i & /* src = "generated/sv2v_out.v:14699.18-14699.57" */ _1234_;
assign _0112_ = instr_ret_spec_i & /* src = "generated/sv2v_out.v:14706.27-14706.63" */ _1234_;
assign icache_enable_o = cpuctrlsts_part_q[0] & /* src = "generated/sv2v_out.v:14910.27-14910.89" */ _1235_;
assign _0113_ = ~ _0265_;
assign _0114_ = ~ mcountinhibit_we;
assign _0286_ = { _0265_, _0265_ } & priv_lvl_d_t0;
assign _0288_ = { mcountinhibit_we, mcountinhibit_we } & { dummy_instr_seed_o_t0[2], dummy_instr_seed_o_t0[0] };
assign _0287_ = { _0113_, _0113_ } & priv_mode_id_o_t0;
assign _0289_ = { _0114_, _0114_ } & { mcountinhibit_t0[2], mcountinhibit_t0[0] };
assign _0784_ = _0286_ | _0287_;
assign _0785_ = _0288_ | _0289_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers  */
/* PC_TAINT_INFO STATE_NAME priv_mode_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) priv_mode_id_o_t0 <= 2'h0;
else priv_mode_id_o_t0 <= _0784_;
reg [1:0] _1372_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers  */
/* PC_TAINT_INFO STATE_NAME _1372_ */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) _1372_ <= 2'h0;
else _1372_ <= _0785_;
assign { mcountinhibit_t0[2], mcountinhibit_t0[0] } = _1372_;
assign _0271_ = csr_access_i_t0 & _1241_;
assign _0274_ = csr_wdata_i_t0 & csr_rdata_o;
assign _0277_ = { irq_software_i_t0, irq_timer_i_t0, irq_external_i_t0, irq_fast_i_t0 } & mie_q;
assign _0280_ = instr_ret_i_t0 & _1234_;
assign _0283_ = cpuctrlsts_part_q_t0[0] & _1235_;
assign illegal_csr_dbg_t0 = debug_mode_i_t0 & dbg_csr;
assign _0272_ = _1242_ & csr_access_i;
assign _0275_ = csr_rdata_o_t0 & _0245_;
assign _0278_ = mie_q_t0 & { irq_software_i, irq_timer_i, irq_external_i, irq_fast_i };
assign _0281_ = mcountinhibit_t0[2] & instr_ret_i;
assign _0284_ = _1236_ & cpuctrlsts_part_q[0];
assign _0273_ = csr_access_i_t0 & _1242_;
assign _0276_ = csr_wdata_i_t0 & csr_rdata_o_t0;
assign _0279_ = { irq_software_i_t0, irq_timer_i_t0, irq_external_i_t0, irq_fast_i_t0 } & mie_q_t0;
assign _0282_ = instr_ret_i_t0 & mcountinhibit_t0[2];
assign _0285_ = cpuctrlsts_part_q_t0[0] & _1236_;
assign _0779_ = _0271_ | _0272_;
assign _0780_ = _0274_ | _0275_;
assign _0781_ = _0277_ | _0278_;
assign _0782_ = _0280_ | _0281_;
assign _0783_ = _0283_ | _0284_;
assign illegal_csr_insn_o_t0 = _0779_ | _0273_;
assign _0107_ = _0780_ | _0276_;
assign irqs_o_t0 = _0781_ | _0279_;
assign _0111_ = _0782_ | _0282_;
assign icache_enable_o_t0 = _0783_ | _0285_;
/* src = "generated/sv2v_out.v:14299.2-14303.29" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers  */
/* PC_TAINT_INFO STATE_NAME priv_mode_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) priv_mode_id_o <= 2'h3;
else if (_0265_) priv_mode_id_o <= priv_lvl_d;
reg [1:0] _1400_;
/* src = "generated/sv2v_out.v:14761.2-14765.39" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers  */
/* PC_TAINT_INFO STATE_NAME _1400_ */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) _1400_ <= 2'h0;
else if (mcountinhibit_we) _1400_ <= { dummy_instr_seed_o[2], dummy_instr_seed_o[0] };
assign { mcountinhibit[2], mcountinhibit[0] } = _1400_;
assign _0115_ = ~ { _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_ };
assign _0116_ = ~ { _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_ };
assign _0117_ = ~ _1294_;
assign _0119_ = ~ _1301_;
assign _0121_ = ~ _0253_;
assign _0122_ = ~ _1304_;
assign _0124_ = ~ _1302_;
assign _0125_ = ~ _0768_;
assign _0126_ = ~ _0254_;
assign _0127_ = ~ _0255_;
assign _0128_ = ~ _1297_;
assign _0129_ = ~ _0769_;
assign _0120_ = ~ _0767_;
assign _0133_ = ~ _0770_;
assign _0136_ = ~ _0771_;
assign _0141_ = ~ { _1299_, _1299_, _1299_ };
assign _0142_ = ~ { _1301_, _1301_, _1301_ };
assign _0143_ = ~ { _0767_, _0767_, _0767_ };
assign _0144_ = ~ { _0256_, _0256_, _0256_ };
assign _0145_ = ~ { _1303_, _1303_, _1303_ };
assign _0146_ = ~ { _1305_, _1305_, _1305_ };
assign _0147_ = ~ { _0770_, _0770_, _0770_ };
assign _0148_ = ~ { _1306_, _1306_, _1306_ };
assign _0149_ = ~ { _0257_, _0257_, _0257_ };
assign _0150_ = ~ { _0259_, _0259_, _0259_ };
assign _0131_ = ~ _0256_;
assign _0138_ = ~ _0258_;
assign _0139_ = ~ { _1297_, _1297_, _1297_ };
assign _0140_ = ~ { _0769_, _0769_, _0769_ };
assign _0151_ = ~ { _1298_, _1298_, _1298_ };
assign _0152_ = ~ { _1300_, _1300_, _1300_ };
assign _0153_ = ~ { _0773_, _0773_, _0773_ };
assign _0155_ = ~ { _0260_, _0260_, _0260_ };
assign _0154_ = ~ { _0774_, _0774_, _0774_ };
assign _0159_ = ~ { _1310_, _1310_, _1310_ };
assign _0160_ = ~ { _0775_, _0775_, _0775_ };
assign _0161_ = ~ { _1291_, _1291_, _1291_ };
assign _0162_ = ~ { _0776_, _0776_, _0776_ };
assign _0163_ = ~ { _0261_, _0261_, _0261_ };
assign _0164_ = ~ { _1346_, _1346_, _1346_ };
assign _0165_ = ~ { _0771_, _0771_, _0771_ };
assign _0166_ = ~ { _0262_, _0262_, _0262_ };
assign _0172_ = ~ _0777_;
assign _0174_ = ~ _0778_;
assign _0175_ = ~ _0263_;
assign _0176_ = ~ _0264_;
assign _0169_ = ~ _1300_;
assign _0132_ = ~ _1305_;
assign _0156_ = ~ { _1294_, _1294_, _1294_ };
assign _0157_ = ~ { _0253_, _0253_, _0253_ };
assign _0178_ = ~ { _1304_, _1304_, _1304_ };
assign _0179_ = ~ { _1302_, _1302_, _1302_ };
assign _0180_ = ~ { _0768_, _0768_, _0768_ };
assign _0181_ = ~ { _0254_, _0254_, _0254_ };
assign _0158_ = ~ { _0255_, _0255_, _0255_ };
assign _0171_ = ~ _0261_;
assign _0134_ = ~ _1306_;
assign _0177_ = ~ _0262_;
assign _0182_ = ~ { _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_ };
assign _0183_ = ~ { _1310_, _1310_, _1310_, _1310_, _1310_, _1310_, _1310_, _1310_, _1310_ };
assign _0184_ = ~ { _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_ };
assign _0185_ = ~ { _1300_, _1300_, _1300_, _1300_, _1300_, _1300_, _1300_, _1300_, _1300_ };
assign _0186_ = ~ { _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_ };
assign _0187_ = ~ { _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_ };
assign _0188_ = ~ { _0261_, _0261_, _0261_, _0261_, _0261_, _0261_, _0261_, _0261_, _0261_ };
assign _0189_ = ~ { _1305_, _1305_, _1305_, _1305_, _1305_, _1305_, _1305_, _1305_, _1305_ };
assign _0190_ = ~ { _0770_, _0770_, _0770_, _0770_, _0770_, _0770_, _0770_, _0770_, _0770_ };
assign _0191_ = ~ { _1306_, _1306_, _1306_, _1306_, _1306_, _1306_, _1306_, _1306_, _1306_ };
assign _0192_ = ~ { _1346_, _1346_, _1346_, _1346_, _1346_, _1346_, _1346_, _1346_, _1346_ };
assign _0193_ = ~ { _0771_, _0771_, _0771_, _0771_, _0771_, _0771_, _0771_, _0771_, _0771_ };
assign _0194_ = ~ { _0257_, _0257_, _0257_, _0257_, _0257_, _0257_, _0257_, _0257_, _0257_ };
assign _0195_ = ~ { _0262_, _0262_, _0262_, _0262_, _0262_, _0262_, _0262_, _0262_, _0262_ };
assign _0168_ = ~ _0775_;
assign _0170_ = ~ _0776_;
assign _0123_ = ~ _1303_;
assign _0135_ = ~ _1292_;
assign _0137_ = ~ _0257_;
assign _0196_ = ~ { _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_ };
assign _0197_ = ~ { _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_, _0270_ };
assign _0167_ = ~ _1310_;
assign _0199_ = ~ { nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i };
assign _0200_ = ~ _1231_;
assign _0201_ = ~ { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
assign _0202_ = ~ { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
assign _0207_ = ~ _1226_;
assign _0206_ = ~ cpuctrlsts_part_q[6];
assign _0210_ = ~ { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i };
assign _0211_ = ~ { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i };
assign _0209_ = ~ { debug_mode_i, debug_mode_i };
assign _0212_ = ~ { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
assign _0213_ = ~ { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
assign _0214_ = ~ { debug_csr_save_i, debug_csr_save_i };
assign _0215_ = ~ { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
assign _0216_ = ~ { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
assign _0217_ = ~ { csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i };
assign _0218_ = ~ { csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i };
assign _0219_ = ~ { csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i };
assign _0204_ = ~ csr_restore_mret_i;
assign _0205_ = ~ csr_restore_dret_i;
assign _0198_ = ~ csr_save_cause_i;
assign _0203_ = ~ { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
assign _0221_ = ~ { csr_save_cause_i, csr_save_cause_i };
assign _0220_ = ~ { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
assign _0222_ = ~ { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
assign _0223_ = ~ { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
assign _0224_ = ~ { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
assign _0225_ = ~ { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
assign _0226_ = ~ { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
assign _0227_ = ~ { nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i };
assign _0228_ = ~ { csr_restore_dret_i, csr_restore_dret_i };
assign _0208_ = ~ debug_mode_i;
assign _0229_ = ~ { _1291_, _1291_, _1291_, _1291_ };
assign _0230_ = ~ { _1292_, _1292_ };
assign _0231_ = ~ { _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_ };
assign _0232_ = ~ { _1291_, _1291_ };
assign _0130_ = ~ _1291_;
assign _0233_ = ~ { _1225_, _1225_ };
assign _0234_ = ~ { _1224_, _1224_ };
assign _0235_ = ~ { _1297_, _1297_, _1297_, _1297_, _1297_, _1297_, _1297_, _1297_ };
assign _0118_ = ~ _1299_;
assign _0237_ = ~ { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int };
assign _0238_ = ~ { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int };
assign _0236_ = ~ csr_we_int;
assign _0239_ = ~ { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int };
assign _0240_ = ~ { csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i };
assign _0241_ = ~ { mstatus_q[1], mstatus_q[1] };
assign _0242_ = ~ { _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_ };
assign _0290_ = _0115_ & _1246_;
assign _0292_ = _0116_ & _0792_;
assign _0294_ = _0117_ & _0794_;
assign _0296_ = _0118_ & dscratch0_q_t0[31];
assign _0298_ = _0119_ & dcsr_q_t0[31];
assign _0300_ = _0120_ & _0800_;
assign _0302_ = _0121_ & _0802_;
assign _0304_ = _0122_ & csr_mepc_o_t0[31];
assign _0306_ = _0123_ & _0806_;
assign _0308_ = _0124_ & mscratch_q_t0[31];
assign _0310_ = _0125_ & _0812_;
assign _0312_ = _0126_ & _0814_;
assign _0314_ = _0127_ & _0816_;
assign _0316_ = _0128_ & _0015_[39];
assign _0318_ = _0129_ & _0820_;
assign _0320_ = _0118_ & dscratch0_q_t0[7];
assign _0322_ = _0130_ & irq_timer_i_t0;
assign _0324_ = _0119_ & _0826_;
assign _0326_ = _0120_ & _0828_;
assign _0328_ = _0131_ & _0830_;
assign _0330_ = _0132_ & csr_mtvec_o_t0[7];
assign _0332_ = _0133_ & _0836_;
assign _0334_ = _0134_ & mie_q_t0[16];
assign _0336_ = _0135_ & _0842_;
assign _0338_ = _0136_ & _0844_;
assign _0340_ = _0137_ & _0846_;
assign _0342_ = _0138_ & _0848_;
assign _0344_ = _0139_ & _0015_[38:36];
assign _0346_ = _0140_ & _0852_;
assign _0348_ = _0141_ & dscratch0_q_t0[6:4];
assign _0350_ = _0142_ & dcsr_q_t0[6:4];
assign _0352_ = _0143_ & _0858_;
assign _0354_ = _0144_ & _0860_;
assign _0356_ = _0145_ & { 2'h0, mcause_q_t0[4] };
assign _0358_ = _0146_ & csr_mtvec_o_t0[6:4];
assign _0360_ = _0147_ & _0866_;
assign _0362_ = _0148_ & hart_id_i_t0[6:4];
assign _0364_ = _0149_ & _0873_;
assign _0366_ = _0150_ & _0875_;
assign _0368_ = _0128_ & _0015_[35];
assign _0370_ = _0129_ & _0879_;
assign _0372_ = _0118_ & dscratch0_q_t0[3];
assign _0374_ = _0130_ & irq_software_i_t0;
assign _0376_ = _0119_ & _0885_;
assign _0378_ = _0120_ & _0887_;
assign _0380_ = _0131_ & _0889_;
assign _0382_ = _0123_ & mcause_q_t0[3];
assign _0384_ = _0132_ & csr_mtvec_o_t0[3];
assign _0386_ = _0133_ & _0895_;
assign _0388_ = _0134_ & mie_q_t0[17];
assign _0390_ = _0135_ & _0901_;
assign _0392_ = _0136_ & _0903_;
assign _0394_ = _0137_ & _0905_;
assign _0396_ = _0138_ & _0907_;
assign _0398_ = _0139_ & _0015_[34:32];
assign _0400_ = _0140_ & _0911_;
assign _0402_ = _0151_ & dscratch1_q_t0[2:0];
assign _0404_ = _0142_ & dcsr_q_t0[2:0];
assign _0406_ = _0152_ & _0917_;
assign _0408_ = _0153_ & _0919_;
assign _0410_ = _0144_ & _0921_;
assign _0412_ = _0145_ & mcause_q_t0[2:0];
assign _0414_ = _0146_ & csr_mtvec_o_t0[2:0];
assign _0416_ = _0147_ & _0927_;
assign _0418_ = _0154_ & _0934_;
assign _0420_ = _0149_ & _0936_;
assign _0422_ = _0155_ & _0938_;
assign _0424_ = _0156_ & _0940_;
assign _0426_ = _0141_ & dscratch0_q_t0[10:8];
assign _0428_ = _0142_ & dcsr_q_t0[10:8];
assign _0430_ = _0143_ & _0946_;
assign _0432_ = _0157_ & _0948_;
assign _0434_ = _0146_ & csr_mtvec_o_t0[10:8];
assign _0436_ = _0147_ & _0954_;
assign _0438_ = _0154_ & _0960_;
assign _0440_ = _0149_ & _0962_;
assign _0442_ = _0158_ & _0964_;
assign _0444_ = _0156_ & _0015_[20:18];
assign _0968_ = _0159_ & dscratch1_q_t0[20:18];
assign _0446_ = _0160_ & _0968_;
assign _0448_ = _0152_ & csr_depc_o_t0[20:18];
assign _0450_ = _0161_ & irq_fast_i_t0[4:2];
assign _0452_ = _0162_ & _0974_;
assign _0454_ = _0163_ & _0976_;
assign _0456_ = _0146_ & csr_mtvec_o_t0[20:18];
assign _0458_ = _0147_ & _0982_;
assign _0460_ = _0148_ & mie_q_t0[4:2];
assign _0990_ = _0164_ & _0988_;
assign _0462_ = _0165_ & _0990_;
assign _0464_ = _0149_ & _0992_;
assign _0466_ = _0166_ & _0994_;
assign _0468_ = _0117_ & _0015_[12];
assign _0998_ = _0167_ & dscratch1_q_t0[12];
assign _0470_ = _0168_ & _0998_;
assign _0472_ = _0169_ & csr_depc_o_t0[12];
assign _0474_ = _0130_ & csr_mtval_o_t0[12];
assign _0476_ = _0170_ & _1004_;
assign _0478_ = _0171_ & _1006_;
assign _1010_ = _0122_ & csr_mepc_o_t0[12];
assign _0480_ = _0124_ & mscratch_q_t0[12];
assign _0482_ = _0172_ & _1012_;
assign _1016_ = _0173_ & mstatus_q_t0[3];
assign _0484_ = _0174_ & _1018_;
assign _0486_ = _0175_ & _1020_;
assign _0488_ = _0176_ & _1022_;
assign _0490_ = _0117_ & _0015_[17];
assign _1026_ = _0167_ & dscratch1_q_t0[17];
assign _0492_ = _0168_ & _1026_;
assign _0494_ = _0169_ & csr_depc_o_t0[17];
assign _0496_ = _0130_ & irq_fast_i_t0[1];
assign _0498_ = _0170_ & _1032_;
assign _0500_ = _0171_ & _1034_;
assign _0502_ = _0132_ & csr_mtvec_o_t0[17];
assign _0504_ = _0133_ & _1040_;
assign _0506_ = _0134_ & mie_q_t0[1];
assign _0508_ = _0135_ & _1046_;
assign _0510_ = _0136_ & _1048_;
assign _0512_ = _0137_ & _1050_;
assign _0514_ = _0177_ & _1052_;
assign _0516_ = _0156_ & _1054_;
assign _0518_ = _0141_ & dscratch0_q_t0[15:13];
assign _0520_ = _0142_ & dcsr_q_t0[15:13];
assign _0522_ = _0143_ & _1060_;
assign _0524_ = _0157_ & _1062_;
assign _1066_ = _0178_ & csr_mepc_o_t0[15:13];
assign _0526_ = _0145_ & _1066_;
assign _0528_ = _0179_ & mscratch_q_t0[15:13];
assign _0530_ = _0180_ & _1072_;
assign _0532_ = _0181_ & _1074_;
assign _0534_ = _0158_ & _1076_;
assign _0536_ = _0117_ & _0015_[16];
assign _1080_ = _0167_ & dscratch1_q_t0[16];
assign _0538_ = _0168_ & _1080_;
assign _0540_ = _0169_ & csr_depc_o_t0[16];
assign _0542_ = _0130_ & irq_fast_i_t0[0];
assign _0544_ = _0170_ & _1086_;
assign _0546_ = _0171_ & _1088_;
assign _0548_ = _0132_ & csr_mtvec_o_t0[16];
assign _0550_ = _0133_ & _1094_;
assign _0552_ = _0134_ & mie_q_t0[0];
assign _0554_ = _0136_ & _1100_;
assign _0556_ = _0137_ & _1102_;
assign _0558_ = _0177_ & _1104_;
assign _0560_ = _0182_ & _0015_[30:22];
assign _1108_ = _0183_ & dscratch1_q_t0[30:22];
assign _0562_ = _0184_ & _1108_;
assign _0564_ = _0185_ & csr_depc_o_t0[30:22];
assign _0566_ = _0186_ & irq_fast_i_t0[14:6];
assign _0568_ = _0187_ & _1114_;
assign _0570_ = _0188_ & _1116_;
assign _0572_ = _0189_ & csr_mtvec_o_t0[30:22];
assign _0574_ = _0190_ & _1122_;
assign _0576_ = _0191_ & mie_q_t0[14:6];
assign _1130_ = _0192_ & _1128_;
assign _0578_ = _0193_ & _1130_;
assign _0580_ = _0194_ & _1132_;
assign _0582_ = _0195_ & _1134_;
assign _0584_ = _0117_ & _0015_[11];
assign _1138_ = _0167_ & dscratch1_q_t0[11];
assign _0586_ = _0168_ & _1138_;
assign _0588_ = _0169_ & csr_depc_o_t0[11];
assign _0590_ = _0130_ & irq_external_i_t0;
assign _0592_ = _0170_ & _1144_;
assign _0594_ = _0171_ & _1146_;
assign _0596_ = _0132_ & csr_mtvec_o_t0[11];
assign _0598_ = _0133_ & _1152_;
assign _0600_ = _0134_ & mie_q_t0[15];
assign _0602_ = _0135_ & _1158_;
assign _0604_ = _0136_ & _1160_;
assign _0606_ = _0137_ & _1162_;
assign _0608_ = _0177_ & _1164_;
assign _0610_ = _0196_ & \mhpmcounter[0]_t0 ;
assign _0015_ = _0197_ & _1166_;
assign _0612_ = _0117_ & _0015_[21];
assign _1170_ = _0167_ & dscratch1_q_t0[21];
assign _0614_ = _0168_ & _1170_;
assign _0616_ = _0169_ & csr_depc_o_t0[21];
assign _0618_ = _0130_ & irq_fast_i_t0[5];
assign _0620_ = _0170_ & _1176_;
assign _0622_ = _0171_ & _1178_;
assign _0624_ = _0132_ & csr_mtvec_o_t0[21];
assign _0626_ = _0133_ & _1184_;
assign _0628_ = _0134_ & mie_q_t0[5];
assign _0630_ = _0135_ & _1190_;
assign _0632_ = _0136_ & _1192_;
assign _0634_ = _0137_ & _1194_;
assign _0636_ = _0177_ & _1196_;
assign _0651_ = _0198_ & _0001_[7];
assign _0653_ = _0199_ & { dummy_instr_seed_o_t0[31:1], 1'h0 };
assign _0103_ = _0200_ & _0011_[1];
assign _0655_ = _0201_ & _0011_[4:2];
assign _0657_ = _0202_ & _1252_;
assign _0659_ = _0203_ & _1254_;
assign _0661_ = _0204_ & _0011_[1];
assign _0663_ = _0205_ & _1256_;
assign _0665_ = _0198_ & _1258_;
assign _0667_ = _0204_ & _0011_[5];
assign _0669_ = _0205_ & _1260_;
assign _0671_ = _0198_ & _1262_;
assign _0099_ = _0206_ & _0001_[7];
assign _0673_ = _0209_ & _0090_;
assign _0675_ = _0210_ & csr_mcause_i_t0;
assign _0677_ = _0211_ & _0030_;
assign _0679_ = _0207_ & _0099_;
assign _0681_ = _0209_ & priv_mode_id_o_t0;
assign _0683_ = _0208_ & mstatus_q_t0[5];
assign _0685_ = _0211_ & csr_mtval_i_t0;
assign _0687_ = _0212_ & { dummy_instr_seed_o_t0[31:1], 1'h0 };
assign _0689_ = _0213_ & _0004_[8:6];
assign _0691_ = _0214_ & _0004_[1:0];
assign _0693_ = _0214_ & _0080_;
assign _0695_ = _0212_ & _0064_;
assign _0697_ = _0215_ & _0057_;
assign _0699_ = _0212_ & _0059_;
assign _0701_ = _0216_ & _0097_;
assign _0703_ = _0217_ & pc_id_i_t0;
assign _0705_ = _0218_ & _1264_;
assign _0707_ = _0219_ & _1266_;
assign _1270_ = _0204_ & _0001_[6];
assign _0709_ = _0205_ & _1270_;
assign _0711_ = _0198_ & _1272_;
assign _0713_ = _0220_ & { dummy_instr_seed_o_t0[31:1], 1'h0 };
assign _0715_ = _0203_ & _0004_[8:6];
assign _0717_ = _0221_ & _0004_[1:0];
assign _0719_ = _0220_ & dummy_instr_seed_o_t0;
assign _0721_ = _0222_ & { 2'h0, dummy_instr_seed_o_t0[4:0] };
assign _0723_ = _0223_ & _1276_;
assign _0725_ = _0224_ & _1278_;
assign _0727_ = _0225_ & { dummy_instr_seed_o_t0[31:1], 1'h0 };
assign _0729_ = _0226_ & _1282_;
assign _0731_ = _0220_ & _1284_;
assign _0733_ = _0227_ & { 2'h0, dummy_instr_seed_o_t0[4:0] };
assign _0735_ = _0228_ & _1288_;
assign priv_lvl_d_t0 = _0221_ & _1290_;
assign _0021_[31:28] = _0229_ & dcsr_q_t0[31:28];
assign _0737_ = _0230_ & mstatus_q_t0[5:4];
assign _0739_ = _0230_ & mstatus_q_t0[3:2];
assign _0741_ = _0130_ & dcsr_q_t0[15];
assign _0021_[14] = _0130_ & dcsr_q_t0[14];
assign _0021_[27:16] = _0231_ & dcsr_q_t0[27:16];
assign _0743_ = _0230_ & mstatus_q_t0[1:0];
assign _0745_ = _0232_ & dcsr_q_t0[1:0];
assign _0021_[5] = _0130_ & dcsr_q_t0[5];
assign _0021_[4] = _0130_ & dcsr_q_t0[4];
assign _0021_[3] = _0130_ & dcsr_q_t0[3];
assign _0747_ = _0130_ & dcsr_q_t0[2];
assign _0749_ = _0232_ & dcsr_q_t0[13:12];
assign _0021_[11] = _0130_ & dcsr_q_t0[11];
assign _0054_ = _0233_ & dummy_instr_seed_o_t0[1:0];
assign _0021_[9] = _0130_ & dcsr_q_t0[9];
assign _0062_ = _0234_ & dummy_instr_seed_o_t0[12:11];
assign _0751_ = _0235_ & cpuctrlsts_part_q_t0;
assign _0021_[10] = _0130_ & dcsr_q_t0[10];
assign _0052_ = _0124_ & csr_mtvec_init_i_t0;
assign _0753_ = _0237_ & cpuctrlsts_part_q_t0;
assign _0755_ = _0238_ & dcsr_q_t0;
assign _0757_ = _0236_ & csr_mtvec_init_i_t0;
assign _0759_ = _0239_ & mstatus_q_t0;
assign _0761_ = _0240_ & { dummy_instr_seed_o_t0[31:8], 8'h00 };
assign _0763_ = _0241_ & priv_mode_id_o_t0;
assign _0765_ = _0242_ & minstret_raw_t0;
assign _0291_ = { _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_, _1220_ } & _0107_;
assign _0293_ = { _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_, _0269_ } & csr_wdata_i_t0;
assign _0794_ = _1296_ & _0015_[31];
assign _0295_ = _1294_ & _0015_[63];
assign _0297_ = _1299_ & dscratch1_q_t0[31];
assign _0299_ = _1301_ & csr_depc_o_t0[31];
assign _0301_ = _0767_ & _0798_;
assign _0303_ = _0253_ & _0796_;
assign _0305_ = _1304_ & _1244_;
assign _0307_ = _1303_ & csr_mtval_o_t0[31];
assign _0309_ = _1302_ & csr_mtvec_o_t0[31];
assign _0812_ = _1311_ & hart_id_i_t0[31];
assign _0311_ = _0768_ & _0810_;
assign _0313_ = _0254_ & _0808_;
assign _0315_ = _0255_ & _0804_;
assign _0317_ = _1297_ & cpuctrlsts_part_q_t0[7];
assign _0820_ = _1296_ & _0015_[7];
assign _0319_ = _0769_ & _0818_;
assign _0321_ = _1299_ & dscratch1_q_t0[7];
assign _0323_ = _1291_ & dcsr_q_t0[7];
assign _0325_ = _1301_ & csr_depc_o_t0[7];
assign _0327_ = _0767_ & _0824_;
assign _0329_ = _0256_ & _0822_;
assign _0834_ = _1303_ & csr_mtval_o_t0[7];
assign _0331_ = _1305_ & csr_mepc_o_t0[7];
assign _0333_ = _0770_ & _0834_;
assign _0335_ = _1306_ & mscratch_q_t0[7];
assign _0842_ = _1311_ & hart_id_i_t0[7];
assign _0337_ = _1292_ & mstatus_q_t0[4];
assign _0339_ = _0771_ & _0840_;
assign _0341_ = _0257_ & _0838_;
assign _0343_ = _0258_ & _0832_;
assign _0345_ = { _1297_, _1297_, _1297_ } & cpuctrlsts_part_q_t0[6:4];
assign _0852_ = { _1296_, _1296_, _1296_ } & _0015_[6:4];
assign _0347_ = { _0769_, _0769_, _0769_ } & _0850_;
assign _0349_ = { _1299_, _1299_, _1299_ } & dscratch1_q_t0[6:4];
assign _0351_ = { _1301_, _1301_, _1301_ } & csr_depc_o_t0[6:4];
assign _0353_ = { _0767_, _0767_, _0767_ } & _0856_;
assign _0355_ = { _0256_, _0256_, _0256_ } & _0854_;
assign _0357_ = { _1303_, _1303_, _1303_ } & csr_mtval_o_t0[6:4];
assign _0359_ = { _1305_, _1305_, _1305_ } & csr_mepc_o_t0[6:4];
assign _0361_ = { _0770_, _0770_, _0770_ } & _0864_;
assign _0363_ = { _1306_, _1306_, _1306_ } & mscratch_q_t0[6:4];
assign _0873_ = { _0772_, _0772_, _0772_ } & _0870_;
assign _0365_ = { _0257_, _0257_, _0257_ } & _0868_;
assign _0367_ = { _0259_, _0259_, _0259_ } & _0862_;
assign _0369_ = _1297_ & cpuctrlsts_part_q_t0[3];
assign _0879_ = _1296_ & _0015_[3];
assign _0371_ = _0769_ & _0877_;
assign _0373_ = _1299_ & dscratch1_q_t0[3];
assign _0375_ = _1291_ & dcsr_q_t0[3];
assign _0377_ = _1301_ & csr_depc_o_t0[3];
assign _0379_ = _0767_ & _0883_;
assign _0381_ = _0256_ & _0881_;
assign _0383_ = _1303_ & csr_mtval_o_t0[3];
assign _0385_ = _1305_ & csr_mepc_o_t0[3];
assign _0387_ = _0770_ & _0893_;
assign _0389_ = _1306_ & mscratch_q_t0[3];
assign _0901_ = _1311_ & hart_id_i_t0[3];
assign _0391_ = _1292_ & mstatus_q_t0[5];
assign _0393_ = _0771_ & _0899_;
assign _0395_ = _0257_ & _0897_;
assign _0397_ = _0258_ & _0891_;
assign _0399_ = { _1297_, _1297_, _1297_ } & cpuctrlsts_part_q_t0[2:0];
assign _0911_ = { _1296_, _1296_, _1296_ } & _0015_[2:0];
assign _0401_ = { _0769_, _0769_, _0769_ } & _0909_;
assign _0403_ = { _1298_, _1298_, _1298_ } & { mcountinhibit_t0[2], 1'h0, mcountinhibit_t0[0] };
assign _0405_ = { _1301_, _1301_, _1301_ } & csr_depc_o_t0[2:0];
assign _0407_ = { _1300_, _1300_, _1300_ } & dscratch0_q_t0[2:0];
assign _0409_ = { _0773_, _0773_, _0773_ } & _0915_;
assign _0411_ = { _0256_, _0256_, _0256_ } & _0913_;
assign _0413_ = { _1303_, _1303_, _1303_ } & csr_mtval_o_t0[2:0];
assign _0415_ = { _1305_, _1305_, _1305_ } & csr_mepc_o_t0[2:0];
assign _0417_ = { _0770_, _0770_, _0770_ } & _0925_;
assign _0931_ = { _1306_, _1306_, _1306_ } & mscratch_q_t0[2:0];
assign _0934_ = { _1311_, _1311_, _1311_ } & hart_id_i_t0[2:0];
assign _0419_ = { _0774_, _0774_, _0774_ } & _0931_;
assign _0421_ = { _0257_, _0257_, _0257_ } & _0929_;
assign _0423_ = { _0260_, _0260_, _0260_ } & _0923_;
assign _0940_ = { _1296_, _1296_, _1296_ } & _0015_[10:8];
assign _0425_ = { _1294_, _1294_, _1294_ } & _0015_[42:40];
assign _0427_ = { _1299_, _1299_, _1299_ } & dscratch1_q_t0[10:8];
assign _0429_ = { _1301_, _1301_, _1301_ } & csr_depc_o_t0[10:8];
assign _0431_ = { _0767_, _0767_, _0767_ } & _0944_;
assign _0433_ = { _0253_, _0253_, _0253_ } & _0942_;
assign _0952_ = { _1303_, _1303_, _1303_ } & csr_mtval_o_t0[10:8];
assign _0435_ = { _1305_, _1305_, _1305_ } & csr_mepc_o_t0[10:8];
assign _0437_ = { _0770_, _0770_, _0770_ } & _0952_;
assign _0958_ = { _1306_, _1306_, _1306_ } & mscratch_q_t0[10:8];
assign _0960_ = { _1311_, _1311_, _1311_ } & hart_id_i_t0[10:8];
assign _0439_ = { _0774_, _0774_, _0774_ } & _0958_;
assign _0441_ = { _0257_, _0257_, _0257_ } & _0956_;
assign _0443_ = { _0255_, _0255_, _0255_ } & _0950_;
assign _0445_ = { _1294_, _1294_, _1294_ } & _0015_[52:50];
assign _0447_ = { _0775_, _0775_, _0775_ } & _0966_;
assign _0449_ = { _1300_, _1300_, _1300_ } & dscratch0_q_t0[20:18];
assign _0451_ = { _1291_, _1291_, _1291_ } & dcsr_q_t0[20:18];
assign _0453_ = { _0776_, _0776_, _0776_ } & _0972_;
assign _0455_ = { _0261_, _0261_, _0261_ } & _0970_;
assign _0980_ = { _1303_, _1303_, _1303_ } & csr_mtval_o_t0[20:18];
assign _0457_ = { _1305_, _1305_, _1305_ } & csr_mepc_o_t0[20:18];
assign _0459_ = { _0770_, _0770_, _0770_ } & _0980_;
assign _0461_ = { _1306_, _1306_, _1306_ } & mscratch_q_t0[20:18];
assign _0988_ = { _1311_, _1311_, _1311_ } & hart_id_i_t0[20:18];
assign _0463_ = { _0771_, _0771_, _0771_ } & _0986_;
assign _0465_ = { _0257_, _0257_, _0257_ } & _0984_;
assign _0467_ = { _0262_, _0262_, _0262_ } & _0978_;
assign _0469_ = _1294_ & _0015_[44];
assign _0471_ = _0775_ & _0996_;
assign _0473_ = _1300_ & dscratch0_q_t0[12];
assign _0475_ = _1291_ & dcsr_q_t0[12];
assign _0477_ = _0776_ & _1002_;
assign _0479_ = _0261_ & _1000_;
assign _0481_ = _1302_ & csr_mtvec_o_t0[12];
assign _0483_ = _0777_ & _1010_;
assign _1018_ = _1311_ & hart_id_i_t0[12];
assign _0485_ = _0778_ & _1016_;
assign _0487_ = _0263_ & _1014_;
assign _0489_ = _0264_ & _1008_;
assign _0491_ = _1294_ & _0015_[49];
assign _0493_ = _0775_ & _1024_;
assign _0495_ = _1300_ & dscratch0_q_t0[17];
assign _0497_ = _1291_ & dcsr_q_t0[17];
assign _0499_ = _0776_ & _1030_;
assign _0501_ = _0261_ & _1028_;
assign _1038_ = _1303_ & csr_mtval_o_t0[17];
assign _0503_ = _1305_ & csr_mepc_o_t0[17];
assign _0505_ = _0770_ & _1038_;
assign _0507_ = _1306_ & mscratch_q_t0[17];
assign _1046_ = _1311_ & hart_id_i_t0[17];
assign _0509_ = _1292_ & mstatus_q_t0[1];
assign _0511_ = _0771_ & _1044_;
assign _0513_ = _0257_ & _1042_;
assign _0515_ = _0262_ & _1036_;
assign _1054_ = { _1296_, _1296_, _1296_ } & _0015_[15:13];
assign _0517_ = { _1294_, _1294_, _1294_ } & _0015_[47:45];
assign _0519_ = { _1299_, _1299_, _1299_ } & dscratch1_q_t0[15:13];
assign _0521_ = { _1301_, _1301_, _1301_ } & csr_depc_o_t0[15:13];
assign _0523_ = { _0767_, _0767_, _0767_ } & _1058_;
assign _0525_ = { _0253_, _0253_, _0253_ } & _1056_;
assign _0527_ = { _1303_, _1303_, _1303_ } & csr_mtval_o_t0[15:13];
assign _0529_ = { _1302_, _1302_, _1302_ } & csr_mtvec_o_t0[15:13];
assign _1072_ = { _1311_, _1311_, _1311_ } & hart_id_i_t0[15:13];
assign _0531_ = { _0768_, _0768_, _0768_ } & _1070_;
assign _0533_ = { _0254_, _0254_, _0254_ } & _1068_;
assign _0535_ = { _0255_, _0255_, _0255_ } & _1064_;
assign _0537_ = _1294_ & _0015_[48];
assign _0539_ = _0775_ & _1078_;
assign _0541_ = _1300_ & dscratch0_q_t0[16];
assign _0543_ = _1291_ & dcsr_q_t0[16];
assign _0545_ = _0776_ & _1084_;
assign _0547_ = _0261_ & _1082_;
assign _1092_ = _1303_ & csr_mtval_o_t0[16];
assign _0549_ = _1305_ & csr_mepc_o_t0[16];
assign _0551_ = _0770_ & _1092_;
assign _0553_ = _1306_ & mscratch_q_t0[16];
assign _1100_ = _1311_ & hart_id_i_t0[16];
assign _0555_ = _0771_ & _1098_;
assign _0557_ = _0257_ & _1096_;
assign _0559_ = _0262_ & _1090_;
assign _0561_ = { _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_ } & _0015_[62:54];
assign _0563_ = { _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_ } & _1106_;
assign _0565_ = { _1300_, _1300_, _1300_, _1300_, _1300_, _1300_, _1300_, _1300_, _1300_ } & dscratch0_q_t0[30:22];
assign _0567_ = { _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_, _1291_ } & dcsr_q_t0[30:22];
assign _0569_ = { _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_ } & _1112_;
assign _0571_ = { _0261_, _0261_, _0261_, _0261_, _0261_, _0261_, _0261_, _0261_, _0261_ } & _1110_;
assign _1120_ = { _1303_, _1303_, _1303_, _1303_, _1303_, _1303_, _1303_, _1303_, _1303_ } & csr_mtval_o_t0[30:22];
assign _0573_ = { _1305_, _1305_, _1305_, _1305_, _1305_, _1305_, _1305_, _1305_, _1305_ } & csr_mepc_o_t0[30:22];
assign _0575_ = { _0770_, _0770_, _0770_, _0770_, _0770_, _0770_, _0770_, _0770_, _0770_ } & _1120_;
assign _0577_ = { _1306_, _1306_, _1306_, _1306_, _1306_, _1306_, _1306_, _1306_, _1306_ } & mscratch_q_t0[30:22];
assign _1128_ = { _1311_, _1311_, _1311_, _1311_, _1311_, _1311_, _1311_, _1311_, _1311_ } & hart_id_i_t0[30:22];
assign _0579_ = { _0771_, _0771_, _0771_, _0771_, _0771_, _0771_, _0771_, _0771_, _0771_ } & _1126_;
assign _0581_ = { _0257_, _0257_, _0257_, _0257_, _0257_, _0257_, _0257_, _0257_, _0257_ } & _1124_;
assign _0583_ = { _0262_, _0262_, _0262_, _0262_, _0262_, _0262_, _0262_, _0262_, _0262_ } & _1118_;
assign _0585_ = _1294_ & _0015_[43];
assign _0587_ = _0775_ & _1136_;
assign _0589_ = _1300_ & dscratch0_q_t0[11];
assign _0591_ = _1291_ & dcsr_q_t0[11];
assign _0593_ = _0776_ & _1142_;
assign _0595_ = _0261_ & _1140_;
assign _1150_ = _1303_ & csr_mtval_o_t0[11];
assign _0597_ = _1305_ & csr_mepc_o_t0[11];
assign _0599_ = _0770_ & _1150_;
assign _0601_ = _1306_ & mscratch_q_t0[11];
assign _1158_ = _1311_ & hart_id_i_t0[11];
assign _0603_ = _1292_ & mstatus_q_t0[2];
assign _0605_ = _0771_ & _1156_;
assign _0607_ = _0257_ & _1154_;
assign _0609_ = _0262_ & _1148_;
assign _0611_ = { _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_, _1343_ } & \mhpmcounter[2]_t0 ;
assign _0613_ = _1294_ & _0015_[53];
assign _0615_ = _0775_ & _1168_;
assign _0617_ = _1300_ & dscratch0_q_t0[21];
assign _0619_ = _1291_ & dcsr_q_t0[21];
assign _0621_ = _0776_ & _1174_;
assign _0623_ = _0261_ & _1172_;
assign _1182_ = _1303_ & csr_mtval_o_t0[21];
assign _0625_ = _1305_ & csr_mepc_o_t0[21];
assign _0627_ = _0770_ & _1182_;
assign _0629_ = _1306_ & mscratch_q_t0[21];
assign _1190_ = _1311_ & hart_id_i_t0[21];
assign _0631_ = _1292_ & mstatus_q_t0[0];
assign _0633_ = _0771_ & _1188_;
assign _0635_ = _0257_ & _1186_;
assign _0637_ = _0262_ & _1180_;
assign _0652_ = csr_save_cause_i & _0066_[1];
assign _0654_ = { nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i } & mstack_epc_q_t0;
assign _0105_[1:0] = { nmi_mode_i, nmi_mode_i } & mstack_q_t0[1:0];
assign _0105_[2] = nmi_mode_i & mstack_q_t0[2];
assign _0656_ = { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i } & _0105_;
assign _0658_ = { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i } & _0011_[4:2];
assign _0660_ = { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i } & _0086_[2:0];
assign _0662_ = csr_restore_mret_i & _0103_;
assign _0664_ = csr_restore_dret_i & _0011_[1];
assign _0666_ = csr_save_cause_i & _0011_[1];
assign _0668_ = csr_restore_mret_i & mstatus_q_t0[4];
assign _0670_ = csr_restore_dret_i & _0011_[5];
assign _0672_ = csr_save_cause_i & _0086_[3];
assign _0090_[0] = _1226_ & _0001_[6];
assign _0674_ = { debug_mode_i, debug_mode_i } & _0001_[7:6];
assign _0676_ = { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i } & { 2'h0, dummy_instr_seed_o_t0[4:0] };
assign _0678_ = { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i } & { dummy_instr_seed_o_t0[31:1], 1'h0 };
assign _0680_ = _1226_ & _0001_[7];
assign _0682_ = { debug_mode_i, debug_mode_i } & _0011_[3:2];
assign _0684_ = debug_mode_i & _0011_[4];
assign _0686_ = { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i } & dummy_instr_seed_o_t0;
assign _0688_ = { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i } & _0030_;
assign _0690_ = { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i } & debug_cause_i_t0;
assign _0692_ = { debug_csr_save_i, debug_csr_save_i } & priv_mode_id_o_t0;
assign _0694_ = { debug_csr_save_i, debug_csr_save_i } & _0001_[7:6];
assign _0696_ = { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i } & dummy_instr_seed_o_t0;
assign _0698_ = { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i } & { 2'h0, dummy_instr_seed_o_t0[4:0] };
assign _0700_ = { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i } & { dummy_instr_seed_o_t0[31:1], 1'h0 };
assign _0702_ = { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i } & _0011_[5:2];
assign _0704_ = { csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i } & pc_wb_i_t0;
assign _0706_ = { csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i } & pc_id_i_t0;
assign _0708_ = { csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i } & pc_if_i_t0;
assign _0710_ = csr_restore_dret_i & _0001_[6];
assign _0712_ = csr_save_cause_i & _0066_[0];
assign _0714_ = { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i } & _0024_;
assign _0716_ = { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i } & _0101_;
assign _0718_ = { csr_save_cause_i, csr_save_cause_i } & _0093_;
assign _0720_ = { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i } & _0049_;
assign _0722_ = { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i } & _0072_;
assign _0724_ = { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i } & { 2'h0, dummy_instr_seed_o_t0[4:0] };
assign _0726_ = { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i } & _0032_;
assign _0728_ = { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i } & _0075_;
assign _0730_ = { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i } & { dummy_instr_seed_o_t0[31:1], 1'h0 };
assign _0732_ = { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i } & _0036_;
assign _0734_ = { nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i } & mstack_cause_q_t0;
assign _1288_ = { csr_restore_mret_i, csr_restore_mret_i } & mstatus_q_t0[3:2];
assign _0736_ = { csr_restore_dret_i, csr_restore_dret_i } & dcsr_q_t0[1:0];
assign _0097_[3] = debug_mode_i & _0011_[5];
assign _0738_ = { _1292_, _1292_ } & { dummy_instr_seed_o_t0[3], dummy_instr_seed_o_t0[7] };
assign _0740_ = { _1292_, _1292_ } & _0062_;
assign _0742_ = _1291_ & dummy_instr_seed_o_t0[15];
assign _0744_ = { _1292_, _1292_ } & { dummy_instr_seed_o_t0[17], dummy_instr_seed_o_t0[21] };
assign _0746_ = { _1291_, _1291_ } & _0054_;
assign _0748_ = _1291_ & dummy_instr_seed_o_t0[2];
assign _0750_ = { _1291_, _1291_ } & dummy_instr_seed_o_t0[13:12];
assign _0752_ = { _1297_, _1297_, _1297_, _1297_, _1297_, _1297_, _1297_, _1297_ } & { dummy_instr_seed_o_t0[7:1], 1'h0 };
assign _0041_ = { _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_, _1294_ } & _1238_;
assign _0039_ = { _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_, _1296_ } & _1238_;
assign _0754_ = { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int } & _0018_;
assign mhpmcounterh_we_t0 = { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int } & _0041_;
assign mhpmcounter_we_t0 = { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int } & _0039_;
assign _0756_ = { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int } & { _0021_[31:9], dcsr_q_t0[8:6], _0021_[5:0] };
assign _0758_ = csr_we_int & _0052_;
assign _0760_ = { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int } & _0046_;
assign _0762_ = { csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i } & { boot_addr_i_t0[31:8], 8'h00 };
assign _0764_ = { mstatus_q[1], mstatus_q[1] } & mstatus_q_t0[3:2];
assign _0766_ = { _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_, _0112_ } & minstret_next_t0;
assign _0792_ = _0290_ | _0291_;
assign dummy_instr_seed_o_t0 = _0292_ | _0293_;
assign _0796_ = _0294_ | _0295_;
assign _0798_ = _0296_ | _0297_;
assign _0800_ = _0298_ | _0299_;
assign _0802_ = _0300_ | _0301_;
assign _0804_ = _0302_ | _0303_;
assign _0806_ = _0304_ | _0305_;
assign _0808_ = _0306_ | _0307_;
assign _0810_ = _0308_ | _0309_;
assign _0814_ = _0310_ | _0311_;
assign _0816_ = _0312_ | _0313_;
assign csr_rdata_o_t0[31] = _0314_ | _0315_;
assign _0818_ = _0316_ | _0317_;
assign _0822_ = _0318_ | _0319_;
assign _0824_ = _0320_ | _0321_;
assign _0826_ = _0322_ | _0323_;
assign _0828_ = _0324_ | _0325_;
assign _0830_ = _0326_ | _0327_;
assign _0832_ = _0328_ | _0329_;
assign _0836_ = _0330_ | _0331_;
assign _0838_ = _0332_ | _0333_;
assign _0840_ = _0334_ | _0335_;
assign _0844_ = _0336_ | _0337_;
assign _0846_ = _0338_ | _0339_;
assign _0848_ = _0340_ | _0341_;
assign csr_rdata_o_t0[7] = _0342_ | _0343_;
assign _0850_ = _0344_ | _0345_;
assign _0854_ = _0346_ | _0347_;
assign _0856_ = _0348_ | _0349_;
assign _0858_ = _0350_ | _0351_;
assign _0860_ = _0352_ | _0353_;
assign _0862_ = _0354_ | _0355_;
assign _0864_ = _0356_ | _0357_;
assign _0866_ = _0358_ | _0359_;
assign _0868_ = _0360_ | _0361_;
assign _0870_ = _0362_ | _0363_;
assign _0875_ = _0364_ | _0365_;
assign csr_rdata_o_t0[6:4] = _0366_ | _0367_;
assign _0877_ = _0368_ | _0369_;
assign _0881_ = _0370_ | _0371_;
assign _0883_ = _0372_ | _0373_;
assign _0885_ = _0374_ | _0375_;
assign _0887_ = _0376_ | _0377_;
assign _0889_ = _0378_ | _0379_;
assign _0891_ = _0380_ | _0381_;
assign _0893_ = _0382_ | _0383_;
assign _0895_ = _0384_ | _0385_;
assign _0897_ = _0386_ | _0387_;
assign _0899_ = _0388_ | _0389_;
assign _0903_ = _0390_ | _0391_;
assign _0905_ = _0392_ | _0393_;
assign _0907_ = _0394_ | _0395_;
assign csr_rdata_o_t0[3] = _0396_ | _0397_;
assign _0909_ = _0398_ | _0399_;
assign _0913_ = _0400_ | _0401_;
assign _0915_ = _0402_ | _0403_;
assign _0917_ = _0404_ | _0405_;
assign _0919_ = _0406_ | _0407_;
assign _0921_ = _0408_ | _0409_;
assign _0923_ = _0410_ | _0411_;
assign _0925_ = _0412_ | _0413_;
assign _0927_ = _0414_ | _0415_;
assign _0929_ = _0416_ | _0417_;
assign _0936_ = _0418_ | _0419_;
assign _0938_ = _0420_ | _0421_;
assign csr_rdata_o_t0[2:0] = _0422_ | _0423_;
assign _0942_ = _0424_ | _0425_;
assign _0944_ = _0426_ | _0427_;
assign _0946_ = _0428_ | _0429_;
assign _0948_ = _0430_ | _0431_;
assign _0950_ = _0432_ | _0433_;
assign _0954_ = _0434_ | _0435_;
assign _0956_ = _0436_ | _0437_;
assign _0962_ = _0438_ | _0439_;
assign _0964_ = _0440_ | _0441_;
assign csr_rdata_o_t0[10:8] = _0442_ | _0443_;
assign _0966_ = _0444_ | _0445_;
assign _0970_ = _0446_ | _0447_;
assign _0972_ = _0448_ | _0449_;
assign _0974_ = _0450_ | _0451_;
assign _0976_ = _0452_ | _0453_;
assign _0978_ = _0454_ | _0455_;
assign _0982_ = _0456_ | _0457_;
assign _0984_ = _0458_ | _0459_;
assign _0986_ = _0460_ | _0461_;
assign _0992_ = _0462_ | _0463_;
assign _0994_ = _0464_ | _0465_;
assign csr_rdata_o_t0[20:18] = _0466_ | _0467_;
assign _0996_ = _0468_ | _0469_;
assign _1000_ = _0470_ | _0471_;
assign _1002_ = _0472_ | _0473_;
assign _1004_ = _0474_ | _0475_;
assign _1006_ = _0476_ | _0477_;
assign _1008_ = _0478_ | _0479_;
assign _1012_ = _0480_ | _0481_;
assign _1014_ = _0482_ | _0483_;
assign _1020_ = _0484_ | _0485_;
assign _1022_ = _0486_ | _0487_;
assign csr_rdata_o_t0[12] = _0488_ | _0489_;
assign _1024_ = _0490_ | _0491_;
assign _1028_ = _0492_ | _0493_;
assign _1030_ = _0494_ | _0495_;
assign _1032_ = _0496_ | _0497_;
assign _1034_ = _0498_ | _0499_;
assign _1036_ = _0500_ | _0501_;
assign _1040_ = _0502_ | _0503_;
assign _1042_ = _0504_ | _0505_;
assign _1044_ = _0506_ | _0507_;
assign _1048_ = _0508_ | _0509_;
assign _1050_ = _0510_ | _0511_;
assign _1052_ = _0512_ | _0513_;
assign csr_rdata_o_t0[17] = _0514_ | _0515_;
assign _1056_ = _0516_ | _0517_;
assign _1058_ = _0518_ | _0519_;
assign _1060_ = _0520_ | _0521_;
assign _1062_ = _0522_ | _0523_;
assign _1064_ = _0524_ | _0525_;
assign _1068_ = _0526_ | _0527_;
assign _1070_ = _0528_ | _0529_;
assign _1074_ = _0530_ | _0531_;
assign _1076_ = _0532_ | _0533_;
assign csr_rdata_o_t0[15:13] = _0534_ | _0535_;
assign _1078_ = _0536_ | _0537_;
assign _1082_ = _0538_ | _0539_;
assign _1084_ = _0540_ | _0541_;
assign _1086_ = _0542_ | _0543_;
assign _1088_ = _0544_ | _0545_;
assign _1090_ = _0546_ | _0547_;
assign _1094_ = _0548_ | _0549_;
assign _1096_ = _0550_ | _0551_;
assign _1098_ = _0552_ | _0553_;
assign _1102_ = _0554_ | _0555_;
assign _1104_ = _0556_ | _0557_;
assign csr_rdata_o_t0[16] = _0558_ | _0559_;
assign _1106_ = _0560_ | _0561_;
assign _1110_ = _0562_ | _0563_;
assign _1112_ = _0564_ | _0565_;
assign _1114_ = _0566_ | _0567_;
assign _1116_ = _0568_ | _0569_;
assign _1118_ = _0570_ | _0571_;
assign _1122_ = _0572_ | _0573_;
assign _1124_ = _0574_ | _0575_;
assign _1126_ = _0576_ | _0577_;
assign _1132_ = _0578_ | _0579_;
assign _1134_ = _0580_ | _0581_;
assign csr_rdata_o_t0[30:22] = _0582_ | _0583_;
assign _1136_ = _0584_ | _0585_;
assign _1140_ = _0586_ | _0587_;
assign _1142_ = _0588_ | _0589_;
assign _1144_ = _0590_ | _0591_;
assign _1146_ = _0592_ | _0593_;
assign _1148_ = _0594_ | _0595_;
assign _1152_ = _0596_ | _0597_;
assign _1154_ = _0598_ | _0599_;
assign _1156_ = _0600_ | _0601_;
assign _1160_ = _0602_ | _0603_;
assign _1162_ = _0604_ | _0605_;
assign _1164_ = _0606_ | _0607_;
assign csr_rdata_o_t0[11] = _0608_ | _0609_;
assign _1166_ = _0610_ | _0611_;
assign _1168_ = _0612_ | _0613_;
assign _1172_ = _0614_ | _0615_;
assign _1174_ = _0616_ | _0617_;
assign _1176_ = _0618_ | _0619_;
assign _1178_ = _0620_ | _0621_;
assign _1180_ = _0622_ | _0623_;
assign _1184_ = _0624_ | _0625_;
assign _1186_ = _0626_ | _0627_;
assign _1188_ = _0628_ | _0629_;
assign _1192_ = _0630_ | _0631_;
assign _1194_ = _0632_ | _0633_;
assign _1196_ = _0634_ | _0635_;
assign csr_rdata_o_t0[21] = _0636_ | _0637_;
assign cpuctrlsts_part_d_t0[7] = _0651_ | _0652_;
assign _0075_ = _0653_ | _0654_;
assign _1252_ = _0655_ | _0656_;
assign _1254_ = _0657_ | _0658_;
assign mstatus_d_t0[4:2] = _0659_ | _0660_;
assign _1256_ = _0661_ | _0662_;
assign _1258_ = _0663_ | _0664_;
assign mstatus_d_t0[1] = _0665_ | _0666_;
assign _1260_ = _0667_ | _0668_;
assign _1262_ = _0669_ | _0670_;
assign mstatus_d_t0[5] = _0671_ | _0672_;
assign _0080_ = _0673_ | _0674_;
assign _0057_ = _0675_ | _0676_;
assign _0059_ = _0677_ | _0678_;
assign _0090_[1] = _0679_ | _0680_;
assign _0097_[1:0] = _0681_ | _0682_;
assign _0097_[2] = _0683_ | _0684_;
assign _0064_ = _0685_ | _0686_;
assign _0024_ = _0687_ | _0688_;
assign _0101_ = _0689_ | _0690_;
assign _0093_ = _0691_ | _0692_;
assign _0066_ = _0693_ | _0694_;
assign _0049_ = _0695_ | _0696_;
assign _0032_ = _0697_ | _0698_;
assign _0036_ = _0699_ | _0700_;
assign _0086_ = _0701_ | _0702_;
assign _1264_ = _0703_ | _0704_;
assign _1266_ = _0705_ | _0706_;
assign _0030_ = _0707_ | _0708_;
assign _1272_ = _0709_ | _0710_;
assign cpuctrlsts_part_d_t0[6] = _0711_ | _0712_;
assign depc_d_t0 = _0713_ | _0714_;
assign dcsr_d_t0[8:6] = _0715_ | _0716_;
assign dcsr_d_t0[1:0] = _0717_ | _0718_;
assign mtval_d_t0 = _0719_ | _0720_;
assign _1276_ = _0721_ | _0722_;
assign _1278_ = _0723_ | _0724_;
assign mcause_d_t0 = _0725_ | _0726_;
assign _1282_ = _0727_ | _0728_;
assign _1284_ = _0729_ | _0730_;
assign mepc_d_t0 = _0731_ | _0732_;
assign _0072_ = _0733_ | _0734_;
assign _1290_ = _0735_ | _0736_;
assign _0046_[5:4] = _0737_ | _0738_;
assign _0046_[3:2] = _0739_ | _0740_;
assign _0021_[15] = _0741_ | _0742_;
assign _0046_[1:0] = _0743_ | _0744_;
assign _0021_[1:0] = _0745_ | _0746_;
assign _0021_[2] = _0747_ | _0748_;
assign _0021_[13:12] = _0749_ | _0750_;
assign _0018_ = _0751_ | _0752_;
assign { _0001_[7:6], cpuctrlsts_part_d_t0[5:0] } = _0753_ | _0754_;
assign { dcsr_d_t0[31:9], _0004_[8:6], dcsr_d_t0[5:2], _0004_[1:0] } = _0755_ | _0756_;
assign mtvec_en_t0 = _0757_ | _0758_;
assign { _0011_[5:1], mstatus_d_t0[0] } = _0759_ | _0760_;
assign mtvec_d_t0 = _0761_ | _0762_;
assign priv_mode_lsu_o_t0 = _0763_ | _0764_;
assign \mhpmcounter[2]_t0  = _0765_ | _0766_;
assign _0265_ = | { csr_save_cause_i, csr_restore_dret_i, csr_restore_mret_i };
assign _0266_ = | { _1352_, _1351_, _1350_, _1349_, _1348_, _1347_, _1346_, _1313_, _1312_, _1311_, _1309_, _1307_, _1306_, _1305_, _1304_, _1303_, _1302_, _1301_, _1300_, _1299_, _1298_, _1297_, _1295_, _1293_, _1292_, _1291_, _1223_, _1217_, _1216_, _1215_, _1214_, _1213_, _1212_, _1211_, _1210_, _1209_, _1208_, _1207_, _1206_, _1205_, _1204_, _1203_, _1202_, _1201_, _1200_, _1199_, _1198_ };
assign _0267_ = | { _1345_, _1344_, _1343_, _1342_, _1341_, _1340_, _1339_, _1338_, _1337_, _1336_, _1335_, _1334_, _1333_, _1332_, _1331_, _1330_, _1329_, _1328_, _1327_, _1326_, _1325_, _1324_, _1323_, _1322_, _1321_, _1320_, _1319_, _1318_, _1317_, _1316_, _1315_, _1314_ };
assign _0268_ = | { _1301_, _1300_, _1299_, _1291_ };
assign _0269_ = | { _1222_, _1250_ };
assign _0270_ = | { _1344_, _1342_, _1341_, _1340_, _1339_, _1338_, _1337_, _1336_, _1335_, _1334_, _1333_, _1332_, _1331_, _1330_, _1329_, _1328_, _1327_, _1326_, _1325_, _1324_, _1323_, _1322_, _1321_, _1320_, _1319_, _1318_, _1317_, _1316_, _1315_, _1314_ };
assign _0173_ = ~ _1346_;
assign _0243_ = ~ _1240_;
assign _0244_ = ~ mcause_q[5];
assign _0245_ = ~ csr_wdata_i;
assign _0246_ = ~ mstatus_err;
assign _0247_ = ~ _1248_;
assign _0248_ = ~ mcause_q[6];
assign _0249_ = ~ csr_rdata_o;
assign _0250_ = ~ debug_mode_entering_i;
assign _0251_ = ~ mtvec_err;
assign _0252_ = ~ cpuctrlsts_part_err;
assign _0638_ = mcause_q_t0[5] & _0248_;
assign _0641_ = csr_wdata_i_t0 & _0249_;
assign _0642_ = debug_mode_i_t0 & _0250_;
assign _0645_ = mstatus_err_t0 & _0251_;
assign _0648_ = _1249_ & _0252_;
assign _1242_ = illegal_csr_dbg_t0 & _0243_;
assign _0639_ = mcause_q_t0[6] & _0244_;
assign _0643_ = debug_mode_entering_i_t0 & _0208_;
assign _0646_ = mtvec_err_t0 & _0246_;
assign _0649_ = cpuctrlsts_part_err_t0 & _0247_;
assign _0640_ = mcause_q_t0[5] & mcause_q_t0[6];
assign _0644_ = debug_mode_i_t0 & debug_mode_entering_i_t0;
assign _0647_ = mstatus_err_t0 & mtvec_err_t0;
assign _0650_ = _1249_ & cpuctrlsts_part_err_t0;
assign _0786_ = _0638_ | _0639_;
assign _0787_ = _0641_ | _0275_;
assign _0788_ = _0642_ | _0643_;
assign _0789_ = _0645_ | _0646_;
assign _0790_ = _0648_ | _0649_;
assign _1244_ = _0786_ | _0640_;
assign _1246_ = _0787_ | _0276_;
assign _1236_ = _0788_ | _0644_;
assign _1249_ = _0789_ | _0647_;
assign csr_shadow_err_o_t0 = _0790_ | _0650_;
assign _0772_ = _1311_ | _1306_;
assign _0769_ = _1294_ | _1297_;
assign _0773_ = _1299_ | _1298_;
assign _0774_ = _1346_ | _1306_;
assign _0777_ = _1305_ | _1304_;
assign _0778_ = _1292_ | _1346_;
assign _0767_ = _1300_ | _1299_;
assign _0768_ = _1306_ | _1302_;
assign _0775_ = _1296_ | _1294_;
assign _0776_ = _1301_ | _1300_;
assign _0770_ = _1304_ | _1303_;
assign _0771_ = _1307_ | _1306_;
assign _0259_ = | { _1309_, _1301_, _1295_, _1291_, _0767_, _0769_ };
assign _0258_ = | { _1312_, _1309_, _1301_, _1295_, _1291_, _0767_, _0769_ };
assign _0256_ = | { _1309_, _1295_, _0769_ };
assign _0260_ = | { _0773_, _1309_, _1301_, _1300_, _1295_, _1291_, _0769_ };
assign _0263_ = | { _1306_, _1302_, _0777_ };
assign _0264_ = | { _0775_, _0776_, _1309_, _1303_, _1299_, _1291_ };
assign _0262_ = | { _0775_, _0776_, _1312_, _1309_, _1299_, _1291_ };
assign _0253_ = | { _1309_, _1295_, _1293_ };
assign _0254_ = | { _1305_, _1304_, _1303_ };
assign _0255_ = | { _1309_, _1301_, _1295_, _1293_, _1291_, _0767_ };
assign _0261_ = | { _0775_, _1309_, _1299_ };
assign _0257_ = | { _1305_, _1302_, _0770_ };
assign _0791_ = _1220_ ? _0106_ : _1245_;
assign dummy_instr_seed_o = _0269_ ? csr_wdata_i : _0791_;
assign _0793_ = _1296_ ? _0014_[31] : _0016_[31];
assign _0795_ = _1294_ ? _0014_[63] : _0793_;
assign _0797_ = _1299_ ? dscratch1_q[31] : dscratch0_q[31];
assign _0799_ = _1301_ ? csr_depc_o[31] : dcsr_q[31];
assign _0801_ = _0767_ ? _0797_ : _0799_;
assign _0803_ = _0253_ ? _0795_ : _0801_;
assign _0805_ = _1304_ ? _1243_ : csr_mepc_o[31];
assign _0807_ = _1303_ ? csr_mtval_o[31] : _0805_;
assign _0809_ = _1302_ ? csr_mtvec_o[31] : mscratch_q[31];
assign _0811_ = _1311_ ? hart_id_i[31] : 1'h0;
assign _0813_ = _0768_ ? _0809_ : _0811_;
assign _0815_ = _0254_ ? _0807_ : _0813_;
assign csr_rdata_o[31] = _0255_ ? _0803_ : _0815_;
assign _0817_ = _1297_ ? cpuctrlsts_part_q[7] : _0014_[39];
assign _0819_ = _1296_ ? _0014_[7] : _0016_[7];
assign _0821_ = _0769_ ? _0817_ : _0819_;
assign _0823_ = _1299_ ? dscratch1_q[7] : dscratch0_q[7];
assign _0825_ = _1291_ ? dcsr_q[7] : irq_timer_i;
assign _0827_ = _1301_ ? csr_depc_o[7] : _0825_;
assign _0829_ = _0767_ ? _0823_ : _0827_;
assign _0831_ = _0256_ ? _0821_ : _0829_;
assign _0833_ = _1303_ ? csr_mtval_o[7] : _1353_[2];
assign _0835_ = _1305_ ? csr_mepc_o[7] : csr_mtvec_o[7];
assign _0837_ = _0770_ ? _0833_ : _0835_;
assign _0839_ = _1306_ ? mscratch_q[7] : mie_q[16];
assign _0841_ = _1311_ ? hart_id_i[7] : 1'h0;
assign _0843_ = _1292_ ? mstatus_q[4] : _0841_;
assign _0845_ = _0771_ ? _0839_ : _0843_;
assign _0847_ = _0257_ ? _0837_ : _0845_;
assign csr_rdata_o[7] = _0258_ ? _0831_ : _0847_;
assign _0849_ = _1297_ ? cpuctrlsts_part_q[6:4] : _0014_[38:36];
assign _0851_ = _1296_ ? _0014_[6:4] : _0016_[6:4];
assign _0853_ = _0769_ ? _0849_ : _0851_;
assign _0855_ = _1299_ ? dscratch1_q[6:4] : dscratch0_q[6:4];
assign _0857_ = _1301_ ? csr_depc_o[6:4] : dcsr_q[6:4];
assign _0859_ = _0767_ ? _0855_ : _0857_;
assign _0861_ = _0256_ ? _0853_ : _0859_;
assign _0863_ = _1303_ ? csr_mtval_o[6:4] : { _1353_[1:0], mcause_q[4] };
assign _0865_ = _1305_ ? csr_mepc_o[6:4] : csr_mtvec_o[6:4];
assign _0867_ = _0770_ ? _0863_ : _0865_;
assign _0869_ = _1306_ ? mscratch_q[6:4] : hart_id_i[6:4];
assign _0871_ = _1313_ ? 3'h1 : 3'h0;
assign _0872_ = _0772_ ? _0869_ : _0871_;
assign _0874_ = _0257_ ? _0867_ : _0872_;
assign csr_rdata_o[6:4] = _0259_ ? _0861_ : _0874_;
assign _0876_ = _1297_ ? cpuctrlsts_part_q[3] : _0014_[35];
assign _0878_ = _1296_ ? _0014_[3] : _0016_[3];
assign _0880_ = _0769_ ? _0876_ : _0878_;
assign _0882_ = _1299_ ? dscratch1_q[3] : dscratch0_q[3];
assign _0884_ = _1291_ ? dcsr_q[3] : irq_software_i;
assign _0886_ = _1301_ ? csr_depc_o[3] : _0884_;
assign _0888_ = _0767_ ? _0882_ : _0886_;
assign _0890_ = _0256_ ? _0880_ : _0888_;
assign _0892_ = _1303_ ? csr_mtval_o[3] : mcause_q[3];
assign _0894_ = _1305_ ? csr_mepc_o[3] : csr_mtvec_o[3];
assign _0896_ = _0770_ ? _0892_ : _0894_;
assign _0898_ = _1306_ ? mscratch_q[3] : mie_q[17];
assign _0900_ = _1311_ ? hart_id_i[3] : 1'h0;
assign _0902_ = _1292_ ? mstatus_q[5] : _0900_;
assign _0904_ = _0771_ ? _0898_ : _0902_;
assign _0906_ = _0257_ ? _0896_ : _0904_;
assign csr_rdata_o[3] = _0258_ ? _0890_ : _0906_;
assign _0908_ = _1297_ ? cpuctrlsts_part_q[2:0] : _0014_[34:32];
assign _0910_ = _1296_ ? _0014_[2:0] : _0016_[2:0];
assign _0912_ = _0769_ ? _0908_ : _0910_;
assign _0914_ = _1298_ ? { mcountinhibit[2], 1'h0, mcountinhibit[0] } : dscratch1_q[2:0];
assign _0916_ = _1301_ ? csr_depc_o[2:0] : dcsr_q[2:0];
assign _0918_ = _1300_ ? dscratch0_q[2:0] : _0916_;
assign _0920_ = _0773_ ? _0914_ : _0918_;
assign _0922_ = _0256_ ? _0912_ : _0920_;
assign _0924_ = _1303_ ? csr_mtval_o[2:0] : mcause_q[2:0];
assign _0926_ = _1305_ ? csr_mepc_o[2:0] : csr_mtvec_o[2:0];
assign _0928_ = _0770_ ? _0924_ : _0926_;
assign _0930_ = _1306_ ? mscratch_q[2:0] : 3'h4;
assign _0932_ = _1313_ ? 3'h6 : 3'h0;
assign _0933_ = _1311_ ? hart_id_i[2:0] : _0932_;
assign _0935_ = _0774_ ? _0930_ : _0933_;
assign _0937_ = _0257_ ? _0928_ : _0935_;
assign csr_rdata_o[2:0] = _0260_ ? _0922_ : _0937_;
assign _0939_ = _1296_ ? _0014_[10:8] : _0016_[10:8];
assign _0941_ = _1294_ ? _0014_[42:40] : _0939_;
assign _0943_ = _1299_ ? dscratch1_q[10:8] : dscratch0_q[10:8];
assign _0945_ = _1301_ ? csr_depc_o[10:8] : dcsr_q[10:8];
assign _0947_ = _0767_ ? _0943_ : _0945_;
assign _0949_ = _0253_ ? _0941_ : _0947_;
assign _0951_ = _1303_ ? csr_mtval_o[10:8] : _1353_[5:3];
assign _0953_ = _1305_ ? csr_mepc_o[10:8] : csr_mtvec_o[10:8];
assign _0955_ = _0770_ ? _0951_ : _0953_;
assign _0957_ = _1306_ ? mscratch_q[10:8] : 3'h1;
assign _0959_ = _1311_ ? hart_id_i[10:8] : 3'h0;
assign _0961_ = _0774_ ? _0957_ : _0959_;
assign _0963_ = _0257_ ? _0955_ : _0961_;
assign csr_rdata_o[10:8] = _0255_ ? _0949_ : _0963_;
assign _0965_ = _1294_ ? _0014_[52:50] : _0014_[20:18];
assign _0967_ = _1310_ ? _0016_[20:18] : dscratch1_q[20:18];
assign _0969_ = _0775_ ? _0965_ : _0967_;
assign _0971_ = _1300_ ? dscratch0_q[20:18] : csr_depc_o[20:18];
assign _0973_ = _1291_ ? dcsr_q[20:18] : irq_fast_i[4:2];
assign _0975_ = _0776_ ? _0971_ : _0973_;
assign _0977_ = _0261_ ? _0969_ : _0975_;
assign _0979_ = _1303_ ? csr_mtval_o[20:18] : _1353_[15:13];
assign _0981_ = _1305_ ? csr_mepc_o[20:18] : csr_mtvec_o[20:18];
assign _0983_ = _0770_ ? _0979_ : _0981_;
assign _0985_ = _1306_ ? mscratch_q[20:18] : mie_q[4:2];
assign _0987_ = _1311_ ? hart_id_i[20:18] : 3'h0;
assign _0989_ = _1346_ ? 3'h4 : _0987_;
assign _0991_ = _0771_ ? _0985_ : _0989_;
assign _0993_ = _0257_ ? _0983_ : _0991_;
assign csr_rdata_o[20:18] = _0262_ ? _0977_ : _0993_;
assign _0995_ = _1294_ ? _0014_[44] : _0014_[12];
assign _0997_ = _1310_ ? _0016_[12] : dscratch1_q[12];
assign _0999_ = _0775_ ? _0995_ : _0997_;
assign _1001_ = _1300_ ? dscratch0_q[12] : csr_depc_o[12];
assign _1003_ = _1291_ ? dcsr_q[12] : csr_mtval_o[12];
assign _1005_ = _0776_ ? _1001_ : _1003_;
assign _1007_ = _0261_ ? _0999_ : _1005_;
assign _1009_ = _1304_ ? _1353_[7] : csr_mepc_o[12];
assign _1011_ = _1302_ ? csr_mtvec_o[12] : mscratch_q[12];
assign _1013_ = _0777_ ? _1009_ : _1011_;
assign _1015_ = _1346_ ? 1'h1 : mstatus_q[3];
assign _1017_ = _1311_ ? hart_id_i[12] : 1'h0;
assign _1019_ = _0778_ ? _1015_ : _1017_;
assign _1021_ = _0263_ ? _1013_ : _1019_;
assign csr_rdata_o[12] = _0264_ ? _1007_ : _1021_;
assign _1023_ = _1294_ ? _0014_[49] : _0014_[17];
assign _1025_ = _1310_ ? _0016_[17] : dscratch1_q[17];
assign _1027_ = _0775_ ? _1023_ : _1025_;
assign _1029_ = _1300_ ? dscratch0_q[17] : csr_depc_o[17];
assign _1031_ = _1291_ ? dcsr_q[17] : irq_fast_i[1];
assign _1033_ = _0776_ ? _1029_ : _1031_;
assign _1035_ = _0261_ ? _1027_ : _1033_;
assign _1037_ = _1303_ ? csr_mtval_o[17] : _1353_[12];
assign _1039_ = _1305_ ? csr_mepc_o[17] : csr_mtvec_o[17];
assign _1041_ = _0770_ ? _1037_ : _1039_;
assign _1043_ = _1306_ ? mscratch_q[17] : mie_q[1];
assign _1045_ = _1311_ ? hart_id_i[17] : 1'h0;
assign _1047_ = _1292_ ? mstatus_q[1] : _1045_;
assign _1049_ = _0771_ ? _1043_ : _1047_;
assign _1051_ = _0257_ ? _1041_ : _1049_;
assign csr_rdata_o[17] = _0262_ ? _1035_ : _1051_;
assign _1053_ = _1296_ ? _0014_[15:13] : _0016_[15:13];
assign _1055_ = _1294_ ? _0014_[47:45] : _1053_;
assign _1057_ = _1299_ ? dscratch1_q[15:13] : dscratch0_q[15:13];
assign _1059_ = _1301_ ? csr_depc_o[15:13] : dcsr_q[15:13];
assign _1061_ = _0767_ ? _1057_ : _1059_;
assign _1063_ = _0253_ ? _1055_ : _1061_;
assign _1065_ = _1304_ ? _1353_[10:8] : csr_mepc_o[15:13];
assign _1067_ = _1303_ ? csr_mtval_o[15:13] : _1065_;
assign _1069_ = _1302_ ? csr_mtvec_o[15:13] : mscratch_q[15:13];
assign _1071_ = _1311_ ? hart_id_i[15:13] : 3'h0;
assign _1073_ = _0768_ ? _1069_ : _1071_;
assign _1075_ = _0254_ ? _1067_ : _1073_;
assign csr_rdata_o[15:13] = _0255_ ? _1063_ : _1075_;
assign _1077_ = _1294_ ? _0014_[48] : _0014_[16];
assign _1079_ = _1310_ ? _0016_[16] : dscratch1_q[16];
assign _1081_ = _0775_ ? _1077_ : _1079_;
assign _1083_ = _1300_ ? dscratch0_q[16] : csr_depc_o[16];
assign _1085_ = _1291_ ? dcsr_q[16] : irq_fast_i[0];
assign _1087_ = _0776_ ? _1083_ : _1085_;
assign _1089_ = _0261_ ? _1081_ : _1087_;
assign _1091_ = _1303_ ? csr_mtval_o[16] : _1353_[11];
assign _1093_ = _1305_ ? csr_mepc_o[16] : csr_mtvec_o[16];
assign _1095_ = _0770_ ? _1091_ : _1093_;
assign _1097_ = _1306_ ? mscratch_q[16] : mie_q[0];
assign _1099_ = _1311_ ? hart_id_i[16] : 1'h0;
assign _1101_ = _0771_ ? _1097_ : _1099_;
assign _1103_ = _0257_ ? _1095_ : _1101_;
assign csr_rdata_o[16] = _0262_ ? _1089_ : _1103_;
assign _1105_ = _1294_ ? _0014_[62:54] : _0014_[30:22];
assign _1107_ = _1310_ ? _0016_[30:22] : dscratch1_q[30:22];
assign _1109_ = _0775_ ? _1105_ : _1107_;
assign _1111_ = _1300_ ? dscratch0_q[30:22] : csr_depc_o[30:22];
assign _1113_ = _1291_ ? dcsr_q[30:22] : irq_fast_i[14:6];
assign _1115_ = _0776_ ? _1111_ : _1113_;
assign _1117_ = _0261_ ? _1109_ : _1115_;
assign _1119_ = _1303_ ? csr_mtval_o[30:22] : _1353_[25:17];
assign _1121_ = _1305_ ? csr_mepc_o[30:22] : csr_mtvec_o[30:22];
assign _1123_ = _0770_ ? _1119_ : _1121_;
assign _1125_ = _1306_ ? mscratch_q[30:22] : mie_q[14:6];
assign _1127_ = _1311_ ? hart_id_i[30:22] : 9'h000;
assign _1129_ = _1346_ ? 9'h100 : _1127_;
assign _1131_ = _0771_ ? _1125_ : _1129_;
assign _1133_ = _0257_ ? _1123_ : _1131_;
assign csr_rdata_o[30:22] = _0262_ ? _1117_ : _1133_;
assign _1135_ = _1294_ ? _0014_[43] : _0014_[11];
assign _1137_ = _1310_ ? _0016_[11] : dscratch1_q[11];
assign _1139_ = _0775_ ? _1135_ : _1137_;
assign _1141_ = _1300_ ? dscratch0_q[11] : csr_depc_o[11];
assign _1143_ = _1291_ ? dcsr_q[11] : irq_external_i;
assign _1145_ = _0776_ ? _1141_ : _1143_;
assign _1147_ = _0261_ ? _1139_ : _1145_;
assign _1149_ = _1303_ ? csr_mtval_o[11] : _1353_[6];
assign _1151_ = _1305_ ? csr_mepc_o[11] : csr_mtvec_o[11];
assign _1153_ = _0770_ ? _1149_ : _1151_;
assign _1155_ = _1306_ ? mscratch_q[11] : mie_q[15];
assign _1157_ = _1311_ ? hart_id_i[11] : 1'h0;
assign _1159_ = _1292_ ? mstatus_q[2] : _1157_;
assign _1161_ = _0771_ ? _1155_ : _1159_;
assign _1163_ = _0257_ ? _1153_ : _1161_;
assign csr_rdata_o[11] = _0262_ ? _1147_ : _1163_;
assign _1165_ = _1343_ ? \mhpmcounter[2]  : \mhpmcounter[0] ;
assign _0014_ = _0270_ ? 64'h0000000000000000 : _1165_;
assign _1167_ = _1294_ ? _0014_[53] : _0014_[21];
assign _1169_ = _1310_ ? _0016_[21] : dscratch1_q[21];
assign _1171_ = _0775_ ? _1167_ : _1169_;
assign _1173_ = _1300_ ? dscratch0_q[21] : csr_depc_o[21];
assign _1175_ = _1291_ ? dcsr_q[21] : irq_fast_i[5];
assign _1177_ = _0776_ ? _1173_ : _1175_;
assign _1179_ = _0261_ ? _1171_ : _1177_;
assign _1181_ = _1303_ ? csr_mtval_o[21] : _1353_[16];
assign _1183_ = _1305_ ? csr_mepc_o[21] : csr_mtvec_o[21];
assign _1185_ = _0770_ ? _1181_ : _1183_;
assign _1187_ = _1306_ ? mscratch_q[21] : mie_q[5];
assign _1189_ = _1311_ ? hart_id_i[21] : 1'h0;
assign _1191_ = _1292_ ? mstatus_q[0] : _1189_;
assign _1193_ = _0771_ ? _1187_ : _1191_;
assign _1195_ = _0257_ ? _1185_ : _1193_;
assign csr_rdata_o[21] = _0262_ ? _1179_ : _1195_;
assign _1238_ = 1'h0 >> _1232_;
assign _1197_ = csr_addr_i[11:10] == /* src = "generated/sv2v_out.v:14000.30-14000.54" */ 2'h3;
assign _1218_ = dummy_instr_seed_o[31:30] == /* src = "generated/sv2v_out.v:14169.46-14169.75" */ 2'h2;
assign _1219_ = dummy_instr_seed_o[31:30] == /* src = "generated/sv2v_out.v:14169.15-14169.44" */ 2'h3;
assign illegal_csr_priv = csr_addr_i[9:8] > /* src = "generated/sv2v_out.v:13999.28-13999.56" */ priv_mode_id_o;
assign illegal_csr_write = _1197_ && /* src = "generated/sv2v_out.v:14000.29-14000.65" */ csr_wr;
assign _1224_ = _1227_ && /* src = "generated/sv2v_out.v:14196.10-14196.66" */ _1228_;
assign _1225_ = _1229_ && /* src = "generated/sv2v_out.v:14208.10-14208.60" */ _1230_;
assign dummy_instr_seed_en_o = csr_we_int && /* src = "generated/sv2v_out.v:14866.35-14866.70" */ _1223_;
assign _1226_ = csr_mcause_i[5] || /* src = "generated/sv2v_out.v:14263.12-14263.38" */ csr_mcause_i[6];
assign _1227_ = dummy_instr_seed_o[12:11] != /* src = "generated/sv2v_out.v:14196.11-14196.35" */ 2'h3;
assign _1228_ = | /* src = "generated/sv2v_out.v:14196.41-14196.65" */ dummy_instr_seed_o[12:11];
assign _1229_ = dummy_instr_seed_o[1:0] != /* src = "generated/sv2v_out.v:14208.11-14208.32" */ 2'h3;
assign _1230_ = | /* src = "generated/sv2v_out.v:14208.38-14208.59" */ dummy_instr_seed_o[1:0];
assign _1231_ = mstatus_q[3:2] != /* src = "generated/sv2v_out.v:14278.9-14278.33" */ 2'h3;
assign _1232_ = - /* src = "generated/sv2v_out.v:0.0-0.0" */ $signed({ 27'h0000000, csr_addr_i[4:0] });
assign _1233_ = ~ /* src = "generated/sv2v_out.v:14315.47-14315.66" */ illegal_csr_insn_o;
assign _0109_ = ~ /* src = "generated/sv2v_out.v:14687.40-14687.57" */ mcountinhibit[0];
assign _1234_ = ~ /* src = "generated/sv2v_out.v:14706.46-14706.63" */ mcountinhibit[2];
assign _1235_ = ~ /* src = "generated/sv2v_out.v:14910.50-14910.89" */ _1247_;
assign _1239_ = illegal_csr | /* src = "generated/sv2v_out.v:14001.48-14001.79" */ illegal_csr_write;
assign _1240_ = _1239_ | /* src = "generated/sv2v_out.v:14001.47-14001.99" */ illegal_csr_priv;
assign _1241_ = _1240_ | /* src = "generated/sv2v_out.v:14001.46-14001.118" */ illegal_csr_dbg;
assign _1243_ = mcause_q[5] | /* src = "generated/sv2v_out.v:14056.30-14056.55" */ mcause_q[6];
assign _1245_ = csr_wdata_i | /* src = "generated/sv2v_out.v:14309.26-14309.51" */ csr_rdata_o;
assign _1247_ = debug_mode_i | /* src = "generated/sv2v_out.v:14910.52-14910.88" */ debug_mode_entering_i;
assign _1248_ = mstatus_err | /* src = "generated/sv2v_out.v:14923.31-14923.54" */ mtvec_err;
assign csr_shadow_err_o = _1248_ | /* src = "generated/sv2v_out.v:14923.29-14923.92" */ cpuctrlsts_part_err;
assign _1250_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14307.3-14313.10" */ csr_op_i;
assign _1220_ = csr_op_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14307.3-14313.10" */ 2'h3;
assign _1221_ = csr_op_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14307.3-14313.10" */ 2'h2;
assign _1222_ = csr_op_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14307.3-14313.10" */ 2'h1;
assign cpuctrlsts_part_d[7] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0065_[1] : _0000_[7];
assign _0094_ = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14282.9-14282.19|generated/sv2v_out.v:14282.5-14293.8" */ 1'h1 : _0008_;
assign _0074_ = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14282.9-14282.19|generated/sv2v_out.v:14282.5-14293.8" */ mstack_epc_q : { dummy_instr_seed_o[31:1], 1'h0 };
assign _0095_ = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14282.9-14282.19|generated/sv2v_out.v:14282.5-14293.8" */ 1'h1 : _0009_;
assign _0104_[1:0] = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14282.9-14282.19|generated/sv2v_out.v:14282.5-14293.8" */ mstack_q[1:0] : 2'h0;
assign _0104_[2] = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14282.9-14282.19|generated/sv2v_out.v:14282.5-14293.8" */ mstack_q[2] : 1'h1;
assign _0102_ = _1231_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14278.9-14278.33|generated/sv2v_out.v:14278.5-14279.26" */ 1'h0 : _0010_[1];
assign _1251_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0104_ : _0010_[4:2];
assign _1253_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0010_[4:2] : _1251_;
assign mstatus_d[4:2] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0085_[2:0] : _1253_;
assign _1255_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0102_ : _0010_[1];
assign _1257_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0010_[1] : _1255_;
assign mstatus_d[1] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0010_[1] : _1257_;
assign _1259_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ mstatus_q[4] : _0010_[5];
assign _1261_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0010_[5] : _1259_;
assign mstatus_d[5] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0085_[3] : _1261_;
assign _0082_ = cpuctrlsts_part_q[6] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14266.11-14266.31|generated/sv2v_out.v:14266.7-14269.10" */ 1'h1 : 1'h0;
assign _0089_[0] = _1226_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14263.10-14263.39|generated/sv2v_out.v:14263.6-14270.9" */ _0000_[6] : 1'h1;
assign _0070_ = _1226_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14263.10-14263.39|generated/sv2v_out.v:14263.6-14270.9" */ 1'h0 : _0082_;
assign _0098_ = cpuctrlsts_part_q[6] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14266.11-14266.31|generated/sv2v_out.v:14266.7-14269.10" */ 1'h1 : _0000_[7];
assign _0091_ = _1226_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14263.10-14263.39|generated/sv2v_out.v:14263.6-14270.9" */ _0002_ : 1'h1;
assign _0081_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14251.14-14251.27|generated/sv2v_out.v:14251.10-14271.8" */ _0002_ : _0091_;
assign _0079_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14251.14-14251.27|generated/sv2v_out.v:14251.10-14271.8" */ _0000_[7:6] : _0089_;
assign _0055_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14251.14-14251.27|generated/sv2v_out.v:14251.10-14271.8" */ 1'h0 : _0070_;
assign _0060_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14251.14-14251.27|generated/sv2v_out.v:14251.10-14271.8" */ 1'h0 : 1'h1;
assign _0056_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14251.14-14251.27|generated/sv2v_out.v:14251.10-14271.8" */ { _1219_, _1218_, dummy_instr_seed_o[4:0] } : csr_mcause_i;
assign _0083_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14251.14-14251.27|generated/sv2v_out.v:14251.10-14271.8" */ _0008_ : 1'h1;
assign _0058_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14251.14-14251.27|generated/sv2v_out.v:14251.10-14271.8" */ { dummy_instr_seed_o[31:1], 1'h0 } : _0029_;
assign _0084_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14251.14-14251.27|generated/sv2v_out.v:14251.10-14271.8" */ _0009_ : 1'h1;
assign _0089_[1] = _1226_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14263.10-14263.39|generated/sv2v_out.v:14263.6-14270.9" */ _0000_[7] : _0098_;
assign _0096_[1:0] = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14251.14-14251.27|generated/sv2v_out.v:14251.10-14271.8" */ _0010_[3:2] : priv_mode_id_o;
assign _0096_[2] = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14251.14-14251.27|generated/sv2v_out.v:14251.10-14271.8" */ _0010_[4] : mstatus_q[5];
assign _0087_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14251.14-14251.27|generated/sv2v_out.v:14251.10-14271.8" */ _0012_ : 1'h1;
assign _0063_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14251.14-14251.27|generated/sv2v_out.v:14251.10-14271.8" */ dummy_instr_seed_o : csr_mtval_i;
assign _0088_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14251.14-14251.27|generated/sv2v_out.v:14251.10-14271.8" */ _0013_ : 1'h1;
assign _0069_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ 1'h1 : _0006_;
assign _0023_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ _0029_ : { dummy_instr_seed_o[31:1], 1'h0 };
assign _0068_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ 1'h1 : _0005_;
assign _0100_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ debug_cause_i : _0003_[8:6];
assign _0092_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ priv_mode_id_o : _0003_[1:0];
assign _0067_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ _0002_ : _0081_;
assign _0065_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ _0000_[7:6] : _0079_;
assign _0044_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ 1'h0 : _0060_;
assign _0078_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ _0013_ : _0088_;
assign _0048_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ dummy_instr_seed_o : _0063_;
assign _0073_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ _0008_ : _0083_;
assign _0031_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ { _1219_, _1218_, dummy_instr_seed_o[4:0] } : _0056_;
assign _0076_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ _0009_ : _0084_;
assign _0035_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ { dummy_instr_seed_o[31:1], 1'h0 } : _0058_;
assign _0077_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ _0012_ : _0087_;
assign _0085_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ _0010_[5:2] : _0096_;
assign _0026_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14244.9-14244.25|generated/sv2v_out.v:14244.5-14271.8" */ 1'h0 : _0055_;
assign _1263_ = csr_save_wb_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14236.5-14242.12" */ pc_wb_i : pc_id_i;
assign _1265_ = csr_save_id_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14236.5-14242.12" */ pc_id_i : _1263_;
assign _0029_ = csr_save_if_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14236.5-14242.12" */ pc_if_i : _1265_;
assign _1267_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ 1'h1 : _0002_;
assign _1268_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0002_ : _1267_;
assign cpuctrlsts_part_we = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0067_ : _1268_;
assign _1269_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ 1'h0 : _0000_[6];
assign _1271_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0000_[6] : _1269_;
assign cpuctrlsts_part_d[6] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0065_[0] : _1271_;
assign mstack_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0044_ : 1'h0;
assign depc_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0069_ : _0006_;
assign depc_d = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0023_ : { dummy_instr_seed_o[31:1], 1'h0 };
assign dcsr_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0068_ : _0005_;
assign dcsr_d[8:6] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0100_ : _0003_[8:6];
assign dcsr_d[1:0] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0092_ : _0003_[1:0];
assign mtval_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0078_ : _0013_;
assign mtval_d = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0048_ : dummy_instr_seed_o;
assign _1273_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0094_ : _0008_;
assign _1274_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0008_ : _1273_;
assign mcause_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0073_ : _1274_;
assign _1275_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0071_ : { _1219_, _1218_, dummy_instr_seed_o[4:0] };
assign _1277_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ { _1219_, _1218_, dummy_instr_seed_o[4:0] } : _1275_;
assign mcause_d = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0031_ : _1277_;
assign _1279_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0095_ : _0009_;
assign _1280_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0009_ : _1279_;
assign mepc_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0076_ : _1280_;
assign _1281_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0074_ : { dummy_instr_seed_o[31:1], 1'h0 };
assign _1283_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ { dummy_instr_seed_o[31:1], 1'h0 } : _1281_;
assign mepc_d = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0035_ : _1283_;
assign _1285_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ 1'h1 : _0012_;
assign _1286_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0012_ : _1285_;
assign mstatus_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0077_ : _1286_;
assign _0071_ = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14282.9-14282.19|generated/sv2v_out.v:14282.5-14293.8" */ mstack_cause_q : { _1219_, _1218_, dummy_instr_seed_o[4:0] };
assign double_fault_seen_o = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ _0026_ : 1'h0;
assign _1287_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ mstatus_q[3:2] : 2'hx;
assign _1289_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ dcsr_q[1:0] : _1287_;
assign priv_lvl_d = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14234.3-14297.10" */ 2'h3 : _1289_;
assign _0096_[3] = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14251.14-14251.27|generated/sv2v_out.v:14251.10-14271.8" */ _0010_[5] : 1'h0;
assign _0020_[31:28] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 4'h4 : dcsr_q[31:28];
assign _0045_[5:4] = _1292_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ { dummy_instr_seed_o[3], dummy_instr_seed_o[7] } : mstatus_q[5:4];
assign _0045_[3:2] = _1292_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ _0061_ : mstatus_q[3:2];
assign _0020_[15] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ dummy_instr_seed_o[15] : dcsr_q[15];
assign _0020_[14] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h0 : dcsr_q[14];
assign _0020_[27:16] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 12'h000 : dcsr_q[27:16];
assign _0045_[1:0] = _1292_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ { dummy_instr_seed_o[17], dummy_instr_seed_o[21] } : mstatus_q[1:0];
assign _0020_[1:0] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ _0053_ : dcsr_q[1:0];
assign _0020_[5] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h0 : dcsr_q[5];
assign _0020_[4] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h0 : dcsr_q[4];
assign _0020_[3] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h0 : dcsr_q[3];
assign _0020_[2] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ dummy_instr_seed_o[2] : dcsr_q[2];
assign _0020_[13:12] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ dummy_instr_seed_o[13:12] : dcsr_q[13:12];
assign _0020_[11] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h0 : dcsr_q[11];
assign _0053_ = _1225_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14208.10-14208.60|generated/sv2v_out.v:14208.6-14209.28" */ 2'h0 : dummy_instr_seed_o[1:0];
assign _0020_[9] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h0 : dcsr_q[9];
assign _0061_ = _1224_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14196.10-14196.66|generated/sv2v_out.v:14196.6-14197.31" */ 2'h0 : dummy_instr_seed_o[12:11];
assign _0047_ = _1292_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h1 : 1'h0;
assign _1296_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ _1295_;
assign _0019_ = _1297_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h1 : 1'h0;
assign _0017_ = _1297_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ { dummy_instr_seed_o[7:1], 1'h0 } : cpuctrlsts_part_q;
assign _0040_ = _1294_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ _1237_ : 32'd0;
assign _0038_ = _1296_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ _1237_ : 32'd0;
assign _0034_ = _1298_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h1 : 1'h0;
assign _0028_ = _1299_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h1 : 1'h0;
assign _0027_ = _1300_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h1 : 1'h0;
assign _0025_ = _1301_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h1 : 1'h0;
assign _0022_ = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h1 : 1'h0;
assign _0020_[10] = _1291_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h0 : dcsr_q[10];
assign _0051_ = _1302_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h1 : csr_mtvec_init_i;
assign _0050_ = _1303_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h1 : 1'h0;
assign _0033_ = _1304_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h1 : 1'h0;
assign _0037_ = _1305_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h1 : 1'h0;
assign _0043_ = _1306_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h1 : 1'h0;
assign _0042_ = _1307_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14192.4-14233.11" */ 1'h1 : 1'h0;
assign _0002_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0019_ : 1'h0;
assign { _0000_[7:6], cpuctrlsts_part_d[5:0] } = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0017_ : cpuctrlsts_part_q;
assign mhpmcounterh_we = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0040_ : 32'd0;
assign mhpmcounter_we = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0038_ : 32'd0;
assign mcountinhibit_we = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0034_ : 1'h0;
assign dscratch1_en = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0028_ : 1'h0;
assign dscratch0_en = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0027_ : 1'h0;
assign _0006_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0025_ : 1'h0;
assign _0005_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0022_ : 1'h0;
assign { dcsr_d[31:9], _0003_[8:6], dcsr_d[5:2], _0003_[1:0] } = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ { _0020_[31:9], dcsr_q[8:6], _0020_[5:0] } : dcsr_q;
assign mtvec_en = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0051_ : csr_mtvec_init_i;
assign _0013_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0050_ : 1'h0;
assign _0008_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0033_ : 1'h0;
assign _0009_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0037_ : 1'h0;
assign mscratch_en = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0043_ : 1'h0;
assign mie_en = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0042_ : 1'h0;
assign _0012_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0047_ : 1'h0;
assign { _0010_[5:1], mstatus_d[0] } = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14191.7-14191.17|generated/sv2v_out.v:14191.3-14233.11" */ _0045_ : mstatus_q;
assign illegal_csr = _1308_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14152.8-14152.429|generated/sv2v_out.v:14152.4-14153.24" */ 1'h1 : _0007_;
assign _0016_ = _0267_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 32'd0 : 32'hxxxxxxxx;
assign _1294_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ _1293_;
assign _1298_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h320;
assign _1313_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hf12;
assign _1310_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ _1309_;
assign _1346_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h301;
assign _1314_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1f;
assign _1315_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1e;
assign _1316_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1d;
assign _1317_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1c;
assign _1318_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1b;
assign _1319_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1a;
assign _1320_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h19;
assign _1321_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h18;
assign _1322_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h17;
assign _1323_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h16;
assign _1324_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h15;
assign _1325_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h14;
assign _1326_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h13;
assign _1327_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h12;
assign _1328_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h11;
assign _1329_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h10;
assign _1330_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0f;
assign _1331_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0e;
assign _1332_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0d;
assign _1333_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0c;
assign _1334_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0b;
assign _1335_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0a;
assign _1336_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h09;
assign _1337_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h08;
assign _1338_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h07;
assign _1339_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h06;
assign _1340_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h05;
assign _1341_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h04;
assign _1342_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h03;
assign _1343_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h02;
assign _1344_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h01;
assign _1345_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ csr_addr_i[4:0];
assign _1299_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h7b3;
assign _1300_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h7b2;
assign _1301_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h7b1;
assign _1291_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h7b0;
assign _1198_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3bf;
assign _1199_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3be;
assign _1200_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3bd;
assign _1201_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3bc;
assign _1202_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3bb;
assign _1203_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3ba;
assign _1204_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3b9;
assign _1205_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3b8;
assign _1206_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3b7;
assign _1207_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3b6;
assign _1208_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3b5;
assign _1209_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3b4;
assign _1210_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3b3;
assign _1211_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3b2;
assign _1212_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3b1;
assign _1213_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3b0;
assign _1214_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3a3;
assign _1215_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3a2;
assign _1216_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3a1;
assign _1217_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h3a0;
assign _1312_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h344;
assign _1303_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h343;
assign _1304_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h342;
assign _1305_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h341;
assign _1302_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h305;
assign _1306_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h340;
assign _1307_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h304;
assign _1292_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h300;
assign _1311_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hf14;
assign _1295_[1] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb02;
assign _1295_[10] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb0b;
assign _1295_[11] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb0c;
assign _1295_[12] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb0d;
assign _1295_[13] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb0e;
assign _1295_[14] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb0f;
assign _1295_[15] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb10;
assign _1295_[16] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb11;
assign _1295_[17] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb12;
assign _1295_[18] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb13;
assign _1295_[19] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb14;
assign _1295_[2] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb03;
assign _1295_[20] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb15;
assign _1295_[21] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb16;
assign _1295_[22] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb17;
assign _1295_[23] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb18;
assign _1295_[24] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb19;
assign _1295_[25] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb1a;
assign _1295_[26] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb1b;
assign _1295_[27] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb1c;
assign _1295_[28] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb1d;
assign _1295_[29] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb1e;
assign _1295_[3] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb04;
assign _1295_[30] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb1f;
assign _1295_[4] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb05;
assign _1295_[5] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb06;
assign _1295_[6] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb07;
assign _1295_[7] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb08;
assign _1295_[8] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb09;
assign _1295_[9] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb0a;
assign _1309_[0] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h323;
assign _1309_[1] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h324;
assign _1309_[10] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h32d;
assign _1309_[11] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h32e;
assign _1309_[12] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h32f;
assign _1309_[13] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h330;
assign _1309_[14] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h331;
assign _1309_[15] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h332;
assign _1309_[16] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h333;
assign _1309_[17] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h334;
assign _1309_[18] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h335;
assign _1309_[19] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h336;
assign _1309_[2] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h325;
assign _1309_[20] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h337;
assign _1309_[21] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h338;
assign _1309_[22] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h339;
assign _1309_[23] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h33a;
assign _1309_[24] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h33b;
assign _1309_[25] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h33c;
assign _1309_[26] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h33d;
assign _1309_[27] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h33e;
assign _1309_[28] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h33f;
assign _1309_[3] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h326;
assign _1309_[4] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h327;
assign _1309_[5] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h328;
assign _1309_[6] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h329;
assign _1309_[7] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h32a;
assign _1309_[8] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h32b;
assign _1309_[9] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h32c;
assign _0007_ = _0266_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 1'h0 : 1'h1;
assign _1223_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h7c1;
assign _1297_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h7c0;
assign _1293_[0] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb80;
assign _1293_[1] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb82;
assign _1293_[10] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb8b;
assign _1293_[11] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb8c;
assign _1293_[12] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb8d;
assign _1293_[13] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb8e;
assign _1293_[14] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb8f;
assign _1293_[15] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb90;
assign _1293_[16] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb91;
assign _1293_[17] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb92;
assign _1293_[18] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb93;
assign _1293_[19] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb94;
assign _1293_[2] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb83;
assign _1293_[20] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb95;
assign _1293_[21] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb96;
assign _1293_[22] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb97;
assign _1293_[23] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb98;
assign _1293_[24] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb99;
assign _1293_[25] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb9a;
assign _1293_[26] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb9b;
assign _1293_[27] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb9c;
assign _1293_[28] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb9d;
assign _1293_[29] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb9e;
assign _1293_[3] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb84;
assign _1293_[30] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb9f;
assign _1293_[4] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb85;
assign _1293_[5] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb86;
assign _1293_[6] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb87;
assign _1293_[7] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb88;
assign _1293_[8] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb89;
assign _1293_[9] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb8a;
assign _1295_[0] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hb00;
assign _1347_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h306;
assign _1348_[0] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h30a;
assign _1348_[1] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h31a;
assign _1349_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'h310;
assign _1350_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hf15;
assign _1351_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hf13;
assign _1352_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 12'hf11;
assign dbg_csr = _0268_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14028.3-14150.10" */ 1'h1 : 1'h0;
assign _1308_ = | /* src = "generated/sv2v_out.v:14152.8-14152.429" */ { _1217_, _1216_, _1215_, _1214_, _1213_, _1212_, _1211_, _1210_, _1209_, _1208_, _1207_, _1206_, _1205_, _1204_, _1203_, _1202_, _1201_, _1200_, _1199_, _1198_ };
assign csr_wr = | /* src = "generated/sv2v_out.v:14314.18-14314.73" */ { _1222_, _1221_, _1220_ };
assign irq_pending_o = | /* src = "generated/sv2v_out.v:14327.25-14327.32" */ irqs_o;
assign _1237_ = $signed(_1232_) < 0 ? 1'h1 << - _1232_ : 1'h1 >> _1232_;
assign _1353_ = mcause_q[6] ? /* src = "generated/sv2v_out.v:14056.58-14056.116" */ 26'h3ffffff : 26'h0000000;
assign mtvec_d = csr_mtvec_init_i ? /* src = "generated/sv2v_out.v:14173.14-14173.112" */ { boot_addr_i[31:8], 8'h01 } : { dummy_instr_seed_o[31:8], 8'h01 };
assign priv_mode_lsu_o = mstatus_q[1] ? /* src = "generated/sv2v_out.v:14305.28-14305.71" */ mstatus_q[3:2] : priv_mode_id_o;
assign \mhpmcounter[2]  = _0112_ ? /* src = "generated/sv2v_out.v:14706.27-14706.94" */ minstret_next : minstret_raw;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14684.36-14692.3" */
\$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000  mcycle_counter_i (
.clk_i(clk_i),
.counter_inc_i(_0109_),
.counter_inc_i_t0(mcountinhibit_t0[0]),
.counter_val_i(dummy_instr_seed_o),
.counter_val_i_t0(dummy_instr_seed_o_t0),
.counter_val_o(\mhpmcounter[0] ),
.counter_val_o_t0(\mhpmcounter[0]_t0 ),
.counter_we_i(mhpmcounter_we[0]),
.counter_we_i_t0(mhpmcounter_we_t0[0]),
.counterh_we_i(mhpmcounterh_we[0]),
.counterh_we_i_t0(mhpmcounterh_we_t0[0]),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14696.4-14705.3" */
\$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter  minstret_counter_i (
.clk_i(clk_i),
.counter_inc_i(_0110_),
.counter_inc_i_t0(_0111_),
.counter_val_i(dummy_instr_seed_o),
.counter_val_i_t0(dummy_instr_seed_o_t0),
.counter_val_o(minstret_raw),
.counter_val_o_t0(minstret_raw_t0),
.counter_val_upd_o(minstret_next),
.counter_val_upd_o_t0(minstret_next_t0),
.counter_we_i(mhpmcounter_we[2]),
.counter_we_i_t0(mhpmcounter_we_t0[2]),
.counterh_we_i(mhpmcounterh_we[2]),
.counterh_we_i_t0(mhpmcounterh_we_t0[2]),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14915.4-14922.3" */
\$paramod$a088b13b9337f1e1fba58a671f47d7c7701ffa49\ibex_csr  u_cpuctrlsts_part_csr (
.clk_i(clk_i),
.rd_data_o(cpuctrlsts_part_q),
.rd_data_o_t0(cpuctrlsts_part_q_t0),
.rd_error_o(cpuctrlsts_part_err),
.rd_error_o_t0(cpuctrlsts_part_err_t0),
.rst_ni(rst_ni),
.wr_data_i(cpuctrlsts_part_d),
.wr_data_i_t0(cpuctrlsts_part_d_t0),
.wr_en_i(cpuctrlsts_part_we),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14417.4-14423.3" */
\$paramod$9a435d8f6db004a67362aa9a56f32ea481a74dbe\ibex_csr  u_dcsr_csr (
.clk_i(clk_i),
.rd_data_o(dcsr_q),
.rd_data_o_t0(dcsr_q_t0),
.rst_ni(rst_ni),
.wr_data_i(dcsr_d),
.wr_data_i_t0(dcsr_d_t0),
.wr_en_i(dcsr_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14428.4-14434.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_depc_csr (
.clk_i(clk_i),
.rd_data_o(csr_depc_o),
.rd_data_o_t0(csr_depc_o_t0),
.rst_ni(rst_ni),
.wr_data_i(depc_d),
.wr_data_i_t0(depc_d_t0),
.wr_en_i(depc_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14439.4-14445.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_dscratch0_csr (
.clk_i(clk_i),
.rd_data_o(dscratch0_q),
.rd_data_o_t0(dscratch0_q_t0),
.rst_ni(rst_ni),
.wr_data_i(dummy_instr_seed_o),
.wr_data_i_t0(dummy_instr_seed_o_t0),
.wr_en_i(dscratch0_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14450.4-14456.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_dscratch1_csr (
.clk_i(clk_i),
.rd_data_o(dscratch1_q),
.rd_data_o_t0(dscratch1_q_t0),
.rst_ni(rst_ni),
.wr_data_i(dummy_instr_seed_o),
.wr_data_i_t0(dummy_instr_seed_o_t0),
.wr_en_i(dscratch1_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14382.4-14388.3" */
\$paramod$34601000fe8707ce2501f5ed778e152043201712\ibex_csr  u_mcause_csr (
.clk_i(clk_i),
.rd_data_o(mcause_q),
.rd_data_o_t0(mcause_q_t0),
.rst_ni(rst_ni),
.wr_data_i(mcause_d),
.wr_data_i_t0(mcause_d_t0),
.wr_en_i(mcause_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14345.4-14351.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_mepc_csr (
.clk_i(clk_i),
.rd_data_o(csr_mepc_o),
.rd_data_o_t0(csr_mepc_o_t0),
.rst_ni(rst_ni),
.wr_data_i(mepc_d),
.wr_data_i_t0(mepc_d_t0),
.wr_en_i(mepc_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14360.4-14366.3" */
\$paramod$e55993a14b1fbc43320d549f521b710ed37596c6\ibex_csr  u_mie_csr (
.clk_i(clk_i),
.rd_data_o(mie_q),
.rd_data_o_t0(mie_q_t0),
.rst_ni(rst_ni),
.wr_data_i({ dummy_instr_seed_o[3], dummy_instr_seed_o[7], dummy_instr_seed_o[11], dummy_instr_seed_o[30:16] }),
.wr_data_i_t0({ dummy_instr_seed_o_t0[3], dummy_instr_seed_o_t0[7], dummy_instr_seed_o_t0[11], dummy_instr_seed_o_t0[30:16] }),
.wr_en_i(mie_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14371.4-14377.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_mscratch_csr (
.clk_i(clk_i),
.rd_data_o(mscratch_q),
.rd_data_o_t0(mscratch_q_t0),
.rst_ni(rst_ni),
.wr_data_i(dummy_instr_seed_o),
.wr_data_i_t0(dummy_instr_seed_o_t0),
.wr_en_i(mscratch_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14484.4-14490.3" */
\$paramod$34601000fe8707ce2501f5ed778e152043201712\ibex_csr  u_mstack_cause_csr (
.clk_i(clk_i),
.rd_data_o(mstack_cause_q),
.rd_data_o_t0(mstack_cause_q_t0),
.rst_ni(rst_ni),
.wr_data_i(mcause_q),
.wr_data_i_t0(mcause_q_t0),
.wr_en_i(mstack_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14462.4-14468.3" */
\$paramod$410b37fbfbfa994790f1902c150d2be939cadb3b\ibex_csr  u_mstack_csr (
.clk_i(clk_i),
.rd_data_o(mstack_q),
.rd_data_o_t0(mstack_q_t0),
.rst_ni(rst_ni),
.wr_data_i(mstatus_q[4:2]),
.wr_data_i_t0(mstatus_q_t0[4:2]),
.wr_en_i(mstack_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14473.4-14479.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_mstack_epc_csr (
.clk_i(clk_i),
.rd_data_o(mstack_epc_q),
.rd_data_o_t0(mstack_epc_q_t0),
.rst_ni(rst_ni),
.wr_data_i(csr_mepc_o),
.wr_data_i_t0(csr_mepc_o_t0),
.wr_en_i(mstack_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14333.4-14340.3" */
\$paramod$5714e31d82f2b8816750797f158ebea69a089104\ibex_csr  u_mstatus_csr (
.clk_i(clk_i),
.rd_data_o(mstatus_q),
.rd_data_o_t0(mstatus_q_t0),
.rd_error_o(mstatus_err),
.rd_error_o_t0(mstatus_err_t0),
.rst_ni(rst_ni),
.wr_data_i(mstatus_d),
.wr_data_i_t0(mstatus_d_t0),
.wr_en_i(mstatus_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14393.4-14399.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_mtval_csr (
.clk_i(clk_i),
.rd_data_o(csr_mtval_o),
.rd_data_o_t0(csr_mtval_o_t0),
.rst_ni(rst_ni),
.wr_data_i(mtval_d),
.wr_data_i_t0(mtval_d_t0),
.wr_en_i(mtval_en),
.wr_en_i_t0(1'h0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14404.4-14411.3" */
\$paramod$4f46e25470a27719ee9ca03cee1a0827eff766f7\ibex_csr  u_mtvec_csr (
.clk_i(clk_i),
.rd_data_o(csr_mtvec_o),
.rd_data_o_t0(csr_mtvec_o_t0),
.rd_error_o(mtvec_err),
.rd_error_o_t0(mtvec_err_t0),
.rst_ni(rst_ni),
.wr_data_i(mtvec_d),
.wr_data_i_t0(mtvec_d_t0),
.wr_en_i(mtvec_en),
.wr_en_i_t0(mtvec_en_t0)
);
assign _0000_[5:0] = cpuctrlsts_part_d[5:0];
assign _0001_[5:0] = cpuctrlsts_part_d_t0[5:0];
assign { _0003_[31:9], _0003_[5:2] } = { dcsr_d[31:9], dcsr_d[5:2] };
assign { _0004_[31:9], _0004_[5:2] } = { dcsr_d_t0[31:9], dcsr_d_t0[5:2] };
assign _0010_[0] = mstatus_d[0];
assign _0011_[0] = mstatus_d_t0[0];
assign _0020_[8:6] = dcsr_q[8:6];
assign _0021_[8:6] = dcsr_q_t0[8:6];
assign csr_mstatus_mie_o = mstatus_q[5];
assign csr_mstatus_mie_o_t0 = mstatus_q_t0[5];
assign csr_mstatus_tw_o = mstatus_q[0];
assign csr_mstatus_tw_o_t0 = mstatus_q_t0[0];
assign csr_pmp_addr_o = 136'h0000000000000000000000000000000000;
assign csr_pmp_addr_o_t0 = 136'h0000000000000000000000000000000000;
assign csr_pmp_cfg_o = 24'h000000;
assign csr_pmp_cfg_o_t0 = 24'h000000;
assign csr_pmp_mseccfg_o = 3'h0;
assign csr_pmp_mseccfg_o_t0 = 3'h0;
assign data_ind_timing_o = cpuctrlsts_part_q[1];
assign data_ind_timing_o_t0 = cpuctrlsts_part_q_t0[1];
assign debug_ebreakm_o = dcsr_q[15];
assign debug_ebreakm_o_t0 = dcsr_q_t0[15];
assign debug_ebreaku_o = dcsr_q[12];
assign debug_ebreaku_o_t0 = dcsr_q_t0[12];
assign debug_single_step_o = dcsr_q[2];
assign debug_single_step_o_t0 = dcsr_q_t0[2];
assign double_fault_seen_o_t0 = 1'h0;
assign dummy_instr_en_o = cpuctrlsts_part_q[2];
assign dummy_instr_en_o_t0 = cpuctrlsts_part_q_t0[2];
assign dummy_instr_mask_o = cpuctrlsts_part_q[5:3];
assign dummy_instr_mask_o_t0 = cpuctrlsts_part_q_t0[5:3];
assign dummy_instr_seed_en_o_t0 = 1'h0;
assign irq_pending_o_t0 = 1'h0;
assign { mcountinhibit[31:3], mcountinhibit[1] } = 30'h00000000;
assign { mcountinhibit_t0[31:3], mcountinhibit_t0[1] } = 30'h00000000;
assign trigger_match_o = 1'h0;
assign trigger_match_o_t0 = 1'h0;
endmodule

module \$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter (clk_i, rst_ni, counter_inc_i, counterh_we_i, counter_we_i, counter_val_i, counter_val_o, counter_val_upd_o, counter_inc_i_t0, counter_val_i_t0, counter_val_o_t0, counter_val_upd_o_t0, counter_we_i_t0, counterh_we_i_t0);
/* src = "generated/sv2v_out.v:13678.2-13692.5" */
wire [63:0] _00_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13678.2-13692.5" */
wire [63:0] _01_;
wire [63:0] _02_;
wire _03_;
wire _04_;
wire [63:0] _05_;
wire [31:0] _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire [63:0] _12_;
wire [31:0] _13_;
wire [31:0] _14_;
wire [31:0] _15_;
wire [31:0] _16_;
wire [63:0] _17_;
wire [63:0] _18_;
wire [63:0] _19_;
wire [31:0] _20_;
wire [31:0] _21_;
wire [63:0] _22_;
wire [63:0] _23_;
wire [63:0] _24_;
/* src = "generated/sv2v_out.v:13664.13-13664.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:13676.27-13676.36" */
wire [63:0] counter_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13676.27-13676.36" */
wire [63:0] counter_d_t0;
/* src = "generated/sv2v_out.v:13666.13-13666.26" */
input counter_inc_i;
wire counter_inc_i;
/* cellift = 32'd1 */
input counter_inc_i_t0;
wire counter_inc_i_t0;
/* src = "generated/sv2v_out.v:13674.13-13674.25" */
wire [63:0] counter_load;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13674.13-13674.25" */
wire [63:0] counter_load_t0;
/* src = "generated/sv2v_out.v:13669.20-13669.33" */
input [31:0] counter_val_i;
wire [31:0] counter_val_i;
/* cellift = 32'd1 */
input [31:0] counter_val_i_t0;
wire [31:0] counter_val_i_t0;
/* src = "generated/sv2v_out.v:13670.21-13670.34" */
output [63:0] counter_val_o;
reg [63:0] counter_val_o;
/* cellift = 32'd1 */
output [63:0] counter_val_o_t0;
reg [63:0] counter_val_o_t0;
/* src = "generated/sv2v_out.v:13671.21-13671.38" */
output [63:0] counter_val_upd_o;
wire [63:0] counter_val_upd_o;
/* cellift = 32'd1 */
output [63:0] counter_val_upd_o_t0;
wire [63:0] counter_val_upd_o_t0;
/* src = "generated/sv2v_out.v:13668.13-13668.25" */
input counter_we_i;
wire counter_we_i;
/* cellift = 32'd1 */
input counter_we_i_t0;
wire counter_we_i_t0;
/* src = "generated/sv2v_out.v:13667.13-13667.26" */
input counterh_we_i;
wire counterh_we_i;
/* cellift = 32'd1 */
input counterh_we_i_t0;
wire counterh_we_i_t0;
/* src = "generated/sv2v_out.v:13665.13-13665.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:13675.6-13675.8" */
wire we;
assign counter_val_upd_o = counter_val_o + /* src = "generated/sv2v_out.v:13677.23-13677.86" */ 64'h0000000000000001;
assign _02_ = ~ counter_val_o_t0;
assign _12_ = counter_val_o & _02_;
assign _23_ = _12_ + 64'h0000000000000001;
assign _19_ = counter_val_o | counter_val_o_t0;
assign _24_ = _19_ + 64'h0000000000000001;
assign _22_ = _23_ ^ _24_;
assign counter_val_upd_o_t0 = _22_ | counter_val_o_t0;
assign _03_ = ~ _10_;
assign _04_ = ~ _11_;
assign _13_ = { _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_ } & counter_d_t0[63:32];
assign _15_ = { _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_ } & counter_d_t0[31:0];
assign _14_ = { _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_ } & counter_val_o_t0[63:32];
assign _16_ = { _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_ } & counter_val_o_t0[31:0];
assign _20_ = _13_ | _14_;
assign _21_ = _15_ | _16_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter  */
/* PC_TAINT_INFO STATE_NAME counter_val_o_t0[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o_t0[63:32] <= 32'd0;
else counter_val_o_t0[63:32] <= _20_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter  */
/* PC_TAINT_INFO STATE_NAME counter_val_o_t0[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o_t0[31:0] <= 32'd0;
else counter_val_o_t0[31:0] <= _21_;
/* src = "generated/sv2v_out.v:13694.2-13698.27" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter  */
/* PC_TAINT_INFO STATE_NAME counter_val_o[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o[63:32] <= 32'd0;
else if (_10_) counter_val_o[63:32] <= counter_d[63:32];
/* src = "generated/sv2v_out.v:13694.2-13698.27" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter  */
/* PC_TAINT_INFO STATE_NAME counter_val_o[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o[31:0] <= 32'd0;
else if (_11_) counter_val_o[31:0] <= counter_d[31:0];
assign _05_ = ~ { we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we };
assign _06_ = ~ { counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i };
assign _17_ = _05_ & _01_;
assign counter_load_t0[31:0] = _06_ & counter_val_i_t0;
assign _01_ = { counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i } & counter_val_upd_o_t0;
assign _18_ = { we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we } & counter_load_t0;
assign counter_load_t0[63:32] = { counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i } & counter_val_i_t0;
assign counter_d_t0 = _17_ | _18_;
assign _07_ = | { we, counter_inc_i };
assign _08_ = { we, counterh_we_i } != 2'h2;
assign _09_ = { we, counterh_we_i } != 2'h3;
assign _10_ = & { _08_, _07_ };
assign _11_ = & { _07_, _09_ };
assign we = counter_we_i | /* src = "generated/sv2v_out.v:13679.8-13679.36" */ counterh_we_i;
assign _00_ = counter_inc_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13688.12-13688.25|generated/sv2v_out.v:13688.8-13691.44" */ counter_val_upd_o : 64'hxxxxxxxxxxxxxxxx;
assign counter_d = we ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13686.7-13686.9|generated/sv2v_out.v:13686.3-13691.44" */ counter_load : _00_;
assign counter_load[63:32] = counterh_we_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13682.7-13682.20|generated/sv2v_out.v:13682.3-13685.6" */ counter_val_i : 32'hxxxxxxxx;
assign counter_load[31:0] = counterh_we_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13682.7-13682.20|generated/sv2v_out.v:13682.3-13685.6" */ 32'hxxxxxxxx : counter_val_i;
endmodule

module \$paramod$e55993a14b1fbc43320d549f521b710ed37596c6\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _0_;
wire [17:0] _1_;
wire [17:0] _2_;
wire [17:0] _3_;
/* src = "generated/sv2v_out.v:14936.13-14936.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14940.28-14940.37" */
output [17:0] rd_data_o;
reg [17:0] rd_data_o;
/* cellift = 32'd1 */
output [17:0] rd_data_o_t0;
reg [17:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14941.14-14941.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14937.13-14937.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14938.27-14938.36" */
input [17:0] wr_data_i;
wire [17:0] wr_data_i;
/* cellift = 32'd1 */
input [17:0] wr_data_i_t0;
wire [17:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14939.13-14939.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _0_ = ~ wr_en_i;
assign _1_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _2_ = { _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_, _0_ } & rd_data_o_t0;
assign _3_ = _1_ | _2_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$e55993a14b1fbc43320d549f521b710ed37596c6\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 18'h00000;
else rd_data_o_t0 <= _3_;
/* src = "generated/sv2v_out.v:14943.2-14947.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$e55993a14b1fbc43320d549f521b710ed37596c6\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 18'h00000;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage (clk_i, rst_ni, boot_addr_i, req_i, instr_req_o, instr_addr_o, instr_gnt_i, instr_rvalid_i, instr_rdata_i, instr_bus_err_i, instr_intg_err_o, ic_tag_req_o, ic_tag_write_o, ic_tag_addr_o, ic_tag_wdata_o, ic_tag_rdata_i, ic_data_req_o, ic_data_write_o, ic_data_addr_o, ic_data_wdata_o, ic_data_rdata_i
, ic_scr_key_valid_i, ic_scr_key_req_o, instr_valid_id_o, instr_new_id_o, instr_rdata_id_o, instr_rdata_alu_id_o, instr_rdata_c_id_o, instr_is_compressed_id_o, instr_bp_taken_o, instr_fetch_err_o, instr_fetch_err_plus2_o, illegal_c_insn_id_o, dummy_instr_id_o, pc_if_o, pc_id_o, pmp_err_if_i, pmp_err_if_plus2_i, instr_valid_clear_i, pc_set_i, pc_mux_i, nt_branch_mispredict_i
, nt_branch_addr_i, exc_pc_mux_i, exc_cause, dummy_instr_en_i, dummy_instr_mask_i, dummy_instr_seed_en_i, dummy_instr_seed_i, icache_enable_i, icache_inval_i, icache_ecc_error_o, branch_target_ex_i, csr_mepc_i, csr_depc_i, csr_mtvec_i, csr_mtvec_init_o, id_in_ready_i, pc_mismatch_alert_o, if_busy_o, pmp_err_if_plus2_i_t0, pmp_err_if_i_t0, pc_set_i_t0
, pc_mux_i_t0, pc_mismatch_alert_o_t0, pc_if_o_t0, pc_id_o_t0, nt_branch_mispredict_i_t0, nt_branch_addr_i_t0, instr_valid_id_o_t0, instr_valid_clear_i_t0, instr_rdata_id_o_t0, instr_rdata_c_id_o_t0, instr_rdata_alu_id_o_t0, instr_new_id_o_t0, instr_is_compressed_id_o_t0, instr_intg_err_o_t0, instr_fetch_err_plus2_o_t0, instr_fetch_err_o_t0, instr_bus_err_i_t0, instr_bp_taken_o_t0, illegal_c_insn_id_o_t0, if_busy_o_t0, icache_inval_i_t0
, icache_enable_i_t0, icache_ecc_error_o_t0, ic_tag_write_o_t0, ic_tag_wdata_o_t0, ic_tag_req_o_t0, ic_tag_rdata_i_t0, ic_tag_addr_o_t0, ic_scr_key_valid_i_t0, ic_scr_key_req_o_t0, ic_data_write_o_t0, ic_data_wdata_o_t0, ic_data_req_o_t0, ic_data_rdata_i_t0, ic_data_addr_o_t0, exc_pc_mux_i_t0, exc_cause_t0, dummy_instr_id_o_t0, csr_mtvec_init_o_t0, csr_mtvec_i_t0, csr_mepc_i_t0, csr_depc_i_t0
, branch_target_ex_i_t0, boot_addr_i_t0, id_in_ready_i_t0, dummy_instr_seed_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_mask_i_t0, dummy_instr_en_i_t0, req_i_t0, instr_rvalid_i_t0, instr_req_o_t0, instr_rdata_i_t0, instr_gnt_i_t0, instr_addr_o_t0);
/* src = "generated/sv2v_out.v:18161.45-18161.84" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18161.45-18161.84" */
wire _001_;
/* src = "generated/sv2v_out.v:18161.44-18161.106" */
wire _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18161.44-18161.106" */
wire _003_;
/* src = "generated/sv2v_out.v:18167.12-18167.36" */
wire _004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18167.12-18167.36" */
wire _005_;
/* src = "generated/sv2v_out.v:18222.29-18222.73" */
wire _006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18222.29-18222.73" */
wire _007_;
/* src = "generated/sv2v_out.v:18222.78-18222.117" */
wire _008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18222.78-18222.117" */
wire _009_;
/* src = "generated/sv2v_out.v:18278.32-18278.81" */
wire _010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18278.32-18278.81" */
wire _011_;
/* src = "generated/sv2v_out.v:18278.31-18278.98" */
wire _012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18278.31-18278.98" */
wire _013_;
/* src = "generated/sv2v_out.v:18316.29-18316.61" */
wire _014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18316.29-18316.61" */
wire _015_;
/* src = "generated/sv2v_out.v:18316.28-18316.79" */
wire _016_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18316.28-18316.79" */
wire _017_;
/* src = "generated/sv2v_out.v:18317.34-18317.69" */
wire _018_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18317.34-18317.69" */
wire _019_;
/* src = "generated/sv2v_out.v:18317.33-18317.91" */
wire _020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18317.33-18317.91" */
wire _021_;
/* src = "generated/sv2v_out.v:18353.35-18353.81" */
wire _022_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18353.35-18353.81" */
wire _023_;
/* src = "generated/sv2v_out.v:18354.43-18354.87" */
wire _024_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18354.43-18354.87" */
wire _025_;
/* src = "generated/sv2v_out.v:18359.26-18359.60" */
wire _026_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18359.26-18359.60" */
wire _027_;
wire [31:0] _028_;
wire _029_;
wire _030_;
wire [31:0] _031_;
wire [31:0] _032_;
wire [31:0] _033_;
wire [31:0] _034_;
wire [31:0] _035_;
wire [31:0] _036_;
wire [31:0] _037_;
wire [4:0] _038_;
wire [31:0] _039_;
wire [31:0] _040_;
wire _041_;
wire [31:0] _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire [31:0] _061_;
wire [31:0] _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire [31:0] _129_;
wire [31:0] _130_;
wire [31:0] _131_;
wire [31:0] _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire [31:0] _137_;
wire [31:0] _138_;
wire [15:0] _139_;
wire [15:0] _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire [31:0] _149_;
wire [31:0] _150_;
wire _151_;
wire _152_;
wire [31:0] _153_;
wire [31:0] _154_;
wire [31:0] _155_;
wire [31:0] _156_;
wire [31:0] _157_;
wire [31:0] _158_;
wire [31:0] _159_;
wire [31:0] _160_;
wire [31:0] _161_;
wire [31:0] _162_;
wire [31:0] _163_;
wire [31:0] _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire [31:0] _190_;
wire [31:0] _191_;
wire [31:0] _192_;
wire [31:0] _193_;
wire [31:0] _194_;
wire [31:0] _195_;
wire [31:0] _196_;
wire [31:0] _197_;
wire _198_;
wire _199_;
wire _200_;
wire [31:0] _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire [31:0] _224_;
wire [31:0] _225_;
wire _226_;
wire _227_;
wire [31:0] _228_;
wire [15:0] _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire [31:0] _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire [31:0] _245_;
wire [31:0] _246_;
wire [31:0] _247_;
wire [31:0] _248_;
/* cellift = 32'd1 */
wire [31:0] _249_;
wire [31:0] _250_;
/* cellift = 32'd1 */
wire [31:0] _251_;
wire [31:0] _252_;
/* cellift = 32'd1 */
wire [31:0] _253_;
wire [31:0] _254_;
/* cellift = 32'd1 */
wire [31:0] _255_;
wire [31:0] _256_;
wire [31:0] _257_;
/* cellift = 32'd1 */
wire [31:0] _258_;
/* src = "generated/sv2v_out.v:18046.29-18046.45" */
wire _259_;
/* src = "generated/sv2v_out.v:18034.28-18034.82" */
wire _260_;
/* src = "generated/sv2v_out.v:18034.73-18034.82" */
wire _261_;
/* src = "generated/sv2v_out.v:18289.53-18289.88" */
wire _262_;
/* src = "generated/sv2v_out.v:18161.64-18161.84" */
wire _263_;
/* src = "generated/sv2v_out.v:18167.26-18167.36" */
wire _264_;
/* src = "generated/sv2v_out.v:18222.97-18222.117" */
wire _265_;
/* src = "generated/sv2v_out.v:18278.85-18278.98" */
wire _266_;
/* src = "generated/sv2v_out.v:18316.65-18316.79" */
wire _267_;
/* src = "generated/sv2v_out.v:18163.31-18163.113" */
wire _268_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18163.31-18163.113" */
wire _269_;
/* src = "generated/sv2v_out.v:18278.33-18278.66" */
wire _270_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18278.33-18278.66" */
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire _276_;
wire _277_;
wire _278_;
wire _279_;
/* src = "generated/sv2v_out.v:17917.20-17917.31" */
input [31:0] boot_addr_i;
wire [31:0] boot_addr_i;
/* cellift = 32'd1 */
input [31:0] boot_addr_i_t0;
wire [31:0] boot_addr_i_t0;
/* src = "generated/sv2v_out.v:17982.7-17982.17" */
wire branch_req;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17982.7-17982.17" */
wire branch_req_t0;
/* src = "generated/sv2v_out.v:17967.20-17967.38" */
input [31:0] branch_target_ex_i;
wire [31:0] branch_target_ex_i;
/* cellift = 32'd1 */
input [31:0] branch_target_ex_i_t0;
wire [31:0] branch_target_ex_i_t0;
/* src = "generated/sv2v_out.v:17915.13-17915.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:17969.20-17969.30" */
input [31:0] csr_depc_i;
wire [31:0] csr_depc_i;
/* cellift = 32'd1 */
input [31:0] csr_depc_i_t0;
wire [31:0] csr_depc_i_t0;
/* src = "generated/sv2v_out.v:17968.20-17968.30" */
input [31:0] csr_mepc_i;
wire [31:0] csr_mepc_i;
/* cellift = 32'd1 */
input [31:0] csr_mepc_i_t0;
wire [31:0] csr_mepc_i_t0;
/* src = "generated/sv2v_out.v:17970.20-17970.31" */
input [31:0] csr_mtvec_i;
wire [31:0] csr_mtvec_i;
/* cellift = 32'd1 */
input [31:0] csr_mtvec_i_t0;
wire [31:0] csr_mtvec_i_t0;
/* src = "generated/sv2v_out.v:17971.14-17971.30" */
output csr_mtvec_init_o;
wire csr_mtvec_init_o;
/* cellift = 32'd1 */
output csr_mtvec_init_o_t0;
wire csr_mtvec_init_o_t0;
/* src = "generated/sv2v_out.v:17960.13-17960.29" */
input dummy_instr_en_i;
wire dummy_instr_en_i;
/* cellift = 32'd1 */
input dummy_instr_en_i_t0;
wire dummy_instr_en_i_t0;
/* src = "generated/sv2v_out.v:17948.13-17948.29" */
output dummy_instr_id_o;
reg dummy_instr_id_o;
/* cellift = 32'd1 */
output dummy_instr_id_o_t0;
reg dummy_instr_id_o_t0;
/* src = "generated/sv2v_out.v:17961.19-17961.37" */
input [2:0] dummy_instr_mask_i;
wire [2:0] dummy_instr_mask_i;
/* cellift = 32'd1 */
input [2:0] dummy_instr_mask_i_t0;
wire [2:0] dummy_instr_mask_i_t0;
/* src = "generated/sv2v_out.v:17962.13-17962.34" */
input dummy_instr_seed_en_i;
wire dummy_instr_seed_en_i;
/* cellift = 32'd1 */
input dummy_instr_seed_en_i_t0;
wire dummy_instr_seed_en_i_t0;
/* src = "generated/sv2v_out.v:17963.20-17963.38" */
input [31:0] dummy_instr_seed_i;
wire [31:0] dummy_instr_seed_i;
/* cellift = 32'd1 */
input [31:0] dummy_instr_seed_i_t0;
wire [31:0] dummy_instr_seed_i_t0;
/* src = "generated/sv2v_out.v:17959.19-17959.28" */
input [6:0] exc_cause;
wire [6:0] exc_cause;
/* cellift = 32'd1 */
input [6:0] exc_cause_t0;
wire [6:0] exc_cause_t0;
/* src = "generated/sv2v_out.v:18004.13-18004.19" */
wire [31:0] exc_pc;
/* src = "generated/sv2v_out.v:17958.19-17958.31" */
input [1:0] exc_pc_mux_i;
wire [1:0] exc_pc_mux_i;
/* cellift = 32'd1 */
input [1:0] exc_pc_mux_i_t0;
wire [1:0] exc_pc_mux_i_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18004.13-18004.19" */
wire [31:0] exc_pc_t0;
/* src = "generated/sv2v_out.v:17991.14-17991.24" */
wire [31:0] fetch_addr;
/* src = "generated/sv2v_out.v:17983.13-17983.25" */
/* unused_bits = "0" */
wire [31:0] fetch_addr_n;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17983.13-17983.25" */
/* unused_bits = "0" */
wire [31:0] fetch_addr_n_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17991.14-17991.24" */
wire [31:0] fetch_addr_t0;
/* src = "generated/sv2v_out.v:17992.7-17992.16" */
wire fetch_err;
/* src = "generated/sv2v_out.v:17993.7-17993.22" */
wire fetch_err_plus2;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17993.7-17993.22" */
wire fetch_err_plus2_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17992.7-17992.16" */
wire fetch_err_t0;
/* src = "generated/sv2v_out.v:17990.14-17990.25" */
wire [31:0] fetch_rdata;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17990.14-17990.25" */
wire [31:0] fetch_rdata_t0;
/* src = "generated/sv2v_out.v:17989.7-17989.18" */
wire fetch_ready;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17989.7-17989.18" */
wire fetch_ready_t0;
/* src = "generated/sv2v_out.v:17988.7-17988.18" */
wire fetch_valid;
/* src = "generated/sv2v_out.v:17987.7-17987.22" */
wire fetch_valid_raw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17987.7-17987.22" */
wire fetch_valid_raw_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17988.7-17988.18" */
wire fetch_valid_t0;
/* src = "generated/sv2v_out.v:18302.9-18302.25" */
wire \g_branch_predictor.instr_bp_taken_d ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18302.9-18302.25" */
wire \g_branch_predictor.instr_bp_taken_d_t0 ;
/* src = "generated/sv2v_out.v:18296.15-18296.32" */
reg [31:0] \g_branch_predictor.instr_skid_addr_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18296.15-18296.32" */
reg [31:0] \g_branch_predictor.instr_skid_addr_q_t0 ;
/* src = "generated/sv2v_out.v:18297.8-18297.29" */
reg \g_branch_predictor.instr_skid_bp_taken_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18297.8-18297.29" */
reg \g_branch_predictor.instr_skid_bp_taken_q_t0 ;
/* src = "generated/sv2v_out.v:18295.15-18295.32" */
reg [31:0] \g_branch_predictor.instr_skid_data_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18295.15-18295.32" */
reg [31:0] \g_branch_predictor.instr_skid_data_q_t0 ;
/* src = "generated/sv2v_out.v:18300.9-18300.22" */
wire \g_branch_predictor.instr_skid_en ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18300.9-18300.22" */
wire \g_branch_predictor.instr_skid_en_t0 ;
/* src = "generated/sv2v_out.v:18299.9-18299.27" */
wire \g_branch_predictor.instr_skid_valid_d ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18299.9-18299.27" */
wire \g_branch_predictor.instr_skid_valid_d_t0 ;
/* src = "generated/sv2v_out.v:18298.8-18298.26" */
reg \g_branch_predictor.instr_skid_valid_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18298.8-18298.26" */
reg \g_branch_predictor.instr_skid_valid_q_t0 ;
/* src = "generated/sv2v_out.v:18303.9-18303.33" */
wire \g_branch_predictor.predict_branch_taken_raw ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18303.9-18303.33" */
wire \g_branch_predictor.predict_branch_taken_raw_t0 ;
/* src = "generated/sv2v_out.v:18049.15-18049.22" */
wire [1:0] \g_mem_ecc.ecc_err ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18049.15-18049.22" */
/* unused_bits = "0 1" */
wire [1:0] \g_mem_ecc.ecc_err_t0 ;
/* src = "generated/sv2v_out.v:18050.30-18050.45" */
wire [38:0] \g_mem_ecc.instr_rdata_buf ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18050.30-18050.45" */
wire [38:0] \g_mem_ecc.instr_rdata_buf_t0 ;
/* src = "generated/sv2v_out.v:18274.16-18274.36" */
wire [31:0] \g_secure_pc.prev_instr_addr_incr ;
/* src = "generated/sv2v_out.v:18275.16-18275.40" */
wire [31:0] \g_secure_pc.prev_instr_addr_incr_buf ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18275.16-18275.40" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] \g_secure_pc.prev_instr_addr_incr_buf_t0 ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18274.16-18274.36" */
wire [31:0] \g_secure_pc.prev_instr_addr_incr_t0 ;
/* src = "generated/sv2v_out.v:18277.9-18277.25" */
wire \g_secure_pc.prev_instr_seq_d ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18277.9-18277.25" */
wire \g_secure_pc.prev_instr_seq_d_t0 ;
/* src = "generated/sv2v_out.v:18276.8-18276.24" */
reg \g_secure_pc.prev_instr_seq_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18276.8-18276.24" */
reg \g_secure_pc.prev_instr_seq_q_t0 ;
/* src = "generated/sv2v_out.v:18176.16-18176.32" */
wire [31:0] \gen_dummy_instr.dummy_instr_data ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18176.16-18176.32" */
wire [31:0] \gen_dummy_instr.dummy_instr_data_t0 ;
/* src = "generated/sv2v_out.v:18175.9-18175.27" */
wire \gen_dummy_instr.insert_dummy_instr ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18175.9-18175.27" */
wire \gen_dummy_instr.insert_dummy_instr_t0 ;
/* src = "generated/sv2v_out.v:17933.42-17933.56" */
output [7:0] ic_data_addr_o;
wire [7:0] ic_data_addr_o;
/* cellift = 32'd1 */
output [7:0] ic_data_addr_o_t0;
wire [7:0] ic_data_addr_o_t0;
/* src = "generated/sv2v_out.v:17935.58-17935.73" */
input [127:0] ic_data_rdata_i;
wire [127:0] ic_data_rdata_i;
/* cellift = 32'd1 */
input [127:0] ic_data_rdata_i_t0;
wire [127:0] ic_data_rdata_i_t0;
/* src = "generated/sv2v_out.v:17931.20-17931.33" */
output [1:0] ic_data_req_o;
wire [1:0] ic_data_req_o;
/* cellift = 32'd1 */
output [1:0] ic_data_req_o_t0;
wire [1:0] ic_data_req_o_t0;
/* src = "generated/sv2v_out.v:17934.34-17934.49" */
output [63:0] ic_data_wdata_o;
wire [63:0] ic_data_wdata_o;
/* cellift = 32'd1 */
output [63:0] ic_data_wdata_o_t0;
wire [63:0] ic_data_wdata_o_t0;
/* src = "generated/sv2v_out.v:17932.14-17932.29" */
output ic_data_write_o;
wire ic_data_write_o;
/* cellift = 32'd1 */
output ic_data_write_o_t0;
wire ic_data_write_o_t0;
/* src = "generated/sv2v_out.v:17937.14-17937.30" */
output ic_scr_key_req_o;
wire ic_scr_key_req_o;
/* cellift = 32'd1 */
output ic_scr_key_req_o_t0;
wire ic_scr_key_req_o_t0;
/* src = "generated/sv2v_out.v:17936.13-17936.31" */
input ic_scr_key_valid_i;
wire ic_scr_key_valid_i;
/* cellift = 32'd1 */
input ic_scr_key_valid_i_t0;
wire ic_scr_key_valid_i_t0;
/* src = "generated/sv2v_out.v:17928.42-17928.55" */
output [7:0] ic_tag_addr_o;
wire [7:0] ic_tag_addr_o;
/* cellift = 32'd1 */
output [7:0] ic_tag_addr_o_t0;
wire [7:0] ic_tag_addr_o_t0;
/* src = "generated/sv2v_out.v:17930.57-17930.71" */
input [43:0] ic_tag_rdata_i;
wire [43:0] ic_tag_rdata_i;
/* cellift = 32'd1 */
input [43:0] ic_tag_rdata_i_t0;
wire [43:0] ic_tag_rdata_i_t0;
/* src = "generated/sv2v_out.v:17926.20-17926.32" */
output [1:0] ic_tag_req_o;
wire [1:0] ic_tag_req_o;
/* cellift = 32'd1 */
output [1:0] ic_tag_req_o_t0;
wire [1:0] ic_tag_req_o_t0;
/* src = "generated/sv2v_out.v:17929.33-17929.47" */
output [21:0] ic_tag_wdata_o;
wire [21:0] ic_tag_wdata_o;
/* cellift = 32'd1 */
output [21:0] ic_tag_wdata_o_t0;
wire [21:0] ic_tag_wdata_o_t0;
/* src = "generated/sv2v_out.v:17927.14-17927.28" */
output ic_tag_write_o;
wire ic_tag_write_o;
/* cellift = 32'd1 */
output ic_tag_write_o_t0;
wire ic_tag_write_o_t0;
/* src = "generated/sv2v_out.v:17966.14-17966.32" */
output icache_ecc_error_o;
wire icache_ecc_error_o;
/* cellift = 32'd1 */
output icache_ecc_error_o_t0;
wire icache_ecc_error_o_t0;
/* src = "generated/sv2v_out.v:17964.13-17964.28" */
input icache_enable_i;
wire icache_enable_i;
/* cellift = 32'd1 */
input icache_enable_i_t0;
wire icache_enable_i_t0;
/* src = "generated/sv2v_out.v:17965.13-17965.27" */
input icache_inval_i;
wire icache_inval_i;
/* cellift = 32'd1 */
input icache_inval_i_t0;
wire icache_inval_i_t0;
/* src = "generated/sv2v_out.v:17972.13-17972.26" */
input id_in_ready_i;
wire id_in_ready_i;
/* cellift = 32'd1 */
input id_in_ready_i_t0;
wire id_in_ready_i_t0;
/* src = "generated/sv2v_out.v:17974.14-17974.23" */
output if_busy_o;
wire if_busy_o;
/* cellift = 32'd1 */
output if_busy_o_t0;
wire if_busy_o_t0;
/* src = "generated/sv2v_out.v:18005.7-18005.24" */
wire if_id_pipe_reg_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18005.7-18005.24" */
wire if_id_pipe_reg_we_t0;
/* src = "generated/sv2v_out.v:18000.7-18000.23" */
wire if_instr_bus_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18000.7-18000.23" */
wire if_instr_bus_err_t0;
/* src = "generated/sv2v_out.v:18002.7-18002.19" */
wire if_instr_err;
/* src = "generated/sv2v_out.v:18003.7-18003.25" */
wire if_instr_err_plus2;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18003.7-18003.25" */
wire if_instr_err_plus2_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18002.7-18002.19" */
wire if_instr_err_t0;
/* src = "generated/sv2v_out.v:18001.7-18001.23" */
wire if_instr_pmp_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18001.7-18001.23" */
wire if_instr_pmp_err_t0;
/* src = "generated/sv2v_out.v:17998.14-17998.28" */
wire [31:0] if_instr_rdata;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17998.14-17998.28" */
wire [31:0] if_instr_rdata_t0;
/* src = "generated/sv2v_out.v:17997.7-17997.21" */
wire if_instr_valid;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17997.7-17997.21" */
wire if_instr_valid_t0;
/* src = "generated/sv2v_out.v:17995.7-17995.21" */
wire illegal_c_insn;
/* src = "generated/sv2v_out.v:17947.13-17947.32" */
output illegal_c_insn_id_o;
reg illegal_c_insn_id_o;
/* cellift = 32'd1 */
output illegal_c_insn_id_o_t0;
reg illegal_c_insn_id_o_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17995.7-17995.21" */
wire illegal_c_insn_t0;
/* src = "generated/sv2v_out.v:18009.7-18009.26" */
wire illegal_c_instr_out;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18009.7-18009.26" */
wire illegal_c_instr_out_t0;
/* src = "generated/sv2v_out.v:17920.21-17920.33" */
output [31:0] instr_addr_o;
wire [31:0] instr_addr_o;
/* cellift = 32'd1 */
output [31:0] instr_addr_o_t0;
wire [31:0] instr_addr_o_t0;
/* src = "generated/sv2v_out.v:17944.14-17944.30" */
output instr_bp_taken_o;
reg instr_bp_taken_o;
/* cellift = 32'd1 */
output instr_bp_taken_o_t0;
reg instr_bp_taken_o_t0;
/* src = "generated/sv2v_out.v:17924.13-17924.28" */
input instr_bus_err_i;
wire instr_bus_err_i;
/* cellift = 32'd1 */
input instr_bus_err_i_t0;
wire instr_bus_err_i_t0;
/* src = "generated/sv2v_out.v:17994.14-17994.32" */
wire [31:0] instr_decompressed;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17994.14-17994.32" */
wire [31:0] instr_decompressed_t0;
/* src = "generated/sv2v_out.v:17979.7-17979.16" */
wire instr_err;
/* src = "generated/sv2v_out.v:18010.7-18010.20" */
wire instr_err_out;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18010.7-18010.20" */
wire instr_err_out_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17979.7-17979.16" */
wire instr_err_t0;
/* src = "generated/sv2v_out.v:17945.13-17945.30" */
output instr_fetch_err_o;
reg instr_fetch_err_o;
/* cellift = 32'd1 */
output instr_fetch_err_o_t0;
reg instr_fetch_err_o_t0;
/* src = "generated/sv2v_out.v:17946.13-17946.36" */
output instr_fetch_err_plus2_o;
reg instr_fetch_err_plus2_o;
/* cellift = 32'd1 */
output instr_fetch_err_plus2_o_t0;
reg instr_fetch_err_plus2_o_t0;
/* src = "generated/sv2v_out.v:17921.13-17921.24" */
input instr_gnt_i;
wire instr_gnt_i;
/* cellift = 32'd1 */
input instr_gnt_i_t0;
wire instr_gnt_i_t0;
/* src = "generated/sv2v_out.v:17980.7-17980.21" */
wire instr_intg_err;
/* src = "generated/sv2v_out.v:17925.14-17925.30" */
output instr_intg_err_o;
wire instr_intg_err_o;
/* cellift = 32'd1 */
output instr_intg_err_o_t0;
wire instr_intg_err_o_t0;
/* src = "generated/sv2v_out.v:17996.7-17996.26" */
wire instr_is_compressed;
/* src = "generated/sv2v_out.v:17943.13-17943.37" */
output instr_is_compressed_id_o;
reg instr_is_compressed_id_o;
/* cellift = 32'd1 */
output instr_is_compressed_id_o_t0;
reg instr_is_compressed_id_o_t0;
/* src = "generated/sv2v_out.v:18008.7-18008.30" */
wire instr_is_compressed_out;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18008.7-18008.30" */
wire instr_is_compressed_out_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17996.7-17996.26" */
wire instr_is_compressed_t0;
/* src = "generated/sv2v_out.v:17939.14-17939.28" */
output instr_new_id_o;
reg instr_new_id_o;
/* cellift = 32'd1 */
output instr_new_id_o_t0;
reg instr_new_id_o_t0;
/* src = "generated/sv2v_out.v:18007.14-18007.23" */
wire [31:0] instr_out;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18007.14-18007.23" */
wire [31:0] instr_out_t0;
/* src = "generated/sv2v_out.v:17941.20-17941.40" */
output [31:0] instr_rdata_alu_id_o;
reg [31:0] instr_rdata_alu_id_o;
/* cellift = 32'd1 */
output [31:0] instr_rdata_alu_id_o_t0;
reg [31:0] instr_rdata_alu_id_o_t0;
/* src = "generated/sv2v_out.v:17942.20-17942.38" */
output [15:0] instr_rdata_c_id_o;
reg [15:0] instr_rdata_c_id_o;
/* cellift = 32'd1 */
output [15:0] instr_rdata_c_id_o_t0;
reg [15:0] instr_rdata_c_id_o_t0;
/* src = "generated/sv2v_out.v:17923.34-17923.47" */
input [38:0] instr_rdata_i;
wire [38:0] instr_rdata_i;
/* cellift = 32'd1 */
input [38:0] instr_rdata_i_t0;
wire [38:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:17940.20-17940.36" */
output [31:0] instr_rdata_id_o;
wire [31:0] instr_rdata_id_o;
/* cellift = 32'd1 */
output [31:0] instr_rdata_id_o_t0;
wire [31:0] instr_rdata_id_o_t0;
/* src = "generated/sv2v_out.v:17919.14-17919.25" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:17922.13-17922.27" */
input instr_rvalid_i;
wire instr_rvalid_i;
/* cellift = 32'd1 */
input instr_rvalid_i_t0;
wire instr_rvalid_i_t0;
/* src = "generated/sv2v_out.v:17953.13-17953.32" */
input instr_valid_clear_i;
wire instr_valid_clear_i;
/* cellift = 32'd1 */
input instr_valid_clear_i_t0;
wire instr_valid_clear_i_t0;
/* src = "generated/sv2v_out.v:17975.7-17975.23" */
wire instr_valid_id_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17975.7-17975.23" */
wire instr_valid_id_d_t0;
/* src = "generated/sv2v_out.v:17938.14-17938.30" */
output instr_valid_id_o;
reg instr_valid_id_o;
/* cellift = 32'd1 */
output instr_valid_id_o_t0;
reg instr_valid_id_o_t0;
/* src = "generated/sv2v_out.v:18013.12-18013.19" */
wire [4:0] irq_vec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18013.12-18013.19" */
wire [4:0] irq_vec_t0;
/* src = "generated/sv2v_out.v:17957.20-17957.36" */
input [31:0] nt_branch_addr_i;
wire [31:0] nt_branch_addr_i;
/* cellift = 32'd1 */
input [31:0] nt_branch_addr_i_t0;
wire [31:0] nt_branch_addr_i_t0;
/* src = "generated/sv2v_out.v:17956.13-17956.35" */
input nt_branch_mispredict_i;
wire nt_branch_mispredict_i;
/* cellift = 32'd1 */
input nt_branch_mispredict_i_t0;
wire nt_branch_mispredict_i_t0;
/* src = "generated/sv2v_out.v:17950.20-17950.27" */
output [31:0] pc_id_o;
reg [31:0] pc_id_o;
/* cellift = 32'd1 */
output [31:0] pc_id_o_t0;
reg [31:0] pc_id_o_t0;
/* src = "generated/sv2v_out.v:17949.21-17949.28" */
output [31:0] pc_if_o;
wire [31:0] pc_if_o;
/* cellift = 32'd1 */
output [31:0] pc_if_o_t0;
wire [31:0] pc_if_o_t0;
/* src = "generated/sv2v_out.v:17973.14-17973.33" */
output pc_mismatch_alert_o;
wire pc_mismatch_alert_o;
/* cellift = 32'd1 */
output pc_mismatch_alert_o_t0;
wire pc_mismatch_alert_o_t0;
/* src = "generated/sv2v_out.v:17955.19-17955.27" */
input [2:0] pc_mux_i;
wire [2:0] pc_mux_i;
/* cellift = 32'd1 */
input [2:0] pc_mux_i_t0;
wire [2:0] pc_mux_i_t0;
/* src = "generated/sv2v_out.v:18014.13-18014.28" */
wire [2:0] pc_mux_internal;
/* src = "generated/sv2v_out.v:17954.13-17954.21" */
input pc_set_i;
wire pc_set_i;
/* cellift = 32'd1 */
input pc_set_i_t0;
wire pc_set_i_t0;
/* src = "generated/sv2v_out.v:17951.13-17951.25" */
input pmp_err_if_i;
wire pmp_err_if_i;
/* cellift = 32'd1 */
input pmp_err_if_i_t0;
wire pmp_err_if_i_t0;
/* src = "generated/sv2v_out.v:17952.13-17952.31" */
input pmp_err_if_plus2_i;
wire pmp_err_if_plus2_i;
/* cellift = 32'd1 */
input pmp_err_if_plus2_i_t0;
wire pmp_err_if_plus2_i_t0;
/* src = "generated/sv2v_out.v:18012.14-18012.31" */
wire [31:0] predict_branch_pc;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18012.14-18012.31" */
wire [31:0] predict_branch_pc_t0;
/* src = "generated/sv2v_out.v:18011.7-18011.27" */
wire predict_branch_taken;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18011.7-18011.27" */
wire predict_branch_taken_t0;
/* src = "generated/sv2v_out.v:17986.14-17986.27" */
wire [31:0] prefetch_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17986.14-17986.27" */
wire [31:0] prefetch_addr_t0;
/* src = "generated/sv2v_out.v:17985.7-17985.22" */
wire prefetch_branch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17985.7-17985.22" */
wire prefetch_branch_t0;
/* src = "generated/sv2v_out.v:17918.13-17918.18" */
input req_i;
wire req_i;
/* cellift = 32'd1 */
input req_i_t0;
wire req_i_t0;
/* src = "generated/sv2v_out.v:17916.13-17916.19" */
input rst_ni;
wire rst_ni;
assign \g_secure_pc.prev_instr_addr_incr  = pc_id_o + /* src = "generated/sv2v_out.v:18284.34-18284.86" */ _062_;
assign csr_mtvec_init_o = _259_ & /* src = "generated/sv2v_out.v:18046.28-18046.57" */ pc_set_i;
assign instr_intg_err_o = instr_intg_err & /* src = "generated/sv2v_out.v:18066.28-18066.59" */ instr_rvalid_i;
assign fetch_valid = fetch_valid_raw & /* src = "generated/sv2v_out.v:18069.23-18069.64" */ _054_;
assign _000_ = pc_if_o[1] & /* src = "generated/sv2v_out.v:18163.33-18163.72" */ _263_;
assign _002_ = _000_ & /* src = "generated/sv2v_out.v:18163.32-18163.94" */ pmp_err_if_plus2_i;
assign if_instr_err_plus2 = _268_ & /* src = "generated/sv2v_out.v:18163.30-18163.130" */ _047_;
assign _004_ = fetch_valid & /* src = "generated/sv2v_out.v:18167.12-18167.36" */ _264_;
assign _006_ = if_id_pipe_reg_we & /* src = "generated/sv2v_out.v:18222.29-18222.73" */ _046_;
assign _008_ = instr_valid_id_o & /* src = "generated/sv2v_out.v:18222.78-18222.117" */ _265_;
assign if_id_pipe_reg_we = if_instr_valid & /* src = "generated/sv2v_out.v:18223.26-18223.56" */ id_in_ready_i;
assign _010_ = _270_ & /* src = "generated/sv2v_out.v:18278.32-18278.81" */ _045_;
assign _012_ = _010_ & /* src = "generated/sv2v_out.v:18278.31-18278.98" */ _266_;
assign \g_secure_pc.prev_instr_seq_d  = _012_ & /* src = "generated/sv2v_out.v:18278.30-18278.120" */ _041_;
assign pc_mismatch_alert_o = \g_secure_pc.prev_instr_seq_q  & /* src = "generated/sv2v_out.v:18289.33-18289.89" */ _262_;
assign \g_branch_predictor.instr_skid_en  = _016_ & /* src = "generated/sv2v_out.v:18316.27-18316.102" */ _043_;
assign _014_ = predict_branch_taken & /* src = "generated/sv2v_out.v:18316.29-18316.61" */ _046_;
assign _016_ = _014_ & /* src = "generated/sv2v_out.v:18316.28-18316.79" */ _267_;
assign _018_ = \g_branch_predictor.instr_skid_valid_q  & /* src = "generated/sv2v_out.v:18317.34-18317.69" */ _267_;
assign _020_ = _018_ & /* src = "generated/sv2v_out.v:18317.33-18317.91" */ _041_;
assign _022_ = \g_branch_predictor.predict_branch_taken_raw  & /* src = "generated/sv2v_out.v:18353.35-18353.81" */ _043_;
assign predict_branch_taken = _022_ & /* src = "generated/sv2v_out.v:18353.34-18353.95" */ _264_;
assign _024_ = \g_branch_predictor.instr_skid_valid_q  & /* src = "generated/sv2v_out.v:18354.43-18354.87" */ _054_;
assign if_instr_bus_err = _043_ & /* src = "generated/sv2v_out.v:18357.30-18357.61" */ fetch_err;
assign _026_ = id_in_ready_i & /* src = "generated/sv2v_out.v:18359.26-18359.60" */ _041_;
assign fetch_ready = _026_ & /* src = "generated/sv2v_out.v:18359.25-18359.83" */ _043_;
assign _028_ = ~ pc_id_o_t0;
assign _061_ = pc_id_o & _028_;
assign _246_ = _061_ + _062_;
assign _201_ = pc_id_o | pc_id_o_t0;
assign _247_ = _201_ + _062_;
assign _245_ = _246_ ^ _247_;
assign \g_secure_pc.prev_instr_addr_incr_t0  = _245_ | pc_id_o_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME \g_branch_predictor.instr_skid_valid_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_branch_predictor.instr_skid_valid_q_t0  <= 1'h0;
else \g_branch_predictor.instr_skid_valid_q_t0  <= \g_branch_predictor.instr_skid_valid_d_t0 ;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME \g_secure_pc.prev_instr_seq_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_secure_pc.prev_instr_seq_q_t0  <= 1'h0;
else \g_secure_pc.prev_instr_seq_q_t0  <= \g_secure_pc.prev_instr_seq_d_t0 ;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_valid_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_valid_id_o_t0 <= 1'h0;
else instr_valid_id_o_t0 <= instr_valid_id_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_new_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_new_id_o_t0 <= 1'h0;
else instr_new_id_o_t0 <= if_id_pipe_reg_we_t0;
assign _029_ = ~ \g_branch_predictor.instr_skid_en ;
assign _030_ = ~ if_id_pipe_reg_we;
assign _129_ = { \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en  } & fetch_rdata_t0;
assign _131_ = { \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en , \g_branch_predictor.instr_skid_en  } & fetch_addr_t0;
assign _133_ = \g_branch_predictor.instr_skid_en  & predict_branch_taken_t0;
assign _135_ = if_id_pipe_reg_we & \g_branch_predictor.instr_bp_taken_d_t0 ;
assign _137_ = { if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we } & instr_out_t0;
assign _139_ = { if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we } & if_instr_rdata_t0[15:0];
assign _141_ = if_id_pipe_reg_we & instr_is_compressed_out_t0;
assign _143_ = if_id_pipe_reg_we & instr_err_out_t0;
assign _145_ = if_id_pipe_reg_we & if_instr_err_plus2_t0;
assign _147_ = if_id_pipe_reg_we & illegal_c_instr_out_t0;
assign _149_ = { if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we } & pc_if_o_t0;
assign _151_ = if_id_pipe_reg_we & \gen_dummy_instr.insert_dummy_instr_t0 ;
assign _130_ = { _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_ } & \g_branch_predictor.instr_skid_data_q_t0 ;
assign _132_ = { _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_ } & \g_branch_predictor.instr_skid_addr_q_t0 ;
assign _134_ = _029_ & \g_branch_predictor.instr_skid_bp_taken_q_t0 ;
assign _136_ = _030_ & instr_bp_taken_o_t0;
assign _138_ = { _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_ } & instr_rdata_alu_id_o_t0;
assign _140_ = { _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_ } & instr_rdata_c_id_o_t0;
assign _142_ = _030_ & instr_is_compressed_id_o_t0;
assign _144_ = _030_ & instr_fetch_err_o_t0;
assign _146_ = _030_ & instr_fetch_err_plus2_o_t0;
assign _148_ = _030_ & illegal_c_insn_id_o_t0;
assign _150_ = { _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_ } & pc_id_o_t0;
assign _152_ = _030_ & dummy_instr_id_o_t0;
assign _224_ = _129_ | _130_;
assign _225_ = _131_ | _132_;
assign _226_ = _133_ | _134_;
assign _227_ = _135_ | _136_;
assign _228_ = _137_ | _138_;
assign _229_ = _139_ | _140_;
assign _230_ = _141_ | _142_;
assign _231_ = _143_ | _144_;
assign _232_ = _145_ | _146_;
assign _233_ = _147_ | _148_;
assign _234_ = _149_ | _150_;
assign _235_ = _151_ | _152_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME \g_branch_predictor.instr_skid_data_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_branch_predictor.instr_skid_data_q_t0  <= 32'd0;
else \g_branch_predictor.instr_skid_data_q_t0  <= _224_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME \g_branch_predictor.instr_skid_addr_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_branch_predictor.instr_skid_addr_q_t0  <= 32'd0;
else \g_branch_predictor.instr_skid_addr_q_t0  <= _225_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME \g_branch_predictor.instr_skid_bp_taken_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_branch_predictor.instr_skid_bp_taken_q_t0  <= 1'h0;
else \g_branch_predictor.instr_skid_bp_taken_q_t0  <= _226_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_bp_taken_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_bp_taken_o_t0 <= 1'h0;
else instr_bp_taken_o_t0 <= _227_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_rdata_alu_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_rdata_alu_id_o_t0 <= 32'd0;
else instr_rdata_alu_id_o_t0 <= _228_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_rdata_c_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_rdata_c_id_o_t0 <= 16'h0000;
else instr_rdata_c_id_o_t0 <= _229_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_is_compressed_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_is_compressed_id_o_t0 <= 1'h0;
else instr_is_compressed_id_o_t0 <= _230_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_fetch_err_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_fetch_err_o_t0 <= 1'h0;
else instr_fetch_err_o_t0 <= _231_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_fetch_err_plus2_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_fetch_err_plus2_o_t0 <= 1'h0;
else instr_fetch_err_plus2_o_t0 <= _232_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME illegal_c_insn_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) illegal_c_insn_id_o_t0 <= 1'h0;
else illegal_c_insn_id_o_t0 <= _233_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME pc_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) pc_id_o_t0 <= 32'd0;
else pc_id_o_t0 <= _234_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME dummy_instr_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_instr_id_o_t0 <= 1'h0;
else dummy_instr_id_o_t0 <= _235_;
assign _063_ = fetch_valid_raw_t0 & _054_;
assign _066_ = pc_if_o_t0[1] & _263_;
assign _069_ = _001_ & pmp_err_if_plus2_i;
assign _072_ = _269_ & _047_;
assign _075_ = fetch_valid_t0 & _264_;
assign _078_ = if_id_pipe_reg_we_t0 & _046_;
assign _081_ = instr_valid_id_o_t0 & _265_;
assign _084_ = if_instr_valid_t0 & id_in_ready_i;
assign _087_ = _271_ & _045_;
assign _090_ = _011_ & _266_;
assign _093_ = _013_ & _041_;
assign pc_mismatch_alert_o_t0 = \g_secure_pc.prev_instr_seq_q_t0  & _262_;
assign _096_ = _017_ & _043_;
assign _099_ = predict_branch_taken_t0 & _046_;
assign _102_ = _015_ & _267_;
assign _105_ = \g_branch_predictor.instr_skid_valid_q_t0  & _267_;
assign _108_ = _019_ & _041_;
assign _111_ = \g_branch_predictor.predict_branch_taken_raw_t0  & _043_;
assign _114_ = _023_ & _264_;
assign _117_ = \g_branch_predictor.instr_skid_valid_q_t0  & _054_;
assign _120_ = \g_branch_predictor.instr_skid_valid_q_t0  & fetch_err;
assign _123_ = id_in_ready_i_t0 & _041_;
assign _126_ = _027_ & _043_;
assign csr_mtvec_init_o_t0 = pc_set_i_t0 & _259_;
assign instr_intg_err_o_t0 = instr_rvalid_i_t0 & instr_intg_err;
assign _064_ = nt_branch_mispredict_i_t0 & fetch_valid_raw;
assign _067_ = instr_is_compressed_t0 & pc_if_o[1];
assign _070_ = pmp_err_if_plus2_i_t0 & _000_;
assign _073_ = pmp_err_if_i_t0 & _268_;
assign _076_ = fetch_err_t0 & fetch_valid;
assign _079_ = pc_set_i_t0 & if_id_pipe_reg_we;
assign _082_ = instr_valid_clear_i_t0 & instr_valid_id_o;
assign _085_ = id_in_ready_i_t0 & if_instr_valid;
assign _088_ = branch_req_t0 & _270_;
assign _091_ = if_instr_err_t0 & _010_;
assign _094_ = \gen_dummy_instr.insert_dummy_instr_t0  & _012_;
assign _097_ = \g_branch_predictor.instr_skid_valid_q_t0  & _016_;
assign _100_ = pc_set_i_t0 & predict_branch_taken;
assign _103_ = id_in_ready_i_t0 & _014_;
assign _106_ = id_in_ready_i_t0 & \g_branch_predictor.instr_skid_valid_q ;
assign _109_ = \gen_dummy_instr.insert_dummy_instr_t0  & _018_;
assign _112_ = \g_branch_predictor.instr_skid_valid_q_t0  & \g_branch_predictor.predict_branch_taken_raw ;
assign _115_ = fetch_err_t0 & _022_;
assign _118_ = nt_branch_mispredict_i_t0 & \g_branch_predictor.instr_skid_valid_q ;
assign _121_ = fetch_err_t0 & _043_;
assign _124_ = \gen_dummy_instr.insert_dummy_instr_t0  & id_in_ready_i;
assign _127_ = \g_branch_predictor.instr_skid_valid_q_t0  & _026_;
assign _065_ = fetch_valid_raw_t0 & nt_branch_mispredict_i_t0;
assign _068_ = pc_if_o_t0[1] & instr_is_compressed_t0;
assign _071_ = _001_ & pmp_err_if_plus2_i_t0;
assign _074_ = _269_ & pmp_err_if_i_t0;
assign _077_ = fetch_valid_t0 & fetch_err_t0;
assign _080_ = if_id_pipe_reg_we_t0 & pc_set_i_t0;
assign _083_ = instr_valid_id_o_t0 & instr_valid_clear_i_t0;
assign _086_ = if_instr_valid_t0 & id_in_ready_i_t0;
assign _089_ = _271_ & branch_req_t0;
assign _092_ = _011_ & if_instr_err_t0;
assign _095_ = _013_ & \gen_dummy_instr.insert_dummy_instr_t0 ;
assign _098_ = _017_ & \g_branch_predictor.instr_skid_valid_q_t0 ;
assign _101_ = predict_branch_taken_t0 & pc_set_i_t0;
assign _104_ = _015_ & id_in_ready_i_t0;
assign _107_ = \g_branch_predictor.instr_skid_valid_q_t0  & id_in_ready_i_t0;
assign _110_ = _019_ & \gen_dummy_instr.insert_dummy_instr_t0 ;
assign _113_ = \g_branch_predictor.predict_branch_taken_raw_t0  & \g_branch_predictor.instr_skid_valid_q_t0 ;
assign _116_ = _023_ & fetch_err_t0;
assign _119_ = \g_branch_predictor.instr_skid_valid_q_t0  & nt_branch_mispredict_i_t0;
assign _122_ = \g_branch_predictor.instr_skid_valid_q_t0  & fetch_err_t0;
assign _125_ = id_in_ready_i_t0 & \gen_dummy_instr.insert_dummy_instr_t0 ;
assign _128_ = _027_ & \g_branch_predictor.instr_skid_valid_q_t0 ;
assign _202_ = _063_ | _064_;
assign _203_ = _066_ | _067_;
assign _204_ = _069_ | _070_;
assign _205_ = _072_ | _073_;
assign _206_ = _075_ | _076_;
assign _207_ = _078_ | _079_;
assign _208_ = _081_ | _082_;
assign _209_ = _084_ | _085_;
assign _210_ = _087_ | _088_;
assign _211_ = _090_ | _091_;
assign _212_ = _093_ | _094_;
assign _213_ = _096_ | _097_;
assign _214_ = _099_ | _100_;
assign _215_ = _102_ | _103_;
assign _216_ = _105_ | _106_;
assign _217_ = _108_ | _109_;
assign _218_ = _111_ | _112_;
assign _219_ = _114_ | _115_;
assign _220_ = _117_ | _118_;
assign _221_ = _120_ | _121_;
assign _222_ = _123_ | _124_;
assign _223_ = _126_ | _127_;
assign fetch_valid_t0 = _202_ | _065_;
assign _001_ = _203_ | _068_;
assign _003_ = _204_ | _071_;
assign if_instr_err_plus2_t0 = _205_ | _074_;
assign _005_ = _206_ | _077_;
assign _007_ = _207_ | _080_;
assign _009_ = _208_ | _083_;
assign if_id_pipe_reg_we_t0 = _209_ | _086_;
assign _011_ = _210_ | _089_;
assign _013_ = _211_ | _092_;
assign \g_secure_pc.prev_instr_seq_d_t0  = _212_ | _095_;
assign \g_branch_predictor.instr_skid_en_t0  = _213_ | _098_;
assign _015_ = _214_ | _101_;
assign _017_ = _215_ | _104_;
assign _019_ = _216_ | _107_;
assign _021_ = _217_ | _110_;
assign _023_ = _218_ | _113_;
assign predict_branch_taken_t0 = _219_ | _116_;
assign _025_ = _220_ | _119_;
assign if_instr_bus_err_t0 = _221_ | _122_;
assign _027_ = _222_ | _125_;
assign fetch_ready_t0 = _223_ | _128_;
/* src = "generated/sv2v_out.v:18324.5-18334.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME \g_branch_predictor.instr_skid_data_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_branch_predictor.instr_skid_data_q  <= 32'd0;
else if (\g_branch_predictor.instr_skid_en ) \g_branch_predictor.instr_skid_data_q  <= fetch_rdata;
/* src = "generated/sv2v_out.v:18324.5-18334.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME \g_branch_predictor.instr_skid_addr_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_branch_predictor.instr_skid_addr_q  <= 32'd0;
else if (\g_branch_predictor.instr_skid_en ) \g_branch_predictor.instr_skid_addr_q  <= fetch_addr;
/* src = "generated/sv2v_out.v:18324.5-18334.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME \g_branch_predictor.instr_skid_bp_taken_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_branch_predictor.instr_skid_bp_taken_q  <= 1'h0;
else if (\g_branch_predictor.instr_skid_en ) \g_branch_predictor.instr_skid_bp_taken_q  <= predict_branch_taken;
/* src = "generated/sv2v_out.v:18305.5-18309.44" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_bp_taken_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_bp_taken_o <= 1'h0;
else if (if_id_pipe_reg_we) instr_bp_taken_o <= \g_branch_predictor.instr_bp_taken_d ;
/* src = "generated/sv2v_out.v:18238.4-18258.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_rdata_alu_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_rdata_alu_id_o <= 32'd0;
else if (if_id_pipe_reg_we) instr_rdata_alu_id_o <= instr_out;
/* src = "generated/sv2v_out.v:18238.4-18258.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_rdata_c_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_rdata_c_id_o <= 16'h0000;
else if (if_id_pipe_reg_we) instr_rdata_c_id_o <= if_instr_rdata[15:0];
/* src = "generated/sv2v_out.v:18238.4-18258.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_is_compressed_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_is_compressed_id_o <= 1'h0;
else if (if_id_pipe_reg_we) instr_is_compressed_id_o <= instr_is_compressed_out;
/* src = "generated/sv2v_out.v:18238.4-18258.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_fetch_err_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_fetch_err_o <= 1'h0;
else if (if_id_pipe_reg_we) instr_fetch_err_o <= instr_err_out;
/* src = "generated/sv2v_out.v:18238.4-18258.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_fetch_err_plus2_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_fetch_err_plus2_o <= 1'h0;
else if (if_id_pipe_reg_we) instr_fetch_err_plus2_o <= if_instr_err_plus2;
/* src = "generated/sv2v_out.v:18238.4-18258.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME illegal_c_insn_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) illegal_c_insn_id_o <= 1'h0;
else if (if_id_pipe_reg_we) illegal_c_insn_id_o <= illegal_c_instr_out;
/* src = "generated/sv2v_out.v:18238.4-18258.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME pc_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) pc_id_o <= 32'd0;
else if (if_id_pipe_reg_we) pc_id_o <= pc_if_o;
/* src = "generated/sv2v_out.v:18197.4-18201.45" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME dummy_instr_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_instr_id_o <= 1'h0;
else if (if_id_pipe_reg_we) dummy_instr_id_o <= \gen_dummy_instr.insert_dummy_instr ;
assign _031_ = ~ { _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_ };
assign _032_ = ~ { _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_ };
assign _033_ = ~ { _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_ };
assign _034_ = ~ { _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_ };
assign _035_ = ~ { _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_ };
assign _036_ = ~ { _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_ };
assign _037_ = ~ { _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_, _200_ };
assign _038_ = ~ { exc_cause[6], exc_cause[6], exc_cause[6], exc_cause[6], exc_cause[6] };
assign _039_ = ~ { branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req };
assign _040_ = ~ { \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr  };
assign _041_ = ~ \gen_dummy_instr.insert_dummy_instr ;
assign _042_ = ~ { \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q  };
assign _043_ = ~ \g_branch_predictor.instr_skid_valid_q ;
assign _153_ = _031_ & csr_mepc_i_t0;
assign _155_ = _032_ & _249_;
assign _157_ = _033_ & { boot_addr_i_t0[31:8], 8'h00 };
assign _159_ = _034_ & _253_;
assign _161_ = _035_ & _255_;
assign _163_ = _036_ & { csr_mtvec_i_t0[31:8], 8'h00 };
assign exc_pc_t0 = _037_ & _258_;
assign irq_vec_t0 = _038_ & exc_cause_t0[4:0];
assign _190_ = _039_ & nt_branch_addr_i_t0;
assign _192_ = _040_ & instr_decompressed_t0;
assign instr_is_compressed_out_t0 = _041_ & instr_is_compressed_t0;
assign illegal_c_instr_out_t0 = _041_ & illegal_c_insn_t0;
assign instr_err_out_t0 = _041_ & if_instr_err_t0;
assign _194_ = _042_ & fetch_rdata_t0;
assign _196_ = _042_ & fetch_addr_t0;
assign _198_ = _043_ & predict_branch_taken_t0;
assign _154_ = { _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_, _273_ } & csr_depc_i_t0;
assign _156_ = { _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_, _272_ } & predict_branch_pc_t0;
assign _158_ = { _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_ } & branch_target_ex_i_t0;
assign _160_ = { _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_ } & exc_pc_t0;
assign _162_ = { _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_, _060_ } & _251_;
assign _164_ = { _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_ } & { csr_mtvec_i_t0[31:8], 1'h0, irq_vec_t0, 2'h0 };
assign _191_ = { branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req, branch_req } & { fetch_addr_n_t0[31:1], 1'h0 };
assign _193_ = { \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr  } & \gen_dummy_instr.dummy_instr_data_t0 ;
assign _195_ = { \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q  } & \g_branch_predictor.instr_skid_data_q_t0 ;
assign _197_ = { \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q , \g_branch_predictor.instr_skid_valid_q  } & \g_branch_predictor.instr_skid_addr_q_t0 ;
assign _199_ = \g_branch_predictor.instr_skid_valid_q  & \g_branch_predictor.instr_skid_bp_taken_q_t0 ;
assign _249_ = _153_ | _154_;
assign _251_ = _155_ | _156_;
assign _253_ = _157_ | _158_;
assign _255_ = _159_ | _160_;
assign fetch_addr_n_t0 = _161_ | _162_;
assign _258_ = _163_ | _164_;
assign prefetch_addr_t0 = _190_ | _191_;
assign instr_out_t0 = _192_ | _193_;
assign if_instr_rdata_t0 = _194_ | _195_;
assign pc_if_o_t0 = _196_ | _197_;
assign \g_branch_predictor.instr_bp_taken_d_t0  = _198_ | _199_;
assign _044_ = ~ instr_intg_err;
assign _045_ = ~ branch_req;
assign _046_ = ~ pc_set_i;
assign _047_ = ~ pmp_err_if_i;
assign _048_ = ~ if_instr_bus_err;
assign _049_ = ~ _002_;
assign _050_ = ~ _006_;
assign _051_ = ~ \g_secure_pc.prev_instr_seq_q ;
assign _052_ = ~ _020_;
assign _053_ = ~ fetch_valid;
assign _054_ = ~ nt_branch_mispredict_i;
assign _055_ = ~ predict_branch_taken;
assign _056_ = ~ if_instr_pmp_err;
assign _057_ = ~ fetch_err_plus2;
assign _058_ = ~ _008_;
assign _059_ = ~ _024_;
assign _165_ = branch_req_t0 & _054_;
assign _168_ = pc_set_i_t0 & _055_;
assign _169_ = pmp_err_if_i_t0 & _049_;
assign _172_ = if_instr_bus_err_t0 & _056_;
assign _175_ = _003_ & _057_;
assign _178_ = _007_ & _058_;
assign _181_ = \g_secure_pc.prev_instr_seq_q_t0  & _030_;
assign _184_ = _021_ & _029_;
assign _187_ = fetch_valid_t0 & _059_;
assign instr_err_t0 = instr_bus_err_i_t0 & _044_;
assign _166_ = nt_branch_mispredict_i_t0 & _045_;
assign _170_ = _003_ & _047_;
assign _173_ = if_instr_pmp_err_t0 & _048_;
assign _176_ = fetch_err_plus2_t0 & _049_;
assign _179_ = _009_ & _050_;
assign _182_ = if_id_pipe_reg_we_t0 & _051_;
assign _185_ = \g_branch_predictor.instr_skid_en_t0  & _052_;
assign _188_ = _025_ & _053_;
assign _167_ = branch_req_t0 & nt_branch_mispredict_i_t0;
assign _171_ = pmp_err_if_i_t0 & _003_;
assign _174_ = if_instr_bus_err_t0 & if_instr_pmp_err_t0;
assign _177_ = _003_ & fetch_err_plus2_t0;
assign _180_ = _007_ & _009_;
assign _183_ = \g_secure_pc.prev_instr_seq_q_t0  & if_id_pipe_reg_we_t0;
assign _186_ = _021_ & \g_branch_predictor.instr_skid_en_t0 ;
assign _189_ = fetch_valid_t0 & _025_;
assign _236_ = _165_ | _166_;
assign _237_ = _168_ | _099_;
assign _238_ = _169_ | _170_;
assign _239_ = _172_ | _173_;
assign _240_ = _175_ | _176_;
assign _241_ = _178_ | _179_;
assign _242_ = _181_ | _182_;
assign _243_ = _184_ | _185_;
assign _244_ = _187_ | _188_;
assign prefetch_branch_t0 = _236_ | _167_;
assign branch_req_t0 = _237_ | _101_;
assign if_instr_pmp_err_t0 = _238_ | _171_;
assign if_instr_err_t0 = _239_ | _174_;
assign _269_ = _240_ | _177_;
assign instr_valid_id_d_t0 = _241_ | _180_;
assign _271_ = _242_ | _183_;
assign \g_branch_predictor.instr_skid_valid_d_t0  = _243_ | _186_;
assign if_instr_valid_t0 = _244_ | _189_;
assign _200_ = _278_ | _277_;
assign _060_ = | { _274_, _273_, _272_ };
assign _248_ = _273_ ? csr_depc_i : csr_mepc_i;
assign _250_ = _272_ ? predict_branch_pc : _248_;
assign _252_ = _276_ ? branch_target_ex_i : { boot_addr_i[31:8], 8'h80 };
assign _254_ = _275_ ? exc_pc : _252_;
assign fetch_addr_n = _060_ ? _250_ : _254_;
assign _256_ = _277_ ? 32'd437323784 : 32'd437323776;
assign _257_ = _279_ ? { csr_mtvec_i[31:8], 1'h0, irq_vec, 2'h0 } : { csr_mtvec_i[31:8], 8'h00 };
assign exc_pc = _200_ ? _256_ : _257_;
assign _259_ = ! /* src = "generated/sv2v_out.v:18046.29-18046.45" */ pc_mux_i;
assign _260_ = predict_branch_taken && /* src = "generated/sv2v_out.v:18034.28-18034.82" */ _261_;
assign _261_ = ! /* src = "generated/sv2v_out.v:18034.73-18034.82" */ pc_set_i;
assign _262_ = pc_if_o != /* src = "generated/sv2v_out.v:18289.53-18289.88" */ \g_secure_pc.prev_instr_addr_incr_buf ;
assign _263_ = ~ /* src = "generated/sv2v_out.v:18163.52-18163.72" */ instr_is_compressed;
assign _265_ = ~ /* src = "generated/sv2v_out.v:18222.97-18222.117" */ instr_valid_clear_i;
assign _266_ = ~ /* src = "generated/sv2v_out.v:18278.85-18278.98" */ if_instr_err;
assign _267_ = ~ /* src = "generated/sv2v_out.v:18317.55-18317.69" */ id_in_ready_i;
assign _264_ = ~ /* src = "generated/sv2v_out.v:18353.85-18353.95" */ fetch_err;
assign instr_err = instr_intg_err | /* src = "generated/sv2v_out.v:18065.21-18065.53" */ instr_bus_err_i;
assign prefetch_branch = branch_req | /* src = "generated/sv2v_out.v:18067.27-18067.62" */ nt_branch_mispredict_i;
assign branch_req = pc_set_i | /* src = "generated/sv2v_out.v:18158.22-18158.53" */ predict_branch_taken;
assign if_instr_pmp_err = pmp_err_if_i | /* src = "generated/sv2v_out.v:18161.28-18161.107" */ _002_;
assign if_instr_err = if_instr_bus_err | /* src = "generated/sv2v_out.v:18162.24-18162.59" */ if_instr_pmp_err;
assign _268_ = _002_ | /* src = "generated/sv2v_out.v:18163.31-18163.113" */ fetch_err_plus2;
assign instr_valid_id_d = _006_ | /* src = "generated/sv2v_out.v:18222.28-18222.118" */ _008_;
assign _270_ = \g_secure_pc.prev_instr_seq_q  | /* src = "generated/sv2v_out.v:18278.33-18278.66" */ if_id_pipe_reg_we;
assign \g_branch_predictor.instr_skid_valid_d  = _020_ | /* src = "generated/sv2v_out.v:18317.32-18317.108" */ \g_branch_predictor.instr_skid_en ;
assign if_instr_valid = fetch_valid | /* src = "generated/sv2v_out.v:18354.28-18354.88" */ _024_;
/* src = "generated/sv2v_out.v:18318.4-18322.47" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME \g_branch_predictor.instr_skid_valid_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_branch_predictor.instr_skid_valid_q  <= 1'h0;
else \g_branch_predictor.instr_skid_valid_q  <= \g_branch_predictor.instr_skid_valid_d ;
/* src = "generated/sv2v_out.v:18279.4-18283.43" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME \g_secure_pc.prev_instr_seq_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_secure_pc.prev_instr_seq_q  <= 1'h0;
else \g_secure_pc.prev_instr_seq_q  <= \g_secure_pc.prev_instr_seq_d ;
/* src = "generated/sv2v_out.v:18224.2-18232.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_valid_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_valid_id_o <= 1'h0;
else instr_valid_id_o <= instr_valid_id_d;
/* src = "generated/sv2v_out.v:18224.2-18232.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$fbb75b45794b2f101b0da3ea80b0a23d8e0474ea\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_new_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_new_id_o <= 1'h0;
else instr_new_id_o <= if_id_pipe_reg_we;
assign _272_ = pc_mux_internal == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18036.3-18044.10" */ 3'h5;
assign _273_ = pc_mux_internal == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18036.3-18044.10" */ 3'h4;
assign _274_ = pc_mux_internal == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18036.3-18044.10" */ 3'h3;
assign _275_ = pc_mux_internal == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18036.3-18044.10" */ 3'h2;
assign _276_ = pc_mux_internal == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18036.3-18044.10" */ 3'h1;
assign _277_ = exc_pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18026.3-18032.10" */ 2'h3;
assign _278_ = exc_pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18026.3-18032.10" */ 2'h2;
assign _279_ = exc_pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18026.3-18032.10" */ 2'h1;
assign irq_vec = exc_cause[6] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18024.7-18024.19|generated/sv2v_out.v:18024.3-18025.43" */ 5'h1f : exc_cause[4:0];
assign instr_intg_err = | /* src = "generated/sv2v_out.v:18059.28-18059.36" */ \g_mem_ecc.ecc_err ;
assign pc_mux_internal = _260_ ? /* src = "generated/sv2v_out.v:18034.28-18034.100" */ 3'h5 : pc_mux_i;
assign prefetch_addr = branch_req ? /* src = "generated/sv2v_out.v:18068.26-18068.84" */ { fetch_addr_n[31:1], 1'h0 } : nt_branch_addr_i;
assign instr_out = \gen_dummy_instr.insert_dummy_instr  ? /* src = "generated/sv2v_out.v:18192.24-18192.82" */ \gen_dummy_instr.dummy_instr_data  : instr_decompressed;
assign instr_is_compressed_out = \gen_dummy_instr.insert_dummy_instr  ? /* src = "generated/sv2v_out.v:18193.38-18193.85" */ 1'h0 : instr_is_compressed;
assign illegal_c_instr_out = \gen_dummy_instr.insert_dummy_instr  ? /* src = "generated/sv2v_out.v:18194.34-18194.76" */ 1'h0 : illegal_c_insn;
assign instr_err_out = \gen_dummy_instr.insert_dummy_instr  ? /* src = "generated/sv2v_out.v:18195.28-18195.68" */ 1'h0 : if_instr_err;
assign _062_ = instr_is_compressed_id_o ? /* src = "generated/sv2v_out.v:18284.45-18284.85" */ 32'd2 : 32'd4;
assign if_instr_rdata = \g_branch_predictor.instr_skid_valid_q  ? /* src = "generated/sv2v_out.v:18355.29-18355.81" */ \g_branch_predictor.instr_skid_data_q  : fetch_rdata;
assign pc_if_o = \g_branch_predictor.instr_skid_valid_q  ? /* src = "generated/sv2v_out.v:18356.28-18356.79" */ \g_branch_predictor.instr_skid_addr_q  : fetch_addr;
assign \g_branch_predictor.instr_bp_taken_d  = \g_branch_predictor.instr_skid_valid_q  ? /* src = "generated/sv2v_out.v:18358.31-18358.96" */ \g_branch_predictor.instr_skid_bp_taken_q  : predict_branch_taken;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18164.26-18172.3" */
ibex_compressed_decoder compressed_decoder_i (
.clk_i(clk_i),
.illegal_instr_o(illegal_c_insn),
.illegal_instr_o_t0(illegal_c_insn_t0),
.instr_i(if_instr_rdata),
.instr_i_t0(if_instr_rdata_t0),
.instr_o(instr_decompressed),
.instr_o_t0(instr_decompressed_t0),
.is_compressed_o(instr_is_compressed),
.is_compressed_o_t0(instr_is_compressed_t0),
.rst_ni(rst_ni),
.valid_i(_004_),
.valid_i_t0(_005_)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18344.24-18352.5" */
ibex_branch_predict \g_branch_predictor.branch_predict_i  (
.clk_i(clk_i),
.fetch_pc_i(fetch_addr),
.fetch_pc_i_t0(fetch_addr_t0),
.fetch_rdata_i(fetch_rdata),
.fetch_rdata_i_t0(fetch_rdata_t0),
.fetch_valid_i(fetch_valid),
.fetch_valid_i_t0(fetch_valid_t0),
.predict_branch_pc_o(predict_branch_pc),
.predict_branch_pc_o_t0(predict_branch_pc_t0),
.predict_branch_taken_o(\g_branch_predictor.predict_branch_taken_raw ),
.predict_branch_taken_o_t0(\g_branch_predictor.predict_branch_taken_raw_t0 ),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18055.30-18058.5" */
prim_secded_inv_39_32_dec \g_mem_ecc.u_instr_intg_dec  (
.data_i(\g_mem_ecc.instr_rdata_buf ),
.data_i_t0(\g_mem_ecc.instr_rdata_buf_t0 ),
.err_o(\g_mem_ecc.ecc_err ),
.err_o_t0(\g_mem_ecc.ecc_err_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18051.37-18054.5" */
\$paramod\prim_buf\Width=32'00000000000000000000000000100111  \g_mem_ecc.u_prim_buf_instr_rdata  (
.in_i(instr_rdata_i),
.in_i_t0(instr_rdata_i_t0),
.out_o(\g_mem_ecc.instr_rdata_buf ),
.out_o_t0(\g_mem_ecc.instr_rdata_buf_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18285.27-18288.5" */
\$paramod\prim_buf\Width=s32'00000000000000000000000000100000  \g_secure_pc.u_prev_instr_addr_incr_buf  (
.in_i(\g_secure_pc.prev_instr_addr_incr ),
.in_i_t0(\g_secure_pc.prev_instr_addr_incr_t0 ),
.out_o(\g_secure_pc.prev_instr_addr_incr_buf ),
.out_o_t0(\g_secure_pc.prev_instr_addr_incr_buf_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18180.6-18191.5" */
\$paramod$501c60d7519704ee720c78ef16ad88cf05835059\ibex_dummy_instr  \gen_dummy_instr.dummy_instr_i  (
.clk_i(clk_i),
.dummy_instr_data_o(\gen_dummy_instr.dummy_instr_data ),
.dummy_instr_data_o_t0(\gen_dummy_instr.dummy_instr_data_t0 ),
.dummy_instr_en_i(dummy_instr_en_i),
.dummy_instr_en_i_t0(dummy_instr_en_i_t0),
.dummy_instr_mask_i(dummy_instr_mask_i),
.dummy_instr_mask_i_t0(dummy_instr_mask_i_t0),
.dummy_instr_seed_en_i(dummy_instr_seed_en_i),
.dummy_instr_seed_en_i_t0(dummy_instr_seed_en_i_t0),
.dummy_instr_seed_i(dummy_instr_seed_i),
.dummy_instr_seed_i_t0(dummy_instr_seed_i_t0),
.fetch_valid_i(fetch_valid),
.fetch_valid_i_t0(fetch_valid_t0),
.id_in_ready_i(id_in_ready_i),
.id_in_ready_i_t0(id_in_ready_i_t0),
.insert_dummy_instr_o(\gen_dummy_instr.insert_dummy_instr ),
.insert_dummy_instr_o_t0(\gen_dummy_instr.insert_dummy_instr_t0 ),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18115.48-18134.5" */
\$paramod\ibex_prefetch_buffer\ResetAll=1'1  \gen_prefetch_buffer.prefetch_buffer_i  (
.addr_i(prefetch_addr),
.addr_i_t0(prefetch_addr_t0),
.addr_o(fetch_addr),
.addr_o_t0(fetch_addr_t0),
.branch_i(prefetch_branch),
.branch_i_t0(prefetch_branch_t0),
.busy_o(if_busy_o),
.busy_o_t0(if_busy_o_t0),
.clk_i(clk_i),
.err_o(fetch_err),
.err_o_t0(fetch_err_t0),
.err_plus2_o(fetch_err_plus2),
.err_plus2_o_t0(fetch_err_plus2_t0),
.instr_addr_o(instr_addr_o),
.instr_addr_o_t0(instr_addr_o_t0),
.instr_err_i(instr_err),
.instr_err_i_t0(instr_err_t0),
.instr_gnt_i(instr_gnt_i),
.instr_gnt_i_t0(instr_gnt_i_t0),
.instr_rdata_i(instr_rdata_i[31:0]),
.instr_rdata_i_t0(instr_rdata_i_t0[31:0]),
.instr_req_o(instr_req_o),
.instr_req_o_t0(instr_req_o_t0),
.instr_rvalid_i(instr_rvalid_i),
.instr_rvalid_i_t0(instr_rvalid_i_t0),
.rdata_o(fetch_rdata),
.rdata_o_t0(fetch_rdata_t0),
.ready_i(fetch_ready),
.ready_i_t0(fetch_ready_t0),
.req_i(req_i),
.req_i_t0(req_i_t0),
.rst_ni(rst_ni),
.valid_o(fetch_valid_raw),
.valid_o_t0(fetch_valid_raw_t0)
);
assign ic_data_addr_o = 8'h00;
assign ic_data_addr_o_t0 = 8'h00;
assign ic_data_req_o = 2'h0;
assign ic_data_req_o_t0 = 2'h0;
assign ic_data_wdata_o = 64'h0000000000000000;
assign ic_data_wdata_o_t0 = 64'h0000000000000000;
assign ic_data_write_o = 1'h0;
assign ic_data_write_o_t0 = 1'h0;
assign ic_scr_key_req_o = 1'h0;
assign ic_scr_key_req_o_t0 = 1'h0;
assign ic_tag_addr_o = 8'h00;
assign ic_tag_addr_o_t0 = 8'h00;
assign ic_tag_req_o = 2'h0;
assign ic_tag_req_o_t0 = 2'h0;
assign ic_tag_wdata_o = 22'h000000;
assign ic_tag_wdata_o_t0 = 22'h000000;
assign ic_tag_write_o = 1'h0;
assign ic_tag_write_o_t0 = 1'h0;
assign icache_ecc_error_o = 1'h0;
assign icache_ecc_error_o_t0 = 1'h0;
assign instr_rdata_id_o = instr_rdata_alu_id_o;
assign instr_rdata_id_o_t0 = instr_rdata_alu_id_o_t0;
endmodule

module \$paramod\ibex_alu\RV32B=s32'00000000000000000000000000000000 (operator_i, operand_a_i, operand_b_i, instr_first_cycle_i, multdiv_operand_a_i, multdiv_operand_b_i, multdiv_sel_i, imd_val_q_i, imd_val_d_o, imd_val_we_o, adder_result_o, adder_result_ext_o, result_o, comparison_result_o, is_equal_result_o, adder_result_ext_o_t0, adder_result_o_t0, comparison_result_o_t0, is_equal_result_o_t0, multdiv_operand_a_i_t0, multdiv_operand_b_i_t0
, multdiv_sel_i_t0, operand_a_i_t0, operand_b_i_t0, result_o_t0, imd_val_d_o_t0, imd_val_q_i_t0, instr_first_cycle_i_t0, imd_val_we_o_t0, operator_i_t0);
/* src = "generated/sv2v_out.v:11462.52-11462.83" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11462.52-11462.83" */
wire _001_;
wire [33:0] _002_;
wire [33:0] _003_;
wire [31:0] _004_;
wire [31:0] _005_;
wire [31:0] _006_;
wire _007_;
wire [31:0] _008_;
wire [31:0] _009_;
wire _010_;
wire [32:0] _011_;
wire [32:0] _012_;
wire [31:0] _013_;
wire [31:0] _014_;
wire [31:0] _015_;
wire _016_;
wire [33:0] _017_;
wire [33:0] _018_;
wire [31:0] _019_;
wire [31:0] _020_;
wire [31:0] _021_;
wire [31:0] _022_;
wire [31:0] _023_;
wire [31:0] _024_;
wire [31:0] _025_;
wire [31:0] _026_;
wire [31:0] _027_;
wire _028_;
wire _029_;
wire [31:0] _030_;
wire [31:0] _031_;
wire [31:0] _032_;
wire [31:0] _033_;
wire [31:0] _034_;
wire [31:0] _035_;
wire _036_;
wire _037_;
wire [32:0] _038_;
wire [32:0] _039_;
wire [32:0] _040_;
wire [32:0] _041_;
wire [32:0] _042_;
wire [32:0] _043_;
wire [31:0] _044_;
wire [31:0] _045_;
wire [31:0] _046_;
wire [31:0] _047_;
wire _048_;
wire _049_;
wire [33:0] _050_;
wire [33:0] _051_;
wire [33:0] _052_;
wire [31:0] _053_;
wire [31:0] _054_;
wire [33:0] _055_;
wire [33:0] _056_;
wire [33:0] _057_;
wire [31:0] _058_;
/* cellift = 32'd1 */
wire [31:0] _059_;
wire [31:0] _060_;
/* cellift = 32'd1 */
wire [31:0] _061_;
wire [31:0] _062_;
/* cellift = 32'd1 */
wire [31:0] _063_;
wire _064_;
/* cellift = 32'd1 */
wire _065_;
wire _066_;
/* src = "generated/sv2v_out.v:11383.23-11383.47" */
wire _067_;
/* src = "generated/sv2v_out.v:11491.23-11491.41" */
wire _068_;
/* src = "generated/sv2v_out.v:11491.46-11491.64" */
wire _069_;
/* src = "generated/sv2v_out.v:11492.24-11492.42" */
wire _070_;
/* src = "generated/sv2v_out.v:11492.47-11492.65" */
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
/* src = "generated/sv2v_out.v:11390.24-11390.33" */
wire _088_;
/* src = "generated/sv2v_out.v:11392.59-11392.76" */
wire _089_;
wire [7:0] _090_;
wire _091_;
wire [4:0] _092_;
wire _093_;
wire [4:0] _094_;
wire _095_;
wire [5:0] _096_;
wire _097_;
wire [31:0] _098_;
/* cellift = 32'd1 */
wire [31:0] _099_;
wire [5:0] _100_;
wire _101_;
wire [3:0] _102_;
wire _103_;
wire _104_;
wire [32:0] _105_;
/* cellift = 32'd1 */
wire [32:0] _106_;
/* src = "generated/sv2v_out.v:11429.27-11429.48" */
/* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] _107_;
/* src = "generated/sv2v_out.v:11382.8-11382.41" */
wire _108_;
/* src = "generated/sv2v_out.v:11385.23-11385.51" */
wire _109_;
/* src = "generated/sv2v_out.v:11330.13-11330.23" */
wire [32:0] adder_in_a;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11330.13-11330.23" */
wire [32:0] adder_in_a_t0;
/* src = "generated/sv2v_out.v:11331.13-11331.23" */
wire [32:0] adder_in_b;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11331.13-11331.23" */
wire [32:0] adder_in_b_t0;
/* src = "generated/sv2v_out.v:11329.6-11329.23" */
wire adder_op_b_negate;
/* src = "generated/sv2v_out.v:11314.21-11314.39" */
output [33:0] adder_result_ext_o;
wire [33:0] adder_result_ext_o;
/* cellift = 32'd1 */
output [33:0] adder_result_ext_o_t0;
wire [33:0] adder_result_ext_o_t0;
/* src = "generated/sv2v_out.v:11313.21-11313.35" */
output [31:0] adder_result_o;
wire [31:0] adder_result_o;
/* cellift = 32'd1 */
output [31:0] adder_result_o_t0;
wire [31:0] adder_result_o_t0;
/* src = "generated/sv2v_out.v:11474.7-11474.18" */
wire bwlogic_and;
/* src = "generated/sv2v_out.v:11477.14-11477.32" */
wire [31:0] bwlogic_and_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11477.14-11477.32" */
wire [31:0] bwlogic_and_result_t0;
/* src = "generated/sv2v_out.v:11473.7-11473.17" */
wire bwlogic_or;
/* src = "generated/sv2v_out.v:11476.14-11476.31" */
wire [31:0] bwlogic_or_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11476.14-11476.31" */
wire [31:0] bwlogic_or_result_t0;
/* src = "generated/sv2v_out.v:11479.13-11479.27" */
wire [31:0] bwlogic_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11479.13-11479.27" */
wire [31:0] bwlogic_result_t0;
/* src = "generated/sv2v_out.v:11478.14-11478.32" */
wire [31:0] bwlogic_xor_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11478.14-11478.32" */
wire [31:0] bwlogic_xor_result_t0;
/* src = "generated/sv2v_out.v:11373.6-11373.16" */
wire cmp_signed;
/* src = "generated/sv2v_out.v:11316.14-11316.33" */
output comparison_result_o;
wire comparison_result_o;
/* cellift = 32'd1 */
output comparison_result_o_t0;
wire comparison_result_o_t0;
/* src = "generated/sv2v_out.v:11311.20-11311.31" */
output [63:0] imd_val_d_o;
wire [63:0] imd_val_d_o;
/* cellift = 32'd1 */
output [63:0] imd_val_d_o_t0;
wire [63:0] imd_val_d_o_t0;
/* src = "generated/sv2v_out.v:11310.20-11310.31" */
input [63:0] imd_val_q_i;
wire [63:0] imd_val_q_i;
/* cellift = 32'd1 */
input [63:0] imd_val_q_i_t0;
wire [63:0] imd_val_q_i_t0;
/* src = "generated/sv2v_out.v:11312.19-11312.31" */
output [1:0] imd_val_we_o;
wire [1:0] imd_val_we_o;
/* cellift = 32'd1 */
output [1:0] imd_val_we_o_t0;
wire [1:0] imd_val_we_o_t0;
/* src = "generated/sv2v_out.v:11306.13-11306.32" */
input instr_first_cycle_i;
wire instr_first_cycle_i;
/* cellift = 32'd1 */
input instr_first_cycle_i_t0;
wire instr_first_cycle_i_t0;
/* src = "generated/sv2v_out.v:11317.14-11317.31" */
output is_equal_result_o;
wire is_equal_result_o;
/* cellift = 32'd1 */
output is_equal_result_o_t0;
wire is_equal_result_o_t0;
/* src = "generated/sv2v_out.v:11372.6-11372.22" */
wire is_greater_equal;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11372.6-11372.22" */
wire is_greater_equal_t0;
/* src = "generated/sv2v_out.v:11307.20-11307.39" */
input [32:0] multdiv_operand_a_i;
wire [32:0] multdiv_operand_a_i;
/* cellift = 32'd1 */
input [32:0] multdiv_operand_a_i_t0;
wire [32:0] multdiv_operand_a_i_t0;
/* src = "generated/sv2v_out.v:11308.20-11308.39" */
input [32:0] multdiv_operand_b_i;
wire [32:0] multdiv_operand_b_i;
/* cellift = 32'd1 */
input [32:0] multdiv_operand_b_i_t0;
wire [32:0] multdiv_operand_b_i_t0;
/* src = "generated/sv2v_out.v:11309.13-11309.26" */
input multdiv_sel_i;
wire multdiv_sel_i;
/* cellift = 32'd1 */
input multdiv_sel_i_t0;
wire multdiv_sel_i_t0;
/* src = "generated/sv2v_out.v:11304.20-11304.31" */
input [31:0] operand_a_i;
wire [31:0] operand_a_i;
/* cellift = 32'd1 */
input [31:0] operand_a_i_t0;
wire [31:0] operand_a_i_t0;
/* src = "generated/sv2v_out.v:11305.20-11305.31" */
input [31:0] operand_b_i;
wire [31:0] operand_b_i;
/* cellift = 32'd1 */
input [31:0] operand_b_i_t0;
wire [31:0] operand_b_i_t0;
/* src = "generated/sv2v_out.v:11319.14-11319.27" */
wire [32:0] operand_b_neg;
/* src = "generated/sv2v_out.v:11303.19-11303.29" */
input [6:0] operator_i;
wire [6:0] operator_i;
/* cellift = 32'd1 */
input [6:0] operator_i_t0;
wire [6:0] operator_i_t0;
/* src = "generated/sv2v_out.v:11315.20-11315.28" */
output [31:0] result_o;
wire [31:0] result_o;
/* cellift = 32'd1 */
output [31:0] result_o_t0;
wire [31:0] result_o_t0;
/* src = "generated/sv2v_out.v:11401.12-11401.21" */
wire [5:0] shift_amt;
/* src = "generated/sv2v_out.v:11402.13-11402.28" */
/* unused_bits = "5" */
wire [5:0] shift_amt_compl;
/* src = "generated/sv2v_out.v:11398.7-11398.18" */
wire shift_arith;
/* src = "generated/sv2v_out.v:11396.6-11396.16" */
wire shift_left;
/* src = "generated/sv2v_out.v:11403.13-11403.26" */
wire [31:0] shift_operand;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11403.13-11403.26" */
wire [31:0] shift_operand_t0;
/* src = "generated/sv2v_out.v:11407.13-11407.25" */
wire [31:0] shift_result;
/* src = "generated/sv2v_out.v:11405.13-11405.29" */
/* unused_bits = "32" */
wire [32:0] shift_result_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11405.13-11405.29" */
/* unused_bits = "32" */
wire [32:0] shift_result_ext_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11407.13-11407.25" */
wire [31:0] shift_result_t0;
assign adder_result_ext_o = { 1'h0, adder_in_a } + /* src = "generated/sv2v_out.v:11368.30-11368.75" */ { 1'h0, adder_in_b };
assign _000_ = shift_arith & /* src = "generated/sv2v_out.v:11462.52-11462.83" */ shift_operand[31];
assign bwlogic_and_result = operand_a_i & /* src = "generated/sv2v_out.v:11489.30-11489.61" */ operand_b_i;
assign _002_ = ~ { 1'h0, adder_in_a_t0 };
assign _003_ = ~ { 1'h0, adder_in_b_t0 };
assign _017_ = { 1'h0, adder_in_a } & _002_;
assign _018_ = { 1'h0, adder_in_b } & _003_;
assign _056_ = _017_ + _018_;
assign _050_ = { 1'h0, adder_in_a } | { 1'h0, adder_in_a_t0 };
assign _051_ = { 1'h0, adder_in_b } | { 1'h0, adder_in_b_t0 };
assign _057_ = _050_ + _051_;
assign _055_ = _056_ ^ _057_;
assign _052_ = _055_ | { 1'h0, adder_in_a_t0 };
assign adder_result_ext_o_t0 = _052_ | { 1'h0, adder_in_b_t0 };
assign _019_ = operand_a_i_t0 & operand_b_i;
assign _001_ = shift_operand_t0[31] & shift_arith;
assign _020_ = operand_b_i_t0 & operand_a_i;
assign _021_ = operand_a_i_t0 & operand_b_i_t0;
assign _053_ = _019_ | _020_;
assign bwlogic_and_result_t0 = _053_ | _021_;
assign _004_ = ~ { _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_ };
assign _005_ = ~ { _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_ };
assign _006_ = ~ { _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_ };
assign _008_ = ~ { bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and };
assign _009_ = ~ { bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or };
assign _010_ = ~ _108_;
assign _011_ = ~ { adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate };
assign _012_ = ~ { multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i };
assign _013_ = ~ { shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left };
assign _022_ = _004_ & shift_result_t0;
assign _024_ = _005_ & _061_;
assign _026_ = _006_ & _063_;
assign _028_ = _007_ & is_greater_equal_t0;
assign _032_ = _008_ & bwlogic_xor_result_t0;
assign _034_ = _009_ & _099_;
assign _036_ = _010_ & adder_result_ext_o_t0[32];
assign _038_ = _011_ & { operand_b_i_t0, 1'h0 };
assign _040_ = _012_ & _106_;
assign _042_ = _012_ & { operand_a_i_t0, 1'h0 };
assign _044_ = _013_ & operand_a_i_t0;
assign _046_ = _013_ & shift_result_ext_t0[31:0];
assign _023_ = { _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_, _091_ } & { 31'h00000000, comparison_result_o_t0 };
assign _061_ = { _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_, _097_ } & bwlogic_result_t0;
assign _025_ = { _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_, _095_ } & adder_result_ext_o_t0[32:1];
assign _027_ = { _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_, _048_ } & _059_;
assign _029_ = _101_ & is_greater_equal_t0;
assign comparison_result_o_t0 = _049_ & _065_;
assign _033_ = { bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and } & bwlogic_and_result_t0;
assign _035_ = { bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or } & bwlogic_or_result_t0;
assign _037_ = _108_ & operand_a_i_t0[31];
assign _039_ = { adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate } & { operand_b_i_t0, 1'h0 };
assign _041_ = { multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i } & multdiv_operand_b_i_t0;
assign _043_ = { multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i } & multdiv_operand_a_i_t0;
assign _045_ = { shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left } & { operand_a_i_t0[0], operand_a_i_t0[1], operand_a_i_t0[2], operand_a_i_t0[3], operand_a_i_t0[4], operand_a_i_t0[5], operand_a_i_t0[6], operand_a_i_t0[7], operand_a_i_t0[8], operand_a_i_t0[9], operand_a_i_t0[10], operand_a_i_t0[11], operand_a_i_t0[12], operand_a_i_t0[13], operand_a_i_t0[14], operand_a_i_t0[15], operand_a_i_t0[16], operand_a_i_t0[17], operand_a_i_t0[18], operand_a_i_t0[19], operand_a_i_t0[20], operand_a_i_t0[21], operand_a_i_t0[22], operand_a_i_t0[23], operand_a_i_t0[24], operand_a_i_t0[25], operand_a_i_t0[26], operand_a_i_t0[27], operand_a_i_t0[28], operand_a_i_t0[29], operand_a_i_t0[30], operand_a_i_t0[31] };
assign _047_ = { shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left } & { shift_result_ext_t0[0], shift_result_ext_t0[1], shift_result_ext_t0[2], shift_result_ext_t0[3], shift_result_ext_t0[4], shift_result_ext_t0[5], shift_result_ext_t0[6], shift_result_ext_t0[7], shift_result_ext_t0[8], shift_result_ext_t0[9], shift_result_ext_t0[10], shift_result_ext_t0[11], shift_result_ext_t0[12], shift_result_ext_t0[13], shift_result_ext_t0[14], shift_result_ext_t0[15], shift_result_ext_t0[16], shift_result_ext_t0[17], shift_result_ext_t0[18], shift_result_ext_t0[19], shift_result_ext_t0[20], shift_result_ext_t0[21], shift_result_ext_t0[22], shift_result_ext_t0[23], shift_result_ext_t0[24], shift_result_ext_t0[25], shift_result_ext_t0[26], shift_result_ext_t0[27], shift_result_ext_t0[28], shift_result_ext_t0[29], shift_result_ext_t0[30], shift_result_ext_t0[31] };
assign _059_ = _022_ | _023_;
assign _063_ = _024_ | _025_;
assign result_o_t0 = _026_ | _027_;
assign _065_ = _028_ | _029_;
assign _099_ = _032_ | _033_;
assign bwlogic_result_t0 = _034_ | _035_;
assign is_greater_equal_t0 = _036_ | _037_;
assign _106_ = _038_ | _039_;
assign adder_in_b_t0 = _040_ | _041_;
assign adder_in_a_t0 = _042_ | _043_;
assign shift_operand_t0 = _044_ | _045_;
assign shift_result_t0 = _046_ | _047_;
assign operand_b_neg = ~ { operand_b_i, 1'h0 };
assign _014_ = ~ operand_a_i;
assign _007_ = ~ _101_;
assign _015_ = ~ operand_b_i;
assign _030_ = operand_a_i_t0 & _015_;
assign _031_ = operand_b_i_t0 & _014_;
assign _054_ = _030_ | _031_;
assign bwlogic_or_result_t0 = _054_ | _021_;
assign _048_ = _093_ | _091_;
assign _049_ = _103_ | _101_;
assign _058_ = _091_ ? { 31'h00000000, comparison_result_o } : shift_result;
assign _060_ = _097_ ? bwlogic_result : 32'd0;
assign _062_ = _095_ ? adder_result_ext_o[32:1] : _060_;
assign result_o = _048_ ? _058_ : _062_;
assign _064_ = _101_ ? _089_ : is_greater_equal;
assign _066_ = _090_[1] ? _088_ : is_equal_result_o;
assign comparison_result_o = _049_ ? _064_ : _066_;
assign shift_result_ext_t0 = { _001_, shift_operand_t0 } >>> shift_amt[4:0];
assign bwlogic_xor_result_t0 = operand_a_i_t0 | operand_b_i_t0;
assign is_equal_result_o = ! /* src = "generated/sv2v_out.v:11379.20-11379.72" */ adder_result_ext_o[32:1];
assign _067_ = ~ /* src = "generated/sv2v_out.v:11383.23-11383.47" */ adder_result_ext_o[32];
assign _016_ = operator_i[5] ? _073_ : _072_;
assign _072_ = operator_i[4] ? _075_ : _074_;
assign _073_ = operator_i[4] ? 1'h0 : _076_;
assign _074_ = operator_i[3] ? 1'h0 : _077_;
assign _075_ = operator_i[3] ? _078_ : 1'h0;
assign _076_ = operator_i[3] ? _080_ : _079_;
assign _077_ = operator_i[2] ? 1'h0 : _081_;
assign _078_ = operator_i[2] ? 1'h1 : _082_;
assign _079_ = operator_i[2] ? 1'h0 : _083_;
assign _080_ = operator_i[2] ? _085_ : _084_;
assign _081_ = operator_i[1] ? 1'h0 : _086_;
assign _084_ = operator_i[1] ? _086_ : 1'h0;
assign _085_ = operator_i[1] ? 1'h0 : _087_;
assign _082_ = operator_i[1] ? 1'h1 : _086_;
assign _083_ = operator_i[1] ? _087_ : 1'h1;
assign _087_ = operator_i[0] ? 1'h0 : 1'h1;
assign _086_ = operator_i[0] ? 1'h1 : 1'h0;
assign _088_ = ~ /* src = "generated/sv2v_out.v:11390.24-11390.33" */ is_equal_result_o;
assign _089_ = ~ /* src = "generated/sv2v_out.v:11392.59-11392.76" */ is_greater_equal;
assign bwlogic_or_result = operand_a_i | /* src = "generated/sv2v_out.v:11488.29-11488.60" */ operand_b_i;
assign bwlogic_or = _068_ | /* src = "generated/sv2v_out.v:11491.22-11491.65" */ _069_;
assign bwlogic_and = _070_ | /* src = "generated/sv2v_out.v:11492.23-11492.66" */ _071_;
assign _091_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ _090_;
assign _090_[0] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ 7'h1d;
assign _093_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ { _092_[4:3], _092_[1:0], shift_arith };
assign _092_[1] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ 7'h09;
assign shift_arith = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ 7'h08;
assign _092_[3] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ 7'h0c;
assign _092_[4] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ 7'h0b;
assign _095_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ _094_;
assign _094_[0] = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ operator_i;
assign _094_[1] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ 7'h01;
assign _094_[2] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ 7'h16;
assign _094_[3] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ 7'h17;
assign _094_[4] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ 7'h18;
assign _097_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ { _096_[1:0], _071_, _070_, _069_, _068_ };
assign _096_[0] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ 7'h02;
assign _096_[1] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ 7'h05;
assign _068_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ 7'h03;
assign _069_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ 7'h06;
assign _070_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ 7'h04;
assign _071_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12023.3-12041.10" */ 7'h07;
assign _098_ = bwlogic_and ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11494.3-11498.10" */ bwlogic_and_result : bwlogic_xor_result;
assign bwlogic_result = bwlogic_or ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11494.3-11498.10" */ bwlogic_or_result : _098_;
assign shift_left = _092_[0] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11437.3-11446.10" */ 1'h1 : 1'h0;
assign _092_[0] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11437.3-11446.10" */ 7'h0a;
assign _101_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11388.3-11394.10" */ { _100_[3:2], _090_[7:4] };
assign _090_[4] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11388.3-11394.10" */ 7'h19;
assign _090_[5] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11388.3-11394.10" */ 7'h1a;
assign _100_[2] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11388.3-11394.10" */ 7'h1f;
assign _100_[3] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11388.3-11394.10" */ 7'h20;
assign _090_[6] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11388.3-11394.10" */ 7'h2b;
assign _090_[7] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11388.3-11394.10" */ 7'h2c;
assign _103_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11388.3-11394.10" */ { _102_[3:2], _090_[3:2] };
assign _090_[3] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11388.3-11394.10" */ 7'h1c;
assign _102_[2] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11388.3-11394.10" */ 7'h21;
assign _102_[3] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11388.3-11394.10" */ 7'h22;
assign _090_[1] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11388.3-11394.10" */ 7'h1e;
assign is_greater_equal = _108_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:11382.7-11382.50|generated/sv2v_out.v:11382.3-11385.52" */ _109_ : _067_;
assign cmp_signed = _104_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11375.3-11378.10" */ 1'h1 : 1'h0;
assign _104_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11375.3-11378.10" */ { _102_[2], _100_[2], _090_[6], _090_[4], _090_[2] };
assign _090_[2] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11375.3-11378.10" */ 7'h1b;
assign _105_ = adder_op_b_negate ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11363.3-11367.10" */ operand_b_neg : { operand_b_i, 1'h0 };
assign adder_in_b = multdiv_sel_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11363.3-11367.10" */ multdiv_operand_b_i : _105_;
assign adder_in_a = multdiv_sel_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11354.3-11360.10" */ multdiv_operand_a_i : { operand_a_i, 1'h1 };
assign adder_op_b_negate = operator_i[6] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:11338.3-11351.10" */ 1'h0 : _016_;
assign shift_result_ext = $signed({ _000_, shift_operand }) >>> /* src = "generated/sv2v_out.v:11462.29-11462.120" */ shift_amt[4:0];
assign { _107_[31:6], shift_amt_compl } = 32'd32 - /* src = "generated/sv2v_out.v:11429.27-11429.48" */ operand_b_i[4:0];
assign shift_amt[4:0] = instr_first_cycle_i ? /* src = "generated/sv2v_out.v:11434.22-11434.195" */ operand_b_i[4:0] : shift_amt_compl[4:0];
assign shift_operand = shift_left ? /* src = "generated/sv2v_out.v:11455.21-11455.61" */ { operand_a_i[0], operand_a_i[1], operand_a_i[2], operand_a_i[3], operand_a_i[4], operand_a_i[5], operand_a_i[6], operand_a_i[7], operand_a_i[8], operand_a_i[9], operand_a_i[10], operand_a_i[11], operand_a_i[12], operand_a_i[13], operand_a_i[14], operand_a_i[15], operand_a_i[16], operand_a_i[17], operand_a_i[18], operand_a_i[19], operand_a_i[20], operand_a_i[21], operand_a_i[22], operand_a_i[23], operand_a_i[24], operand_a_i[25], operand_a_i[26], operand_a_i[27], operand_a_i[28], operand_a_i[29], operand_a_i[30], operand_a_i[31] } : operand_a_i;
assign shift_result = shift_left ? /* src = "generated/sv2v_out.v:11471.19-11471.63" */ { shift_result_ext[0], shift_result_ext[1], shift_result_ext[2], shift_result_ext[3], shift_result_ext[4], shift_result_ext[5], shift_result_ext[6], shift_result_ext[7], shift_result_ext[8], shift_result_ext[9], shift_result_ext[10], shift_result_ext[11], shift_result_ext[12], shift_result_ext[13], shift_result_ext[14], shift_result_ext[15], shift_result_ext[16], shift_result_ext[17], shift_result_ext[18], shift_result_ext[19], shift_result_ext[20], shift_result_ext[21], shift_result_ext[22], shift_result_ext[23], shift_result_ext[24], shift_result_ext[25], shift_result_ext[26], shift_result_ext[27], shift_result_ext[28], shift_result_ext[29], shift_result_ext[30], shift_result_ext[31] } : shift_result_ext[31:0];
assign _108_ = operand_a_i[31] ^ /* src = "generated/sv2v_out.v:11382.8-11382.41" */ operand_b_i[31];
assign _109_ = operand_a_i[31] ^ /* src = "generated/sv2v_out.v:11385.23-11385.51" */ cmp_signed;
assign bwlogic_xor_result = operand_a_i ^ /* src = "generated/sv2v_out.v:11490.30-11490.61" */ operand_b_i;
assign _092_[2] = shift_arith;
assign _096_[5:2] = { _071_, _070_, _069_, _068_ };
assign { _100_[5:4], _100_[1:0] } = _090_[7:4];
assign _102_[1:0] = _090_[3:2];
assign _107_[5:0] = shift_amt_compl;
assign adder_result_o = adder_result_ext_o[32:1];
assign adder_result_o_t0 = adder_result_ext_o_t0[32:1];
assign imd_val_d_o = 64'h0000000000000000;
assign imd_val_d_o_t0 = 64'h0000000000000000;
assign imd_val_we_o = 2'h0;
assign imd_val_we_o_t0 = 2'h0;
assign is_equal_result_o_t0 = 1'h0;
assign shift_amt[5] = 1'h0;
endmodule

module \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1 (clk_i, rst_ni, ctrl_busy_o, illegal_insn_i, ecall_insn_i, mret_insn_i, dret_insn_i, wfi_insn_i, ebrk_insn_i, csr_pipe_flush_i, instr_valid_i, instr_i, instr_compressed_i, instr_is_compressed_i, instr_bp_taken_i, instr_fetch_err_i, instr_fetch_err_plus2_i, pc_id_i, instr_valid_clear_o, id_in_ready_o, controller_run_o
, instr_exec_i, instr_req_o, pc_set_o, pc_mux_o, nt_branch_mispredict_o, exc_pc_mux_o, exc_cause_o, lsu_addr_last_i, load_err_i, store_err_i, mem_resp_intg_err_i, wb_exception_o, id_exception_o, branch_set_i, branch_not_set_i, jump_set_i, csr_mstatus_mie_i, irq_pending_i, irqs_i, irq_nm_ext_i, nmi_mode_o
, debug_req_i, debug_cause_o, debug_csr_save_o, debug_mode_o, debug_mode_entering_o, debug_single_step_i, debug_ebreakm_i, debug_ebreaku_i, trigger_match_i, csr_save_if_o, csr_save_id_o, csr_save_wb_o, csr_restore_mret_id_o, csr_restore_dret_id_o, csr_save_cause_o, csr_mtval_o, priv_mode_i, stall_id_i, stall_wb_i, flush_id_o, ready_wb_i
, perf_jump_o, perf_tbranch_o, wfi_insn_i_t0, wb_exception_o_t0, trigger_match_i_t0, store_err_i_t0, debug_cause_o_t0, debug_csr_save_o_t0, debug_ebreakm_i_t0, debug_ebreaku_i_t0, debug_mode_entering_o_t0, debug_mode_o_t0, debug_req_i_t0, debug_single_step_i_t0, dret_insn_i_t0, ebrk_insn_i_t0, ecall_insn_i_t0, exc_cause_o_t0, exc_pc_mux_o_t0, flush_id_o_t0, id_exception_o_t0
, id_in_ready_o_t0, illegal_insn_i_t0, instr_bp_taken_i_t0, instr_compressed_i_t0, instr_exec_i_t0, instr_fetch_err_i_t0, instr_fetch_err_plus2_i_t0, instr_is_compressed_i_t0, instr_valid_clear_o_t0, instr_valid_i_t0, irq_nm_ext_i_t0, irq_pending_i_t0, irqs_i_t0, jump_set_i_t0, load_err_i_t0, lsu_addr_last_i_t0, mem_resp_intg_err_i_t0, mret_insn_i_t0, nmi_mode_o_t0, nt_branch_mispredict_o_t0, stall_wb_i_t0
, pc_id_i_t0, pc_mux_o_t0, pc_set_o_t0, branch_not_set_i_t0, branch_set_i_t0, controller_run_o_t0, perf_jump_o_t0, csr_mstatus_mie_i_t0, perf_tbranch_o_t0, priv_mode_i_t0, csr_mtval_o_t0, ready_wb_i_t0, csr_pipe_flush_i_t0, stall_id_i_t0, csr_restore_dret_id_o_t0, csr_restore_mret_id_o_t0, csr_save_cause_o_t0, csr_save_id_o_t0, csr_save_if_o_t0, csr_save_wb_o_t0, ctrl_busy_o_t0
, instr_i_t0, instr_req_o_t0);
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [3:0] _000_;
/* src = "generated/sv2v_out.v:12506.2-12514.5" */
wire [3:0] _001_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [3:0] _002_;
/* src = "generated/sv2v_out.v:12506.2-12514.5" */
wire [3:0] _003_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [3:0] _004_;
/* src = "generated/sv2v_out.v:12506.2-12514.5" */
wire [3:0] _005_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [3:0] _006_;
/* src = "generated/sv2v_out.v:12506.2-12514.5" */
wire [3:0] _007_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [3:0] _008_;
/* src = "generated/sv2v_out.v:12506.2-12514.5" */
wire [3:0] _009_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [3:0] _010_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [3:0] _011_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [3:0] _012_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _013_;
/* src = "generated/sv2v_out.v:12506.2-12514.5" */
wire [3:0] _014_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [31:0] _015_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [31:0] _016_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _017_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _018_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _019_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _020_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _021_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _022_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _023_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [3:0] _024_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _025_;
/* src = "generated/sv2v_out.v:12410.4-12429.7" */
wire _026_;
/* src = "generated/sv2v_out.v:12410.4-12429.7" */
wire _027_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [6:0] _028_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [1:0] _029_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _030_;
/* src = "generated/sv2v_out.v:12464.4-12476.7" */
wire _031_;
/* src = "generated/sv2v_out.v:12464.4-12476.7" */
wire _032_;
/* src = "generated/sv2v_out.v:12410.4-12429.7" */
wire _033_;
/* src = "generated/sv2v_out.v:12410.4-12429.7" */
wire _034_;
/* src = "generated/sv2v_out.v:12410.4-12429.7" */
wire _035_;
/* src = "generated/sv2v_out.v:12506.2-12514.5" */
wire [3:0] _036_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _037_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _038_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _039_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [2:0] _040_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _041_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _042_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _043_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _044_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _045_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _046_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _047_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [31:0] _048_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [31:0] _049_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _050_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _051_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _052_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _053_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _054_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _055_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [3:0] _056_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _057_;
/* src = "generated/sv2v_out.v:12410.4-12429.7" */
wire _058_;
/* src = "generated/sv2v_out.v:12410.4-12429.7" */
wire _059_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [6:0] _060_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _061_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _062_;
/* src = "generated/sv2v_out.v:12410.4-12429.7" */
wire _063_;
/* src = "generated/sv2v_out.v:12410.4-12429.7" */
wire _064_;
/* src = "generated/sv2v_out.v:12506.2-12514.5" */
wire [3:0] _065_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _066_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _067_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [2:0] _068_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [31:0] _069_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [31:0] _070_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _071_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _072_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _073_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [3:0] _074_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _075_;
/* src = "generated/sv2v_out.v:12410.4-12429.7" */
wire _076_;
/* src = "generated/sv2v_out.v:12410.4-12429.7" */
wire _077_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [6:0] _078_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _079_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _080_;
/* src = "generated/sv2v_out.v:12410.4-12429.7" */
wire _081_;
/* src = "generated/sv2v_out.v:12506.2-12514.5" */
wire [3:0] _082_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _083_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _084_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [2:0] _085_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _086_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [31:0] _087_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [31:0] _088_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _089_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _090_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [3:0] _091_;
/* src = "generated/sv2v_out.v:12410.4-12429.7" */
wire _092_;
/* src = "generated/sv2v_out.v:12410.4-12429.7" */
wire _093_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [6:0] _094_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _095_;
/* src = "generated/sv2v_out.v:12506.2-12514.5" */
wire [3:0] _096_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _097_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _098_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [31:0] _099_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [31:0] _100_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _101_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _102_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [3:0] _103_;
/* src = "generated/sv2v_out.v:12410.4-12429.7" */
wire _104_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [6:0] _105_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _106_;
/* src = "generated/sv2v_out.v:12506.2-12514.5" */
wire [3:0] _107_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [3:0] _108_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [6:0] _109_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _110_;
/* src = "generated/sv2v_out.v:12506.2-12514.5" */
wire [3:0] _111_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire _112_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [3:0] _113_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [6:0] _114_;
/* src = "generated/sv2v_out.v:12506.2-12514.5" */
wire [3:0] _115_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [3:0] _116_;
/* src = "generated/sv2v_out.v:12539.2-12757.5" */
wire [6:0] _117_;
/* src = "generated/sv2v_out.v:12506.2-12514.5" */
wire [3:0] _118_;
/* src = "generated/sv2v_out.v:12703.49-12703.64" */
wire [31:0] _119_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12703.49-12703.64" */
wire [31:0] _120_;
/* src = "generated/sv2v_out.v:12469.10-12469.38" */
wire _121_;
/* src = "generated/sv2v_out.v:12477.46-12477.108" */
wire _122_;
/* src = "generated/sv2v_out.v:12499.45-12499.80" */
wire _123_;
/* src = "generated/sv2v_out.v:12501.55-12501.86" */
wire _124_;
/* src = "generated/sv2v_out.v:12505.24-12505.60" */
wire _125_;
/* src = "generated/sv2v_out.v:12505.23-12505.75" */
wire _126_;
/* src = "generated/sv2v_out.v:12505.90-12505.117" */
wire _127_;
/* src = "generated/sv2v_out.v:12516.52-12516.86" */
wire _128_;
/* src = "generated/sv2v_out.v:12620.10-12620.45" */
wire _129_;
/* src = "generated/sv2v_out.v:12643.11-12643.37" */
wire _130_;
/* src = "generated/sv2v_out.v:12762.26-12762.43" */
wire _131_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12762.26-12762.43" */
wire _132_;
wire [31:0] _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire [31:0] _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire [31:0] _148_;
wire [31:0] _149_;
wire [31:0] _150_;
wire [31:0] _151_;
wire [31:0] _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire [31:0] _160_;
wire [31:0] _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire [31:0] _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire [31:0] _207_;
wire [31:0] _208_;
wire _209_;
wire _210_;
wire _211_;
wire _212_;
wire [31:0] _213_;
wire [31:0] _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire [31:0] _236_;
wire [31:0] _237_;
wire [31:0] _238_;
wire [31:0] _239_;
wire [31:0] _240_;
wire [31:0] _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire [31:0] _254_;
wire [31:0] _255_;
wire [31:0] _256_;
wire [31:0] _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire [31:0] _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire [31:0] _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire _273_;
wire _274_;
wire _275_;
wire [31:0] _276_;
wire [31:0] _277_;
wire [31:0] _278_;
wire [3:0] _279_;
wire [3:0] _280_;
wire [3:0] _281_;
wire [3:0] _282_;
wire [3:0] _283_;
wire [3:0] _284_;
wire [3:0] _285_;
wire _286_;
wire _287_;
/* cellift = 32'd1 */
wire _288_;
wire _289_;
/* cellift = 32'd1 */
wire _290_;
wire [2:0] _291_;
wire [2:0] _292_;
wire _293_;
wire _294_;
wire _295_;
/* cellift = 32'd1 */
wire _296_;
wire _297_;
wire _298_;
wire [31:0] _299_;
/* cellift = 32'd1 */
wire [31:0] _300_;
wire _301_;
wire _302_;
wire _303_;
wire [6:0] _304_;
wire [1:0] _305_;
wire _306_;
/* src = "generated/sv2v_out.v:12502.30-12502.50" */
wire _307_;
/* src = "generated/sv2v_out.v:12502.72-12502.92" */
wire _308_;
/* src = "generated/sv2v_out.v:12622.9-12622.69" */
wire _309_;
/* src = "generated/sv2v_out.v:12624.10-12624.32" */
wire _310_;
/* src = "generated/sv2v_out.v:12624.9-12624.51" */
wire _311_;
/* src = "generated/sv2v_out.v:12641.10-12641.31" */
wire _312_;
/* src = "generated/sv2v_out.v:12675.9-12675.43" */
wire _313_;
/* src = "generated/sv2v_out.v:12747.38-12747.73" */
wire _314_;
/* src = "generated/sv2v_out.v:12747.9-12747.74" */
wire _315_;
/* src = "generated/sv2v_out.v:12469.25-12469.38" */
wire _316_;
/* src = "generated/sv2v_out.v:12624.10-12624.16" */
wire _317_;
/* src = "generated/sv2v_out.v:12624.20-12624.32" */
wire _318_;
/* src = "generated/sv2v_out.v:12624.37-12624.51" */
wire _319_;
/* src = "generated/sv2v_out.v:12641.20-12641.31" */
wire _320_;
/* src = "generated/sv2v_out.v:12675.30-12675.43" */
wire _321_;
/* src = "generated/sv2v_out.v:12747.36-12747.74" */
wire _322_;
/* src = "generated/sv2v_out.v:12589.12-12589.35" */
wire _323_;
/* src = "generated/sv2v_out.v:12589.11-12589.51" */
wire _324_;
/* src = "generated/sv2v_out.v:12589.10-12589.68" */
wire _325_;
/* src = "generated/sv2v_out.v:12589.9-12589.92" */
wire _326_;
/* src = "generated/sv2v_out.v:12614.9-12614.35" */
wire _327_;
/* src = "generated/sv2v_out.v:12622.10-12622.40" */
wire _328_;
/* src = "generated/sv2v_out.v:12622.46-12622.68" */
wire _329_;
/* src = "generated/sv2v_out.v:12688.10-12688.34" */
wire _330_;
/* src = "generated/sv2v_out.v:12688.9-12688.49" */
wire _331_;
/* src = "generated/sv2v_out.v:12400.44-12400.63" */
wire _332_;
/* src = "generated/sv2v_out.v:12647.15-12647.52" */
wire _333_;
/* src = "generated/sv2v_out.v:12463.39-12463.50" */
wire _334_;
/* src = "generated/sv2v_out.v:12477.80-12477.108" */
wire _335_;
/* src = "generated/sv2v_out.v:12505.40-12505.60" */
wire _336_;
/* src = "generated/sv2v_out.v:12615.36-12615.53" */
wire _337_;
/* src = "generated/sv2v_out.v:12762.35-12762.43" */
wire _338_;
/* src = "generated/sv2v_out.v:12763.31-12763.51" */
wire _339_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12763.31-12763.51" */
wire _340_;
/* src = "generated/sv2v_out.v:12401.24-12401.46" */
wire _341_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12401.24-12401.46" */
wire _342_;
/* src = "generated/sv2v_out.v:12401.23-12401.64" */
wire _343_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12401.23-12401.64" */
wire _344_;
/* src = "generated/sv2v_out.v:12401.22-12401.83" */
wire _345_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12401.22-12401.83" */
wire _346_;
/* src = "generated/sv2v_out.v:12405.35-12405.56" */
wire _347_;
/* src = "generated/sv2v_out.v:12405.34-12405.69" */
wire _348_;
/* src = "generated/sv2v_out.v:12430.29-12430.68" */
wire _349_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12430.29-12430.68" */
wire _350_;
/* src = "generated/sv2v_out.v:12500.36-12500.66" */
wire _351_;
/* src = "generated/sv2v_out.v:12505.80-12505.118" */
wire _352_;
/* src = "generated/sv2v_out.v:12611.10-12611.37" */
wire _353_;
/* src = "generated/sv2v_out.v:12711.12-12711.44" */
wire _354_;
wire _355_;
wire [31:0] _356_;
/* cellift = 32'd1 */
wire [31:0] _357_;
wire [31:0] _358_;
/* cellift = 32'd1 */
wire [31:0] _359_;
wire [31:0] _360_;
/* cellift = 32'd1 */
wire [31:0] _361_;
wire [31:0] _362_;
/* cellift = 32'd1 */
wire [31:0] _363_;
wire [31:0] _364_;
/* cellift = 32'd1 */
wire [31:0] _365_;
wire [6:0] _366_;
wire [6:0] _367_;
wire [6:0] _368_;
wire [6:0] _369_;
wire [6:0] _370_;
wire [3:0] _371_;
wire [3:0] _372_;
wire [3:0] _373_;
wire _374_;
wire _375_;
wire _376_;
wire _377_;
/* cellift = 32'd1 */
wire _378_;
wire _379_;
/* cellift = 32'd1 */
wire _380_;
wire _381_;
/* cellift = 32'd1 */
wire _382_;
wire _383_;
wire _384_;
wire _385_;
wire _386_;
wire _387_;
wire _388_;
wire _389_;
wire _390_;
wire _391_;
/* src = "generated/sv2v_out.v:12502.72-12502.117" */
wire _392_;
/* src = "generated/sv2v_out.v:12516.119-12516.149" */
wire [2:0] _393_;
/* src = "generated/sv2v_out.v:12516.97-12516.150" */
wire [2:0] _394_;
/* src = "generated/sv2v_out.v:12516.52-12516.151" */
wire [2:0] _395_;
/* src = "generated/sv2v_out.v:12642.22-12642.87" */
wire [6:0] _396_;
/* src = "generated/sv2v_out.v:12691.22-12691.48" */
wire [1:0] _397_;
/* src = "generated/sv2v_out.v:12703.23-12703.74" */
wire [31:0] _398_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12703.23-12703.74" */
wire [31:0] _399_;
/* src = "generated/sv2v_out.v:12707.23-12707.99" */
wire [31:0] _400_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12707.23-12707.99" */
wire [31:0] _401_;
/* src = "generated/sv2v_out.v:12709.39-12709.119" */
wire [6:0] _402_;
/* src = "generated/sv2v_out.v:12309.13-12309.29" */
input branch_not_set_i;
wire branch_not_set_i;
/* cellift = 32'd1 */
input branch_not_set_i_t0;
wire branch_not_set_i_t0;
/* src = "generated/sv2v_out.v:12308.13-12308.25" */
input branch_set_i;
wire branch_set_i;
/* cellift = 32'd1 */
input branch_set_i_t0;
wire branch_set_i_t0;
/* src = "generated/sv2v_out.v:12274.13-12274.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:12294.13-12294.29" */
output controller_run_o;
wire controller_run_o;
/* cellift = 32'd1 */
output controller_run_o_t0;
wire controller_run_o_t0;
/* src = "generated/sv2v_out.v:12311.13-12311.30" */
input csr_mstatus_mie_i;
wire csr_mstatus_mie_i;
/* cellift = 32'd1 */
input csr_mstatus_mie_i_t0;
wire csr_mstatus_mie_i_t0;
/* src = "generated/sv2v_out.v:12331.20-12331.31" */
output [31:0] csr_mtval_o;
wire [31:0] csr_mtval_o;
/* cellift = 32'd1 */
output [31:0] csr_mtval_o_t0;
wire [31:0] csr_mtval_o_t0;
/* src = "generated/sv2v_out.v:12389.7-12389.21" */
wire csr_pipe_flush;
/* src = "generated/sv2v_out.v:12283.13-12283.29" */
input csr_pipe_flush_i;
wire csr_pipe_flush_i;
/* cellift = 32'd1 */
input csr_pipe_flush_i_t0;
wire csr_pipe_flush_i_t0;
/* src = "generated/sv2v_out.v:12329.13-12329.34" */
output csr_restore_dret_id_o;
wire csr_restore_dret_id_o;
/* cellift = 32'd1 */
output csr_restore_dret_id_o_t0;
wire csr_restore_dret_id_o_t0;
/* src = "generated/sv2v_out.v:12328.13-12328.34" */
output csr_restore_mret_id_o;
wire csr_restore_mret_id_o;
/* cellift = 32'd1 */
output csr_restore_mret_id_o_t0;
wire csr_restore_mret_id_o_t0;
/* src = "generated/sv2v_out.v:12330.13-12330.29" */
output csr_save_cause_o;
wire csr_save_cause_o;
/* cellift = 32'd1 */
output csr_save_cause_o_t0;
wire csr_save_cause_o_t0;
/* src = "generated/sv2v_out.v:12326.13-12326.26" */
output csr_save_id_o;
wire csr_save_id_o;
/* cellift = 32'd1 */
output csr_save_id_o_t0;
wire csr_save_id_o_t0;
/* src = "generated/sv2v_out.v:12325.13-12325.26" */
output csr_save_if_o;
wire csr_save_if_o;
/* cellift = 32'd1 */
output csr_save_if_o_t0;
wire csr_save_if_o_t0;
/* src = "generated/sv2v_out.v:12327.13-12327.26" */
output csr_save_wb_o;
wire csr_save_wb_o;
/* cellift = 32'd1 */
output csr_save_wb_o_t0;
wire csr_save_wb_o_t0;
/* src = "generated/sv2v_out.v:12276.13-12276.24" */
output ctrl_busy_o;
wire ctrl_busy_o;
/* cellift = 32'd1 */
output ctrl_busy_o_t0;
wire ctrl_busy_o_t0;
/* src = "generated/sv2v_out.v:12339.12-12339.23" */
reg [3:0] ctrl_fsm_cs;
/* src = "generated/sv2v_out.v:12340.12-12340.23" */
wire [3:0] ctrl_fsm_ns;
/* src = "generated/sv2v_out.v:12345.13-12345.26" */
wire [2:0] debug_cause_d;
/* src = "generated/sv2v_out.v:12317.20-12317.33" */
output [2:0] debug_cause_o;
reg [2:0] debug_cause_o;
/* cellift = 32'd1 */
output [2:0] debug_cause_o_t0;
wire [2:0] debug_cause_o_t0;
/* src = "generated/sv2v_out.v:12318.13-12318.29" */
output debug_csr_save_o;
wire debug_csr_save_o;
/* cellift = 32'd1 */
output debug_csr_save_o_t0;
wire debug_csr_save_o_t0;
/* src = "generated/sv2v_out.v:12322.13-12322.28" */
input debug_ebreakm_i;
wire debug_ebreakm_i;
/* cellift = 32'd1 */
input debug_ebreakm_i_t0;
wire debug_ebreakm_i_t0;
/* src = "generated/sv2v_out.v:12323.13-12323.28" */
input debug_ebreaku_i;
wire debug_ebreaku_i;
/* cellift = 32'd1 */
input debug_ebreaku_i_t0;
wire debug_ebreaku_i_t0;
/* src = "generated/sv2v_out.v:12344.6-12344.18" */
wire debug_mode_d;
/* src = "generated/sv2v_out.v:12320.13-12320.34" */
output debug_mode_entering_o;
wire debug_mode_entering_o;
/* cellift = 32'd1 */
output debug_mode_entering_o_t0;
wire debug_mode_entering_o_t0;
/* src = "generated/sv2v_out.v:12319.14-12319.26" */
output debug_mode_o;
reg debug_mode_o;
/* cellift = 32'd1 */
output debug_mode_o_t0;
reg debug_mode_o_t0;
/* src = "generated/sv2v_out.v:12316.13-12316.24" */
input debug_req_i;
wire debug_req_i;
/* cellift = 32'd1 */
input debug_req_i_t0;
wire debug_req_i_t0;
/* src = "generated/sv2v_out.v:12321.13-12321.32" */
input debug_single_step_i;
wire debug_single_step_i;
/* cellift = 32'd1 */
input debug_single_step_i_t0;
wire debug_single_step_i_t0;
/* src = "generated/sv2v_out.v:12369.7-12369.23" */
wire do_single_step_d;
/* src = "generated/sv2v_out.v:12370.6-12370.22" */
reg do_single_step_q;
/* src = "generated/sv2v_out.v:12386.7-12386.16" */
wire dret_insn;
/* src = "generated/sv2v_out.v:12280.13-12280.24" */
input dret_insn_i;
wire dret_insn_i;
/* cellift = 32'd1 */
input dret_insn_i_t0;
wire dret_insn_i_t0;
/* src = "generated/sv2v_out.v:12374.7-12374.24" */
wire ebreak_into_debug;
/* src = "generated/sv2v_out.v:12388.7-12388.16" */
wire ebrk_insn;
/* src = "generated/sv2v_out.v:12282.13-12282.24" */
input ebrk_insn_i;
wire ebrk_insn_i;
/* cellift = 32'd1 */
input ebrk_insn_i_t0;
wire ebrk_insn_i_t0;
/* src = "generated/sv2v_out.v:12358.6-12358.20" */
wire ebrk_insn_prio;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12388.7-12388.16" */
wire ebrk_insn_t0;
/* src = "generated/sv2v_out.v:12384.7-12384.17" */
wire ecall_insn;
/* src = "generated/sv2v_out.v:12278.13-12278.25" */
input ecall_insn_i;
wire ecall_insn_i;
/* cellift = 32'd1 */
input ecall_insn_i_t0;
wire ecall_insn_i_t0;
/* src = "generated/sv2v_out.v:12357.6-12357.21" */
wire ecall_insn_prio;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12384.7-12384.17" */
wire ecall_insn_t0;
/* src = "generated/sv2v_out.v:12373.7-12373.23" */
wire enter_debug_mode;
/* src = "generated/sv2v_out.v:12371.7-12371.30" */
wire enter_debug_mode_prio_d;
/* src = "generated/sv2v_out.v:12372.6-12372.29" */
reg enter_debug_mode_prio_q;
/* src = "generated/sv2v_out.v:12301.19-12301.30" */
output [6:0] exc_cause_o;
wire [6:0] exc_cause_o;
/* cellift = 32'd1 */
output [6:0] exc_cause_o_t0;
wire [6:0] exc_cause_o_t0;
/* src = "generated/sv2v_out.v:12300.19-12300.31" */
output [1:0] exc_pc_mux_o;
wire [1:0] exc_pc_mux_o;
/* cellift = 32'd1 */
output [1:0] exc_pc_mux_o_t0;
wire [1:0] exc_pc_mux_o_t0;
/* src = "generated/sv2v_out.v:12352.7-12352.16" */
wire exc_req_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12352.7-12352.16" */
wire exc_req_d_t0;
/* src = "generated/sv2v_out.v:12365.7-12365.18" */
wire exc_req_lsu;
/* src = "generated/sv2v_out.v:12351.6-12351.15" */
reg exc_req_q;
/* src = "generated/sv2v_out.v:12335.14-12335.24" */
output flush_id_o;
wire flush_id_o;
/* cellift = 32'd1 */
output flush_id_o_t0;
wire flush_id_o_t0;
/* src = "generated/sv2v_out.v:12462.9-12462.21" */
wire \g_intg_irq_int.entering_nmi ;
/* src = "generated/sv2v_out.v:12458.15-12458.39" */
reg [31:0] \g_intg_irq_int.mem_resp_intg_err_addr_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12458.15-12458.39" */
reg [31:0] \g_intg_irq_int.mem_resp_intg_err_addr_q_t0 ;
/* src = "generated/sv2v_out.v:12461.8-12461.35" */
wire \g_intg_irq_int.mem_resp_intg_err_irq_clear ;
/* src = "generated/sv2v_out.v:12457.9-12457.40" */
wire \g_intg_irq_int.mem_resp_intg_err_irq_pending_d ;
/* src = "generated/sv2v_out.v:12456.8-12456.39" */
reg \g_intg_irq_int.mem_resp_intg_err_irq_pending_q ;
/* src = "generated/sv2v_out.v:12460.8-12460.33" */
wire \g_intg_irq_int.mem_resp_intg_err_irq_set ;
/* src = "generated/sv2v_out.v:12362.6-12362.13" */
wire halt_if;
/* src = "generated/sv2v_out.v:12376.7-12376.17" */
wire handle_irq;
/* src = "generated/sv2v_out.v:12307.14-12307.28" */
output id_exception_o;
wire id_exception_o;
/* cellift = 32'd1 */
output id_exception_o_t0;
wire id_exception_o_t0;
/* src = "generated/sv2v_out.v:12293.14-12293.27" */
output id_in_ready_o;
wire id_in_ready_o;
/* cellift = 32'd1 */
output id_in_ready_o_t0;
wire id_in_ready_o_t0;
/* src = "generated/sv2v_out.v:12377.7-12377.20" */
wire id_wb_pending;
/* src = "generated/sv2v_out.v:12354.7-12354.21" */
wire illegal_insn_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12354.7-12354.21" */
wire illegal_insn_d_t0;
/* src = "generated/sv2v_out.v:12277.13-12277.27" */
input illegal_insn_i;
wire illegal_insn_i;
/* cellift = 32'd1 */
input illegal_insn_i_t0;
wire illegal_insn_i_t0;
/* src = "generated/sv2v_out.v:12356.6-12356.23" */
wire illegal_insn_prio;
/* src = "generated/sv2v_out.v:12353.6-12353.20" */
reg illegal_insn_q;
/* src = "generated/sv2v_out.v:12288.13-12288.29" */
input instr_bp_taken_i;
wire instr_bp_taken_i;
/* cellift = 32'd1 */
input instr_bp_taken_i_t0;
wire instr_bp_taken_i_t0;
/* src = "generated/sv2v_out.v:12286.20-12286.38" */
input [15:0] instr_compressed_i;
wire [15:0] instr_compressed_i;
/* cellift = 32'd1 */
input [15:0] instr_compressed_i_t0;
wire [15:0] instr_compressed_i_t0;
/* src = "generated/sv2v_out.v:12295.13-12295.25" */
input instr_exec_i;
wire instr_exec_i;
/* cellift = 32'd1 */
input instr_exec_i_t0;
wire instr_exec_i_t0;
/* src = "generated/sv2v_out.v:12390.7-12390.22" */
wire instr_fetch_err;
/* src = "generated/sv2v_out.v:12289.13-12289.30" */
input instr_fetch_err_i;
wire instr_fetch_err_i;
/* cellift = 32'd1 */
input instr_fetch_err_i_t0;
wire instr_fetch_err_i_t0;
/* src = "generated/sv2v_out.v:12290.13-12290.36" */
input instr_fetch_err_plus2_i;
wire instr_fetch_err_plus2_i;
/* cellift = 32'd1 */
input instr_fetch_err_plus2_i_t0;
wire instr_fetch_err_plus2_i_t0;
/* src = "generated/sv2v_out.v:12355.6-12355.26" */
wire instr_fetch_err_prio;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12390.7-12390.22" */
wire instr_fetch_err_t0;
/* src = "generated/sv2v_out.v:12285.20-12285.27" */
input [31:0] instr_i;
wire [31:0] instr_i;
/* cellift = 32'd1 */
input [31:0] instr_i_t0;
wire [31:0] instr_i_t0;
/* src = "generated/sv2v_out.v:12287.13-12287.34" */
input instr_is_compressed_i;
wire instr_is_compressed_i;
/* cellift = 32'd1 */
input instr_is_compressed_i_t0;
wire instr_is_compressed_i_t0;
/* src = "generated/sv2v_out.v:12296.13-12296.24" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:12292.14-12292.33" */
output instr_valid_clear_o;
wire instr_valid_clear_o;
/* cellift = 32'd1 */
output instr_valid_clear_o_t0;
wire instr_valid_clear_o_t0;
/* src = "generated/sv2v_out.v:12284.13-12284.26" */
input instr_valid_i;
wire instr_valid_i;
/* cellift = 32'd1 */
input instr_valid_i_t0;
wire instr_valid_i_t0;
/* src = "generated/sv2v_out.v:12375.7-12375.18" */
wire irq_enabled;
/* src = "generated/sv2v_out.v:12378.7-12378.13" */
wire irq_nm;
/* src = "generated/sv2v_out.v:12314.13-12314.25" */
input irq_nm_ext_i;
wire irq_nm_ext_i;
/* cellift = 32'd1 */
input irq_nm_ext_i_t0;
wire irq_nm_ext_i_t0;
/* src = "generated/sv2v_out.v:12379.7-12379.17" */
wire irq_nm_int;
/* src = "generated/sv2v_out.v:12312.13-12312.26" */
input irq_pending_i;
wire irq_pending_i;
/* cellift = 32'd1 */
input irq_pending_i_t0;
wire irq_pending_i_t0;
/* src = "generated/sv2v_out.v:12313.20-12313.26" */
input [17:0] irqs_i;
wire [17:0] irqs_i;
/* cellift = 32'd1 */
input [17:0] irqs_i_t0;
wire [17:0] irqs_i_t0;
/* src = "generated/sv2v_out.v:12310.13-12310.23" */
input jump_set_i;
wire jump_set_i;
/* cellift = 32'd1 */
input jump_set_i_t0;
wire jump_set_i_t0;
/* src = "generated/sv2v_out.v:12303.13-12303.23" */
input load_err_i;
wire load_err_i;
/* cellift = 32'd1 */
input load_err_i_t0;
wire load_err_i_t0;
/* src = "generated/sv2v_out.v:12360.6-12360.19" */
wire load_err_prio;
/* src = "generated/sv2v_out.v:12347.6-12347.16" */
reg load_err_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12347.6-12347.16" */
reg load_err_q_t0;
/* src = "generated/sv2v_out.v:12302.20-12302.35" */
input [31:0] lsu_addr_last_i;
wire [31:0] lsu_addr_last_i;
/* cellift = 32'd1 */
input [31:0] lsu_addr_last_i_t0;
wire [31:0] lsu_addr_last_i_t0;
/* src = "generated/sv2v_out.v:12305.13-12305.32" */
input mem_resp_intg_err_i;
wire mem_resp_intg_err_i;
/* cellift = 32'd1 */
input mem_resp_intg_err_i_t0;
wire mem_resp_intg_err_i_t0;
/* src = "generated/sv2v_out.v:12382.12-12382.19" */
wire [3:0] mfip_id;
/* src = "generated/sv2v_out.v:12385.7-12385.16" */
wire mret_insn;
/* src = "generated/sv2v_out.v:12279.13-12279.24" */
input mret_insn_i;
wire mret_insn_i;
/* cellift = 32'd1 */
input mret_insn_i_t0;
wire mret_insn_i_t0;
/* src = "generated/sv2v_out.v:12342.6-12342.16" */
wire nmi_mode_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12342.6-12342.16" */
wire nmi_mode_d_t0;
/* src = "generated/sv2v_out.v:12315.14-12315.24" */
output nmi_mode_o;
reg nmi_mode_o;
/* cellift = 32'd1 */
output nmi_mode_o_t0;
reg nmi_mode_o_t0;
/* src = "generated/sv2v_out.v:12299.13-12299.35" */
output nt_branch_mispredict_o;
wire nt_branch_mispredict_o;
/* cellift = 32'd1 */
output nt_branch_mispredict_o_t0;
wire nt_branch_mispredict_o_t0;
/* src = "generated/sv2v_out.v:12291.20-12291.27" */
input [31:0] pc_id_i;
wire [31:0] pc_id_i;
/* cellift = 32'd1 */
input [31:0] pc_id_i_t0;
wire [31:0] pc_id_i_t0;
/* src = "generated/sv2v_out.v:12298.19-12298.27" */
output [2:0] pc_mux_o;
wire [2:0] pc_mux_o;
/* cellift = 32'd1 */
output [2:0] pc_mux_o_t0;
wire [2:0] pc_mux_o_t0;
/* src = "generated/sv2v_out.v:12297.13-12297.21" */
output pc_set_o;
wire pc_set_o;
/* cellift = 32'd1 */
output pc_set_o_t0;
wire pc_set_o_t0;
/* src = "generated/sv2v_out.v:12337.13-12337.24" */
output perf_jump_o;
wire perf_jump_o;
/* cellift = 32'd1 */
output perf_jump_o_t0;
wire perf_jump_o_t0;
/* src = "generated/sv2v_out.v:12338.13-12338.27" */
output perf_tbranch_o;
wire perf_tbranch_o;
/* cellift = 32'd1 */
output perf_tbranch_o_t0;
wire perf_tbranch_o_t0;
/* src = "generated/sv2v_out.v:12332.19-12332.30" */
input [1:0] priv_mode_i;
wire [1:0] priv_mode_i;
/* cellift = 32'd1 */
input [1:0] priv_mode_i_t0;
wire [1:0] priv_mode_i_t0;
/* src = "generated/sv2v_out.v:12336.13-12336.23" */
input ready_wb_i;
wire ready_wb_i;
/* cellift = 32'd1 */
input ready_wb_i_t0;
wire ready_wb_i_t0;
/* src = "generated/sv2v_out.v:12363.6-12363.15" */
wire retain_id;
/* src = "generated/sv2v_out.v:12275.13-12275.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:12366.7-12366.18" */
wire special_req;
/* src = "generated/sv2v_out.v:12368.7-12368.29" */
wire special_req_flush_only;
/* src = "generated/sv2v_out.v:12367.7-12367.28" */
wire special_req_pc_change;
/* src = "generated/sv2v_out.v:12361.7-12361.12" */
wire stall;
/* src = "generated/sv2v_out.v:12333.13-12333.23" */
input stall_id_i;
wire stall_id_i;
/* cellift = 32'd1 */
input stall_id_i_t0;
wire stall_id_i_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12361.7-12361.12" */
wire stall_t0;
/* src = "generated/sv2v_out.v:12334.13-12334.23" */
input stall_wb_i;
wire stall_wb_i;
/* cellift = 32'd1 */
input stall_wb_i_t0;
wire stall_wb_i_t0;
/* src = "generated/sv2v_out.v:12304.13-12304.24" */
input store_err_i;
wire store_err_i;
/* cellift = 32'd1 */
input store_err_i_t0;
wire store_err_i_t0;
/* src = "generated/sv2v_out.v:12359.6-12359.20" */
wire store_err_prio;
/* src = "generated/sv2v_out.v:12349.6-12349.17" */
reg store_err_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12349.6-12349.17" */
reg store_err_q_t0;
/* src = "generated/sv2v_out.v:12324.13-12324.28" */
input trigger_match_i;
wire trigger_match_i;
/* cellift = 32'd1 */
input trigger_match_i_t0;
wire trigger_match_i_t0;
/* src = "generated/sv2v_out.v:12306.14-12306.28" */
output wb_exception_o;
wire wb_exception_o;
/* cellift = 32'd1 */
output wb_exception_o_t0;
wire wb_exception_o_t0;
/* src = "generated/sv2v_out.v:12387.7-12387.15" */
wire wfi_insn;
/* src = "generated/sv2v_out.v:12281.13-12281.23" */
input wfi_insn_i;
wire wfi_insn_i;
/* cellift = 32'd1 */
input wfi_insn_i_t0;
wire wfi_insn_i_t0;
assign _119_ = pc_id_i + /* src = "generated/sv2v_out.v:12703.49-12703.64" */ 32'd2;
assign ecall_insn = ecall_insn_i & /* src = "generated/sv2v_out.v:12393.22-12393.50" */ instr_valid_i;
assign mret_insn = mret_insn_i & /* src = "generated/sv2v_out.v:12394.21-12394.48" */ instr_valid_i;
assign dret_insn = dret_insn_i & /* src = "generated/sv2v_out.v:12395.21-12395.48" */ instr_valid_i;
assign wfi_insn = wfi_insn_i & /* src = "generated/sv2v_out.v:12396.20-12396.46" */ instr_valid_i;
assign ebrk_insn = ebrk_insn_i & /* src = "generated/sv2v_out.v:12397.21-12397.48" */ instr_valid_i;
assign csr_pipe_flush = csr_pipe_flush_i & /* src = "generated/sv2v_out.v:12398.26-12398.58" */ instr_valid_i;
assign instr_fetch_err = instr_fetch_err_i & /* src = "generated/sv2v_out.v:12399.27-12399.60" */ instr_valid_i;
assign illegal_insn_d = illegal_insn_i & /* src = "generated/sv2v_out.v:12400.26-12400.64" */ _332_;
assign exc_req_d = _345_ & /* src = "generated/sv2v_out.v:12401.21-12401.108" */ _332_;
assign id_exception_o = exc_req_d & /* src = "generated/sv2v_out.v:12403.26-12403.53" */ _173_;
assign \g_intg_irq_int.entering_nmi  = nmi_mode_d & /* src = "generated/sv2v_out.v:12463.26-12463.50" */ _334_;
assign _121_ = \g_intg_irq_int.entering_nmi  & /* src = "generated/sv2v_out.v:12469.10-12469.38" */ _316_;
assign _122_ = \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  & /* src = "generated/sv2v_out.v:12477.46-12477.108" */ _335_;
assign _123_ = _167_ & /* src = "generated/sv2v_out.v:12499.45-12499.80" */ debug_single_step_i;
assign enter_debug_mode_prio_d = _351_ & /* src = "generated/sv2v_out.v:12500.35-12500.83" */ _167_;
assign _124_ = trigger_match_i & /* src = "generated/sv2v_out.v:12501.55-12501.86" */ _167_;
assign _125_ = _167_ & /* src = "generated/sv2v_out.v:12505.24-12505.60" */ _336_;
assign _126_ = _125_ & /* src = "generated/sv2v_out.v:12505.23-12505.75" */ _334_;
assign _127_ = irq_pending_i & /* src = "generated/sv2v_out.v:12505.90-12505.117" */ irq_enabled;
assign handle_irq = _126_ & /* src = "generated/sv2v_out.v:12505.22-12505.119" */ _352_;
assign _128_ = ebrk_insn_prio & /* src = "generated/sv2v_out.v:12516.52-12516.86" */ ebreak_into_debug;
assign _129_ = instr_bp_taken_i & /* src = "generated/sv2v_out.v:12620.10-12620.45" */ branch_not_set_i;
assign _130_ = irq_nm_int & /* src = "generated/sv2v_out.v:12643.11-12643.37" */ _316_;
assign _131_ = _169_ & /* src = "generated/sv2v_out.v:12762.26-12762.43" */ _338_;
assign id_in_ready_o = _131_ & /* src = "generated/sv2v_out.v:12762.25-12762.57" */ _175_;
assign _133_ = ~ pc_id_i_t0;
assign _193_ = pc_id_i & _133_;
assign _277_ = _193_ + 32'd2;
assign _263_ = pc_id_i | pc_id_i_t0;
assign _278_ = _263_ + 32'd2;
assign _276_ = _277_ ^ _278_;
assign _120_ = _276_ | pc_id_i_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME nmi_mode_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) nmi_mode_o_t0 <= 1'h0;
else nmi_mode_o_t0 <= nmi_mode_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME load_err_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) load_err_q_t0 <= 1'h0;
else load_err_q_t0 <= load_err_i_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME store_err_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) store_err_q_t0 <= 1'h0;
else store_err_q_t0 <= store_err_i_t0;
assign _134_ = ~ _185_;
assign _135_ = ~ _187_;
assign _207_ = { _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_, _187_ } & lsu_addr_last_i_t0;
assign _206_ = _134_ & debug_mode_o_t0;
assign _208_ = { _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_, _135_ } & \g_intg_irq_int.mem_resp_intg_err_addr_q_t0 ;
assign _268_ = _207_ | _208_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME debug_mode_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) debug_mode_o_t0 <= 1'h0;
else debug_mode_o_t0 <= _206_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_intg_irq_int.mem_resp_intg_err_addr_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_intg_irq_int.mem_resp_intg_err_addr_q_t0  <= 32'd0;
else \g_intg_irq_int.mem_resp_intg_err_addr_q_t0  <= _268_;
assign _194_ = ecall_insn_i_t0 & instr_valid_i;
assign _197_ = ebrk_insn_i_t0 & instr_valid_i;
assign _200_ = instr_fetch_err_i_t0 & instr_valid_i;
assign illegal_insn_d_t0 = illegal_insn_i_t0 & _332_;
assign exc_req_d_t0 = _346_ & _332_;
assign _203_ = exc_req_d_t0 & _173_;
assign _132_ = stall_t0 & _338_;
assign id_in_ready_o_t0 = _132_ & _175_;
assign _195_ = instr_valid_i_t0 & ecall_insn_i;
assign _198_ = instr_valid_i_t0 & ebrk_insn_i;
assign _201_ = instr_valid_i_t0 & instr_fetch_err_i;
assign _204_ = wb_exception_o_t0 & exc_req_d;
assign _196_ = ecall_insn_i_t0 & instr_valid_i_t0;
assign _199_ = ebrk_insn_i_t0 & instr_valid_i_t0;
assign _202_ = instr_fetch_err_i_t0 & instr_valid_i_t0;
assign _205_ = exc_req_d_t0 & wb_exception_o_t0;
assign _264_ = _194_ | _195_;
assign _265_ = _197_ | _198_;
assign _266_ = _200_ | _201_;
assign _267_ = _203_ | _204_;
assign ecall_insn_t0 = _264_ | _196_;
assign ebrk_insn_t0 = _265_ | _199_;
assign instr_fetch_err_t0 = _266_ | _202_;
assign id_exception_o_t0 = _267_ | _205_;
/* src = "generated/sv2v_out.v:12764.2-12787.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME debug_mode_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) debug_mode_o <= 1'h0;
else if (_185_) debug_mode_o <= debug_mode_d;
/* src = "generated/sv2v_out.v:12764.2-12787.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME ctrl_fsm_cs */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) ctrl_fsm_cs <= 4'h0;
else if (_186_) ctrl_fsm_cs <= ctrl_fsm_ns;
/* src = "generated/sv2v_out.v:12478.4-12486.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_intg_irq_int.mem_resp_intg_err_addr_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_intg_irq_int.mem_resp_intg_err_addr_q  <= 32'd0;
else if (_187_) \g_intg_irq_int.mem_resp_intg_err_addr_q  <= lsu_addr_last_i;
assign _138_ = ~ _260_;
assign _136_ = ~ _355_;
assign _137_ = ~ _384_;
assign _139_ = ~ { _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_ };
assign _140_ = ~ \g_intg_irq_int.mem_resp_intg_err_irq_pending_q ;
assign _141_ = ~ ebrk_insn;
assign _142_ = ~ ecall_insn;
assign _143_ = ~ instr_fetch_err;
assign _144_ = ~ load_err_q;
assign _145_ = ~ store_err_q;
assign _146_ = ~ mret_insn;
assign _147_ = ~ _354_;
assign _148_ = ~ { store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio };
assign _149_ = ~ { ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio };
assign _150_ = ~ { ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio };
assign _151_ = ~ { illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio };
assign _152_ = ~ { instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio };
assign _153_ = ~ ebrk_insn_prio;
assign _155_ = ~ illegal_insn_prio;
assign _154_ = ~ ecall_insn_prio;
assign _156_ = ~ instr_fetch_err_prio;
assign _157_ = ~ _331_;
assign _158_ = ~ _312_;
assign _159_ = ~ handle_irq;
assign _160_ = ~ { instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i };
assign _161_ = ~ { instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i };
assign _290_ = _137_ & _288_;
assign pc_set_o_t0 = _138_ & _290_;
assign _209_ = _137_ & nmi_mode_o_t0;
assign _211_ = _136_ & _296_;
assign _213_ = _139_ & _300_;
assign _098_ = _146_ & nmi_mode_o_t0;
assign _102_ = _147_ & _055_;
assign _236_ = _148_ & _357_;
assign _361_ = _149_ & _359_;
assign _363_ = _150_ & _361_;
assign _238_ = _151_ & _363_;
assign _240_ = _152_ & _365_;
assign _242_ = _153_ & _055_;
assign _244_ = _154_ & _378_;
assign _246_ = _155_ & _380_;
assign _248_ = _156_ & _382_;
assign _250_ = _157_ & _098_;
assign _067_ = _158_ & nmi_mode_o_t0;
assign _252_ = _159_ & nmi_mode_o_t0;
assign _254_ = _160_ & pc_id_i_t0;
assign _256_ = _161_ & instr_i_t0;
assign _288_ = _385_ & _042_;
assign _210_ = _384_ & _038_;
assign _212_ = _355_ & _084_;
assign _300_ = { _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_, _384_ } & _016_;
assign _214_ = { _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_, _355_ } & _088_;
assign csr_save_id_o_t0 = _355_ & _053_;
assign _357_ = { load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio } & lsu_addr_last_i_t0;
assign _237_ = { store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio } & lsu_addr_last_i_t0;
assign _239_ = { illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio } & _401_;
assign _241_ = { instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio } & _399_;
assign _243_ = ebrk_insn_prio & _102_;
assign _245_ = ecall_insn_prio & _055_;
assign _247_ = illegal_insn_prio & _055_;
assign _249_ = instr_fetch_err_prio & _055_;
assign _088_ = { _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_ } & _100_;
assign _053_ = _331_ & _090_;
assign _022_ = _331_ & _055_;
assign _251_ = _331_ & nmi_mode_o_t0;
assign _070_ = { _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_, _130_ } & \g_intg_irq_int.mem_resp_intg_err_addr_q_t0 ;
assign _049_ = { _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_, _312_ } & _070_;
assign _253_ = handle_irq & _067_;
assign _016_ = { handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq } & _049_;
assign _044_ = _327_ & jump_set_i_t0;
assign _046_ = _327_ & branch_set_i_t0;
assign _042_ = _327_ & instr_bp_taken_i_t0;
assign perf_tbranch_o_t0 = _385_ & _046_;
assign perf_jump_o_t0 = _385_ & _044_;
assign csr_save_wb_o_t0 = _355_ & _022_;
assign _255_ = { instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i } & _120_;
assign _257_ = { instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i } & { 16'h0000, instr_compressed_i_t0 };
assign _296_ = _209_ | _210_;
assign nmi_mode_d_t0 = _211_ | _212_;
assign csr_mtval_o_t0 = _213_ | _214_;
assign _359_ = _236_ | _237_;
assign _365_ = _238_ | _239_;
assign _100_ = _240_ | _241_;
assign _378_ = _242_ | _243_;
assign _380_ = _244_ | _245_;
assign _382_ = _246_ | _247_;
assign _090_ = _248_ | _249_;
assign _084_ = _250_ | _251_;
assign _038_ = _252_ | _253_;
assign _399_ = _254_ | _255_;
assign _401_ = _256_ | _257_;
assign _179_ = { _355_, _331_, dret_insn, mret_insn } != 4'h8;
assign _180_ = { _355_, _331_, mret_insn } != 3'h5;
assign _181_ = { _355_, _331_ } != 2'h3;
assign _182_ = | { _177_, _355_ };
assign _183_ = { _386_, id_in_ready_o, handle_irq, enter_debug_mode } != 4'h8;
assign _184_ = { _387_, _326_ } != 2'h2;
assign _185_ = & { _182_, _180_, _179_, _181_ };
assign _186_ = & { _183_, _184_ };
assign _187_ = & { _140_, mem_resp_intg_err_i };
assign _188_ = | { _389_, _387_, _355_ };
assign _190_ = | { _391_, _390_, _388_, _383_ };
assign _191_ = | { _389_, _388_, _387_, _383_ };
assign _189_ = | { _388_, _384_, _383_ };
assign _192_ = | { _390_, _388_, _386_, _385_, _384_, _383_, _355_ };
assign _162_ = ~ _341_;
assign _163_ = ~ _343_;
assign _164_ = ~ store_err_i;
assign _073_ = ~ _054_;
assign _165_ = ~ _349_;
assign _166_ = ~ ready_wb_i;
assign _167_ = ~ debug_mode_o;
assign _168_ = ~ stall_id_i;
assign _169_ = ~ stall;
assign _171_ = ~ illegal_insn_d;
assign _172_ = ~ load_err_i;
assign _173_ = ~ wb_exception_o;
assign _174_ = ~ stall_wb_i;
assign _175_ = ~ retain_id;
assign _176_ = ~ flush_id_o;
assign _215_ = ecall_insn_t0 & _141_;
assign _218_ = _342_ & _171_;
assign _221_ = _344_ & _143_;
assign _224_ = load_err_q_t0 & _145_;
assign _227_ = _055_ & _172_;
assign _230_ = _350_ & _164_;
assign _233_ = stall_id_i_t0 & _174_;
assign _340_ = stall_t0 & _175_;
assign instr_valid_clear_o_t0 = _340_ & _176_;
assign _216_ = ebrk_insn_t0 & _142_;
assign _219_ = illegal_insn_d_t0 & _162_;
assign _222_ = instr_fetch_err_t0 & _163_;
assign _225_ = store_err_q_t0 & _144_;
assign _228_ = load_err_i_t0 & _073_;
assign _231_ = store_err_i_t0 & _165_;
assign _234_ = stall_wb_i_t0 & _168_;
assign _217_ = ecall_insn_t0 & ebrk_insn_t0;
assign _220_ = _342_ & illegal_insn_d_t0;
assign _223_ = _344_ & instr_fetch_err_t0;
assign _226_ = load_err_q_t0 & store_err_q_t0;
assign _229_ = _055_ & load_err_i_t0;
assign _232_ = _350_ & store_err_i_t0;
assign _235_ = stall_id_i_t0 & stall_wb_i_t0;
assign _269_ = _215_ | _216_;
assign _270_ = _218_ | _219_;
assign _271_ = _221_ | _222_;
assign _272_ = _224_ | _225_;
assign _273_ = _227_ | _228_;
assign _274_ = _230_ | _231_;
assign _275_ = _233_ | _234_;
assign _342_ = _269_ | _217_;
assign _344_ = _270_ | _220_;
assign _346_ = _271_ | _223_;
assign _055_ = _272_ | _226_;
assign _350_ = _273_ | _229_;
assign wb_exception_o_t0 = _274_ | _232_;
assign stall_t0 = _275_ | _235_;
assign _177_ = | { _388_, _383_ };
assign _259_ = _389_ | _387_;
assign _260_ = _190_ | _355_;
assign _258_ = _189_ | _355_;
assign _261_ = _385_ | _188_;
assign _262_ = _383_ | _355_;
assign _178_ = | { _386_, _385_, _258_ };
assign _279_ = _355_ ? _012_ : 4'h5;
assign _280_ = _385_ ? _113_ : _091_;
assign _281_ = _258_ ? _279_ : _280_;
assign _282_ = _387_ ? _024_ : 4'h3;
assign _283_ = _391_ ? 4'h1 : 4'h0;
assign _284_ = _390_ ? 4'h4 : _283_;
assign _285_ = _259_ ? _282_ : _284_;
assign ctrl_fsm_ns = _178_ ? _281_ : _285_;
assign _286_ = _355_ ? _086_ : 1'h1;
assign _287_ = _385_ ? _041_ : 1'h0;
assign _289_ = _384_ ? _019_ : _287_;
assign pc_set_o = _260_ ? _286_ : _289_;
assign _291_ = _355_ ? _040_ : 3'h2;
assign _292_ = _385_ ? 3'h1 : 3'h0;
assign pc_mux_o = _258_ ? _291_ : _292_;
assign _293_ = _188_ ? 1'h1 : _095_;
assign _294_ = _386_ ? _062_ : 1'h0;
assign _013_ = _261_ ? _293_ : _294_;
assign debug_mode_d = _355_ ? _025_ : 1'h1;
assign _295_ = _384_ ? _037_ : nmi_mode_o;
assign nmi_mode_d = _355_ ? _083_ : _295_;
assign _297_ = _191_ ? 1'h1 : 1'h0;
assign flush_id_o = _355_ ? _030_ : _297_;
assign _298_ = _388_ ? 1'h1 : 1'h0;
assign debug_csr_save_o = _383_ ? _020_ : _298_;
assign _299_ = _384_ ? _015_ : 32'd0;
assign csr_mtval_o = _355_ ? _087_ : _299_;
assign _301_ = _355_ ? _072_ : _020_;
assign csr_save_if_o = _388_ ? 1'h1 : _302_;
assign csr_save_cause_o = _262_ ? _301_ : csr_save_if_o;
assign _303_ = _383_ ? _020_ : 1'h0;
assign csr_save_id_o = _355_ ? _052_ : _303_;
assign _302_ = _384_ ? _019_ : 1'h0;
assign _304_ = _384_ ? _028_ : 7'h00;
assign exc_cause_o = _355_ ? _109_ : _304_;
assign _305_ = _177_ ? 2'h2 : 2'h1;
assign exc_pc_mux_o = _355_ ? _029_ : _305_;
assign _306_ = _389_ ? 1'h0 : 1'h1;
assign ctrl_busy_o = _387_ ? _023_ : _306_;
assign _308_ = ! /* src = "generated/sv2v_out.v:12504.44-12504.64" */ priv_mode_i;
assign _307_ = priv_mode_i == /* src = "generated/sv2v_out.v:12709.39-12709.59" */ 2'h3;
assign _309_ = _328_ && /* src = "generated/sv2v_out.v:12622.9-12622.69" */ _329_;
assign _310_ = _317_ && /* src = "generated/sv2v_out.v:12624.10-12624.32" */ _318_;
assign _311_ = _310_ && /* src = "generated/sv2v_out.v:12624.9-12624.51" */ _319_;
assign _312_ = irq_nm && /* src = "generated/sv2v_out.v:12641.10-12641.31" */ _320_;
assign _313_ = ebreak_into_debug && /* src = "generated/sv2v_out.v:12675.9-12675.43" */ _321_;
assign _314_ = ebrk_insn_prio && /* src = "generated/sv2v_out.v:12747.38-12747.73" */ ebreak_into_debug;
assign _315_ = enter_debug_mode_prio_q && /* src = "generated/sv2v_out.v:12747.9-12747.74" */ _322_;
assign _316_ = ! /* src = "generated/sv2v_out.v:12469.25-12469.38" */ irq_nm_ext_i;
assign _317_ = ! /* src = "generated/sv2v_out.v:12624.10-12624.16" */ stall;
assign _318_ = ! /* src = "generated/sv2v_out.v:12624.20-12624.32" */ special_req;
assign _319_ = ! /* src = "generated/sv2v_out.v:12624.37-12624.51" */ id_wb_pending;
assign _320_ = ! /* src = "generated/sv2v_out.v:12641.20-12641.31" */ nmi_mode_o;
assign _321_ = ! /* src = "generated/sv2v_out.v:12675.30-12675.43" */ debug_mode_o;
assign _322_ = ! /* src = "generated/sv2v_out.v:12747.36-12747.74" */ _314_;
assign _323_ = irq_nm || /* src = "generated/sv2v_out.v:12589.12-12589.35" */ irq_pending_i;
assign _324_ = _323_ || /* src = "generated/sv2v_out.v:12589.11-12589.51" */ debug_req_i;
assign _325_ = _324_ || /* src = "generated/sv2v_out.v:12589.10-12589.68" */ debug_mode_o;
assign _326_ = _325_ || /* src = "generated/sv2v_out.v:12589.9-12589.92" */ debug_single_step_i;
assign _327_ = branch_set_i || /* src = "generated/sv2v_out.v:12614.9-12614.35" */ jump_set_i;
assign _328_ = enter_debug_mode || /* src = "generated/sv2v_out.v:12622.10-12622.40" */ handle_irq;
assign _329_ = stall || /* src = "generated/sv2v_out.v:12622.46-12622.68" */ id_wb_pending;
assign _330_ = exc_req_q || /* src = "generated/sv2v_out.v:12688.10-12688.34" */ store_err_q;
assign _331_ = _330_ || /* src = "generated/sv2v_out.v:12688.9-12688.49" */ load_err_q;
assign _332_ = ctrl_fsm_cs != /* src = "generated/sv2v_out.v:12401.88-12401.107" */ 4'h6;
assign _333_ = | /* src = "generated/sv2v_out.v:12647.15-12647.52" */ irqs_i[14:0];
assign _334_ = ~ /* src = "generated/sv2v_out.v:12463.39-12463.50" */ nmi_mode_o;
assign _335_ = ~ /* src = "generated/sv2v_out.v:12477.80-12477.108" */ \g_intg_irq_int.mem_resp_intg_err_irq_clear ;
assign _336_ = ~ /* src = "generated/sv2v_out.v:12505.40-12505.60" */ debug_single_step_i;
assign _337_ = ~ /* src = "generated/sv2v_out.v:12615.36-12615.53" */ instr_bp_taken_i;
assign _338_ = ~ /* src = "generated/sv2v_out.v:12762.35-12762.43" */ halt_if;
assign _339_ = ~ /* src = "generated/sv2v_out.v:12763.31-12763.51" */ _170_;
assign _341_ = ecall_insn | /* src = "generated/sv2v_out.v:12401.24-12401.46" */ ebrk_insn;
assign _343_ = _341_ | /* src = "generated/sv2v_out.v:12401.23-12401.64" */ illegal_insn_d;
assign _345_ = _343_ | /* src = "generated/sv2v_out.v:12401.22-12401.83" */ instr_fetch_err;
assign exc_req_lsu = store_err_i | /* src = "generated/sv2v_out.v:12402.23-12402.47" */ load_err_i;
assign special_req_flush_only = wfi_insn | /* src = "generated/sv2v_out.v:12404.34-12404.59" */ csr_pipe_flush;
assign _347_ = mret_insn | /* src = "generated/sv2v_out.v:12405.35-12405.56" */ dret_insn;
assign _348_ = _347_ | /* src = "generated/sv2v_out.v:12405.34-12405.69" */ exc_req_d;
assign special_req_pc_change = _348_ | /* src = "generated/sv2v_out.v:12405.33-12405.84" */ exc_req_lsu;
assign special_req = special_req_pc_change | /* src = "generated/sv2v_out.v:12406.23-12406.69" */ special_req_flush_only;
assign id_wb_pending = instr_valid_i | /* src = "generated/sv2v_out.v:12407.25-12407.52" */ _166_;
assign _054_ = load_err_q | /* src = "generated/sv2v_out.v:12430.30-12430.54" */ store_err_q;
assign _349_ = _054_ | /* src = "generated/sv2v_out.v:12430.29-12430.68" */ load_err_i;
assign wb_exception_o = _349_ | /* src = "generated/sv2v_out.v:12430.28-12430.83" */ store_err_i;
assign \g_intg_irq_int.mem_resp_intg_err_irq_pending_d  = _122_ | /* src = "generated/sv2v_out.v:12477.45-12477.137" */ \g_intg_irq_int.mem_resp_intg_err_irq_set ;
assign irq_nm_int = \g_intg_irq_int.mem_resp_intg_err_irq_set  | /* src = "generated/sv2v_out.v:12487.24-12487.83" */ \g_intg_irq_int.mem_resp_intg_err_irq_pending_q ;
assign _351_ = debug_req_i | /* src = "generated/sv2v_out.v:12500.36-12500.66" */ do_single_step_d;
assign enter_debug_mode = enter_debug_mode_prio_d | /* src = "generated/sv2v_out.v:12501.28-12501.87" */ _124_;
assign irq_nm = irq_nm_ext_i | /* src = "generated/sv2v_out.v:12503.18-12503.43" */ irq_nm_int;
assign irq_enabled = csr_mstatus_mie_i | /* src = "generated/sv2v_out.v:12504.23-12504.65" */ _308_;
assign _352_ = irq_nm | /* src = "generated/sv2v_out.v:12505.80-12505.118" */ _127_;
assign _353_ = ready_wb_i | /* src = "generated/sv2v_out.v:12611.10-12611.37" */ wb_exception_o;
assign _354_ = debug_mode_o | /* src = "generated/sv2v_out.v:12711.12-12711.44" */ ebreak_into_debug;
assign stall = stall_id_i | /* src = "generated/sv2v_out.v:12761.17-12761.40" */ stall_wb_i;
assign _170_ = stall | /* src = "generated/sv2v_out.v:12763.33-12763.50" */ retain_id;
assign instr_valid_clear_o = _339_ | /* src = "generated/sv2v_out.v:12763.31-12763.62" */ flush_id_o;
/* src = "generated/sv2v_out.v:12478.4-12486.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  <= 1'h0;
else \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  <= \g_intg_irq_int.mem_resp_intg_err_irq_pending_d ;
/* src = "generated/sv2v_out.v:12764.2-12787.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME nmi_mode_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) nmi_mode_o <= 1'h0;
else nmi_mode_o <= nmi_mode_d;
/* src = "generated/sv2v_out.v:12764.2-12787.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME load_err_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) load_err_q <= 1'h0;
else load_err_q <= load_err_i;
/* src = "generated/sv2v_out.v:12764.2-12787.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME store_err_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) store_err_q <= 1'h0;
else store_err_q <= store_err_i;
/* src = "generated/sv2v_out.v:12764.2-12787.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME exc_req_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) exc_req_q <= 1'h0;
else exc_req_q <= exc_req_d;
/* src = "generated/sv2v_out.v:12764.2-12787.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME illegal_insn_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) illegal_insn_q <= 1'h0;
else illegal_insn_q <= illegal_insn_d;
/* src = "generated/sv2v_out.v:12764.2-12787.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME do_single_step_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) do_single_step_q <= 1'h0;
else do_single_step_q <= do_single_step_d;
/* src = "generated/sv2v_out.v:12764.2-12787.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME enter_debug_mode_prio_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) enter_debug_mode_prio_q <= 1'h0;
else enter_debug_mode_prio_q <= enter_debug_mode_prio_d;
/* src = "generated/sv2v_out.v:12517.2-12521.35" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'1\BranchPredictor=1'1\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME debug_cause_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) debug_cause_o <= 3'h0;
else debug_cause_o <= debug_cause_d;
assign _032_ = mem_resp_intg_err_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12472.14-12472.33|generated/sv2v_out.v:12472.10-12475.8" */ 1'h1 : 1'h0;
assign _031_ = _121_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12469.10-12469.38|generated/sv2v_out.v:12469.6-12470.42" */ 1'h1 : 1'h0;
assign \g_intg_irq_int.mem_resp_intg_err_irq_clear  = \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12468.9-12468.40|generated/sv2v_out.v:12468.5-12475.8" */ _031_ : 1'h0;
assign \g_intg_irq_int.mem_resp_intg_err_irq_set  = \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12468.9-12468.40|generated/sv2v_out.v:12468.5-12475.8" */ 1'h0 : _032_;
assign _104_ = ebrk_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12427.14-12427.23|generated/sv2v_out.v:12427.10-12428.28" */ 1'h1 : 1'h0;
assign _093_ = ecall_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12425.14-12425.24|generated/sv2v_out.v:12425.10-12428.28" */ 1'h1 : 1'h0;
assign _092_ = ecall_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12425.14-12425.24|generated/sv2v_out.v:12425.10-12428.28" */ 1'h0 : _104_;
assign _081_ = illegal_insn_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12423.14-12423.28|generated/sv2v_out.v:12423.10-12428.28" */ 1'h1 : 1'h0;
assign _076_ = illegal_insn_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12423.14-12423.28|generated/sv2v_out.v:12423.10-12428.28" */ 1'h0 : _092_;
assign _077_ = illegal_insn_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12423.14-12423.28|generated/sv2v_out.v:12423.10-12428.28" */ 1'h0 : _093_;
assign _064_ = instr_fetch_err ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12421.14-12421.29|generated/sv2v_out.v:12421.10-12428.28" */ 1'h1 : 1'h0;
assign _058_ = instr_fetch_err ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12421.14-12421.29|generated/sv2v_out.v:12421.10-12428.28" */ 1'h0 : _076_;
assign _059_ = instr_fetch_err ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12421.14-12421.29|generated/sv2v_out.v:12421.10-12428.28" */ 1'h0 : _077_;
assign _063_ = instr_fetch_err ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12421.14-12421.29|generated/sv2v_out.v:12421.10-12428.28" */ 1'h0 : _081_;
assign _035_ = load_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12419.14-12419.24|generated/sv2v_out.v:12419.10-12428.28" */ 1'h1 : 1'h0;
assign _026_ = load_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12419.14-12419.24|generated/sv2v_out.v:12419.10-12428.28" */ 1'h0 : _058_;
assign _027_ = load_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12419.14-12419.24|generated/sv2v_out.v:12419.10-12428.28" */ 1'h0 : _059_;
assign _033_ = load_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12419.14-12419.24|generated/sv2v_out.v:12419.10-12428.28" */ 1'h0 : _063_;
assign _034_ = load_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12419.14-12419.24|generated/sv2v_out.v:12419.10-12428.28" */ 1'h0 : _064_;
assign store_err_prio = store_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12417.9-12417.20|generated/sv2v_out.v:12417.5-12428.28" */ 1'h1 : 1'h0;
assign load_err_prio = store_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12417.9-12417.20|generated/sv2v_out.v:12417.5-12428.28" */ 1'h0 : _035_;
assign ebrk_insn_prio = store_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12417.9-12417.20|generated/sv2v_out.v:12417.5-12428.28" */ 1'h0 : _026_;
assign ecall_insn_prio = store_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12417.9-12417.20|generated/sv2v_out.v:12417.5-12428.28" */ 1'h0 : _027_;
assign illegal_insn_prio = store_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12417.9-12417.20|generated/sv2v_out.v:12417.5-12428.28" */ 1'h0 : _033_;
assign instr_fetch_err_prio = store_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12417.9-12417.20|generated/sv2v_out.v:12417.5-12428.28" */ 1'h0 : _034_;
assign halt_if = instr_exec_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12755.7-12755.20|generated/sv2v_out.v:12755.3-12756.19" */ _013_ : 1'h1;
assign _012_ = _315_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12747.9-12747.74|generated/sv2v_out.v:12747.5-12748.25" */ 4'h8 : _002_;
assign _011_ = wfi_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12745.14-12745.22|generated/sv2v_out.v:12745.10-12746.25" */ 4'h2 : 4'h5;
assign _075_ = dret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12739.14-12739.23|generated/sv2v_out.v:12739.10-12746.25" */ 1'h0 : 1'hx;
assign _071_ = dret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12739.14-12739.23|generated/sv2v_out.v:12739.10-12746.25" */ 1'h1 : 1'h0;
assign _085_ = dret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12739.14-12739.23|generated/sv2v_out.v:12739.10-12746.25" */ 3'h4 : 3'h0;
assign _010_ = dret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12739.14-12739.23|generated/sv2v_out.v:12739.10-12746.25" */ 4'h5 : _011_;
assign _097_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12732.14-12732.23|generated/sv2v_out.v:12732.10-12746.25" */ 1'h0 : nmi_mode_o;
assign _051_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12732.14-12732.23|generated/sv2v_out.v:12732.10-12746.25" */ 1'h1 : 1'h0;
assign _112_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12732.14-12732.23|generated/sv2v_out.v:12732.10-12746.25" */ 1'h1 : _071_;
assign _068_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12732.14-12732.23|generated/sv2v_out.v:12732.10-12746.25" */ 3'h3 : _085_;
assign _057_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12732.14-12732.23|generated/sv2v_out.v:12732.10-12746.25" */ 1'hx : _075_;
assign _008_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12732.14-12732.23|generated/sv2v_out.v:12732.10-12746.25" */ 4'h5 : _010_;
assign _050_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12732.14-12732.23|generated/sv2v_out.v:12732.10-12746.25" */ 1'h0 : _071_;
assign _006_ = _354_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12711.12-12711.44|generated/sv2v_out.v:12711.8-12719.51" */ 4'h9 : 4'h5;
assign _101_ = _354_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12711.12-12711.44|generated/sv2v_out.v:12711.8-12719.51" */ 1'h0 : _073_;
assign _079_ = _354_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12711.12-12711.44|generated/sv2v_out.v:12711.8-12719.51" */ 1'h0 : 1'h1;
assign _117_ = _354_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12711.12-12711.44|generated/sv2v_out.v:12711.8-12719.51" */ 7'h00 : 7'h03;
assign _356_ = load_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ lsu_addr_last_i : 32'd0;
assign _358_ = store_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ lsu_addr_last_i : _356_;
assign _360_ = ebrk_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ 32'd0 : _358_;
assign _362_ = ecall_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ 32'd0 : _360_;
assign _364_ = illegal_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ _400_ : _362_;
assign _099_ = instr_fetch_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ _398_ : _364_;
assign _366_ = load_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ 7'h05 : 7'h00;
assign _367_ = store_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ 7'h07 : _366_;
assign _368_ = ebrk_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ _117_ : _367_;
assign _369_ = ecall_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ _402_ : _368_;
assign _370_ = illegal_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ 7'h02 : _369_;
assign _114_ = instr_fetch_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ 7'h01 : _370_;
assign _371_ = ebrk_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ _006_ : 4'h5;
assign _372_ = ecall_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ 4'h5 : _371_;
assign _373_ = illegal_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ 4'h5 : _372_;
assign _004_ = instr_fetch_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ 4'h5 : _373_;
assign _377_ = ebrk_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ _101_ : _073_;
assign _379_ = ecall_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ _073_ : _377_;
assign _381_ = illegal_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ _073_ : _379_;
assign _089_ = instr_fetch_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ _073_ : _381_;
assign _374_ = ebrk_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ _079_ : 1'h1;
assign _375_ = ecall_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ 1'h1 : _374_;
assign _376_ = illegal_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ 1'h1 : _375_;
assign _061_ = instr_fetch_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12700.6-12730.13" */ 1'h1 : _376_;
assign _002_ = _331_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12688.9-12688.49|generated/sv2v_out.v:12688.5-12746.25" */ _004_ : _008_;
assign _030_ = _331_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12688.9-12688.49|generated/sv2v_out.v:12688.5-12746.25" */ _061_ : 1'h1;
assign _087_ = _331_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12688.9-12688.49|generated/sv2v_out.v:12688.5-12746.25" */ _099_ : 32'd0;
assign _072_ = _331_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12688.9-12688.49|generated/sv2v_out.v:12688.5-12746.25" */ _061_ : 1'h0;
assign _052_ = _331_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12688.9-12688.49|generated/sv2v_out.v:12688.5-12746.25" */ _089_ : 1'h0;
assign _109_ = _331_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12688.9-12688.49|generated/sv2v_out.v:12688.5-12746.25" */ _114_ : 7'h00;
assign _086_ = _331_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12688.9-12688.49|generated/sv2v_out.v:12688.5-12746.25" */ _061_ : _112_;
assign _021_ = _331_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12688.9-12688.49|generated/sv2v_out.v:12688.5-12746.25" */ _054_ : 1'h0;
assign _029_ = _331_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12688.9-12688.49|generated/sv2v_out.v:12688.5-12746.25" */ _397_ : 2'h1;
assign _040_ = _331_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12688.9-12688.49|generated/sv2v_out.v:12688.5-12746.25" */ 3'h2 : _068_;
assign _025_ = _331_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12688.9-12688.49|generated/sv2v_out.v:12688.5-12746.25" */ 1'hx : _057_;
assign _083_ = _331_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12688.9-12688.49|generated/sv2v_out.v:12688.5-12746.25" */ nmi_mode_o : _097_;
assign _017_ = _331_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12688.9-12688.49|generated/sv2v_out.v:12688.5-12746.25" */ 1'h0 : _050_;
assign _018_ = _331_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12688.9-12688.49|generated/sv2v_out.v:12688.5-12746.25" */ 1'h0 : _051_;
assign _020_ = _313_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12675.9-12675.43|generated/sv2v_out.v:12675.5-12679.8" */ 1'h1 : 1'h0;
assign _105_ = irqs_i[17] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12651.15-12651.25|generated/sv2v_out.v:12651.11-12654.48" */ 7'h23 : 7'h27;
assign _094_ = irqs_i[15] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12649.15-12649.25|generated/sv2v_out.v:12649.11-12654.48" */ 7'h2b : _105_;
assign _078_ = _333_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12647.15-12647.52|generated/sv2v_out.v:12647.11-12654.48" */ { 3'h3, mfip_id } : _094_;
assign _069_ = _130_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12643.11-12643.37|generated/sv2v_out.v:12643.7-12644.39" */ \g_intg_irq_int.mem_resp_intg_err_addr_q  : 32'd0;
assign _066_ = _312_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12641.10-12641.31|generated/sv2v_out.v:12641.6-12654.48" */ 1'h1 : nmi_mode_o;
assign _048_ = _312_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12641.10-12641.31|generated/sv2v_out.v:12641.6-12654.48" */ _069_ : 32'd0;
assign _060_ = _312_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12641.10-12641.31|generated/sv2v_out.v:12641.6-12654.48" */ _396_ : _078_;
assign _037_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12637.9-12637.19|generated/sv2v_out.v:12637.5-12655.8" */ _066_ : nmi_mode_o;
assign _015_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12637.9-12637.19|generated/sv2v_out.v:12637.5-12655.8" */ _048_ : 32'd0;
assign _028_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12637.9-12637.19|generated/sv2v_out.v:12637.5-12655.8" */ _060_ : 7'h00;
assign _019_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12637.9-12637.19|generated/sv2v_out.v:12637.5-12655.8" */ 1'h1 : 1'h0;
assign _110_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12629.15-12629.25|generated/sv2v_out.v:12629.11-12632.9" */ 1'h1 : _080_;
assign _000_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12629.15-12629.25|generated/sv2v_out.v:12629.11-12632.9" */ 4'h7 : _103_;
assign _106_ = enter_debug_mode ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12625.10-12625.26|generated/sv2v_out.v:12625.6-12632.9" */ 1'h1 : _110_;
assign _116_ = enter_debug_mode ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12625.10-12625.26|generated/sv2v_out.v:12625.6-12632.9" */ 4'h8 : _000_;
assign _095_ = _311_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12624.9-12624.51|generated/sv2v_out.v:12624.5-12632.9" */ _106_ : _080_;
assign _113_ = _311_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12624.9-12624.51|generated/sv2v_out.v:12624.5-12632.9" */ _116_ : _103_;
assign _080_ = _309_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12622.9-12622.69|generated/sv2v_out.v:12622.5-12623.21" */ 1'h1 : 1'h0;
assign _039_ = _129_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12620.10-12620.45|generated/sv2v_out.v:12620.6-12621.37" */ 1'h1 : 1'h0;
assign _043_ = _327_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12614.9-12614.35|generated/sv2v_out.v:12614.5-12618.8" */ jump_set_i : 1'h0;
assign _045_ = _327_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12614.9-12614.35|generated/sv2v_out.v:12614.5-12618.8" */ branch_set_i : 1'h0;
assign _041_ = _327_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12614.9-12614.35|generated/sv2v_out.v:12614.5-12618.8" */ _337_ : 1'h0;
assign _108_ = _353_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12611.10-12611.37|generated/sv2v_out.v:12611.6-12612.26" */ 4'h6 : ctrl_fsm_cs;
assign _103_ = special_req ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12609.9-12609.20|generated/sv2v_out.v:12609.5-12613.8" */ _108_ : ctrl_fsm_cs;
assign _047_ = special_req ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12609.9-12609.20|generated/sv2v_out.v:12609.5-12613.8" */ 1'h1 : 1'h0;
assign _062_ = enter_debug_mode ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12601.9-12601.25|generated/sv2v_out.v:12601.5-12604.8" */ 1'h1 : _019_;
assign _091_ = enter_debug_mode ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12601.9-12601.25|generated/sv2v_out.v:12601.5-12604.8" */ 4'h8 : _074_;
assign _074_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12597.9-12597.19|generated/sv2v_out.v:12597.5-12600.8" */ 4'h7 : _056_;
assign _056_ = id_in_ready_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12595.9-12595.22|generated/sv2v_out.v:12595.5-12596.25" */ 4'h5 : 4'hx;
assign _024_ = _326_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12589.9-12589.92|generated/sv2v_out.v:12589.5-12592.25" */ 4'h4 : 4'hx;
assign _023_ = _326_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12589.9-12589.92|generated/sv2v_out.v:12589.5-12592.25" */ 1'h1 : 1'h0;
assign _391_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ ctrl_fsm_cs;
assign instr_req_o = _192_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ 1'h1 : 1'h0;
assign _390_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ 4'h1;
assign retain_id = _385_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ _047_ : 1'h0;
assign _386_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ 4'h4;
assign controller_run_o = _385_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ 1'h1 : 1'h0;
assign _387_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ 4'h3;
assign _389_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ 4'h2;
assign perf_tbranch_o = _385_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ _045_ : 1'h0;
assign perf_jump_o = _385_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ _043_ : 1'h0;
assign _385_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ 4'h5;
assign debug_mode_entering_o = _177_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ 1'h1 : 1'h0;
assign _383_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ 4'h9;
assign _388_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ 4'h8;
assign _355_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ 4'h6;
assign _384_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ 4'h7;
assign csr_restore_dret_id_o = _355_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ _017_ : 1'h0;
assign csr_restore_mret_id_o = _355_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ _018_ : 1'h0;
assign csr_save_wb_o = _355_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ _021_ : 1'h0;
assign nt_branch_mispredict_o = _385_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12565.3-12754.10" */ _039_ : 1'h0;
assign mfip_id = irqs_i[0] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12511.9-12511.22|generated/sv2v_out.v:12511.5-12512.23" */ 4'h0 : _009_;
assign _009_ = irqs_i[1] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12511.9-12511.22|generated/sv2v_out.v:12511.5-12512.23" */ 4'h1 : _007_;
assign _007_ = irqs_i[2] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12511.9-12511.22|generated/sv2v_out.v:12511.5-12512.23" */ 4'h2 : _005_;
assign _005_ = irqs_i[3] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12511.9-12511.22|generated/sv2v_out.v:12511.5-12512.23" */ 4'h3 : _003_;
assign _003_ = irqs_i[4] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12511.9-12511.22|generated/sv2v_out.v:12511.5-12512.23" */ 4'h4 : _001_;
assign _001_ = irqs_i[5] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12511.9-12511.22|generated/sv2v_out.v:12511.5-12512.23" */ 4'h5 : _118_;
assign _118_ = irqs_i[6] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12511.9-12511.22|generated/sv2v_out.v:12511.5-12512.23" */ 4'h6 : _115_;
assign _115_ = irqs_i[7] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12511.9-12511.22|generated/sv2v_out.v:12511.5-12512.23" */ 4'h7 : _111_;
assign _111_ = irqs_i[8] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12511.9-12511.22|generated/sv2v_out.v:12511.5-12512.23" */ 4'h8 : _107_;
assign _107_ = irqs_i[9] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12511.9-12511.22|generated/sv2v_out.v:12511.5-12512.23" */ 4'h9 : _096_;
assign _096_ = irqs_i[10] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12511.9-12511.22|generated/sv2v_out.v:12511.5-12512.23" */ 4'ha : _082_;
assign _082_ = irqs_i[11] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12511.9-12511.22|generated/sv2v_out.v:12511.5-12512.23" */ 4'hb : _065_;
assign _065_ = irqs_i[12] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12511.9-12511.22|generated/sv2v_out.v:12511.5-12512.23" */ 4'hc : _036_;
assign _036_ = irqs_i[13] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12511.9-12511.22|generated/sv2v_out.v:12511.5-12512.23" */ 4'hd : _014_;
assign _014_ = irqs_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12511.9-12511.22|generated/sv2v_out.v:12511.5-12512.23" */ 4'he : 4'h0;
assign do_single_step_d = instr_valid_i ? /* src = "generated/sv2v_out.v:12499.29-12499.99" */ _123_ : do_single_step_q;
assign _392_ = _308_ ? /* src = "generated/sv2v_out.v:12502.72-12502.117" */ debug_ebreaku_i : 1'h0;
assign ebreak_into_debug = _307_ ? /* src = "generated/sv2v_out.v:12502.30-12502.118" */ debug_ebreakm_i : _392_;
assign _393_ = do_single_step_d ? /* src = "generated/sv2v_out.v:12516.119-12516.149" */ 3'h4 : 3'h0;
assign _394_ = debug_req_i ? /* src = "generated/sv2v_out.v:12516.97-12516.150" */ 3'h3 : _393_;
assign _395_ = _128_ ? /* src = "generated/sv2v_out.v:12516.52-12516.151" */ 3'h1 : _394_;
assign debug_cause_d = trigger_match_i ? /* src = "generated/sv2v_out.v:12516.26-12516.152" */ 3'h2 : _395_;
assign _396_ = irq_nm_ext_i ? /* src = "generated/sv2v_out.v:12642.22-12642.87" */ 7'h3f : 7'h40;
assign _397_ = debug_mode_o ? /* src = "generated/sv2v_out.v:12691.22-12691.48" */ 2'h3 : 2'h0;
assign _398_ = instr_fetch_err_plus2_i ? /* src = "generated/sv2v_out.v:12703.23-12703.74" */ _119_ : pc_id_i;
assign _400_ = instr_is_compressed_i ? /* src = "generated/sv2v_out.v:12707.23-12707.99" */ { 16'h0000, instr_compressed_i } : instr_i;
assign _402_ = _307_ ? /* src = "generated/sv2v_out.v:12709.39-12709.119" */ 7'h0b : 7'h08;
assign controller_run_o_t0 = 1'h0;
assign csr_restore_dret_id_o_t0 = 1'h0;
assign csr_restore_mret_id_o_t0 = 1'h0;
assign csr_save_cause_o_t0 = 1'h0;
assign csr_save_if_o_t0 = 1'h0;
assign ctrl_busy_o_t0 = 1'h0;
assign debug_cause_o_t0 = 3'h0;
assign debug_csr_save_o_t0 = 1'h0;
assign debug_mode_entering_o_t0 = 1'h0;
assign exc_cause_o_t0 = 7'h00;
assign exc_pc_mux_o_t0 = 2'h0;
assign flush_id_o_t0 = 1'h0;
assign instr_req_o_t0 = 1'h0;
assign nt_branch_mispredict_o_t0 = 1'h0;
assign pc_mux_o_t0 = 3'h0;
endmodule

module \$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000 (clk_i, rst_ni, counter_inc_i, counterh_we_i, counter_we_i, counter_val_i, counter_val_o, counter_val_upd_o, counter_inc_i_t0, counter_val_i_t0, counter_val_o_t0, counter_val_upd_o_t0, counter_we_i_t0, counterh_we_i_t0);
/* src = "generated/sv2v_out.v:13678.2-13692.5" */
wire [63:0] _00_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13678.2-13692.5" */
wire [63:0] _01_;
wire [63:0] _02_;
wire _03_;
wire _04_;
wire [63:0] _05_;
wire [31:0] _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire [63:0] _12_;
wire [31:0] _13_;
wire [31:0] _14_;
wire [31:0] _15_;
wire [31:0] _16_;
wire [63:0] _17_;
wire [63:0] _18_;
wire [63:0] _19_;
wire [31:0] _20_;
wire [31:0] _21_;
wire [63:0] _22_;
wire [63:0] _23_;
wire [63:0] _24_;
/* src = "generated/sv2v_out.v:13664.13-13664.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:13676.27-13676.36" */
wire [63:0] counter_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13676.27-13676.36" */
wire [63:0] counter_d_t0;
/* src = "generated/sv2v_out.v:13666.13-13666.26" */
input counter_inc_i;
wire counter_inc_i;
/* cellift = 32'd1 */
input counter_inc_i_t0;
wire counter_inc_i_t0;
/* src = "generated/sv2v_out.v:13674.13-13674.25" */
wire [63:0] counter_load;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13674.13-13674.25" */
wire [63:0] counter_load_t0;
/* src = "generated/sv2v_out.v:13673.28-13673.39" */
wire [63:0] counter_upd;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13673.28-13673.39" */
wire [63:0] counter_upd_t0;
/* src = "generated/sv2v_out.v:13669.20-13669.33" */
input [31:0] counter_val_i;
wire [31:0] counter_val_i;
/* cellift = 32'd1 */
input [31:0] counter_val_i_t0;
wire [31:0] counter_val_i_t0;
/* src = "generated/sv2v_out.v:13670.21-13670.34" */
output [63:0] counter_val_o;
reg [63:0] counter_val_o;
/* cellift = 32'd1 */
output [63:0] counter_val_o_t0;
reg [63:0] counter_val_o_t0;
/* src = "generated/sv2v_out.v:13671.21-13671.38" */
output [63:0] counter_val_upd_o;
wire [63:0] counter_val_upd_o;
/* cellift = 32'd1 */
output [63:0] counter_val_upd_o_t0;
wire [63:0] counter_val_upd_o_t0;
/* src = "generated/sv2v_out.v:13668.13-13668.25" */
input counter_we_i;
wire counter_we_i;
/* cellift = 32'd1 */
input counter_we_i_t0;
wire counter_we_i_t0;
/* src = "generated/sv2v_out.v:13667.13-13667.26" */
input counterh_we_i;
wire counterh_we_i;
/* cellift = 32'd1 */
input counterh_we_i_t0;
wire counterh_we_i_t0;
/* src = "generated/sv2v_out.v:13665.13-13665.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:13675.6-13675.8" */
wire we;
assign counter_upd = counter_val_o + /* src = "generated/sv2v_out.v:13677.23-13677.86" */ 64'h0000000000000001;
assign _02_ = ~ counter_val_o_t0;
assign _12_ = counter_val_o & _02_;
assign _23_ = _12_ + 64'h0000000000000001;
assign _19_ = counter_val_o | counter_val_o_t0;
assign _24_ = _19_ + 64'h0000000000000001;
assign _22_ = _23_ ^ _24_;
assign counter_upd_t0 = _22_ | counter_val_o_t0;
assign _03_ = ~ _10_;
assign _04_ = ~ _11_;
assign _13_ = { _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_, _10_ } & counter_d_t0[63:32];
assign _15_ = { _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_, _11_ } & counter_d_t0[31:0];
assign _14_ = { _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_, _03_ } & counter_val_o_t0[63:32];
assign _16_ = { _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_, _04_ } & counter_val_o_t0[31:0];
assign _20_ = _13_ | _14_;
assign _21_ = _15_ | _16_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000  */
/* PC_TAINT_INFO STATE_NAME counter_val_o_t0[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o_t0[63:32] <= 32'd0;
else counter_val_o_t0[63:32] <= _20_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000  */
/* PC_TAINT_INFO STATE_NAME counter_val_o_t0[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o_t0[31:0] <= 32'd0;
else counter_val_o_t0[31:0] <= _21_;
/* src = "generated/sv2v_out.v:13694.2-13698.27" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000  */
/* PC_TAINT_INFO STATE_NAME counter_val_o[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o[63:32] <= 32'd0;
else if (_10_) counter_val_o[63:32] <= counter_d[63:32];
/* src = "generated/sv2v_out.v:13694.2-13698.27" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000  */
/* PC_TAINT_INFO STATE_NAME counter_val_o[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o[31:0] <= 32'd0;
else if (_11_) counter_val_o[31:0] <= counter_d[31:0];
assign _05_ = ~ { we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we };
assign _06_ = ~ { counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i };
assign _17_ = _05_ & _01_;
assign counter_load_t0[31:0] = _06_ & counter_val_i_t0;
assign _01_ = { counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i } & counter_upd_t0;
assign _18_ = { we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we } & counter_load_t0;
assign counter_load_t0[63:32] = { counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i } & counter_val_i_t0;
assign counter_d_t0 = _17_ | _18_;
assign _07_ = | { we, counter_inc_i };
assign _08_ = { we, counterh_we_i } != 2'h2;
assign _09_ = { we, counterh_we_i } != 2'h3;
assign _10_ = & { _07_, _08_ };
assign _11_ = & { _07_, _09_ };
assign we = counter_we_i | /* src = "generated/sv2v_out.v:13679.8-13679.36" */ counterh_we_i;
assign _00_ = counter_inc_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13688.12-13688.25|generated/sv2v_out.v:13688.8-13691.44" */ counter_upd : 64'hxxxxxxxxxxxxxxxx;
assign counter_d = we ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13686.7-13686.9|generated/sv2v_out.v:13686.3-13691.44" */ counter_load : _00_;
assign counter_load[63:32] = counterh_we_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13682.7-13682.20|generated/sv2v_out.v:13682.3-13685.6" */ counter_val_i : 32'hxxxxxxxx;
assign counter_load[31:0] = counterh_we_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13682.7-13682.20|generated/sv2v_out.v:13682.3-13685.6" */ 32'hxxxxxxxx : counter_val_i;
assign counter_val_upd_o = 64'h0000000000000000;
assign counter_val_upd_o_t0 = 64'h0000000000000000;
endmodule

module \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1 (clk_i, rst_ni, clear_i, busy_o, in_valid_i, in_addr_i, in_rdata_i, in_err_i, out_valid_o, out_ready_i, out_addr_o, out_rdata_o, out_err_o, out_err_plus2_o, clear_i_t0, busy_o_t0, out_valid_o_t0, out_ready_i_t0, out_rdata_o_t0, out_err_plus2_o_t0, out_err_o_t0
, out_addr_o_t0, in_valid_i_t0, in_rdata_i_t0, in_err_i_t0, in_addr_i_t0);
/* src = "generated/sv2v_out.v:16192.2-16207.6" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16192.2-16207.6" */
wire _001_;
/* src = "generated/sv2v_out.v:16187.40-16187.75" */
wire _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16187.40-16187.75" */
wire _003_;
/* src = "generated/sv2v_out.v:16187.91-16187.112" */
wire _004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16187.91-16187.112" */
wire _005_;
/* src = "generated/sv2v_out.v:16187.117-16187.168" */
wire _006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16187.117-16187.168" */
wire _007_;
/* src = "generated/sv2v_out.v:16188.35-16188.55" */
wire _008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16188.35-16188.55" */
wire _009_;
/* src = "generated/sv2v_out.v:16188.59-16188.80" */
wire _010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16188.59-16188.80" */
wire _011_;
/* src = "generated/sv2v_out.v:16188.58-16188.93" */
wire _012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16188.58-16188.93" */
wire _013_;
/* src = "generated/sv2v_out.v:16189.48-16189.71" */
wire _014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16189.48-16189.71" */
wire _015_;
/* src = "generated/sv2v_out.v:16208.36-16208.61" */
wire _016_;
/* src = "generated/sv2v_out.v:16239.30-16239.63" */
wire _017_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16239.30-16239.63" */
wire _018_;
/* src = "generated/sv2v_out.v:16239.30-16239.63" */
wire _019_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16239.30-16239.63" */
wire _020_;
/* src = "generated/sv2v_out.v:16242.26-16242.56" */
wire _021_;
/* src = "generated/sv2v_out.v:16242.61-16242.108" */
wire _022_;
/* src = "generated/sv2v_out.v:16242.26-16242.56" */
wire _023_;
/* src = "generated/sv2v_out.v:16242.61-16242.108" */
wire _024_;
wire [30:0] _025_;
wire [30:0] _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire [31:0] _033_;
wire [31:0] _034_;
wire [31:0] _035_;
wire _036_;
wire [30:0] _037_;
wire _038_;
wire [31:0] _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire [30:0] _049_;
wire [30:0] _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire [31:0] _098_;
wire [31:0] _099_;
wire _100_;
wire _101_;
wire [31:0] _102_;
wire [31:0] _103_;
wire _104_;
wire _105_;
wire [31:0] _106_;
wire [31:0] _107_;
wire [30:0] _108_;
wire [30:0] _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire [31:0] _136_;
wire [31:0] _137_;
wire [31:0] _138_;
wire [31:0] _139_;
wire _140_;
wire [31:0] _141_;
wire [31:0] _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire [30:0] _148_;
wire [30:0] _149_;
wire _150_;
wire _151_;
wire [31:0] _152_;
wire [31:0] _153_;
wire [31:0] _154_;
wire [31:0] _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire [30:0] _160_;
wire [30:0] _161_;
wire [30:0] _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire [31:0] _179_;
wire _180_;
wire [31:0] _181_;
wire _182_;
wire [31:0] _183_;
wire [30:0] _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire [30:0] _192_;
wire [30:0] _193_;
wire [30:0] _194_;
/* src = "generated/sv2v_out.v:16190.36-16190.57" */
wire _195_;
/* src = "generated/sv2v_out.v:16191.34-16191.53" */
wire _196_;
/* src = "generated/sv2v_out.v:16190.61-16190.65" */
wire _197_;
/* src = "generated/sv2v_out.v:16210.56-16210.70" */
wire _198_;
/* src = "generated/sv2v_out.v:16229.51-16229.73" */
wire _199_;
/* src = "generated/sv2v_out.v:16187.39-16187.87" */
wire _200_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16187.39-16187.87" */
wire _201_;
/* src = "generated/sv2v_out.v:16187.129-16187.167" */
wire _202_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16187.129-16187.167" */
wire _203_;
/* src = "generated/sv2v_out.v:16187.90-16187.169" */
wire _204_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16187.90-16187.169" */
wire _205_;
/* src = "generated/sv2v_out.v:16229.51-16229.89" */
wire _206_;
/* src = "generated/sv2v_out.v:16177.7-16177.20" */
wire addr_incr_two;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16177.7-16177.20" */
wire addr_incr_two_t0;
/* src = "generated/sv2v_out.v:16175.7-16175.28" */
wire aligned_is_compressed;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16175.7-16175.28" */
wire aligned_is_compressed_t0;
/* src = "generated/sv2v_out.v:16145.31-16145.37" */
output [1:0] busy_o;
wire [1:0] busy_o;
/* cellift = 32'd1 */
output [1:0] busy_o_t0;
wire [1:0] busy_o_t0;
/* src = "generated/sv2v_out.v:16144.13-16144.20" */
input clear_i;
wire clear_i;
/* cellift = 32'd1 */
input clear_i_t0;
wire clear_i_t0;
/* src = "generated/sv2v_out.v:16142.13-16142.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:16166.21-16166.29" */
wire [2:0] entry_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16166.21-16166.29" */
/* unused_bits = "0 1" */
wire [2:0] entry_en_t0;
/* src = "generated/sv2v_out.v:16170.7-16170.10" */
wire err;
/* src = "generated/sv2v_out.v:16159.21-16159.26" */
wire [2:0] err_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16159.21-16159.26" */
wire [2:0] err_d_t0;
/* src = "generated/sv2v_out.v:16172.7-16172.16" */
wire err_plus2;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16172.7-16172.16" */
wire err_plus2_t0;
/* src = "generated/sv2v_out.v:16160.20-16160.25" */
reg [2:0] err_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16160.20-16160.25" */
reg [2:0] err_q_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16170.7-16170.10" */
wire err_t0;
/* src = "generated/sv2v_out.v:16171.7-16171.20" */
wire err_unaligned;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16171.7-16171.20" */
wire err_unaligned_t0;
/* src = "generated/sv2v_out.v:16147.20-16147.29" */
input [31:0] in_addr_i;
wire [31:0] in_addr_i;
/* cellift = 32'd1 */
input [31:0] in_addr_i_t0;
wire [31:0] in_addr_i_t0;
/* src = "generated/sv2v_out.v:16149.13-16149.21" */
input in_err_i;
wire in_err_i;
/* cellift = 32'd1 */
input in_err_i_t0;
wire in_err_i_t0;
/* src = "generated/sv2v_out.v:16148.20-16148.30" */
input [31:0] in_rdata_i;
wire [31:0] in_rdata_i;
/* cellift = 32'd1 */
input [31:0] in_rdata_i_t0;
wire [31:0] in_rdata_i_t0;
/* src = "generated/sv2v_out.v:16146.13-16146.23" */
input in_valid_i;
wire in_valid_i;
/* cellift = 32'd1 */
input in_valid_i_t0;
wire in_valid_i_t0;
/* src = "generated/sv2v_out.v:16179.14-16179.26" */
wire [31:1] instr_addr_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16179.14-16179.26" */
wire [31:1] instr_addr_d_t0;
/* src = "generated/sv2v_out.v:16181.7-16181.20" */
wire instr_addr_en;
/* src = "generated/sv2v_out.v:16178.14-16178.29" */
wire [31:1] instr_addr_next;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16178.14-16178.29" */
wire [31:1] instr_addr_next_t0;
/* src = "generated/sv2v_out.v:16180.13-16180.25" */
reg [31:1] instr_addr_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16180.13-16180.25" */
reg [31:1] instr_addr_q_t0;
/* src = "generated/sv2v_out.v:16163.21-16163.38" */
wire [2:0] lowest_free_entry;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16163.21-16163.38" */
wire [2:0] lowest_free_entry_t0;
/* src = "generated/sv2v_out.v:16152.21-16152.31" */
output [31:0] out_addr_o;
wire [31:0] out_addr_o;
/* cellift = 32'd1 */
output [31:0] out_addr_o_t0;
wire [31:0] out_addr_o_t0;
/* src = "generated/sv2v_out.v:16154.13-16154.22" */
output out_err_o;
wire out_err_o;
/* cellift = 32'd1 */
output out_err_o_t0;
wire out_err_o_t0;
/* src = "generated/sv2v_out.v:16155.13-16155.28" */
output out_err_plus2_o;
wire out_err_plus2_o;
/* cellift = 32'd1 */
output out_err_plus2_o_t0;
wire out_err_plus2_o_t0;
/* src = "generated/sv2v_out.v:16153.20-16153.31" */
output [31:0] out_rdata_o;
wire [31:0] out_rdata_o;
/* cellift = 32'd1 */
output [31:0] out_rdata_o_t0;
wire [31:0] out_rdata_o_t0;
/* src = "generated/sv2v_out.v:16151.13-16151.24" */
input out_ready_i;
wire out_ready_i;
/* cellift = 32'd1 */
input out_ready_i_t0;
wire out_ready_i_t0;
/* src = "generated/sv2v_out.v:16150.13-16150.24" */
output out_valid_o;
wire out_valid_o;
/* cellift = 32'd1 */
output out_valid_o_t0;
wire out_valid_o_t0;
/* src = "generated/sv2v_out.v:16167.7-16167.15" */
wire pop_fifo;
/* src = "generated/sv2v_out.v:16168.14-16168.19" */
wire [31:0] rdata;
/* src = "generated/sv2v_out.v:16157.28-16157.35" */
wire [95:0] rdata_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16157.28-16157.35" */
wire [95:0] rdata_d_t0;
/* src = "generated/sv2v_out.v:16158.27-16158.34" */
reg [95:0] rdata_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16158.27-16158.34" */
reg [95:0] rdata_q_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16168.14-16168.19" */
wire [31:0] rdata_t0;
/* src = "generated/sv2v_out.v:16169.14-16169.29" */
wire [31:0] rdata_unaligned;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16169.14-16169.29" */
wire [31:0] rdata_unaligned_t0;
/* src = "generated/sv2v_out.v:16143.13-16143.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:16176.7-16176.30" */
wire unaligned_is_compressed;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16176.7-16176.30" */
wire unaligned_is_compressed_t0;
/* src = "generated/sv2v_out.v:16173.7-16173.12" */
wire valid;
/* src = "generated/sv2v_out.v:16161.21-16161.28" */
wire [2:0] valid_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16161.21-16161.28" */
wire [2:0] valid_d_t0;
/* src = "generated/sv2v_out.v:16165.21-16165.33" */
wire [2:0] valid_popped;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16165.21-16165.33" */
wire [2:0] valid_popped_t0;
/* src = "generated/sv2v_out.v:16164.21-16164.33" */
wire [2:0] valid_pushed;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16164.21-16164.33" */
wire [2:0] valid_pushed_t0;
/* src = "generated/sv2v_out.v:16162.20-16162.27" */
reg [2:0] valid_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16162.20-16162.27" */
reg [2:0] valid_q_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16173.7-16173.12" */
wire valid_t0;
/* src = "generated/sv2v_out.v:16174.7-16174.22" */
wire valid_unaligned;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16174.7-16174.22" */
wire valid_unaligned_t0;
assign instr_addr_next = instr_addr_q + /* src = "generated/sv2v_out.v:16210.27-16210.86" */ { 29'h00000000, _198_, addr_incr_two };
assign _002_ = err_q[1] & /* src = "generated/sv2v_out.v:16187.40-16187.75" */ _031_;
assign _004_ = valid_q[0] & /* src = "generated/sv2v_out.v:16187.91-16187.112" */ err_q[0];
assign _006_ = in_err_i & /* src = "generated/sv2v_out.v:16187.117-16187.168" */ _202_;
assign _008_ = err_q[1] & /* src = "generated/sv2v_out.v:16188.35-16188.55" */ _047_;
assign _010_ = in_err_i & /* src = "generated/sv2v_out.v:16188.59-16188.80" */ valid_q[0];
assign _012_ = _010_ & /* src = "generated/sv2v_out.v:16188.58-16188.93" */ _047_;
assign _014_ = valid_q[0] & /* src = "generated/sv2v_out.v:16189.48-16189.71" */ in_valid_i;
assign unaligned_is_compressed = _195_ & /* src = "generated/sv2v_out.v:16190.35-16190.65" */ _197_;
assign aligned_is_compressed = _196_ & /* src = "generated/sv2v_out.v:16191.33-16191.61" */ _197_;
assign _016_ = out_ready_i & /* src = "generated/sv2v_out.v:16229.21-16229.46" */ out_valid_o;
assign pop_fifo = _016_ & /* src = "generated/sv2v_out.v:16229.20-16229.90" */ _206_;
assign lowest_free_entry[1] = _036_ & /* src = "generated/sv2v_out.v:16237.35-16237.63" */ valid_q[0];
assign valid_d[0] = valid_popped[0] & /* src = "generated/sv2v_out.v:16241.24-16241.50" */ _043_;
assign valid_d[1] = valid_popped[1] & /* src = "generated/sv2v_out.v:16241.24-16241.50" */ _043_;
assign _021_ = valid_pushed[1] & /* src = "generated/sv2v_out.v:16242.26-16242.56" */ pop_fifo;
assign _017_ = in_valid_i & /* src = "generated/sv2v_out.v:16242.62-16242.95" */ lowest_free_entry[0];
assign _022_ = _017_ & /* src = "generated/sv2v_out.v:16242.61-16242.108" */ _038_;
assign _023_ = valid_pushed[2] & /* src = "generated/sv2v_out.v:16242.26-16242.56" */ pop_fifo;
assign _019_ = in_valid_i & /* src = "generated/sv2v_out.v:16242.62-16242.95" */ lowest_free_entry[1];
assign _024_ = _019_ & /* src = "generated/sv2v_out.v:16242.61-16242.108" */ _038_;
assign lowest_free_entry[2] = _040_ & /* src = "generated/sv2v_out.v:16247.40-16247.80" */ valid_q[1];
assign valid_d[2] = valid_popped[2] & /* src = "generated/sv2v_out.v:16250.30-16250.64" */ _043_;
assign entry_en[2] = in_valid_i & /* src = "generated/sv2v_out.v:16251.31-16251.72" */ lowest_free_entry[2];
assign _025_ = ~ instr_addr_q_t0;
assign _026_ = ~ { 29'h00000000, addr_incr_two_t0, addr_incr_two_t0 };
assign _049_ = instr_addr_q & _025_;
assign _050_ = { 29'h00000000, _198_, addr_incr_two } & _026_;
assign _193_ = _049_ + _050_;
assign _160_ = instr_addr_q | instr_addr_q_t0;
assign _161_ = { 29'h00000000, _198_, addr_incr_two } | { 29'h00000000, addr_incr_two_t0, addr_incr_two_t0 };
assign _194_ = _160_ + _161_;
assign _192_ = _193_ ^ _194_;
assign _162_ = _192_ | instr_addr_q_t0;
assign instr_addr_next_t0 = _162_ | { 29'h00000000, addr_incr_two_t0, addr_incr_two_t0 };
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME valid_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) valid_q_t0 <= 3'h0;
else valid_q_t0 <= valid_d_t0;
assign _027_ = ~ entry_en[2];
assign _028_ = ~ entry_en[1];
assign _029_ = ~ entry_en[0];
assign _030_ = ~ instr_addr_en;
assign _096_ = entry_en[2] & in_err_i_t0;
assign _098_ = { entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2] } & in_rdata_i_t0;
assign _100_ = entry_en[1] & err_d_t0[1];
assign _102_ = { entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1] } & rdata_d_t0[63:32];
assign _104_ = entry_en[0] & err_d_t0[0];
assign _106_ = { entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0] } & rdata_d_t0[31:0];
assign _108_ = { instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en } & instr_addr_d_t0;
assign _097_ = _027_ & err_q_t0[2];
assign _099_ = { _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_ } & rdata_q_t0[95:64];
assign _101_ = _028_ & err_q_t0[1];
assign _103_ = { _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_, _028_ } & rdata_q_t0[63:32];
assign _105_ = _029_ & err_q_t0[0];
assign _107_ = { _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_, _029_ } & rdata_q_t0[31:0];
assign _109_ = { _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_, _030_ } & instr_addr_q_t0;
assign _178_ = _096_ | _097_;
assign _179_ = _098_ | _099_;
assign _180_ = _100_ | _101_;
assign _181_ = _102_ | _103_;
assign _182_ = _104_ | _105_;
assign _183_ = _106_ | _107_;
assign _184_ = _108_ | _109_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q_t0[2] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q_t0[2] <= 1'h0;
else err_q_t0[2] <= _178_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q_t0[95:64] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q_t0[95:64] <= 32'd0;
else rdata_q_t0[95:64] <= _179_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q_t0[1] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q_t0[1] <= 1'h0;
else err_q_t0[1] <= _180_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q_t0[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q_t0[63:32] <= 32'd0;
else rdata_q_t0[63:32] <= _181_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q_t0[0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q_t0[0] <= 1'h0;
else err_q_t0[0] <= _182_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q_t0[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q_t0[31:0] <= 32'd0;
else rdata_q_t0[31:0] <= _183_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME instr_addr_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_addr_q_t0 <= 31'h00000000;
else instr_addr_q_t0 <= _184_;
assign _051_ = err_q_t0[1] & _031_;
assign _054_ = valid_q_t0[0] & err_q[0];
assign _057_ = in_err_i_t0 & _202_;
assign _060_ = err_q_t0[1] & _047_;
assign _063_ = in_err_i_t0 & valid_q[0];
assign _066_ = _011_ & _047_;
assign _069_ = valid_q_t0[0] & in_valid_i;
assign _072_ = valid_q_t0[1] & valid_q[0];
assign _075_ = valid_popped_t0[0] & _043_;
assign _078_ = valid_popped_t0[1] & _043_;
assign _081_ = valid_pushed_t0[1] & pop_fifo;
assign _082_ = in_valid_i_t0 & lowest_free_entry[0];
assign _083_ = valid_pushed_t0[2] & pop_fifo;
assign _084_ = in_valid_i_t0 & lowest_free_entry[1];
assign _087_ = valid_q_t0[2] & valid_q[1];
assign _090_ = valid_popped_t0[2] & _043_;
assign _093_ = in_valid_i_t0 & lowest_free_entry[2];
assign _052_ = unaligned_is_compressed_t0 & err_q[1];
assign _055_ = err_q_t0[0] & valid_q[0];
assign _058_ = _203_ & in_err_i;
assign _061_ = err_q_t0[0] & err_q[1];
assign _064_ = valid_q_t0[0] & in_err_i;
assign _067_ = err_q_t0[0] & _010_;
assign _070_ = in_valid_i_t0 & valid_q[0];
assign unaligned_is_compressed_t0 = err_t0 & _195_;
assign aligned_is_compressed_t0 = err_t0 & _196_;
assign _073_ = valid_q_t0[0] & _036_;
assign _076_ = clear_i_t0 & valid_popped[0];
assign _079_ = clear_i_t0 & valid_popped[1];
assign _085_ = lowest_free_entry_t0[1] & in_valid_i;
assign _088_ = valid_q_t0[1] & _040_;
assign _091_ = clear_i_t0 & valid_popped[2];
assign _094_ = lowest_free_entry_t0[2] & in_valid_i;
assign _053_ = err_q_t0[1] & unaligned_is_compressed_t0;
assign _056_ = valid_q_t0[0] & err_q_t0[0];
assign _059_ = in_err_i_t0 & _203_;
assign _062_ = err_q_t0[1] & err_q_t0[0];
assign _065_ = in_err_i_t0 & valid_q_t0[0];
assign _068_ = _011_ & err_q_t0[0];
assign _071_ = valid_q_t0[0] & in_valid_i_t0;
assign _074_ = valid_q_t0[1] & valid_q_t0[0];
assign _077_ = valid_popped_t0[0] & clear_i_t0;
assign _080_ = valid_popped_t0[1] & clear_i_t0;
assign _086_ = in_valid_i_t0 & lowest_free_entry_t0[1];
assign _089_ = valid_q_t0[2] & valid_q_t0[1];
assign _092_ = valid_popped_t0[2] & clear_i_t0;
assign _095_ = in_valid_i_t0 & lowest_free_entry_t0[2];
assign _163_ = _051_ | _052_;
assign _164_ = _054_ | _055_;
assign _165_ = _057_ | _058_;
assign _166_ = _060_ | _061_;
assign _167_ = _063_ | _064_;
assign _168_ = _066_ | _067_;
assign _169_ = _069_ | _070_;
assign _170_ = _072_ | _073_;
assign _171_ = _075_ | _076_;
assign _172_ = _078_ | _079_;
assign _173_ = _082_ | _069_;
assign _174_ = _084_ | _085_;
assign _175_ = _087_ | _088_;
assign _176_ = _090_ | _091_;
assign _177_ = _093_ | _094_;
assign _003_ = _163_ | _053_;
assign _005_ = _164_ | _056_;
assign _007_ = _165_ | _059_;
assign _009_ = _166_ | _062_;
assign _011_ = _167_ | _065_;
assign _013_ = _168_ | _068_;
assign _015_ = _169_ | _071_;
assign lowest_free_entry_t0[1] = _170_ | _074_;
assign valid_d_t0[0] = _171_ | _077_;
assign valid_d_t0[1] = _172_ | _080_;
assign _018_ = _173_ | _071_;
assign _020_ = _174_ | _086_;
assign lowest_free_entry_t0[2] = _175_ | _089_;
assign valid_d_t0[2] = _176_ | _092_;
assign entry_en_t0[2] = _177_ | _095_;
/* src = "generated/sv2v_out.v:16262.5-16270.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q[2] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q[2] <= 1'h0;
else if (entry_en[2]) err_q[2] <= in_err_i;
/* src = "generated/sv2v_out.v:16262.5-16270.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q[95:64] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q[95:64] <= 32'd0;
else if (entry_en[2]) rdata_q[95:64] <= in_rdata_i;
/* src = "generated/sv2v_out.v:16262.5-16270.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q[1] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q[1] <= 1'h0;
else if (entry_en[1]) err_q[1] <= err_d[1];
/* src = "generated/sv2v_out.v:16262.5-16270.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q[63:32] <= 32'd0;
else if (entry_en[1]) rdata_q[63:32] <= rdata_d[63:32];
/* src = "generated/sv2v_out.v:16262.5-16270.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q[0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q[0] <= 1'h0;
else if (entry_en[0]) err_q[0] <= err_d[0];
/* src = "generated/sv2v_out.v:16262.5-16270.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q[31:0] <= 32'd0;
else if (entry_en[0]) rdata_q[31:0] <= rdata_d[31:0];
/* src = "generated/sv2v_out.v:16214.4-16218.35" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME instr_addr_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_addr_q <= 31'h00000000;
else if (instr_addr_en) instr_addr_q <= instr_addr_d;
assign _031_ = ~ unaligned_is_compressed;
assign _032_ = ~ instr_addr_q[1];
assign _033_ = ~ { instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1] };
assign _034_ = ~ { valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0] };
assign lowest_free_entry[0] = ~ valid_q[0];
assign _035_ = ~ { valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1] };
assign _036_ = ~ valid_q[1];
assign _037_ = ~ { clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i };
assign _038_ = ~ pop_fifo;
assign _039_ = ~ { valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2] };
assign _040_ = ~ valid_q[2];
assign _130_ = _031_ & valid_unaligned_t0;
assign _132_ = _032_ & valid_t0;
assign _134_ = _032_ & err_t0;
assign _136_ = _033_ & rdata_t0;
assign _138_ = _034_ & in_rdata_i_t0;
assign _140_ = lowest_free_entry[0] & in_err_i_t0;
assign _141_ = _035_ & { in_rdata_i_t0[15:0], rdata_t0[31:16] };
assign _143_ = _036_ & _205_;
assign _145_ = _036_ & _013_;
assign valid_unaligned_t0 = _036_ & _015_;
assign _120_ = _032_ & aligned_is_compressed_t0;
assign _148_ = _037_ & instr_addr_next_t0;
assign _150_ = _038_ & valid_pushed_t0[0];
assign _151_ = _038_ & valid_pushed_t0[1];
assign _152_ = _035_ & in_rdata_i_t0;
assign _154_ = _039_ & in_rdata_i_t0;
assign _156_ = _036_ & in_err_i_t0;
assign _158_ = _040_ & in_err_i_t0;
assign valid_popped_t0[2] = _038_ & valid_pushed_t0[2];
assign _131_ = unaligned_is_compressed & valid_t0;
assign _133_ = instr_addr_q[1] & _001_;
assign out_err_plus2_o_t0 = instr_addr_q[1] & err_plus2_t0;
assign _135_ = instr_addr_q[1] & err_unaligned_t0;
assign _137_ = { instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1] } & rdata_unaligned_t0;
assign _139_ = { valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0] } & rdata_q_t0[31:0];
assign _142_ = { valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1] } & { rdata_q_t0[47:32], rdata_t0[31:16] };
assign _144_ = valid_q[1] & _201_;
assign _146_ = valid_q[1] & _009_;
assign _147_ = instr_addr_q[1] & unaligned_is_compressed_t0;
assign _149_ = { clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i } & in_addr_i_t0[31:1];
assign _153_ = { valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1] } & rdata_q_t0[63:32];
assign _155_ = { valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2] } & rdata_q_t0[95:64];
assign _157_ = valid_q[1] & err_q_t0[1];
assign _159_ = valid_q[2] & err_q_t0[2];
assign _001_ = _130_ | _131_;
assign out_valid_o_t0 = _132_ | _133_;
assign out_err_o_t0 = _134_ | _135_;
assign out_rdata_o_t0 = _136_ | _137_;
assign rdata_t0 = _138_ | _139_;
assign err_t0 = _140_ | _055_;
assign rdata_unaligned_t0 = _141_ | _142_;
assign err_unaligned_t0 = _143_ | _144_;
assign err_plus2_t0 = _145_ | _146_;
assign addr_incr_two_t0 = _120_ | _147_;
assign instr_addr_d_t0 = _148_ | _149_;
assign valid_popped_t0[0] = _150_ | _081_;
assign valid_popped_t0[1] = _151_ | _083_;
assign rdata_d_t0[31:0] = _152_ | _153_;
assign rdata_d_t0[63:32] = _154_ | _155_;
assign err_d_t0[0] = _156_ | _157_;
assign err_d_t0[1] = _158_ | _159_;
assign _041_ = ~ _002_;
assign _042_ = ~ _004_;
assign _043_ = ~ clear_i;
assign _044_ = ~ _017_;
assign _045_ = ~ _019_;
assign _046_ = ~ in_valid_i;
assign _047_ = ~ err_q[0];
assign _048_ = ~ _006_;
assign _110_ = valid_q_t0[0] & _046_;
assign _111_ = _003_ & _047_;
assign _114_ = valid_q_t0[0] & unaligned_is_compressed;
assign _117_ = _005_ & _048_;
assign _121_ = _018_ & lowest_free_entry[0];
assign _124_ = _020_ & _036_;
assign _127_ = valid_q_t0[2] & _027_;
assign _112_ = err_q_t0[0] & _041_;
assign _115_ = unaligned_is_compressed_t0 & valid_q[0];
assign _118_ = _007_ & _042_;
assign _122_ = valid_q_t0[0] & _044_;
assign _125_ = valid_q_t0[1] & _045_;
assign _128_ = entry_en_t0[2] & _040_;
assign _113_ = _003_ & err_q_t0[0];
assign _116_ = valid_q_t0[0] & unaligned_is_compressed_t0;
assign _119_ = _005_ & _007_;
assign _123_ = _018_ & valid_q_t0[0];
assign _126_ = _020_ & valid_q_t0[1];
assign _129_ = valid_q_t0[2] & entry_en_t0[2];
assign _185_ = _110_ | _082_;
assign _186_ = _111_ | _112_;
assign _187_ = _114_ | _115_;
assign _188_ = _117_ | _118_;
assign _189_ = _121_ | _122_;
assign _190_ = _124_ | _125_;
assign _191_ = _127_ | _128_;
assign valid_t0 = _185_ | _071_;
assign _201_ = _186_ | _113_;
assign _203_ = _187_ | _116_;
assign _205_ = _188_ | _119_;
assign valid_pushed_t0[0] = _189_ | _123_;
assign valid_pushed_t0[1] = _190_ | _126_;
assign valid_pushed_t0[2] = _191_ | _129_;
assign _195_ = rdata[17:16] != /* src = "generated/sv2v_out.v:16190.36-16190.57" */ 2'h3;
assign _196_ = rdata[1:0] != /* src = "generated/sv2v_out.v:16191.34-16191.53" */ 2'h3;
assign _197_ = ~ /* src = "generated/sv2v_out.v:16191.57-16191.61" */ err;
assign _198_ = ~ /* src = "generated/sv2v_out.v:16210.56-16210.70" */ addr_incr_two;
assign _199_ = ~ /* src = "generated/sv2v_out.v:16229.51-16229.73" */ aligned_is_compressed;
assign valid = valid_q[0] | /* src = "generated/sv2v_out.v:16185.17-16185.40" */ in_valid_i;
assign _200_ = _002_ | /* src = "generated/sv2v_out.v:16187.39-16187.87" */ err_q[0];
assign _202_ = lowest_free_entry[0] | /* src = "generated/sv2v_out.v:16187.129-16187.167" */ _031_;
assign _204_ = _004_ | /* src = "generated/sv2v_out.v:16187.90-16187.169" */ _006_;
assign instr_addr_en = clear_i | /* src = "generated/sv2v_out.v:16208.25-16208.62" */ _016_;
assign _206_ = _199_ | /* src = "generated/sv2v_out.v:16229.51-16229.89" */ instr_addr_q[1];
assign valid_pushed[0] = _017_ | /* src = "generated/sv2v_out.v:16239.29-16239.77" */ valid_q[0];
assign valid_pushed[1] = _019_ | /* src = "generated/sv2v_out.v:16239.29-16239.77" */ valid_q[1];
assign entry_en[0] = _021_ | /* src = "generated/sv2v_out.v:16242.25-16242.109" */ _022_;
assign entry_en[1] = _023_ | /* src = "generated/sv2v_out.v:16242.25-16242.109" */ _024_;
assign valid_pushed[2] = valid_q[2] | /* src = "generated/sv2v_out.v:16248.35-16248.99" */ entry_en[2];
/* src = "generated/sv2v_out.v:16254.2-16258.23" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME valid_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) valid_q <= 3'h0;
else valid_q <= valid_d;
assign _000_ = unaligned_is_compressed ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:16197.8-16197.31|generated/sv2v_out.v:16197.4-16200.35" */ valid : valid_unaligned;
assign out_valid_o = instr_addr_q[1] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:16193.7-16193.20|generated/sv2v_out.v:16193.3-16207.6" */ _000_ : valid;
assign out_err_plus2_o = instr_addr_q[1] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:16193.7-16193.20|generated/sv2v_out.v:16193.3-16207.6" */ err_plus2 : 1'h0;
assign out_err_o = instr_addr_q[1] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:16193.7-16193.20|generated/sv2v_out.v:16193.3-16207.6" */ err_unaligned : err;
assign out_rdata_o = instr_addr_q[1] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:16193.7-16193.20|generated/sv2v_out.v:16193.3-16207.6" */ rdata_unaligned : rdata;
assign rdata = valid_q[0] ? /* src = "generated/sv2v_out.v:16183.18-16183.58" */ rdata_q[31:0] : in_rdata_i;
assign err = valid_q[0] ? /* src = "generated/sv2v_out.v:16184.16-16184.48" */ err_q[0] : in_err_i;
assign rdata_unaligned = valid_q[1] ? /* src = "generated/sv2v_out.v:16186.28-16186.107" */ { rdata_q[47:32], rdata[31:16] } : { in_rdata_i[15:0], rdata[31:16] };
assign err_unaligned = valid_q[1] ? /* src = "generated/sv2v_out.v:16187.26-16187.169" */ _200_ : _204_;
assign err_plus2 = valid_q[1] ? /* src = "generated/sv2v_out.v:16188.22-16188.93" */ _008_ : _012_;
assign valid_unaligned = valid_q[1] ? /* src = "generated/sv2v_out.v:16189.28-16189.71" */ 1'h1 : _014_;
assign addr_incr_two = instr_addr_q[1] ? /* src = "generated/sv2v_out.v:16209.26-16209.91" */ unaligned_is_compressed : aligned_is_compressed;
assign instr_addr_d = clear_i ? /* src = "generated/sv2v_out.v:16211.25-16211.68" */ in_addr_i[31:1] : instr_addr_next;
assign valid_popped[0] = pop_fifo ? /* src = "generated/sv2v_out.v:16240.30-16240.78" */ valid_pushed[1] : valid_pushed[0];
assign valid_popped[1] = pop_fifo ? /* src = "generated/sv2v_out.v:16240.30-16240.78" */ valid_pushed[2] : valid_pushed[1];
assign rdata_d[31:0] = valid_q[1] ? /* src = "generated/sv2v_out.v:16243.34-16243.89" */ rdata_q[63:32] : in_rdata_i;
assign rdata_d[63:32] = valid_q[2] ? /* src = "generated/sv2v_out.v:16243.34-16243.89" */ rdata_q[95:64] : in_rdata_i;
assign err_d[0] = valid_q[1] ? /* src = "generated/sv2v_out.v:16244.23-16244.63" */ err_q[1] : in_err_i;
assign err_d[1] = valid_q[2] ? /* src = "generated/sv2v_out.v:16244.23-16244.63" */ err_q[2] : in_err_i;
assign valid_popped[2] = pop_fifo ? /* src = "generated/sv2v_out.v:16249.36-16249.77" */ 1'h0 : valid_pushed[2];
assign busy_o = valid_q[2:1];
assign busy_o_t0 = valid_q_t0[2:1];
assign err_d[2] = in_err_i;
assign err_d_t0[2] = in_err_i_t0;
assign lowest_free_entry_t0[0] = valid_q_t0[0];
assign out_addr_o = { instr_addr_q, 1'h0 };
assign out_addr_o_t0 = { instr_addr_q_t0, 1'h0 };
assign rdata_d[95:64] = in_rdata_i;
assign rdata_d_t0[95:64] = in_rdata_i_t0;
endmodule

module \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111 (clk_i, rst_ni, data_req_o, data_gnt_i, data_rvalid_i, data_bus_err_i, data_pmp_err_i, data_addr_o, data_we_o, data_be_o, data_wdata_o, data_rdata_i, lsu_we_i, lsu_type_i, lsu_wdata_i, lsu_sign_ext_i, lsu_rdata_o, lsu_rdata_valid_o, lsu_req_i, adder_result_ex_i, addr_incr_req_o
, addr_last_o, lsu_req_done_o, lsu_resp_valid_o, load_err_o, load_resp_intg_err_o, store_err_o, store_resp_intg_err_o, busy_o, perf_load_o, perf_store_o, data_we_o_t0, data_req_o_t0, busy_o_t0, adder_result_ex_i_t0, addr_incr_req_o_t0, addr_last_o_t0, data_addr_o_t0, data_be_o_t0, data_bus_err_i_t0, data_gnt_i_t0, data_pmp_err_i_t0
, data_rdata_i_t0, data_rvalid_i_t0, data_wdata_o_t0, load_err_o_t0, load_resp_intg_err_o_t0, lsu_rdata_o_t0, lsu_rdata_valid_o_t0, lsu_req_done_o_t0, lsu_req_i_t0, lsu_resp_valid_o_t0, lsu_sign_ext_i_t0, lsu_type_i_t0, lsu_wdata_i_t0, lsu_we_i_t0, perf_load_o_t0, perf_store_o_t0, store_err_o_t0, store_resp_intg_err_o_t0);
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _000_;
/* src = "generated/sv2v_out.v:18472.2-18511.10" */
wire [3:0] _001_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _002_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _003_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire [2:0] _004_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _005_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _007_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _008_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _009_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _010_;
/* src = "generated/sv2v_out.v:18576.2-18599.10" */
wire [31:0] _011_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18576.2-18599.10" */
wire [31:0] _012_;
/* src = "generated/sv2v_out.v:18552.2-18575.10" */
wire [31:0] _013_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18552.2-18575.10" */
wire [31:0] _014_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _015_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _016_;
/* src = "generated/sv2v_out.v:18472.2-18511.10" */
wire [3:0] _017_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _018_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire [2:0] _019_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _021_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _022_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _023_;
/* src = "generated/sv2v_out.v:18576.2-18599.10" */
wire [31:0] _024_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18576.2-18599.10" */
wire [31:0] _025_;
/* src = "generated/sv2v_out.v:18552.2-18575.10" */
wire [31:0] _026_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18552.2-18575.10" */
wire [31:0] _027_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _028_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _029_;
/* src = "generated/sv2v_out.v:18472.2-18511.10" */
wire [3:0] _030_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _031_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire [2:0] _032_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _033_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _034_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _035_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _036_;
/* src = "generated/sv2v_out.v:18576.2-18599.10" */
wire [31:0] _037_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18576.2-18599.10" */
wire [31:0] _038_;
/* src = "generated/sv2v_out.v:18552.2-18575.10" */
wire [31:0] _039_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18552.2-18575.10" */
wire [31:0] _040_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _041_;
/* src = "generated/sv2v_out.v:18472.2-18511.10" */
wire [3:0] _042_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _043_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _044_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire [2:0] _045_;
/* src = "generated/sv2v_out.v:18576.2-18599.10" */
wire [31:0] _046_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18576.2-18599.10" */
wire [31:0] _047_;
/* src = "generated/sv2v_out.v:18552.2-18575.10" */
wire [31:0] _048_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18552.2-18575.10" */
wire [31:0] _049_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _050_;
/* src = "generated/sv2v_out.v:18472.2-18511.10" */
wire [3:0] _051_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _052_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire [2:0] _053_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _054_;
/* src = "generated/sv2v_out.v:18472.2-18511.10" */
wire [3:0] _055_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire _056_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire [2:0] _057_;
/* src = "generated/sv2v_out.v:18626.2-18704.5" */
wire [2:0] _058_;
/* src = "generated/sv2v_out.v:18674.20-18674.62" */
wire _059_;
/* src = "generated/sv2v_out.v:18721.32-18721.67" */
wire _060_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18721.32-18721.67" */
wire _061_;
/* src = "generated/sv2v_out.v:18721.31-18721.87" */
wire _062_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18721.31-18721.87" */
wire _063_;
/* src = "generated/sv2v_out.v:18721.30-18721.101" */
wire _064_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18721.30-18721.101" */
wire _065_;
/* src = "generated/sv2v_out.v:18739.23-18739.51" */
wire _066_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18739.23-18739.51" */
wire _067_;
/* src = "generated/sv2v_out.v:18740.24-18740.51" */
wire _068_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18740.24-18740.51" */
wire _069_;
/* src = "generated/sv2v_out.v:18741.33-18741.62" */
wire _070_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18741.33-18741.62" */
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire [31:0] _082_;
wire [31:0] _083_;
wire [31:0] _084_;
wire [31:0] _085_;
wire [31:0] _086_;
wire [31:0] _087_;
wire [31:0] _088_;
wire [31:0] _089_;
wire _090_;
wire _091_;
wire [31:0] _092_;
wire [31:0] _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire [23:0] _143_;
wire [23:0] _144_;
wire [31:0] _145_;
wire [31:0] _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire [31:0] _153_;
wire [31:0] _154_;
wire [31:0] _155_;
wire [31:0] _156_;
wire [31:0] _157_;
wire [31:0] _158_;
wire [31:0] _159_;
wire [31:0] _160_;
wire [31:0] _161_;
wire [31:0] _162_;
wire [31:0] _163_;
wire [31:0] _164_;
wire [31:0] _165_;
wire [31:0] _166_;
wire [31:0] _167_;
wire [31:0] _168_;
wire [31:0] _169_;
wire [31:0] _170_;
wire [31:0] _171_;
wire [31:0] _172_;
wire [31:0] _173_;
wire [31:0] _174_;
wire [31:0] _175_;
wire [31:0] _176_;
wire [31:0] _177_;
wire [31:0] _178_;
wire [31:0] _179_;
wire [31:0] _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire [31:0] _193_;
wire [31:0] _194_;
wire [31:0] _195_;
wire [31:0] _196_;
wire [31:0] _197_;
wire [31:0] _198_;
wire [31:0] _199_;
wire [31:0] _200_;
wire [31:0] _201_;
wire [31:0] _202_;
wire [31:0] _203_;
wire [31:0] _204_;
wire [31:0] _205_;
wire [31:0] _206_;
wire [31:0] _207_;
wire [31:0] _208_;
wire [31:0] _209_;
wire [31:0] _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire _221_;
wire _222_;
wire _223_;
wire _224_;
wire _225_;
wire [23:0] _226_;
wire [31:0] _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire [2:0] _232_;
wire [2:0] _233_;
wire [2:0] _234_;
wire [2:0] _235_;
wire _236_;
/* cellift = 32'd1 */
wire _237_;
wire _238_;
/* cellift = 32'd1 */
wire _239_;
wire _240_;
/* cellift = 32'd1 */
wire _241_;
wire _242_;
wire _243_;
wire _244_;
wire _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
/* cellift = 32'd1 */
wire _250_;
wire [31:0] _251_;
/* cellift = 32'd1 */
wire [31:0] _252_;
wire [31:0] _253_;
/* cellift = 32'd1 */
wire [31:0] _254_;
wire [31:0] _255_;
/* cellift = 32'd1 */
wire [31:0] _256_;
wire [31:0] _257_;
/* cellift = 32'd1 */
wire [31:0] _258_;
wire [31:0] _259_;
/* cellift = 32'd1 */
wire [31:0] _260_;
wire [31:0] _261_;
/* cellift = 32'd1 */
wire [31:0] _262_;
wire [31:0] _263_;
/* cellift = 32'd1 */
wire [31:0] _264_;
wire [31:0] _265_;
/* cellift = 32'd1 */
wire [31:0] _266_;
wire [31:0] _267_;
/* cellift = 32'd1 */
wire [31:0] _268_;
wire [3:0] _269_;
wire [3:0] _270_;
wire [3:0] _271_;
wire [3:0] _272_;
wire [3:0] _273_;
wire [3:0] _274_;
wire [3:0] _275_;
wire [3:0] _276_;
/* src = "generated/sv2v_out.v:18625.37-18625.56" */
wire _277_;
/* src = "generated/sv2v_out.v:18625.90-18625.109" */
wire _278_;
/* src = "generated/sv2v_out.v:18625.115-18625.135" */
wire _279_;
/* src = "generated/sv2v_out.v:18705.63-18705.80" */
wire _280_;
/* src = "generated/sv2v_out.v:18720.59-18720.76" */
wire _281_;
/* src = "generated/sv2v_out.v:18625.36-18625.83" */
wire _282_;
/* src = "generated/sv2v_out.v:18625.89-18625.136" */
wire _283_;
/* src = "generated/sv2v_out.v:18659.9-18659.32" */
wire _284_;
/* src = "generated/sv2v_out.v:18669.9-18669.35" */
wire _285_;
/* src = "generated/sv2v_out.v:18625.62-18625.82" */
wire _286_;
/* src = "generated/sv2v_out.v:18645.20-18645.29" */
wire _287_;
/* src = "generated/sv2v_out.v:18672.21-18672.31" */
wire _288_;
/* src = "generated/sv2v_out.v:18674.33-18674.62" */
wire _289_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18674.33-18674.62" */
wire _290_;
/* src = "generated/sv2v_out.v:18721.71-18721.87" */
wire _291_;
/* src = "generated/sv2v_out.v:18721.105-18721.119" */
wire _292_;
/* src = "generated/sv2v_out.v:18671.18-18671.44" */
wire _293_;
/* src = "generated/sv2v_out.v:18705.27-18705.58" */
wire _294_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18705.27-18705.58" */
wire _295_;
/* src = "generated/sv2v_out.v:18719.28-18719.54" */
wire _296_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18719.28-18719.54" */
wire _297_;
/* src = "generated/sv2v_out.v:18720.29-18720.54" */
wire _298_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18720.29-18720.54" */
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire [1:0] _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire [1:0] _312_;
wire _313_;
/* src = "generated/sv2v_out.v:18651.20-18651.57" */
wire [2:0] _314_;
/* src = "generated/sv2v_out.v:18654.20-18654.57" */
wire [2:0] _315_;
/* src = "generated/sv2v_out.v:18673.19-18673.43" */
wire [2:0] _316_;
/* src = "generated/sv2v_out.v:18428.20-18428.37" */
input [31:0] adder_result_ex_i;
wire [31:0] adder_result_ex_i;
/* cellift = 32'd1 */
input [31:0] adder_result_ex_i_t0;
wire [31:0] adder_result_ex_i_t0;
/* src = "generated/sv2v_out.v:18429.13-18429.28" */
output addr_incr_req_o;
wire addr_incr_req_o;
/* cellift = 32'd1 */
output addr_incr_req_o_t0;
wire addr_incr_req_o_t0;
/* src = "generated/sv2v_out.v:18443.14-18443.25" */
wire [31:0] addr_last_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18443.14-18443.25" */
wire [31:0] addr_last_d_t0;
/* src = "generated/sv2v_out.v:18430.21-18430.32" */
output [31:0] addr_last_o;
reg [31:0] addr_last_o;
/* cellift = 32'd1 */
output [31:0] addr_last_o_t0;
reg [31:0] addr_last_o_t0;
/* src = "generated/sv2v_out.v:18444.6-18444.17" */
wire addr_update;
/* src = "generated/sv2v_out.v:18437.14-18437.20" */
output busy_o;
wire busy_o;
/* cellift = 32'd1 */
output busy_o_t0;
wire busy_o_t0;
/* src = "generated/sv2v_out.v:18409.13-18409.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:18445.6-18445.17" */
wire ctrl_update;
/* src = "generated/sv2v_out.v:18416.21-18416.32" */
output [31:0] data_addr_o;
wire [31:0] data_addr_o;
/* cellift = 32'd1 */
output [31:0] data_addr_o_t0;
wire [31:0] data_addr_o_t0;
/* src = "generated/sv2v_out.v:18418.20-18418.29" */
output [3:0] data_be_o;
wire [3:0] data_be_o;
/* cellift = 32'd1 */
output [3:0] data_be_o_t0;
wire [3:0] data_be_o_t0;
/* src = "generated/sv2v_out.v:18414.13-18414.27" */
input data_bus_err_i;
wire data_bus_err_i;
/* cellift = 32'd1 */
input data_bus_err_i_t0;
wire data_bus_err_i_t0;
/* src = "generated/sv2v_out.v:18412.13-18412.23" */
input data_gnt_i;
wire data_gnt_i;
/* cellift = 32'd1 */
input data_gnt_i_t0;
wire data_gnt_i_t0;
/* src = "generated/sv2v_out.v:18466.7-18466.20" */
wire data_intg_err;
/* src = "generated/sv2v_out.v:18467.7-18467.22" */
wire data_or_pmp_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18467.7-18467.22" */
wire data_or_pmp_err_t0;
/* src = "generated/sv2v_out.v:18415.13-18415.27" */
input data_pmp_err_i;
wire data_pmp_err_i;
/* cellift = 32'd1 */
input data_pmp_err_i_t0;
wire data_pmp_err_i_t0;
/* src = "generated/sv2v_out.v:18420.34-18420.46" */
input [38:0] data_rdata_i;
wire [38:0] data_rdata_i;
/* cellift = 32'd1 */
input [38:0] data_rdata_i_t0;
wire [38:0] data_rdata_i_t0;
/* src = "generated/sv2v_out.v:18411.13-18411.23" */
output data_req_o;
wire data_req_o;
/* cellift = 32'd1 */
output data_req_o_t0;
wire data_req_o_t0;
/* src = "generated/sv2v_out.v:18413.13-18413.26" */
input data_rvalid_i;
wire data_rvalid_i;
/* cellift = 32'd1 */
input data_rvalid_i_t0;
wire data_rvalid_i_t0;
/* src = "generated/sv2v_out.v:18450.6-18450.21" */
reg data_sign_ext_q;
/* src = "generated/sv2v_out.v:18449.12-18449.23" */
reg [1:0] data_type_q;
/* src = "generated/sv2v_out.v:18454.13-18454.23" */
wire [31:0] data_wdata;
/* src = "generated/sv2v_out.v:18419.35-18419.47" */
output [38:0] data_wdata_o;
wire [38:0] data_wdata_o;
/* cellift = 32'd1 */
output [38:0] data_wdata_o_t0;
wire [38:0] data_wdata_o_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18454.13-18454.23" */
wire [31:0] data_wdata_t0;
/* src = "generated/sv2v_out.v:18417.14-18417.23" */
output data_we_o;
wire data_we_o;
/* cellift = 32'd1 */
output data_we_o_t0;
wire data_we_o_t0;
/* src = "generated/sv2v_out.v:18451.6-18451.15" */
reg data_we_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18451.6-18451.15" */
reg data_we_q_t0;
/* src = "generated/sv2v_out.v:18610.30-18610.44" */
wire [38:0] \g_mem_rdata_ecc.data_rdata_buf ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18610.30-18610.44" */
wire [38:0] \g_mem_rdata_ecc.data_rdata_buf_t0 ;
/* src = "generated/sv2v_out.v:18609.15-18609.22" */
wire [1:0] \g_mem_rdata_ecc.ecc_err ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18609.15-18609.22" */
/* unused_bits = "0 1" */
wire [1:0] \g_mem_rdata_ecc.ecc_err_t0 ;
/* src = "generated/sv2v_out.v:18461.6-18461.25" */
wire handle_misaligned_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18461.6-18461.25" */
wire handle_misaligned_d_t0;
/* src = "generated/sv2v_out.v:18460.6-18460.25" */
reg handle_misaligned_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18460.6-18460.25" */
reg handle_misaligned_q_t0;
/* src = "generated/sv2v_out.v:18433.14-18433.24" */
output load_err_o;
wire load_err_o;
/* cellift = 32'd1 */
output load_err_o_t0;
wire load_err_o_t0;
/* src = "generated/sv2v_out.v:18434.14-18434.34" */
output load_resp_intg_err_o;
wire load_resp_intg_err_o;
/* cellift = 32'd1 */
output load_resp_intg_err_o_t0;
wire load_resp_intg_err_o_t0;
/* src = "generated/sv2v_out.v:18468.12-18468.21" */
reg [2:0] ls_fsm_cs;
/* src = "generated/sv2v_out.v:18469.12-18469.21" */
wire [2:0] ls_fsm_ns;
/* src = "generated/sv2v_out.v:18465.6-18465.15" */
wire lsu_err_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18465.6-18465.15" */
wire lsu_err_d_t0;
/* src = "generated/sv2v_out.v:18464.6-18464.15" */
reg lsu_err_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18464.6-18464.15" */
reg lsu_err_q_t0;
/* src = "generated/sv2v_out.v:18425.21-18425.32" */
output [31:0] lsu_rdata_o;
wire [31:0] lsu_rdata_o;
/* cellift = 32'd1 */
output [31:0] lsu_rdata_o_t0;
wire [31:0] lsu_rdata_o_t0;
/* src = "generated/sv2v_out.v:18426.14-18426.31" */
output lsu_rdata_valid_o;
wire lsu_rdata_valid_o;
/* cellift = 32'd1 */
output lsu_rdata_valid_o_t0;
wire lsu_rdata_valid_o_t0;
/* src = "generated/sv2v_out.v:18431.14-18431.28" */
output lsu_req_done_o;
wire lsu_req_done_o;
/* cellift = 32'd1 */
output lsu_req_done_o_t0;
wire lsu_req_done_o_t0;
/* src = "generated/sv2v_out.v:18427.13-18427.22" */
input lsu_req_i;
wire lsu_req_i;
/* cellift = 32'd1 */
input lsu_req_i_t0;
wire lsu_req_i_t0;
/* src = "generated/sv2v_out.v:18432.14-18432.30" */
output lsu_resp_valid_o;
wire lsu_resp_valid_o;
/* cellift = 32'd1 */
output lsu_resp_valid_o_t0;
wire lsu_resp_valid_o_t0;
/* src = "generated/sv2v_out.v:18424.13-18424.27" */
input lsu_sign_ext_i;
wire lsu_sign_ext_i;
/* cellift = 32'd1 */
input lsu_sign_ext_i_t0;
wire lsu_sign_ext_i_t0;
/* src = "generated/sv2v_out.v:18422.19-18422.29" */
input [1:0] lsu_type_i;
wire [1:0] lsu_type_i;
/* cellift = 32'd1 */
input [1:0] lsu_type_i_t0;
wire [1:0] lsu_type_i_t0;
/* src = "generated/sv2v_out.v:18423.20-18423.31" */
input [31:0] lsu_wdata_i;
wire [31:0] lsu_wdata_i;
/* cellift = 32'd1 */
input [31:0] lsu_wdata_i_t0;
wire [31:0] lsu_wdata_i_t0;
/* src = "generated/sv2v_out.v:18421.13-18421.21" */
input lsu_we_i;
wire lsu_we_i;
/* cellift = 32'd1 */
input lsu_we_i_t0;
wire lsu_we_i_t0;
/* src = "generated/sv2v_out.v:18438.13-18438.24" */
output perf_load_o;
wire perf_load_o;
/* cellift = 32'd1 */
output perf_load_o_t0;
wire perf_load_o_t0;
/* src = "generated/sv2v_out.v:18439.13-18439.25" */
output perf_store_o;
wire perf_store_o;
/* cellift = 32'd1 */
output perf_store_o_t0;
wire perf_store_o_t0;
/* src = "generated/sv2v_out.v:18463.6-18463.15" */
wire pmp_err_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18463.6-18463.15" */
wire pmp_err_d_t0;
/* src = "generated/sv2v_out.v:18462.6-18462.15" */
reg pmp_err_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18462.6-18462.15" */
reg pmp_err_q_t0;
/* src = "generated/sv2v_out.v:18458.13-18458.24" */
wire [31:0] rdata_b_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18458.13-18458.24" */
wire [31:0] rdata_b_ext_t0;
/* src = "generated/sv2v_out.v:18457.13-18457.24" */
wire [31:0] rdata_h_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18457.13-18457.24" */
wire [31:0] rdata_h_ext_t0;
/* src = "generated/sv2v_out.v:18448.12-18448.26" */
reg [1:0] rdata_offset_q;
/* src = "generated/sv2v_out.v:18447.13-18447.20" */
reg [31:8] rdata_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18447.13-18447.20" */
reg [31:8] rdata_q_t0;
/* src = "generated/sv2v_out.v:18446.6-18446.18" */
wire rdata_update;
/* src = "generated/sv2v_out.v:18456.13-18456.24" */
wire [31:0] rdata_w_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18456.13-18456.24" */
wire [31:0] rdata_w_ext_t0;
/* src = "generated/sv2v_out.v:18410.13-18410.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:18459.7-18459.30" */
wire split_misaligned_access;
/* src = "generated/sv2v_out.v:18435.14-18435.25" */
output store_err_o;
wire store_err_o;
/* cellift = 32'd1 */
output store_err_o_t0;
wire store_err_o_t0;
/* src = "generated/sv2v_out.v:18436.14-18436.35" */
output store_resp_intg_err_o;
wire store_resp_intg_err_o;
/* cellift = 32'd1 */
output store_resp_intg_err_o_t0;
wire store_resp_intg_err_o_t0;
assign _059_ = data_gnt_i & /* src = "generated/sv2v_out.v:18674.20-18674.62" */ _289_;
assign lsu_req_done_o = _294_ & /* src = "generated/sv2v_out.v:18705.26-18705.81" */ _280_;
assign lsu_resp_valid_o = _298_ & /* src = "generated/sv2v_out.v:18720.28-18720.77" */ _281_;
assign _060_ = _281_ & /* src = "generated/sv2v_out.v:18721.32-18721.67" */ data_rvalid_i;
assign _062_ = _060_ & /* src = "generated/sv2v_out.v:18721.31-18721.87" */ _291_;
assign _064_ = _062_ & /* src = "generated/sv2v_out.v:18721.30-18721.101" */ _288_;
assign lsu_rdata_valid_o = _064_ & /* src = "generated/sv2v_out.v:18721.29-18721.119" */ _292_;
assign _066_ = data_or_pmp_err & /* src = "generated/sv2v_out.v:18739.23-18739.51" */ _288_;
assign load_err_o = _066_ & /* src = "generated/sv2v_out.v:18739.22-18739.71" */ lsu_resp_valid_o;
assign _068_ = data_or_pmp_err & /* src = "generated/sv2v_out.v:18740.24-18740.51" */ data_we_q;
assign store_err_o = _068_ & /* src = "generated/sv2v_out.v:18740.23-18740.71" */ lsu_resp_valid_o;
assign load_resp_intg_err_o = _070_ & /* src = "generated/sv2v_out.v:18741.32-18741.76" */ _288_;
assign _070_ = data_intg_err & /* src = "generated/sv2v_out.v:18742.34-18742.63" */ data_rvalid_i;
assign store_resp_intg_err_o = _070_ & /* src = "generated/sv2v_out.v:18742.33-18742.76" */ data_we_q;
assign _072_ = ~ _110_;
assign _074_ = ~ _111_;
assign _075_ = ~ _112_;
assign _076_ = ~ rdata_update;
assign _077_ = ~ addr_update;
assign _073_ = ~ ctrl_update;
assign _135_ = _110_ & handle_misaligned_d_t0;
assign _137_ = ctrl_update & lsu_we_i_t0;
assign _139_ = _111_ & pmp_err_d_t0;
assign _141_ = _112_ & lsu_err_d_t0;
assign _143_ = { rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update } & data_rdata_i_t0[31:8];
assign _145_ = { addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update } & addr_last_d_t0;
assign _136_ = _072_ & handle_misaligned_q_t0;
assign _138_ = _073_ & data_we_q_t0;
assign _140_ = _074_ & pmp_err_q_t0;
assign _142_ = _075_ & lsu_err_q_t0;
assign _144_ = { _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_, _076_ } & rdata_q_t0;
assign _146_ = { _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_ } & addr_last_o_t0;
assign _222_ = _135_ | _136_;
assign _223_ = _137_ | _138_;
assign _224_ = _139_ | _140_;
assign _225_ = _141_ | _142_;
assign _226_ = _143_ | _144_;
assign _227_ = _145_ | _146_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME handle_misaligned_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) handle_misaligned_q_t0 <= 1'h0;
else handle_misaligned_q_t0 <= _222_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME data_we_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) data_we_q_t0 <= 1'h0;
else data_we_q_t0 <= _223_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME pmp_err_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) pmp_err_q_t0 <= 1'h0;
else pmp_err_q_t0 <= _224_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME lsu_err_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) lsu_err_q_t0 <= 1'h0;
else lsu_err_q_t0 <= _225_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME rdata_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q_t0 <= 24'h000000;
else rdata_q_t0 <= _226_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME addr_last_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) addr_last_o_t0 <= 32'd0;
else addr_last_o_t0 <= _227_;
assign lsu_req_done_o_t0 = _295_ & _280_;
assign lsu_resp_valid_o_t0 = _299_ & _281_;
assign _115_ = _061_ & _291_;
assign _118_ = _063_ & _288_;
assign lsu_rdata_valid_o_t0 = _065_ & _292_;
assign _121_ = data_or_pmp_err_t0 & _288_;
assign _124_ = _067_ & lsu_resp_valid_o;
assign _127_ = data_or_pmp_err_t0 & data_we_q;
assign _128_ = _069_ & lsu_resp_valid_o;
assign _131_ = _071_ & _288_;
assign _134_ = _071_ & data_we_q;
assign _061_ = data_rvalid_i_t0 & _281_;
assign _116_ = data_or_pmp_err_t0 & _060_;
assign _119_ = data_we_q_t0 & _062_;
assign _125_ = lsu_resp_valid_o_t0 & _066_;
assign _122_ = data_we_q_t0 & data_or_pmp_err;
assign _129_ = lsu_resp_valid_o_t0 & _068_;
assign _071_ = data_rvalid_i_t0 & data_intg_err;
assign _132_ = data_we_q_t0 & _070_;
assign _117_ = _061_ & data_or_pmp_err_t0;
assign _120_ = _063_ & data_we_q_t0;
assign _126_ = _067_ & lsu_resp_valid_o_t0;
assign _123_ = data_or_pmp_err_t0 & data_we_q_t0;
assign _130_ = _069_ & lsu_resp_valid_o_t0;
assign _133_ = _071_ & data_we_q_t0;
assign _214_ = _115_ | _116_;
assign _215_ = _118_ | _119_;
assign _216_ = _121_ | _122_;
assign _217_ = _124_ | _125_;
assign _218_ = _127_ | _122_;
assign _219_ = _128_ | _129_;
assign _220_ = _131_ | _132_;
assign _221_ = _134_ | _132_;
assign _063_ = _214_ | _117_;
assign _065_ = _215_ | _120_;
assign _067_ = _216_ | _123_;
assign load_err_o_t0 = _217_ | _126_;
assign _069_ = _218_ | _123_;
assign store_err_o_t0 = _219_ | _130_;
assign load_resp_intg_err_o_t0 = _220_ | _133_;
assign store_resp_intg_err_o_t0 = _221_ | _133_;
/* src = "generated/sv2v_out.v:18706.2-18718.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME handle_misaligned_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) handle_misaligned_q <= 1'h0;
else if (_110_) handle_misaligned_q <= handle_misaligned_d;
/* src = "generated/sv2v_out.v:18525.2-18537.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME data_we_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) data_we_q <= 1'h0;
else if (ctrl_update) data_we_q <= lsu_we_i;
/* src = "generated/sv2v_out.v:18706.2-18718.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME pmp_err_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) pmp_err_q <= 1'h0;
else if (_111_) pmp_err_q <= pmp_err_d;
/* src = "generated/sv2v_out.v:18706.2-18718.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME lsu_err_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) lsu_err_q <= 1'h0;
else if (_112_) lsu_err_q <= lsu_err_d;
/* src = "generated/sv2v_out.v:18520.2-18524.34" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME rdata_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q <= 24'h000000;
else if (rdata_update) rdata_q <= data_rdata_i[31:8];
/* src = "generated/sv2v_out.v:18539.2-18543.31" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME addr_last_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) addr_last_o <= 32'd0;
else if (addr_update) addr_last_o <= addr_last_d;
/* src = "generated/sv2v_out.v:18525.2-18537.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME rdata_offset_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_offset_q <= 2'h0;
else if (ctrl_update) rdata_offset_q <= adder_result_ex_i[1:0];
/* src = "generated/sv2v_out.v:18525.2-18537.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME data_type_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) data_type_q <= 2'h0;
else if (ctrl_update) data_type_q <= lsu_type_i;
/* src = "generated/sv2v_out.v:18525.2-18537.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME data_sign_ext_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) data_sign_ext_q <= 1'h0;
else if (ctrl_update) data_sign_ext_q <= lsu_sign_ext_i;
assign _078_ = ~ _302_;
assign _079_ = ~ _300_;
assign _080_ = ~ _301_;
assign _081_ = ~ _099_;
assign _082_ = ~ { _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_ };
assign _083_ = ~ { _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_ };
assign _084_ = ~ { _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_ };
assign _085_ = ~ { _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_ };
assign _086_ = ~ { _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_ };
assign _087_ = ~ { _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_ };
assign _088_ = ~ { _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_ };
assign _089_ = ~ { _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_ };
assign _090_ = ~ data_rvalid_i;
assign _091_ = ~ data_gnt_i;
assign _092_ = ~ { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q };
assign _093_ = ~ { addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o };
assign _147_ = _079_ & _237_;
assign _149_ = _078_ & _010_;
assign _151_ = _079_ & _239_;
assign _241_ = _080_ & _044_;
assign addr_incr_req_o_t0 = _081_ & _250_;
assign _153_ = _082_ & rdata_w_ext_t0;
assign _155_ = _083_ & _252_;
assign _157_ = _084_ & _038_;
assign _159_ = _085_ & _012_;
assign _161_ = _086_ & _256_;
assign _163_ = _084_ & _040_;
assign _165_ = _085_ & _014_;
assign _167_ = _086_ & _260_;
assign _169_ = _084_ & { data_rdata_i_t0[15:0], rdata_q_t0[31:16] };
assign _171_ = _085_ & data_rdata_i_t0[31:0];
assign _173_ = _086_ & _264_;
assign _175_ = _087_ & { lsu_wdata_i_t0[15:0], lsu_wdata_i_t0[31:16] };
assign _177_ = _088_ & lsu_wdata_i_t0;
assign _179_ = _089_ & _268_;
assign _193_ = _092_ & { 24'h000000, data_rdata_i_t0[31:24] };
assign _195_ = _092_ & { 24'h000000, data_rdata_i_t0[23:16] };
assign _197_ = _092_ & { 24'h000000, data_rdata_i_t0[15:8] };
assign _199_ = _092_ & { 24'h000000, data_rdata_i_t0[7:0] };
assign _201_ = _092_ & { 16'h0000, data_rdata_i_t0[7:0], rdata_q_t0[31:24] };
assign _203_ = _092_ & { 16'h0000, data_rdata_i_t0[31:16] };
assign _205_ = _092_ & { 16'h0000, data_rdata_i_t0[23:8] };
assign _207_ = _092_ & { 16'h0000, data_rdata_i_t0[15:0] };
assign _209_ = _093_ & adder_result_ex_i_t0;
assign _237_ = _302_ & _021_;
assign _148_ = _300_ & _034_;
assign _150_ = _302_ & _023_;
assign _152_ = _300_ & _036_;
assign handle_misaligned_d_t0 = _211_ & _241_;
assign _250_ = _301_ & handle_misaligned_q_t0;
assign _154_ = { _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_, _306_ } & rdata_h_ext_t0;
assign _156_ = { _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_, _305_ } & rdata_b_ext_t0;
assign _158_ = { _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_ } & _047_;
assign _160_ = { _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_ } & _025_;
assign _162_ = { _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_ } & _254_;
assign _164_ = { _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_ } & _049_;
assign _166_ = { _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_ } & _027_;
assign _168_ = { _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_ } & _258_;
assign _170_ = { _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_, _307_ } & { data_rdata_i_t0[23:0], rdata_q_t0[31:24] };
assign _172_ = { _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_, _309_ } & { data_rdata_i_t0[7:0], rdata_q_t0 };
assign _174_ = { _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_, _212_ } & _262_;
assign _176_ = { _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_, _279_ } & { lsu_wdata_i_t0[7:0], lsu_wdata_i_t0[31:8] };
assign _178_ = { _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_, _311_ } & { lsu_wdata_i_t0[23:0], lsu_wdata_i_t0[31:24] };
assign _180_ = { _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_, _213_ } & _266_;
assign _034_ = data_rvalid_i & data_bus_err_i_t0;
assign _036_ = data_rvalid_i & data_pmp_err_i_t0;
assign _044_ = _285_ & data_gnt_i_t0;
assign _021_ = _285_ & _290_;
assign _023_ = _285_ & data_pmp_err_i_t0;
assign _007_ = lsu_req_i & lsu_we_i_t0;
assign _010_ = lsu_req_i & data_pmp_err_i_t0;
assign perf_load_o_t0 = _281_ & _007_;
assign _194_ = { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q } & { data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31:24] };
assign _196_ = { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q } & { data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23:16] };
assign _198_ = { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q } & { data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15:8] };
assign _200_ = { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q } & { data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7:0] };
assign _202_ = { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q } & { data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7:0], rdata_q_t0[31:24] };
assign _204_ = { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q } & { data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31:16] };
assign _206_ = { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q } & { data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23:8] };
assign _208_ = { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q } & { data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15:0] };
assign _210_ = { addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o } & { adder_result_ex_i_t0[31:2], 2'h0 };
assign lsu_err_d_t0 = _147_ | _148_;
assign _239_ = _149_ | _150_;
assign pmp_err_d_t0 = _151_ | _152_;
assign _252_ = _153_ | _154_;
assign lsu_rdata_o_t0 = _155_ | _156_;
assign _254_ = _157_ | _158_;
assign _256_ = _159_ | _160_;
assign rdata_b_ext_t0 = _161_ | _162_;
assign _258_ = _163_ | _164_;
assign _260_ = _165_ | _166_;
assign rdata_h_ext_t0 = _167_ | _168_;
assign _262_ = _169_ | _170_;
assign _264_ = _171_ | _172_;
assign rdata_w_ext_t0 = _173_ | _174_;
assign _266_ = _175_ | _176_;
assign _268_ = _177_ | _178_;
assign data_wdata_t0 = _179_ | _180_;
assign _047_ = _193_ | _194_;
assign _038_ = _195_ | _196_;
assign _025_ = _197_ | _198_;
assign _012_ = _199_ | _200_;
assign _049_ = _201_ | _202_;
assign _040_ = _203_ | _204_;
assign _027_ = _205_ | _206_;
assign _014_ = _207_ | _208_;
assign addr_last_d_t0 = _209_ | _210_;
assign _101_ = { _281_, lsu_req_i, data_gnt_i } != 3'h6;
assign _102_ = { _302_, _285_, data_gnt_i } != 3'h4;
assign _103_ = { _281_, lsu_req_i } != 2'h2;
assign _104_ = { _303_, _284_ } != 2'h2;
assign _105_ = { _301_, _284_ } != 2'h2;
assign _106_ = | { _302_, _301_, _281_, _303_ };
assign _107_ = { _300_, data_rvalid_i } != 2'h2;
assign _108_ = { _302_, _285_ } != 2'h2;
assign _109_ = | { _302_, _300_, _281_ };
assign _110_ = & { _102_, _101_, _103_, _104_, _106_, _105_ };
assign _111_ = & { _108_, _107_, _109_ };
assign _112_ = & { _103_, _108_, _107_, _109_ };
assign _113_ = | { _303_, _302_, _301_ };
assign _114_ = | { _303_, _301_ };
assign _094_ = ~ data_bus_err_i;
assign _095_ = ~ lsu_err_q;
assign _096_ = ~ _296_;
assign _097_ = ~ pmp_err_q;
assign _098_ = ~ busy_o;
assign _181_ = data_bus_err_i_t0 & _097_;
assign _295_ = lsu_req_i_t0 & _098_;
assign _184_ = lsu_err_q_t0 & _094_;
assign _187_ = _297_ & _097_;
assign _190_ = data_rvalid_i_t0 & _097_;
assign _182_ = pmp_err_q_t0 & _094_;
assign _185_ = data_bus_err_i_t0 & _095_;
assign _188_ = pmp_err_q_t0 & _096_;
assign _191_ = pmp_err_q_t0 & _090_;
assign _183_ = data_bus_err_i_t0 & pmp_err_q_t0;
assign _186_ = lsu_err_q_t0 & data_bus_err_i_t0;
assign _189_ = _297_ & pmp_err_q_t0;
assign _192_ = data_rvalid_i_t0 & pmp_err_q_t0;
assign _228_ = _181_ | _182_;
assign _229_ = _184_ | _185_;
assign _230_ = _187_ | _188_;
assign _231_ = _190_ | _191_;
assign _290_ = _228_ | _183_;
assign _297_ = _229_ | _186_;
assign data_or_pmp_err_t0 = _230_ | _189_;
assign _299_ = _231_ | _192_;
assign _099_ = | { _302_, _300_ };
assign _100_ = | { _302_, _301_, _300_ };
assign _211_ = _302_ | _301_;
assign _212_ = _308_ | _307_;
assign _213_ = _310_ | _279_;
assign _232_ = _301_ ? _057_ : _045_;
assign _233_ = _300_ ? _058_ : _232_;
assign _234_ = _281_ ? _004_ : 3'h0;
assign _235_ = _303_ ? _032_ : _234_;
assign ls_fsm_ns = _100_ ? _233_ : _235_;
assign _236_ = _302_ ? _020_ : _005_;
assign lsu_err_d = _300_ ? _033_ : _236_;
assign _238_ = _302_ ? _022_ : _009_;
assign pmp_err_d = _300_ ? _035_ : _238_;
assign _240_ = _301_ ? _056_ : _043_;
assign _242_ = _303_ ? _031_ : _003_;
assign handle_misaligned_d = _211_ ? _240_ : _242_;
assign ctrl_update = _114_ ? _029_ : _243_;
assign _244_ = _301_ ? _050_ : _041_;
assign _245_ = _300_ ? _054_ : _244_;
assign _243_ = _281_ ? _000_ : 1'h0;
assign _246_ = _303_ ? _029_ : _243_;
assign addr_update = _100_ ? _245_ : _246_;
assign _247_ = _281_ ? _002_ : 1'h0;
assign data_req_o = _113_ ? 1'h1 : _247_;
assign _248_ = _302_ ? _015_ : 1'h0;
assign rdata_update = _300_ ? _028_ : _248_;
assign _249_ = _301_ ? handle_misaligned_q : 1'h0;
assign addr_incr_req_o = _099_ ? 1'h1 : _249_;
assign _251_ = _306_ ? rdata_h_ext : rdata_w_ext;
assign lsu_rdata_o = _305_ ? rdata_b_ext : _251_;
assign _253_ = _307_ ? _046_ : _037_;
assign _255_ = _309_ ? _024_ : _011_;
assign rdata_b_ext = _212_ ? _253_ : _255_;
assign _257_ = _307_ ? _048_ : _039_;
assign _259_ = _309_ ? _026_ : _013_;
assign rdata_h_ext = _212_ ? _257_ : _259_;
assign _261_ = _307_ ? { data_rdata_i[23:0], rdata_q[31:24] } : { data_rdata_i[15:0], rdata_q[31:16] };
assign _263_ = _309_ ? { data_rdata_i[7:0], rdata_q } : data_rdata_i[31:0];
assign rdata_w_ext = _212_ ? _261_ : _263_;
assign _265_ = _279_ ? { lsu_wdata_i[7:0], lsu_wdata_i[31:8] } : { lsu_wdata_i[15:0], lsu_wdata_i[31:16] };
assign _267_ = _311_ ? { lsu_wdata_i[23:0], lsu_wdata_i[31:24] } : lsu_wdata_i;
assign data_wdata = _213_ ? _265_ : _267_;
assign _269_ = _279_ ? 4'h8 : 4'h4;
assign _270_ = _311_ ? 4'h2 : 4'h1;
assign _055_ = _213_ ? _269_ : _270_;
assign _272_ = _311_ ? 4'h6 : 4'h3;
assign _051_ = _213_ ? _271_ : _272_;
assign _273_ = _279_ ? 4'h7 : 4'h3;
assign _274_ = _311_ ? 4'h1 : 4'h0;
assign _030_ = _213_ ? _273_ : _274_;
assign _271_ = _279_ ? 4'h8 : 4'hc;
assign _275_ = _311_ ? 4'he : 4'hf;
assign _017_ = _213_ ? _271_ : _275_;
assign _276_ = _278_ ? _042_ : _001_;
assign data_be_o = _313_ ? _055_ : _276_;
assign _280_ = ! /* src = "generated/sv2v_out.v:18705.63-18705.80" */ ls_fsm_ns;
assign _282_ = _277_ && /* src = "generated/sv2v_out.v:18625.36-18625.83" */ _286_;
assign _283_ = _278_ && /* src = "generated/sv2v_out.v:18625.89-18625.136" */ _279_;
assign split_misaligned_access = _282_ || /* src = "generated/sv2v_out.v:18625.35-18625.137" */ _283_;
assign _285_ = data_rvalid_i || /* src = "generated/sv2v_out.v:18669.9-18669.35" */ pmp_err_q;
assign _284_ = data_gnt_i || /* src = "generated/sv2v_out.v:18685.9-18685.32" */ pmp_err_q;
assign _286_ = | /* src = "generated/sv2v_out.v:18625.62-18625.82" */ adder_result_ex_i[1:0];
assign busy_o = | /* src = "generated/sv2v_out.v:18743.18-18743.35" */ ls_fsm_cs;
assign _287_ = ~ /* src = "generated/sv2v_out.v:18645.20-18645.29" */ lsu_we_i;
assign _289_ = ~ /* src = "generated/sv2v_out.v:18674.33-18674.62" */ _293_;
assign _291_ = ~ /* src = "generated/sv2v_out.v:18721.71-18721.87" */ data_or_pmp_err;
assign _292_ = ~ /* src = "generated/sv2v_out.v:18721.105-18721.119" */ data_intg_err;
assign _288_ = ~ /* src = "generated/sv2v_out.v:18741.66-18741.76" */ data_we_q;
assign _293_ = data_bus_err_i | /* src = "generated/sv2v_out.v:18674.35-18674.61" */ pmp_err_q;
assign _294_ = lsu_req_i | /* src = "generated/sv2v_out.v:18705.27-18705.58" */ busy_o;
assign _296_ = lsu_err_q | /* src = "generated/sv2v_out.v:18719.28-18719.54" */ data_bus_err_i;
assign data_or_pmp_err = _296_ | /* src = "generated/sv2v_out.v:18719.27-18719.67" */ pmp_err_q;
assign _298_ = data_rvalid_i | /* src = "generated/sv2v_out.v:18720.29-18720.54" */ pmp_err_q;
/* src = "generated/sv2v_out.v:18706.2-18718.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME ls_fsm_cs */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) ls_fsm_cs <= 3'h0;
else ls_fsm_cs <= ls_fsm_ns;
assign _058_ = data_rvalid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18694.9-18694.22|generated/sv2v_out.v:18694.5-18700.8" */ 3'h0 : ls_fsm_cs;
assign _028_ = data_rvalid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18694.9-18694.22|generated/sv2v_out.v:18694.5-18700.8" */ _288_ : 1'h0;
assign _054_ = data_rvalid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18694.9-18694.22|generated/sv2v_out.v:18694.5-18700.8" */ _094_ : 1'h0;
assign _033_ = data_rvalid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18694.9-18694.22|generated/sv2v_out.v:18694.5-18700.8" */ data_bus_err_i : 1'hx;
assign _035_ = data_rvalid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18694.9-18694.22|generated/sv2v_out.v:18694.5-18700.8" */ data_pmp_err_i : 1'hx;
assign _056_ = _284_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18685.9-18685.32|generated/sv2v_out.v:18685.5-18690.8" */ 1'h0 : 1'hx;
assign _057_ = _284_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18685.9-18685.32|generated/sv2v_out.v:18685.5-18690.8" */ 3'h0 : ls_fsm_cs;
assign _050_ = _284_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18685.9-18685.32|generated/sv2v_out.v:18685.5-18690.8" */ _095_ : 1'h0;
assign _052_ = data_gnt_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18677.14-18677.24|generated/sv2v_out.v:18677.10-18680.8" */ 1'h0 : 1'hx;
assign _053_ = data_gnt_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18677.14-18677.24|generated/sv2v_out.v:18677.10-18680.8" */ 3'h4 : ls_fsm_cs;
assign _043_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18669.9-18669.35|generated/sv2v_out.v:18669.5-18680.8" */ _091_ : _052_;
assign _041_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18669.9-18669.35|generated/sv2v_out.v:18669.5-18680.8" */ _059_ : 1'h0;
assign _045_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18669.9-18669.35|generated/sv2v_out.v:18669.5-18680.8" */ _316_ : _053_;
assign _015_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18669.9-18669.35|generated/sv2v_out.v:18669.5-18680.8" */ _288_ : 1'h0;
assign _020_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18669.9-18669.35|generated/sv2v_out.v:18669.5-18680.8" */ _293_ : 1'hx;
assign _022_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18669.9-18669.35|generated/sv2v_out.v:18669.5-18680.8" */ data_pmp_err_i : 1'hx;
assign _032_ = _284_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18659.9-18659.32|generated/sv2v_out.v:18659.5-18664.8" */ 3'h2 : ls_fsm_cs;
assign _031_ = _284_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18659.9-18659.32|generated/sv2v_out.v:18659.5-18664.8" */ 1'h1 : 1'hx;
assign _029_ = _284_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18659.9-18659.32|generated/sv2v_out.v:18659.5-18664.8" */ 1'h1 : 1'h0;
assign _019_ = data_gnt_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18647.10-18647.20|generated/sv2v_out.v:18647.6-18654.59" */ _314_ : _315_;
assign _018_ = data_gnt_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18647.10-18647.20|generated/sv2v_out.v:18647.6-18654.59" */ split_misaligned_access : 1'hx;
assign _016_ = data_gnt_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18647.10-18647.20|generated/sv2v_out.v:18647.6-18654.59" */ 1'h1 : 1'h0;
assign _004_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18641.9-18641.18|generated/sv2v_out.v:18641.5-18655.8" */ _019_ : ls_fsm_cs;
assign _003_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18641.9-18641.18|generated/sv2v_out.v:18641.5-18655.8" */ _018_ : 1'hx;
assign _000_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18641.9-18641.18|generated/sv2v_out.v:18641.5-18655.8" */ _016_ : 1'h0;
assign _008_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18641.9-18641.18|generated/sv2v_out.v:18641.5-18655.8" */ lsu_we_i : 1'h0;
assign _006_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18641.9-18641.18|generated/sv2v_out.v:18641.5-18655.8" */ _287_ : 1'h0;
assign _005_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18641.9-18641.18|generated/sv2v_out.v:18641.5-18655.8" */ 1'h0 : 1'hx;
assign _009_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18641.9-18641.18|generated/sv2v_out.v:18641.5-18655.8" */ data_pmp_err_i : 1'h0;
assign _002_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18641.9-18641.18|generated/sv2v_out.v:18641.5-18655.8" */ 1'h1 : 1'h0;
assign perf_store_o = _281_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18638.3-18703.10" */ _008_ : 1'h0;
assign perf_load_o = _281_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18638.3-18703.10" */ _006_ : 1'h0;
assign _303_ = ls_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18638.3-18703.10" */ 3'h1;
assign _281_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18638.3-18703.10" */ ls_fsm_cs;
assign _300_ = ls_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18638.3-18703.10" */ 3'h4;
assign _301_ = ls_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18638.3-18703.10" */ 3'h3;
assign _302_ = ls_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18638.3-18703.10" */ 3'h2;
assign _305_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18601.3-18606.10" */ _304_;
assign _304_[0] = data_type_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18601.3-18606.10" */ 2'h2;
assign _304_[1] = data_type_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18601.3-18606.10" */ 2'h3;
assign _306_ = data_type_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18601.3-18606.10" */ 2'h1;
assign _046_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18594.9-18594.25|generated/sv2v_out.v:18594.5-18597.67" */ { data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31:24] } : { 24'h000000, data_rdata_i[31:24] };
assign _037_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18589.9-18589.25|generated/sv2v_out.v:18589.5-18592.67" */ { data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23:16] } : { 24'h000000, data_rdata_i[23:16] };
assign _024_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18584.9-18584.25|generated/sv2v_out.v:18584.5-18587.66" */ { data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15:8] } : { 24'h000000, data_rdata_i[15:8] };
assign _011_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18579.9-18579.25|generated/sv2v_out.v:18579.5-18582.64" */ { data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7:0] } : { 24'h000000, data_rdata_i[7:0] };
assign _048_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18570.9-18570.25|generated/sv2v_out.v:18570.5-18573.80" */ { data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7:0], rdata_q[31:24] } : { 16'h0000, data_rdata_i[7:0], rdata_q[31:24] };
assign _039_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18565.9-18565.25|generated/sv2v_out.v:18565.5-18568.67" */ { data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31:16] } : { 16'h0000, data_rdata_i[31:16] };
assign _026_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18560.9-18560.25|generated/sv2v_out.v:18560.5-18563.66" */ { data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23:8] } : { 16'h0000, data_rdata_i[23:8] };
assign _013_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18555.9-18555.25|generated/sv2v_out.v:18555.5-18558.66" */ { data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15:0] } : { 16'h0000, data_rdata_i[15:0] };
assign _307_ = rdata_offset_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18545.3-18551.10" */ 2'h3;
assign _308_ = rdata_offset_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18545.3-18551.10" */ 2'h2;
assign _309_ = rdata_offset_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18545.3-18551.10" */ 2'h1;
assign _313_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18473.3-18511.10" */ _312_;
assign _042_ = handle_misaligned_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18492.9-18492.29|generated/sv2v_out.v:18492.5-18501.24" */ 4'h1 : _051_;
assign _279_ = adder_result_ex_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18476.6-18482.13" */ 2'h3;
assign _310_ = adder_result_ex_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18476.6-18482.13" */ 2'h2;
assign _311_ = adder_result_ex_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18476.6-18482.13" */ 2'h1;
assign _001_ = handle_misaligned_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18475.9-18475.29|generated/sv2v_out.v:18475.5-18490.13" */ _030_ : _017_;
assign _312_[0] = lsu_type_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18473.3-18511.10" */ 2'h2;
assign _312_[1] = lsu_type_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18473.3-18511.10" */ 2'h3;
assign _278_ = lsu_type_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18473.3-18511.10" */ 2'h1;
assign _277_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18473.3-18511.10" */ lsu_type_i;
assign data_intg_err = | /* src = "generated/sv2v_out.v:18619.27-18619.35" */ \g_mem_rdata_ecc.ecc_err ;
assign addr_last_d = addr_incr_req_o ? /* src = "generated/sv2v_out.v:18538.24-18538.73" */ { adder_result_ex_i[31:2], 2'h0 } : adder_result_ex_i;
assign _314_ = split_misaligned_access ? /* src = "generated/sv2v_out.v:18651.20-18651.57" */ 3'h2 : 3'h0;
assign _315_ = split_misaligned_access ? /* src = "generated/sv2v_out.v:18654.20-18654.57" */ 3'h1 : 3'h3;
assign _316_ = data_gnt_i ? /* src = "generated/sv2v_out.v:18673.19-18673.43" */ 3'h0 : 3'h3;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18615.30-18618.5" */
prim_secded_inv_39_32_dec \g_mem_rdata_ecc.u_data_intg_dec  (
.data_i(\g_mem_rdata_ecc.data_rdata_buf ),
.data_i_t0(\g_mem_rdata_ecc.data_rdata_buf_t0 ),
.err_o(\g_mem_rdata_ecc.ecc_err ),
.err_o_t0(\g_mem_rdata_ecc.ecc_err_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18611.37-18614.5" */
\$paramod\prim_buf\Width=32'00000000000000000000000000100111  \g_mem_rdata_ecc.u_prim_buf_instr_rdata  (
.in_i(data_rdata_i),
.in_i_t0(data_rdata_i_t0),
.out_o(\g_mem_rdata_ecc.data_rdata_buf ),
.out_o_t0(\g_mem_rdata_ecc.data_rdata_buf_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18729.30-18732.5" */
prim_secded_inv_39_32_enc \g_mem_wdata_ecc.u_data_gen  (
.data_i(data_wdata),
.data_i_t0(data_wdata_t0),
.data_o(data_wdata_o),
.data_o_t0(data_wdata_o_t0)
);
assign busy_o_t0 = 1'h0;
assign data_addr_o = { adder_result_ex_i[31:2], 2'h0 };
assign data_addr_o_t0 = { adder_result_ex_i_t0[31:2], 2'h0 };
assign data_be_o_t0 = 4'h0;
assign data_req_o_t0 = 1'h0;
assign data_we_o = lsu_we_i;
assign data_we_o_t0 = lsu_we_i_t0;
assign perf_store_o_t0 = perf_load_o_t0;
endmodule

module \$paramod\ibex_prefetch_buffer\ResetAll=1'1 (clk_i, rst_ni, req_i, branch_i, addr_i, ready_i, valid_o, rdata_o, addr_o, err_o, err_plus2_o, instr_req_o, instr_gnt_i, instr_addr_o, instr_rdata_i, instr_err_i, instr_rvalid_i, busy_o, busy_o_t0, valid_o_t0, req_i_t0
, ready_i_t0, rdata_o_t0, instr_rvalid_i_t0, instr_req_o_t0, instr_rdata_i_t0, instr_gnt_i_t0, instr_err_i_t0, instr_addr_o_t0, err_plus2_o_t0, branch_i_t0, addr_o_t0, addr_i_t0, err_o_t0);
/* src = "generated/sv2v_out.v:20024.26-20024.57" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20024.26-20024.57" */
wire _001_;
/* src = "generated/sv2v_out.v:20028.27-20028.55" */
wire _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20028.27-20028.55" */
wire _003_;
/* src = "generated/sv2v_out.v:20065.38-20065.61" */
wire _004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20065.38-20065.61" */
wire _005_;
/* src = "generated/sv2v_out.v:20066.36-20066.77" */
wire _006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20066.36-20066.77" */
wire _007_;
/* src = "generated/sv2v_out.v:20066.82-20066.115" */
wire _008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20066.82-20066.115" */
wire _009_;
/* src = "generated/sv2v_out.v:20069.38-20069.92" */
wire _010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20069.38-20069.92" */
wire _011_;
/* src = "generated/sv2v_out.v:20070.36-20070.108" */
wire _012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20070.36-20070.108" */
wire _013_;
/* src = "generated/sv2v_out.v:20070.113-20070.146" */
wire _014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20070.113-20070.146" */
wire _015_;
wire [31:0] _016_;
wire [31:0] _017_;
wire _018_;
wire _019_;
wire _020_;
wire [31:0] _021_;
wire [31:0] _022_;
wire [1:0] _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire [31:0] _043_;
wire [31:0] _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire [31:0] _079_;
wire [31:0] _080_;
wire [1:0] _081_;
wire [1:0] _082_;
wire [29:0] _083_;
wire [29:0] _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire [31:0] _106_;
wire [31:0] _107_;
wire [31:0] _108_;
wire [31:0] _109_;
wire [31:0] _110_;
wire [1:0] _111_;
wire [1:0] _112_;
wire [1:0] _113_;
wire [1:0] _114_;
wire [31:0] _115_;
wire [31:0] _116_;
wire [31:0] _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire [31:0] _130_;
wire [1:0] _131_;
wire [29:0] _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire [31:0] _141_;
wire [31:0] _142_;
wire [31:0] _143_;
/* src = "generated/sv2v_out.v:20026.35-20026.47" */
wire _144_;
/* src = "generated/sv2v_out.v:20004.25-20004.58" */
wire [1:0] _145_;
/* src = "generated/sv2v_out.v:20024.35-20024.56" */
wire _146_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20024.35-20024.56" */
wire _147_;
/* src = "generated/sv2v_out.v:20027.40-20027.64" */
wire _148_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20027.40-20027.64" */
wire _149_;
/* src = "generated/sv2v_out.v:20066.35-20066.116" */
wire _150_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20066.35-20066.116" */
wire _151_;
/* src = "generated/sv2v_out.v:20070.35-20070.147" */
wire _152_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20070.35-20070.147" */
wire _153_;
/* src = "generated/sv2v_out.v:19996.18-19996.38" */
wire _154_;
/* src = "generated/sv2v_out.v:20045.25-20045.72" */
wire [31:0] _155_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20045.25-20045.72" */
wire [31:0] _156_;
/* src = "generated/sv2v_out.v:20060.54-20060.86" */
wire [31:0] _157_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20060.54-20060.86" */
wire [31:0] _158_;
/* src = "generated/sv2v_out.v:19955.20-19955.26" */
input [31:0] addr_i;
wire [31:0] addr_i;
/* cellift = 32'd1 */
input [31:0] addr_i_t0;
wire [31:0] addr_i_t0;
/* src = "generated/sv2v_out.v:19959.21-19959.27" */
output [31:0] addr_o;
wire [31:0] addr_o;
/* cellift = 32'd1 */
output [31:0] addr_o_t0;
wire [31:0] addr_o_t0;
/* src = "generated/sv2v_out.v:19979.13-19979.29" */
wire [1:0] branch_discard_n;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19979.13-19979.29" */
wire [1:0] branch_discard_n_t0;
/* src = "generated/sv2v_out.v:19981.12-19981.28" */
reg [1:0] branch_discard_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19981.12-19981.28" */
reg [1:0] branch_discard_q_t0;
/* src = "generated/sv2v_out.v:19980.13-19980.29" */
wire [1:0] branch_discard_s;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19980.13-19980.29" */
wire [1:0] branch_discard_s_t0;
/* src = "generated/sv2v_out.v:19954.13-19954.21" */
input branch_i;
wire branch_i;
/* cellift = 32'd1 */
input branch_i_t0;
wire branch_i_t0;
/* src = "generated/sv2v_out.v:19968.14-19968.20" */
output busy_o;
wire busy_o;
/* cellift = 32'd1 */
output busy_o_t0;
wire busy_o_t0;
/* src = "generated/sv2v_out.v:19951.13-19951.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:19974.7-19974.20" */
wire discard_req_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19974.7-19974.20" */
wire discard_req_d_t0;
/* src = "generated/sv2v_out.v:19975.6-19975.19" */
reg discard_req_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19975.6-19975.19" */
reg discard_req_q_t0;
/* src = "generated/sv2v_out.v:19960.14-19960.19" */
output err_o;
wire err_o;
/* cellift = 32'd1 */
output err_o_t0;
wire err_o_t0;
/* src = "generated/sv2v_out.v:19961.14-19961.25" */
output err_plus2_o;
wire err_plus2_o;
/* cellift = 32'd1 */
output err_plus2_o_t0;
wire err_plus2_o_t0;
/* src = "generated/sv2v_out.v:19986.14-19986.26" */
wire [31:0] fetch_addr_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19986.14-19986.26" */
wire [31:0] fetch_addr_d_t0;
/* src = "generated/sv2v_out.v:19988.7-19988.20" */
wire fetch_addr_en;
/* src = "generated/sv2v_out.v:19987.13-19987.25" */
reg [31:0] fetch_addr_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19987.13-19987.25" */
reg [31:0] fetch_addr_q_t0;
/* src = "generated/sv2v_out.v:19995.13-19995.22" */
wire [1:0] fifo_busy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19995.13-19995.22" */
/* unused_bits = "0 1" */
wire [1:0] fifo_busy_t0;
/* src = "generated/sv2v_out.v:19993.7-19993.17" */
wire fifo_ready;
/* src = "generated/sv2v_out.v:19991.7-19991.17" */
wire fifo_valid;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19991.7-19991.17" */
wire fifo_valid_t0;
/* src = "generated/sv2v_out.v:19989.14-19989.24" */
/* unused_bits = "0 1" */
wire [31:0] instr_addr;
/* src = "generated/sv2v_out.v:19964.21-19964.33" */
output [31:0] instr_addr_o;
wire [31:0] instr_addr_o;
/* cellift = 32'd1 */
output [31:0] instr_addr_o_t0;
wire [31:0] instr_addr_o_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19989.14-19989.24" */
/* unused_bits = "0 1" */
wire [31:0] instr_addr_t0;
/* src = "generated/sv2v_out.v:19966.13-19966.24" */
input instr_err_i;
wire instr_err_i;
/* cellift = 32'd1 */
input instr_err_i_t0;
wire instr_err_i_t0;
/* src = "generated/sv2v_out.v:19963.13-19963.24" */
input instr_gnt_i;
wire instr_gnt_i;
/* cellift = 32'd1 */
input instr_gnt_i_t0;
wire instr_gnt_i_t0;
/* src = "generated/sv2v_out.v:19965.20-19965.33" */
input [31:0] instr_rdata_i;
wire [31:0] instr_rdata_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_i_t0;
wire [31:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:19962.14-19962.25" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:19967.13-19967.27" */
input instr_rvalid_i;
wire instr_rvalid_i;
/* cellift = 32'd1 */
input instr_rvalid_i_t0;
wire instr_rvalid_i_t0;
/* src = "generated/sv2v_out.v:19958.21-19958.28" */
output [31:0] rdata_o;
wire [31:0] rdata_o;
/* cellift = 32'd1 */
output [31:0] rdata_o_t0;
wire [31:0] rdata_o_t0;
/* src = "generated/sv2v_out.v:19976.13-19976.32" */
wire [1:0] rdata_outstanding_n;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19976.13-19976.32" */
wire [1:0] rdata_outstanding_n_t0;
/* src = "generated/sv2v_out.v:19978.12-19978.31" */
reg [1:0] rdata_outstanding_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19978.12-19978.31" */
reg [1:0] rdata_outstanding_q_t0;
/* src = "generated/sv2v_out.v:19977.13-19977.32" */
wire [1:0] rdata_outstanding_s;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19977.13-19977.32" */
wire [1:0] rdata_outstanding_s_t0;
/* src = "generated/sv2v_out.v:19956.13-19956.20" */
input ready_i;
wire ready_i;
/* cellift = 32'd1 */
input ready_i_t0;
wire ready_i_t0;
/* src = "generated/sv2v_out.v:19953.13-19953.18" */
input req_i;
wire req_i;
/* cellift = 32'd1 */
input req_i_t0;
wire req_i_t0;
/* src = "generated/sv2v_out.v:19952.13-19952.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:19985.7-19985.21" */
wire stored_addr_en;
/* src = "generated/sv2v_out.v:19984.13-19984.26" */
reg [31:0] stored_addr_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19984.13-19984.26" */
reg [31:0] stored_addr_q_t0;
/* src = "generated/sv2v_out.v:19970.7-19970.20" */
wire valid_new_req;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19970.7-19970.20" */
wire valid_new_req_t0;
/* src = "generated/sv2v_out.v:19957.14-19957.21" */
output valid_o;
wire valid_o;
/* cellift = 32'd1 */
output valid_o_t0;
wire valid_o_t0;
/* src = "generated/sv2v_out.v:19972.7-19972.18" */
wire valid_req_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19972.7-19972.18" */
wire valid_req_d_t0;
/* src = "generated/sv2v_out.v:19973.6-19973.17" */
reg valid_req_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19973.6-19973.17" */
reg valid_req_q_t0;
assign fetch_addr_d = _155_ + /* src = "generated/sv2v_out.v:20045.24-20045.126" */ { 29'h00000000, _002_, 2'h0 };
assign _000_ = req_i & /* src = "generated/sv2v_out.v:20024.26-20024.57" */ _146_;
assign valid_new_req = _000_ & /* src = "generated/sv2v_out.v:20024.25-20024.84" */ _039_;
assign valid_req_d = instr_req_o & /* src = "generated/sv2v_out.v:20026.23-20026.47" */ _144_;
assign discard_req_d = valid_req_q & /* src = "generated/sv2v_out.v:20027.25-20027.65" */ _148_;
assign stored_addr_en = _002_ & /* src = "generated/sv2v_out.v:20028.26-20028.71" */ _144_;
assign _002_ = valid_new_req & /* src = "generated/sv2v_out.v:20045.90-20045.118" */ _024_;
assign _008_ = branch_i & /* src = "generated/sv2v_out.v:20066.82-20066.115" */ rdata_outstanding_q[0];
assign _010_ = _004_ & /* src = "generated/sv2v_out.v:20069.38-20069.92" */ rdata_outstanding_q[0];
assign _004_ = instr_req_o & /* src = "generated/sv2v_out.v:20070.38-20070.61" */ instr_gnt_i;
assign _006_ = _004_ & /* src = "generated/sv2v_out.v:20070.37-20070.78" */ discard_req_d;
assign _012_ = _006_ & /* src = "generated/sv2v_out.v:20070.36-20070.108" */ rdata_outstanding_q[0];
assign _014_ = branch_i & /* src = "generated/sv2v_out.v:20070.113-20070.146" */ rdata_outstanding_q[1];
assign fifo_valid = instr_rvalid_i & /* src = "generated/sv2v_out.v:20076.22-20076.59" */ _038_;
assign _016_ = ~ _156_;
assign _017_ = ~ { 29'h00000000, _003_, 2'h0 };
assign _043_ = _155_ & _016_;
assign _044_ = { 29'h00000000, _002_, 2'h0 } & _017_;
assign _142_ = _043_ + _044_;
assign _115_ = _155_ | _156_;
assign _116_ = { 29'h00000000, _002_, 2'h0 } | { 29'h00000000, _003_, 2'h0 };
assign _143_ = _115_ + _116_;
assign _141_ = _142_ ^ _143_;
assign _117_ = _141_ | _156_;
assign fetch_addr_d_t0 = _117_ | { 29'h00000000, _003_, 2'h0 };
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME valid_req_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) valid_req_q_t0 <= 1'h0;
else valid_req_q_t0 <= valid_req_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME discard_req_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) discard_req_q_t0 <= 1'h0;
else discard_req_q_t0 <= discard_req_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_outstanding_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_outstanding_q_t0 <= 2'h0;
else rdata_outstanding_q_t0 <= rdata_outstanding_s_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME branch_discard_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_discard_q_t0 <= 2'h0;
else branch_discard_q_t0 <= branch_discard_s_t0;
assign _018_ = ~ fetch_addr_en;
assign _019_ = ~ _042_;
assign _020_ = ~ stored_addr_en;
assign _079_ = { fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en } & fetch_addr_d_t0;
assign _081_ = { _042_, _042_ } & _158_[1:0];
assign _083_ = { stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en } & instr_addr_t0[31:2];
assign _080_ = { _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_ } & fetch_addr_q_t0;
assign _082_ = { _019_, _019_ } & stored_addr_q_t0[1:0];
assign _084_ = { _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_ } & stored_addr_q_t0[31:2];
assign _130_ = _079_ | _080_;
assign _131_ = _081_ | _082_;
assign _132_ = _083_ | _084_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME fetch_addr_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) fetch_addr_q_t0 <= 32'd0;
else fetch_addr_q_t0 <= _130_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME stored_addr_q_t0[1:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) stored_addr_q_t0[1:0] <= 2'h0;
else stored_addr_q_t0[1:0] <= _131_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME stored_addr_q_t0[31:2] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) stored_addr_q_t0[31:2] <= 30'h00000000;
else stored_addr_q_t0[31:2] <= _132_;
assign _045_ = req_i_t0 & _146_;
assign _048_ = _001_ & _039_;
assign _051_ = instr_req_o_t0 & _144_;
assign _054_ = valid_req_q_t0 & _148_;
assign _057_ = valid_new_req_t0 & _024_;
assign _060_ = branch_i_t0 & rdata_outstanding_q[0];
assign _063_ = _005_ & rdata_outstanding_q[0];
assign _066_ = instr_req_o_t0 & instr_gnt_i;
assign _067_ = _005_ & discard_req_d;
assign _070_ = _007_ & rdata_outstanding_q[0];
assign _073_ = branch_i_t0 & rdata_outstanding_q[1];
assign _076_ = instr_rvalid_i_t0 & _038_;
assign _046_ = _147_ & req_i;
assign _049_ = rdata_outstanding_q_t0[1] & _000_;
assign _052_ = instr_gnt_i_t0 & instr_req_o;
assign _055_ = _149_ & valid_req_q;
assign _058_ = valid_req_q_t0 & valid_new_req;
assign _061_ = rdata_outstanding_q_t0[0] & branch_i;
assign _064_ = rdata_outstanding_q_t0[0] & _004_;
assign _068_ = discard_req_d_t0 & _004_;
assign _071_ = rdata_outstanding_q_t0[0] & _006_;
assign _074_ = rdata_outstanding_q_t0[1] & branch_i;
assign _077_ = branch_discard_q_t0[0] & instr_rvalid_i;
assign _047_ = req_i_t0 & _147_;
assign _050_ = _001_ & rdata_outstanding_q_t0[1];
assign _053_ = instr_req_o_t0 & instr_gnt_i_t0;
assign _056_ = valid_req_q_t0 & _149_;
assign _059_ = valid_new_req_t0 & valid_req_q_t0;
assign _062_ = branch_i_t0 & rdata_outstanding_q_t0[0];
assign _065_ = _005_ & rdata_outstanding_q_t0[0];
assign _069_ = _005_ & discard_req_d_t0;
assign _072_ = _007_ & rdata_outstanding_q_t0[0];
assign _075_ = branch_i_t0 & rdata_outstanding_q_t0[1];
assign _078_ = instr_rvalid_i_t0 & branch_discard_q_t0[0];
assign _118_ = _045_ | _046_;
assign _119_ = _048_ | _049_;
assign _120_ = _051_ | _052_;
assign _121_ = _054_ | _055_;
assign _122_ = _057_ | _058_;
assign _123_ = _060_ | _061_;
assign _124_ = _063_ | _064_;
assign _125_ = _066_ | _052_;
assign _126_ = _067_ | _068_;
assign _127_ = _070_ | _071_;
assign _128_ = _073_ | _074_;
assign _129_ = _076_ | _077_;
assign _001_ = _118_ | _047_;
assign valid_new_req_t0 = _119_ | _050_;
assign valid_req_d_t0 = _120_ | _053_;
assign discard_req_d_t0 = _121_ | _056_;
assign _003_ = _122_ | _059_;
assign _009_ = _123_ | _062_;
assign _011_ = _124_ | _065_;
assign _005_ = _125_ | _053_;
assign _007_ = _126_ | _069_;
assign _013_ = _127_ | _072_;
assign _015_ = _128_ | _075_;
assign fifo_valid_t0 = _129_ | _078_;
/* src = "generated/sv2v_out.v:20048.4-20052.35" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME fetch_addr_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) fetch_addr_q <= 32'd0;
else if (fetch_addr_en) fetch_addr_q <= fetch_addr_d;
/* src = "generated/sv2v_out.v:20032.4-20036.37" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME stored_addr_q[1:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) stored_addr_q[1:0] <= 2'h0;
else if (_042_) stored_addr_q[1:0] <= _157_[1:0];
/* src = "generated/sv2v_out.v:20032.4-20036.37" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME stored_addr_q[31:2] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) stored_addr_q[31:2] <= 30'h00000000;
else if (stored_addr_en) stored_addr_q[31:2] <= instr_addr[31:2];
assign _021_ = ~ { branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i };
assign _022_ = ~ { valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q };
assign _023_ = ~ { instr_rvalid_i, instr_rvalid_i };
assign _106_ = _021_ & { fetch_addr_q_t0[31:2], 2'h0 };
assign _108_ = _021_ & fetch_addr_q_t0;
assign _109_ = _022_ & _158_;
assign _111_ = _023_ & rdata_outstanding_n_t0;
assign _113_ = _023_ & branch_discard_n_t0;
assign _107_ = { branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i } & addr_i_t0;
assign _110_ = { valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q } & stored_addr_q_t0;
assign _112_ = { instr_rvalid_i, instr_rvalid_i } & { 1'h0, rdata_outstanding_n_t0[1] };
assign _114_ = { instr_rvalid_i, instr_rvalid_i } & { 1'h0, branch_discard_n_t0[1] };
assign _156_ = _106_ | _107_;
assign _158_ = _108_ | _107_;
assign instr_addr_t0 = _109_ | _110_;
assign rdata_outstanding_s_t0 = _111_ | _112_;
assign branch_discard_s_t0 = _113_ | _114_;
assign _024_ = ~ valid_req_q;
assign _042_ = & { _024_, stored_addr_en };
assign _025_ = ~ _154_;
assign _027_ = ~ branch_i;
assign _028_ = ~ _004_;
assign _029_ = ~ _006_;
assign _030_ = ~ _150_;
assign _031_ = ~ _010_;
assign _032_ = ~ _012_;
assign _033_ = ~ _152_;
assign _034_ = ~ valid_new_req;
assign _035_ = ~ discard_req_q;
assign _036_ = ~ rdata_outstanding_q[0];
assign _037_ = ~ _008_;
assign _038_ = ~ branch_discard_q[0];
assign _039_ = ~ rdata_outstanding_q[1];
assign _040_ = ~ _014_;
assign _041_ = ~ branch_discard_q[1];
assign _085_ = valid_req_q_t0 & _034_;
assign _086_ = branch_i_t0 & _035_;
assign _089_ = _005_ & _036_;
assign _091_ = _007_ & _037_;
assign _094_ = _151_ & _038_;
assign _097_ = _011_ & _039_;
assign _100_ = _013_ & _040_;
assign _103_ = _153_ & _041_;
assign busy_o_t0 = instr_req_o_t0 & _025_;
assign _147_ = branch_i_t0 & _026_;
assign _087_ = discard_req_q_t0 & _027_;
assign _090_ = rdata_outstanding_q_t0[0] & _028_;
assign _092_ = _009_ & _029_;
assign _095_ = branch_discard_q_t0[0] & _030_;
assign _098_ = rdata_outstanding_q_t0[1] & _031_;
assign _101_ = _015_ & _032_;
assign _104_ = branch_discard_q_t0[1] & _033_;
assign _088_ = branch_i_t0 & discard_req_q_t0;
assign _093_ = _007_ & _009_;
assign _096_ = _151_ & branch_discard_q_t0[0];
assign _099_ = _011_ & rdata_outstanding_q_t0[1];
assign _102_ = _013_ & _015_;
assign _105_ = _153_ & branch_discard_q_t0[1];
assign _133_ = _085_ | _057_;
assign _134_ = _086_ | _087_;
assign _135_ = _089_ | _090_;
assign _136_ = _091_ | _092_;
assign _137_ = _094_ | _095_;
assign _138_ = _097_ | _098_;
assign _139_ = _100_ | _101_;
assign _140_ = _103_ | _104_;
assign instr_req_o_t0 = _133_ | _059_;
assign _149_ = _134_ | _088_;
assign rdata_outstanding_n_t0[0] = _135_ | _065_;
assign _151_ = _136_ | _093_;
assign branch_discard_n_t0[0] = _137_ | _096_;
assign rdata_outstanding_n_t0[1] = _138_ | _099_;
assign _153_ = _139_ | _102_;
assign branch_discard_n_t0[1] = _140_ | _105_;
assign fifo_ready = ! /* src = "generated/sv2v_out.v:0.0-0.0" */ _026_;
assign _144_ = ~ /* src = "generated/sv2v_out.v:20028.59-20028.71" */ instr_gnt_i;
assign busy_o = _154_ | /* src = "generated/sv2v_out.v:19996.18-19996.52" */ instr_req_o;
assign _145_ = fifo_busy | /* src = "generated/sv2v_out.v:20004.25-20004.58" */ { rdata_outstanding_q[0], rdata_outstanding_q[1] };
assign _146_ = fifo_ready | /* src = "generated/sv2v_out.v:20024.35-20024.56" */ branch_i;
assign instr_req_o = valid_req_q | /* src = "generated/sv2v_out.v:20025.21-20025.48" */ valid_new_req;
assign _148_ = branch_i | /* src = "generated/sv2v_out.v:20027.40-20027.64" */ discard_req_q;
assign fetch_addr_en = branch_i | /* src = "generated/sv2v_out.v:20044.25-20044.66" */ _002_;
assign rdata_outstanding_n[0] = _004_ | /* src = "generated/sv2v_out.v:20065.37-20065.87" */ rdata_outstanding_q[0];
assign _150_ = _006_ | /* src = "generated/sv2v_out.v:20066.35-20066.116" */ _008_;
assign branch_discard_n[0] = _150_ | /* src = "generated/sv2v_out.v:20066.34-20066.139" */ branch_discard_q[0];
assign rdata_outstanding_n[1] = _010_ | /* src = "generated/sv2v_out.v:20069.37-20069.118" */ rdata_outstanding_q[1];
assign _152_ = _012_ | /* src = "generated/sv2v_out.v:20070.35-20070.147" */ _014_;
assign branch_discard_n[1] = _152_ | /* src = "generated/sv2v_out.v:20070.34-20070.170" */ branch_discard_q[1];
/* src = "generated/sv2v_out.v:20078.2-20090.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME valid_req_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) valid_req_q <= 1'h0;
else valid_req_q <= valid_req_d;
/* src = "generated/sv2v_out.v:20078.2-20090.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME discard_req_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) discard_req_q <= 1'h0;
else discard_req_q <= discard_req_d;
/* src = "generated/sv2v_out.v:20078.2-20090.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_outstanding_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_outstanding_q <= 2'h0;
else rdata_outstanding_q <= rdata_outstanding_s;
/* src = "generated/sv2v_out.v:20078.2-20090.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME branch_discard_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_discard_q <= 2'h0;
else branch_discard_q <= branch_discard_s;
assign _026_ = & /* src = "generated/sv2v_out.v:20004.22-20004.59" */ _145_;
assign _154_ = | /* src = "generated/sv2v_out.v:19996.18-19996.38" */ rdata_outstanding_q;
assign _155_ = branch_i ? /* src = "generated/sv2v_out.v:20045.25-20045.72" */ addr_i : { fetch_addr_q[31:2], 2'h0 };
assign _157_ = branch_i ? /* src = "generated/sv2v_out.v:20060.54-20060.86" */ addr_i : fetch_addr_q;
assign instr_addr = valid_req_q ? /* src = "generated/sv2v_out.v:20060.23-20060.87" */ stored_addr_q : _157_;
assign rdata_outstanding_s = instr_rvalid_i ? /* src = "generated/sv2v_out.v:20074.32-20074.103" */ { 1'h0, rdata_outstanding_n[1] } : rdata_outstanding_n;
assign branch_discard_s = instr_rvalid_i ? /* src = "generated/sv2v_out.v:20075.29-20075.94" */ { 1'h0, branch_discard_n[1] } : branch_discard_n;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20008.4-20023.3" */
\$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  fifo_i (
.busy_o(fifo_busy),
.busy_o_t0(fifo_busy_t0),
.clear_i(branch_i),
.clear_i_t0(branch_i_t0),
.clk_i(clk_i),
.in_addr_i(addr_i),
.in_addr_i_t0(addr_i_t0),
.in_err_i(instr_err_i),
.in_err_i_t0(instr_err_i_t0),
.in_rdata_i(instr_rdata_i),
.in_rdata_i_t0(instr_rdata_i_t0),
.in_valid_i(fifo_valid),
.in_valid_i_t0(fifo_valid_t0),
.out_addr_o(addr_o),
.out_addr_o_t0(addr_o_t0),
.out_err_o(err_o),
.out_err_o_t0(err_o_t0),
.out_err_plus2_o(err_plus2_o),
.out_err_plus2_o_t0(err_plus2_o_t0),
.out_rdata_o(rdata_o),
.out_rdata_o_t0(rdata_o_t0),
.out_ready_i(ready_i),
.out_ready_i_t0(ready_i_t0),
.out_valid_o(valid_o),
.out_valid_o_t0(valid_o_t0),
.rst_ni(rst_ni)
);
assign instr_addr_o = { instr_addr[31:2], 2'h0 };
assign instr_addr_o_t0 = { instr_addr_t0[31:2], 2'h0 };
endmodule

module \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1 (clk_i, rst_ni, en_wb_i, instr_type_wb_i, pc_id_i, instr_is_compressed_id_i, instr_perf_count_id_i, ready_wb_o, rf_write_wb_o, outstanding_load_wb_o, outstanding_store_wb_o, pc_wb_o, perf_instr_ret_wb_o, perf_instr_ret_compressed_wb_o, perf_instr_ret_wb_spec_o, perf_instr_ret_compressed_wb_spec_o, rf_waddr_id_i, rf_wdata_id_i, rf_we_id_i, dummy_instr_id_i, rf_wdata_lsu_i
, rf_we_lsu_i, rf_wdata_fwd_wb_o, rf_waddr_wb_o, rf_wdata_wb_o, rf_we_wb_o, dummy_instr_wb_o, lsu_resp_valid_i, lsu_resp_err_i, instr_done_wb_o, pc_id_i_t0, lsu_resp_valid_i_t0, dummy_instr_id_i_t0, dummy_instr_wb_o_t0, en_wb_i_t0, instr_done_wb_o_t0, instr_is_compressed_id_i_t0, instr_perf_count_id_i_t0, instr_type_wb_i_t0, lsu_resp_err_i_t0, outstanding_load_wb_o_t0, outstanding_store_wb_o_t0
, pc_wb_o_t0, perf_instr_ret_compressed_wb_o_t0, perf_instr_ret_compressed_wb_spec_o_t0, perf_instr_ret_wb_o_t0, perf_instr_ret_wb_spec_o_t0, ready_wb_o_t0, rf_waddr_id_i_t0, rf_waddr_wb_o_t0, rf_wdata_fwd_wb_o_t0, rf_wdata_id_i_t0, rf_wdata_lsu_i_t0, rf_wdata_wb_o_t0, rf_we_id_i_t0, rf_we_lsu_i_t0, rf_we_wb_o_t0, rf_write_wb_o_t0);
/* src = "generated/sv2v_out.v:21025.25-21025.45" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21025.25-21025.45" */
wire _001_;
/* src = "generated/sv2v_out.v:21025.50-21025.71" */
wire _002_;
/* src = "generated/sv2v_out.v:21076.34-21076.62" */
wire _003_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21076.34-21076.62" */
wire _004_;
/* src = "generated/sv2v_out.v:21076.68-21076.101" */
wire _005_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21076.68-21076.101" */
wire _006_;
/* src = "generated/sv2v_out.v:21132.26-21132.75" */
wire [31:0] _007_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21132.26-21132.75" */
wire [31:0] _008_;
/* src = "generated/sv2v_out.v:21132.80-21132.129" */
wire [31:0] _009_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21132.80-21132.129" */
wire [31:0] _010_;
wire _011_;
wire _012_;
wire _013_;
wire [31:0] _014_;
wire _015_;
wire _016_;
wire _017_;
wire [31:0] _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire [31:0] _050_;
wire [31:0] _051_;
wire [31:0] _052_;
wire [31:0] _053_;
wire [31:0] _054_;
wire [31:0] _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire [31:0] _060_;
wire [31:0] _061_;
wire _062_;
wire _063_;
wire [4:0] _064_;
wire [4:0] _065_;
wire [31:0] _066_;
wire [31:0] _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire [31:0] _073_;
wire [31:0] _074_;
wire [31:0] _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire [31:0] _087_;
wire [31:0] _088_;
wire _089_;
wire _090_;
wire [31:0] _091_;
wire _092_;
wire [4:0] _093_;
wire [31:0] _094_;
wire _095_;
wire _096_;
wire [31:0] _097_;
/* src = "generated/sv2v_out.v:21026.22-21026.45" */
wire _098_;
/* src = "generated/sv2v_out.v:21069.55-21069.78" */
wire _099_;
/* src = "generated/sv2v_out.v:21071.50-21071.73" */
wire _100_;
/* src = "generated/sv2v_out.v:21068.24-21068.35" */
wire _101_;
/* src = "generated/sv2v_out.v:21076.66-21076.102" */
wire _102_;
/* src = "generated/sv2v_out.v:21069.41-21069.79" */
wire _103_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21069.41-21069.79" */
wire _104_;
/* src = "generated/sv2v_out.v:20981.13-20981.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:21000.13-21000.29" */
input dummy_instr_id_i;
wire dummy_instr_id_i;
/* cellift = 32'd1 */
input dummy_instr_id_i_t0;
wire dummy_instr_id_i_t0;
/* src = "generated/sv2v_out.v:21007.14-21007.30" */
output dummy_instr_wb_o;
reg dummy_instr_wb_o;
/* cellift = 32'd1 */
output dummy_instr_wb_o_t0;
reg dummy_instr_wb_o_t0;
/* src = "generated/sv2v_out.v:20983.13-20983.20" */
input en_wb_i;
wire en_wb_i;
/* cellift = 32'd1 */
input en_wb_i_t0;
wire en_wb_i_t0;
/* src = "generated/sv2v_out.v:21016.8-21016.18" */
reg \g_writeback_stage.rf_we_wb_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21016.8-21016.18" */
reg \g_writeback_stage.rf_we_wb_q_t0 ;
/* src = "generated/sv2v_out.v:21021.8-21021.23" */
reg \g_writeback_stage.wb_compressed_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21021.8-21021.23" */
reg \g_writeback_stage.wb_compressed_q_t0 ;
/* src = "generated/sv2v_out.v:21018.9-21018.16" */
wire \g_writeback_stage.wb_done ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21018.9-21018.16" */
wire \g_writeback_stage.wb_done_t0 ;
/* src = "generated/sv2v_out.v:21023.14-21023.29" */
reg [1:0] \g_writeback_stage.wb_instr_type_q ;
/* src = "generated/sv2v_out.v:21024.9-21024.19" */
wire \g_writeback_stage.wb_valid_d ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21024.9-21024.19" */
wire \g_writeback_stage.wb_valid_d_t0 ;
/* src = "generated/sv2v_out.v:21019.8-21019.18" */
reg \g_writeback_stage.wb_valid_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21019.8-21019.18" */
reg \g_writeback_stage.wb_valid_q_t0 ;
/* src = "generated/sv2v_out.v:21010.14-21010.29" */
output instr_done_wb_o;
wire instr_done_wb_o;
/* cellift = 32'd1 */
output instr_done_wb_o_t0;
wire instr_done_wb_o_t0;
/* src = "generated/sv2v_out.v:20986.13-20986.37" */
input instr_is_compressed_id_i;
wire instr_is_compressed_id_i;
/* cellift = 32'd1 */
input instr_is_compressed_id_i_t0;
wire instr_is_compressed_id_i_t0;
/* src = "generated/sv2v_out.v:20987.13-20987.34" */
input instr_perf_count_id_i;
wire instr_perf_count_id_i;
/* cellift = 32'd1 */
input instr_perf_count_id_i_t0;
wire instr_perf_count_id_i_t0;
/* src = "generated/sv2v_out.v:20984.19-20984.34" */
input [1:0] instr_type_wb_i;
wire [1:0] instr_type_wb_i;
/* cellift = 32'd1 */
input [1:0] instr_type_wb_i_t0;
wire [1:0] instr_type_wb_i_t0;
/* src = "generated/sv2v_out.v:21009.13-21009.27" */
input lsu_resp_err_i;
wire lsu_resp_err_i;
/* cellift = 32'd1 */
input lsu_resp_err_i_t0;
wire lsu_resp_err_i_t0;
/* src = "generated/sv2v_out.v:21008.13-21008.29" */
input lsu_resp_valid_i;
wire lsu_resp_valid_i;
/* cellift = 32'd1 */
input lsu_resp_valid_i_t0;
wire lsu_resp_valid_i_t0;
/* src = "generated/sv2v_out.v:20990.14-20990.35" */
output outstanding_load_wb_o;
wire outstanding_load_wb_o;
/* cellift = 32'd1 */
output outstanding_load_wb_o_t0;
wire outstanding_load_wb_o_t0;
/* src = "generated/sv2v_out.v:20991.14-20991.36" */
output outstanding_store_wb_o;
wire outstanding_store_wb_o;
/* cellift = 32'd1 */
output outstanding_store_wb_o_t0;
wire outstanding_store_wb_o_t0;
/* src = "generated/sv2v_out.v:20985.20-20985.27" */
input [31:0] pc_id_i;
wire [31:0] pc_id_i;
/* cellift = 32'd1 */
input [31:0] pc_id_i_t0;
wire [31:0] pc_id_i_t0;
/* src = "generated/sv2v_out.v:20992.21-20992.28" */
output [31:0] pc_wb_o;
reg [31:0] pc_wb_o;
/* cellift = 32'd1 */
output [31:0] pc_wb_o_t0;
reg [31:0] pc_wb_o_t0;
/* src = "generated/sv2v_out.v:20994.14-20994.44" */
output perf_instr_ret_compressed_wb_o;
wire perf_instr_ret_compressed_wb_o;
/* cellift = 32'd1 */
output perf_instr_ret_compressed_wb_o_t0;
wire perf_instr_ret_compressed_wb_o_t0;
/* src = "generated/sv2v_out.v:20996.14-20996.49" */
output perf_instr_ret_compressed_wb_spec_o;
wire perf_instr_ret_compressed_wb_spec_o;
/* cellift = 32'd1 */
output perf_instr_ret_compressed_wb_spec_o_t0;
wire perf_instr_ret_compressed_wb_spec_o_t0;
/* src = "generated/sv2v_out.v:20993.14-20993.33" */
output perf_instr_ret_wb_o;
wire perf_instr_ret_wb_o;
/* cellift = 32'd1 */
output perf_instr_ret_wb_o_t0;
wire perf_instr_ret_wb_o_t0;
/* src = "generated/sv2v_out.v:20995.14-20995.38" */
output perf_instr_ret_wb_spec_o;
reg perf_instr_ret_wb_spec_o;
/* cellift = 32'd1 */
output perf_instr_ret_wb_spec_o_t0;
reg perf_instr_ret_wb_spec_o_t0;
/* src = "generated/sv2v_out.v:20988.14-20988.24" */
output ready_wb_o;
wire ready_wb_o;
/* cellift = 32'd1 */
output ready_wb_o_t0;
wire ready_wb_o_t0;
/* src = "generated/sv2v_out.v:20997.19-20997.32" */
input [4:0] rf_waddr_id_i;
wire [4:0] rf_waddr_id_i;
/* cellift = 32'd1 */
input [4:0] rf_waddr_id_i_t0;
wire [4:0] rf_waddr_id_i_t0;
/* src = "generated/sv2v_out.v:21004.20-21004.33" */
output [4:0] rf_waddr_wb_o;
reg [4:0] rf_waddr_wb_o;
/* cellift = 32'd1 */
output [4:0] rf_waddr_wb_o_t0;
reg [4:0] rf_waddr_wb_o_t0;
/* src = "generated/sv2v_out.v:21003.21-21003.38" */
output [31:0] rf_wdata_fwd_wb_o;
reg [31:0] rf_wdata_fwd_wb_o;
/* cellift = 32'd1 */
output [31:0] rf_wdata_fwd_wb_o_t0;
reg [31:0] rf_wdata_fwd_wb_o_t0;
/* src = "generated/sv2v_out.v:20998.20-20998.33" */
input [31:0] rf_wdata_id_i;
wire [31:0] rf_wdata_id_i;
/* cellift = 32'd1 */
input [31:0] rf_wdata_id_i_t0;
wire [31:0] rf_wdata_id_i_t0;
/* src = "generated/sv2v_out.v:21001.20-21001.34" */
input [31:0] rf_wdata_lsu_i;
wire [31:0] rf_wdata_lsu_i;
/* cellift = 32'd1 */
input [31:0] rf_wdata_lsu_i_t0;
wire [31:0] rf_wdata_lsu_i_t0;
/* src = "generated/sv2v_out.v:21012.13-21012.31" */
wire [1:0] rf_wdata_wb_mux_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21012.13-21012.31" */
wire [1:0] rf_wdata_wb_mux_we_t0;
/* src = "generated/sv2v_out.v:21005.21-21005.34" */
output [31:0] rf_wdata_wb_o;
wire [31:0] rf_wdata_wb_o;
/* cellift = 32'd1 */
output [31:0] rf_wdata_wb_o_t0;
wire [31:0] rf_wdata_wb_o_t0;
/* src = "generated/sv2v_out.v:20999.13-20999.23" */
input rf_we_id_i;
wire rf_we_id_i;
/* cellift = 32'd1 */
input rf_we_id_i_t0;
wire rf_we_id_i_t0;
/* src = "generated/sv2v_out.v:21002.13-21002.24" */
input rf_we_lsu_i;
wire rf_we_lsu_i;
/* cellift = 32'd1 */
input rf_we_lsu_i_t0;
wire rf_we_lsu_i_t0;
/* src = "generated/sv2v_out.v:21006.14-21006.24" */
output rf_we_wb_o;
wire rf_we_wb_o;
/* cellift = 32'd1 */
output rf_we_wb_o_t0;
wire rf_we_wb_o_t0;
/* src = "generated/sv2v_out.v:20989.14-20989.27" */
output rf_write_wb_o;
wire rf_write_wb_o;
/* cellift = 32'd1 */
output rf_write_wb_o_t0;
wire rf_write_wb_o_t0;
/* src = "generated/sv2v_out.v:20982.13-20982.19" */
input rst_ni;
wire rst_ni;
assign _000_ = en_wb_i & /* src = "generated/sv2v_out.v:21025.25-21025.45" */ ready_wb_o;
assign _002_ = \g_writeback_stage.wb_valid_q  & /* src = "generated/sv2v_out.v:21025.50-21025.71" */ _016_;
assign rf_wdata_wb_mux_we[0] = \g_writeback_stage.rf_we_wb_q  & /* src = "generated/sv2v_out.v:21067.35-21067.58" */ \g_writeback_stage.wb_valid_q ;
assign rf_write_wb_o = \g_writeback_stage.wb_valid_q  & /* src = "generated/sv2v_out.v:21069.27-21069.80" */ _103_;
assign outstanding_load_wb_o = \g_writeback_stage.wb_valid_q  & /* src = "generated/sv2v_out.v:21070.35-21070.73" */ _099_;
assign outstanding_store_wb_o = \g_writeback_stage.wb_valid_q  & /* src = "generated/sv2v_out.v:21071.36-21071.74" */ _100_;
assign instr_done_wb_o = \g_writeback_stage.wb_valid_q  & /* src = "generated/sv2v_out.v:21073.29-21073.49" */ \g_writeback_stage.wb_done ;
assign perf_instr_ret_compressed_wb_spec_o = perf_instr_ret_wb_spec_o & /* src = "generated/sv2v_out.v:21075.49-21075.91" */ \g_writeback_stage.wb_compressed_q ;
assign _003_ = instr_done_wb_o & /* src = "generated/sv2v_out.v:21076.34-21076.62" */ perf_instr_ret_wb_spec_o;
assign _005_ = lsu_resp_valid_i & /* src = "generated/sv2v_out.v:21076.68-21076.101" */ lsu_resp_err_i;
assign perf_instr_ret_wb_o = _003_ & /* src = "generated/sv2v_out.v:21076.33-21076.102" */ _102_;
assign perf_instr_ret_compressed_wb_o = perf_instr_ret_wb_o & /* src = "generated/sv2v_out.v:21077.44-21077.81" */ \g_writeback_stage.wb_compressed_q ;
assign rf_wdata_wb_mux_we[1] = outstanding_load_wb_o & /* src = "generated/sv2v_out.v:21079.35-21079.70" */ rf_we_lsu_i;
assign _007_ = { rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0] } & /* src = "generated/sv2v_out.v:21132.26-21132.75" */ rf_wdata_fwd_wb_o;
assign _009_ = { rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1] } & /* src = "generated/sv2v_out.v:21132.80-21132.129" */ rf_wdata_lsu_i;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_writeback_stage.wb_valid_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_writeback_stage.wb_valid_q_t0  <= 1'h0;
else \g_writeback_stage.wb_valid_q_t0  <= \g_writeback_stage.wb_valid_d_t0 ;
assign _011_ = ~ en_wb_i;
assign _056_ = en_wb_i & instr_perf_count_id_i_t0;
assign _058_ = en_wb_i & dummy_instr_id_i_t0;
assign _060_ = { en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i } & rf_wdata_id_i_t0;
assign _062_ = en_wb_i & rf_we_id_i_t0;
assign _064_ = { en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i } & rf_waddr_id_i_t0;
assign _066_ = { en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i, en_wb_i } & pc_id_i_t0;
assign _068_ = en_wb_i & instr_is_compressed_id_i_t0;
assign _057_ = _011_ & perf_instr_ret_wb_spec_o_t0;
assign _059_ = _011_ & dummy_instr_wb_o_t0;
assign _061_ = { _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_ } & rf_wdata_fwd_wb_o_t0;
assign _063_ = _011_ & \g_writeback_stage.rf_we_wb_q_t0 ;
assign _065_ = { _011_, _011_, _011_, _011_, _011_ } & rf_waddr_wb_o_t0;
assign _067_ = { _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_ } & pc_wb_o_t0;
assign _069_ = _011_ & \g_writeback_stage.wb_compressed_q_t0 ;
assign _089_ = _056_ | _057_;
assign _090_ = _058_ | _059_;
assign _091_ = _060_ | _061_;
assign _092_ = _062_ | _063_;
assign _093_ = _064_ | _065_;
assign _094_ = _066_ | _067_;
assign _095_ = _068_ | _069_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME perf_instr_ret_wb_spec_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) perf_instr_ret_wb_spec_o_t0 <= 1'h0;
else perf_instr_ret_wb_spec_o_t0 <= _089_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME dummy_instr_wb_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_instr_wb_o_t0 <= 1'h0;
else dummy_instr_wb_o_t0 <= _090_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME rf_wdata_fwd_wb_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rf_wdata_fwd_wb_o_t0 <= 32'd0;
else rf_wdata_fwd_wb_o_t0 <= _091_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_writeback_stage.rf_we_wb_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_writeback_stage.rf_we_wb_q_t0  <= 1'h0;
else \g_writeback_stage.rf_we_wb_q_t0  <= _092_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME rf_waddr_wb_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rf_waddr_wb_o_t0 <= 5'h00;
else rf_waddr_wb_o_t0 <= _093_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME pc_wb_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) pc_wb_o_t0 <= 32'd0;
else pc_wb_o_t0 <= _094_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_writeback_stage.wb_compressed_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_writeback_stage.wb_compressed_q_t0  <= 1'h0;
else \g_writeback_stage.wb_compressed_q_t0  <= _095_;
assign _019_ = en_wb_i_t0 & ready_wb_o;
assign _022_ = \g_writeback_stage.wb_valid_q_t0  & _016_;
assign _025_ = \g_writeback_stage.rf_we_wb_q_t0  & \g_writeback_stage.wb_valid_q ;
assign _028_ = \g_writeback_stage.wb_valid_q_t0  & _103_;
assign outstanding_load_wb_o_t0 = \g_writeback_stage.wb_valid_q_t0  & _099_;
assign outstanding_store_wb_o_t0 = \g_writeback_stage.wb_valid_q_t0  & _100_;
assign _031_ = \g_writeback_stage.wb_valid_q_t0  & \g_writeback_stage.wb_done ;
assign _032_ = perf_instr_ret_wb_spec_o_t0 & \g_writeback_stage.wb_compressed_q ;
assign _035_ = instr_done_wb_o_t0 & perf_instr_ret_wb_spec_o;
assign _038_ = lsu_resp_valid_i_t0 & lsu_resp_err_i;
assign _041_ = _004_ & _102_;
assign _044_ = perf_instr_ret_wb_o_t0 & \g_writeback_stage.wb_compressed_q ;
assign _047_ = outstanding_load_wb_o_t0 & rf_we_lsu_i;
assign _050_ = { rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0] } & rf_wdata_fwd_wb_o;
assign _053_ = { rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1] } & rf_wdata_lsu_i;
assign _020_ = ready_wb_o_t0 & en_wb_i;
assign _023_ = \g_writeback_stage.wb_done_t0  & \g_writeback_stage.wb_valid_q ;
assign _026_ = \g_writeback_stage.wb_valid_q_t0  & \g_writeback_stage.rf_we_wb_q ;
assign _029_ = _104_ & \g_writeback_stage.wb_valid_q ;
assign _033_ = \g_writeback_stage.wb_compressed_q_t0  & perf_instr_ret_wb_spec_o;
assign _036_ = perf_instr_ret_wb_spec_o_t0 & instr_done_wb_o;
assign _039_ = lsu_resp_err_i_t0 & lsu_resp_valid_i;
assign _042_ = _006_ & _003_;
assign _045_ = \g_writeback_stage.wb_compressed_q_t0  & perf_instr_ret_wb_o;
assign _048_ = rf_we_lsu_i_t0 & outstanding_load_wb_o;
assign _051_ = rf_wdata_fwd_wb_o_t0 & { rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0], rf_wdata_wb_mux_we[0] };
assign _054_ = rf_wdata_lsu_i_t0 & { rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1], rf_wdata_wb_mux_we[1] };
assign _021_ = en_wb_i_t0 & ready_wb_o_t0;
assign _024_ = \g_writeback_stage.wb_valid_q_t0  & \g_writeback_stage.wb_done_t0 ;
assign _027_ = \g_writeback_stage.rf_we_wb_q_t0  & \g_writeback_stage.wb_valid_q_t0 ;
assign _030_ = \g_writeback_stage.wb_valid_q_t0  & _104_;
assign _034_ = perf_instr_ret_wb_spec_o_t0 & \g_writeback_stage.wb_compressed_q_t0 ;
assign _037_ = instr_done_wb_o_t0 & perf_instr_ret_wb_spec_o_t0;
assign _040_ = lsu_resp_valid_i_t0 & lsu_resp_err_i_t0;
assign _043_ = _004_ & _006_;
assign _046_ = perf_instr_ret_wb_o_t0 & \g_writeback_stage.wb_compressed_q_t0 ;
assign _049_ = outstanding_load_wb_o_t0 & rf_we_lsu_i_t0;
assign _052_ = { rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0], rf_wdata_wb_mux_we_t0[0] } & rf_wdata_fwd_wb_o_t0;
assign _055_ = { rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1], rf_wdata_wb_mux_we_t0[1] } & rf_wdata_lsu_i_t0;
assign _076_ = _019_ | _020_;
assign _077_ = _022_ | _023_;
assign _078_ = _025_ | _026_;
assign _079_ = _028_ | _029_;
assign _080_ = _031_ | _023_;
assign _081_ = _032_ | _033_;
assign _082_ = _035_ | _036_;
assign _083_ = _038_ | _039_;
assign _084_ = _041_ | _042_;
assign _085_ = _044_ | _045_;
assign _086_ = _047_ | _048_;
assign _087_ = _050_ | _051_;
assign _088_ = _053_ | _054_;
assign _001_ = _076_ | _021_;
assign ready_wb_o_t0 = _077_ | _024_;
assign rf_wdata_wb_mux_we_t0[0] = _078_ | _027_;
assign rf_write_wb_o_t0 = _079_ | _030_;
assign instr_done_wb_o_t0 = _080_ | _024_;
assign perf_instr_ret_compressed_wb_spec_o_t0 = _081_ | _034_;
assign _004_ = _082_ | _037_;
assign _006_ = _083_ | _040_;
assign perf_instr_ret_wb_o_t0 = _084_ | _043_;
assign perf_instr_ret_compressed_wb_o_t0 = _085_ | _046_;
assign rf_wdata_wb_mux_we_t0[1] = _086_ | _049_;
assign _008_ = _087_ | _052_;
assign _010_ = _088_ | _055_;
/* src = "generated/sv2v_out.v:21033.5-21051.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME perf_instr_ret_wb_spec_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) perf_instr_ret_wb_spec_o <= 1'h0;
else if (en_wb_i) perf_instr_ret_wb_spec_o <= instr_perf_count_id_i;
/* src = "generated/sv2v_out.v:21033.5-21051.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_writeback_stage.wb_instr_type_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_writeback_stage.wb_instr_type_q  <= 2'h0;
else if (en_wb_i) \g_writeback_stage.wb_instr_type_q  <= instr_type_wb_i;
/* src = "generated/sv2v_out.v:21083.6-21087.45" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME dummy_instr_wb_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_instr_wb_o <= 1'h0;
else if (en_wb_i) dummy_instr_wb_o <= dummy_instr_id_i;
/* src = "generated/sv2v_out.v:21033.5-21051.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME rf_wdata_fwd_wb_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rf_wdata_fwd_wb_o <= 32'd0;
else if (en_wb_i) rf_wdata_fwd_wb_o <= rf_wdata_id_i;
/* src = "generated/sv2v_out.v:21033.5-21051.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_writeback_stage.rf_we_wb_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_writeback_stage.rf_we_wb_q  <= 1'h0;
else if (en_wb_i) \g_writeback_stage.rf_we_wb_q  <= rf_we_id_i;
/* src = "generated/sv2v_out.v:21033.5-21051.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME rf_waddr_wb_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rf_waddr_wb_o <= 5'h00;
else if (en_wb_i) rf_waddr_wb_o <= rf_waddr_id_i;
/* src = "generated/sv2v_out.v:21033.5-21051.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME pc_wb_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) pc_wb_o <= 32'd0;
else if (en_wb_i) pc_wb_o <= pc_id_i;
/* src = "generated/sv2v_out.v:21033.5-21051.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_writeback_stage.wb_compressed_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_writeback_stage.wb_compressed_q  <= 1'h0;
else if (en_wb_i) \g_writeback_stage.wb_compressed_q  <= instr_is_compressed_id_i;
assign _012_ = ~ _000_;
assign _013_ = ~ _098_;
assign _014_ = ~ _007_;
assign _015_ = ~ _002_;
assign _016_ = ~ \g_writeback_stage.wb_done ;
assign _017_ = ~ _099_;
assign _018_ = ~ _009_;
assign _070_ = _001_ & _015_;
assign _104_ = \g_writeback_stage.rf_we_wb_q_t0  & _017_;
assign _073_ = _008_ & _018_;
assign _071_ = ready_wb_o_t0 & _012_;
assign \g_writeback_stage.wb_done_t0  = lsu_resp_valid_i_t0 & _013_;
assign _074_ = _010_ & _014_;
assign _072_ = _001_ & ready_wb_o_t0;
assign _075_ = _008_ & _010_;
assign _096_ = _070_ | _071_;
assign _097_ = _073_ | _074_;
assign \g_writeback_stage.wb_valid_d_t0  = _096_ | _072_;
assign rf_wdata_wb_o_t0 = _097_ | _075_;
assign _098_ = \g_writeback_stage.wb_instr_type_q  == /* src = "generated/sv2v_out.v:21026.22-21026.45" */ 2'h2;
assign _099_ = ! /* src = "generated/sv2v_out.v:21070.49-21070.72" */ \g_writeback_stage.wb_instr_type_q ;
assign _100_ = \g_writeback_stage.wb_instr_type_q  == /* src = "generated/sv2v_out.v:21071.50-21071.73" */ 2'h1;
assign _101_ = ~ /* src = "generated/sv2v_out.v:21068.24-21068.35" */ \g_writeback_stage.wb_valid_q ;
assign _102_ = ~ /* src = "generated/sv2v_out.v:21076.66-21076.102" */ _005_;
assign \g_writeback_stage.wb_valid_d  = _000_ | /* src = "generated/sv2v_out.v:21025.24-21025.72" */ _002_;
assign \g_writeback_stage.wb_done  = _098_ | /* src = "generated/sv2v_out.v:21026.21-21026.65" */ lsu_resp_valid_i;
assign ready_wb_o = _101_ | /* src = "generated/sv2v_out.v:21068.24-21068.45" */ \g_writeback_stage.wb_done ;
assign _103_ = \g_writeback_stage.rf_we_wb_q  | /* src = "generated/sv2v_out.v:21069.41-21069.79" */ _099_;
assign rf_wdata_wb_o = _007_ | /* src = "generated/sv2v_out.v:21132.25-21132.130" */ _009_;
/* src = "generated/sv2v_out.v:21027.4-21031.31" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'1\DummyInstructions=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_writeback_stage.wb_valid_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_writeback_stage.wb_valid_q  <= 1'h0;
else \g_writeback_stage.wb_valid_q  <= \g_writeback_stage.wb_valid_d ;
assign rf_we_wb_o = | /* src = "generated/sv2v_out.v:21133.22-21133.41" */ rf_wdata_wb_mux_we;
assign rf_we_wb_o_t0 = 1'h0;
endmodule

module \$paramod\prim_buf\Width=32'00000000000000000000000000001100 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23080.22-23080.26" */
input [11:0] in_i;
wire [11:0] in_i;
/* cellift = 32'd1 */
input [11:0] in_i_t0;
wire [11:0] in_i_t0;
/* src = "generated/sv2v_out.v:23081.28-23081.33" */
output [11:0] out_o;
wire [11:0] out_o;
/* cellift = 32'd1 */
output [11:0] out_o_t0;
wire [11:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23091.38-23094.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000001100  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_buf\Width=32'00000000000000000000000000100000 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23080.22-23080.26" */
input [31:0] in_i;
wire [31:0] in_i;
/* cellift = 32'd1 */
input [31:0] in_i_t0;
wire [31:0] in_i_t0;
/* src = "generated/sv2v_out.v:23081.28-23081.33" */
output [31:0] out_o;
wire [31:0] out_o;
/* cellift = 32'd1 */
output [31:0] out_o_t0;
wire [31:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23091.38-23094.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000100000  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_buf\Width=32'00000000000000000000000000100111 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23080.22-23080.26" */
input [38:0] in_i;
wire [38:0] in_i;
/* cellift = 32'd1 */
input [38:0] in_i_t0;
wire [38:0] in_i_t0;
/* src = "generated/sv2v_out.v:23081.28-23081.33" */
output [38:0] out_o;
wire [38:0] out_o;
/* cellift = 32'd1 */
output [38:0] out_o_t0;
wire [38:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23091.38-23094.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000100111  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_buf\Width=s32'00000000000000000000000000000100 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23080.22-23080.26" */
input [3:0] in_i;
wire [3:0] in_i;
/* cellift = 32'd1 */
input [3:0] in_i_t0;
wire [3:0] in_i_t0;
/* src = "generated/sv2v_out.v:23081.28-23081.33" */
output [3:0] out_o;
wire [3:0] out_o;
/* cellift = 32'd1 */
output [3:0] out_o_t0;
wire [3:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23091.38-23094.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000000100  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_buf\Width=s32'00000000000000000000000000000111 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23080.22-23080.26" */
input [6:0] in_i;
wire [6:0] in_i;
/* cellift = 32'd1 */
input [6:0] in_i_t0;
wire [6:0] in_i_t0;
/* src = "generated/sv2v_out.v:23081.28-23081.33" */
output [6:0] out_o;
wire [6:0] out_o;
/* cellift = 32'd1 */
output [6:0] out_o_t0;
wire [6:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23091.38-23094.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000000111  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_buf\Width=s32'00000000000000000000000000100000 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23080.22-23080.26" */
input [31:0] in_i;
wire [31:0] in_i;
/* cellift = 32'd1 */
input [31:0] in_i_t0;
wire [31:0] in_i_t0;
/* src = "generated/sv2v_out.v:23081.28-23081.33" */
output [31:0] out_o;
wire [31:0] out_o;
/* cellift = 32'd1 */
output [31:0] out_o_t0;
wire [31:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23091.38-23094.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000100000  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_generic_buf\Width=s32'00000000000000000000000000000100 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:24927.22-24927.26" */
input [3:0] in_i;
wire [3:0] in_i;
/* cellift = 32'd1 */
input [3:0] in_i_t0;
wire [3:0] in_i_t0;
/* src = "generated/sv2v_out.v:24929.21-24929.24" */
wire [3:0] inv;
/* src = "generated/sv2v_out.v:24928.28-24928.33" */
output [3:0] out_o;
wire [3:0] out_o;
/* cellift = 32'd1 */
output [3:0] out_o_t0;
wire [3:0] out_o_t0;
assign inv = ~ /* src = "generated/sv2v_out.v:24930.15-24930.20" */ in_i;
assign out_o = ~ /* src = "generated/sv2v_out.v:24931.17-24931.21" */ inv;
assign out_o_t0 = in_i_t0;
endmodule

module \$paramod\prim_generic_buf\Width=s32'00000000000000000000000000000111 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:24927.22-24927.26" */
input [6:0] in_i;
wire [6:0] in_i;
/* cellift = 32'd1 */
input [6:0] in_i_t0;
wire [6:0] in_i_t0;
/* src = "generated/sv2v_out.v:24929.21-24929.24" */
wire [6:0] inv;
/* src = "generated/sv2v_out.v:24928.28-24928.33" */
output [6:0] out_o;
wire [6:0] out_o;
/* cellift = 32'd1 */
output [6:0] out_o_t0;
wire [6:0] out_o_t0;
assign inv = ~ /* src = "generated/sv2v_out.v:24930.15-24930.20" */ in_i;
assign out_o = ~ /* src = "generated/sv2v_out.v:24931.17-24931.21" */ inv;
assign out_o_t0 = in_i_t0;
endmodule

module \$paramod\prim_generic_buf\Width=s32'00000000000000000000000000001100 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:24927.22-24927.26" */
input [11:0] in_i;
wire [11:0] in_i;
/* cellift = 32'd1 */
input [11:0] in_i_t0;
wire [11:0] in_i_t0;
/* src = "generated/sv2v_out.v:24929.21-24929.24" */
wire [11:0] inv;
/* src = "generated/sv2v_out.v:24928.28-24928.33" */
output [11:0] out_o;
wire [11:0] out_o;
/* cellift = 32'd1 */
output [11:0] out_o_t0;
wire [11:0] out_o_t0;
assign inv = ~ /* src = "generated/sv2v_out.v:24930.15-24930.20" */ in_i;
assign out_o = ~ /* src = "generated/sv2v_out.v:24931.17-24931.21" */ inv;
assign out_o_t0 = in_i_t0;
endmodule

module \$paramod\prim_generic_buf\Width=s32'00000000000000000000000000100000 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:24927.22-24927.26" */
input [31:0] in_i;
wire [31:0] in_i;
/* cellift = 32'd1 */
input [31:0] in_i_t0;
wire [31:0] in_i_t0;
/* src = "generated/sv2v_out.v:24929.21-24929.24" */
wire [31:0] inv;
/* src = "generated/sv2v_out.v:24928.28-24928.33" */
output [31:0] out_o;
wire [31:0] out_o;
/* cellift = 32'd1 */
output [31:0] out_o_t0;
wire [31:0] out_o_t0;
assign inv = ~ /* src = "generated/sv2v_out.v:24930.15-24930.20" */ in_i;
assign out_o = ~ /* src = "generated/sv2v_out.v:24931.17-24931.21" */ inv;
assign out_o_t0 = in_i_t0;
endmodule

module \$paramod\prim_generic_buf\Width=s32'00000000000000000000000000100111 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:24927.22-24927.26" */
input [38:0] in_i;
wire [38:0] in_i;
/* cellift = 32'd1 */
input [38:0] in_i_t0;
wire [38:0] in_i_t0;
/* src = "generated/sv2v_out.v:24929.21-24929.24" */
wire [38:0] inv;
/* src = "generated/sv2v_out.v:24928.28-24928.33" */
output [38:0] out_o;
wire [38:0] out_o;
/* cellift = 32'd1 */
output [38:0] out_o_t0;
wire [38:0] out_o_t0;
assign inv = ~ /* src = "generated/sv2v_out.v:24930.15-24930.20" */ in_i;
assign out_o = ~ /* src = "generated/sv2v_out.v:24931.17-24931.21" */ inv;
assign out_o_t0 = in_i_t0;
endmodule

module ibex_branch_predict(clk_i, rst_ni, fetch_rdata_i, fetch_pc_i, fetch_valid_i, predict_branch_taken_o, predict_branch_pc_o, predict_branch_taken_o_t0, predict_branch_pc_o_t0, fetch_valid_i_t0, fetch_rdata_i_t0, fetch_pc_i_t0);
/* src = "generated/sv2v_out.v:12093.26-12093.50" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12093.26-12093.50" */
wire _001_;
/* src = "generated/sv2v_out.v:12093.55-12093.81" */
wire _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12093.55-12093.81" */
wire _003_;
wire [31:0] _004_;
wire [31:0] _005_;
wire [31:0] _006_;
wire [31:0] _007_;
wire [31:0] _008_;
wire [31:0] _009_;
wire _010_;
wire _011_;
wire _012_;
wire [31:0] _013_;
wire [31:0] _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire [31:0] _021_;
wire [31:0] _022_;
wire [31:0] _023_;
wire [31:0] _024_;
wire [31:0] _025_;
wire [31:0] _026_;
wire [31:0] _027_;
wire [31:0] _028_;
wire [31:0] _029_;
wire [31:0] _030_;
wire [31:0] _031_;
wire _032_;
wire _033_;
wire [31:0] _034_;
wire [31:0] _035_;
wire [31:0] _036_;
/* src = "generated/sv2v_out.v:12080.21-12080.40" */
wire _037_;
/* src = "generated/sv2v_out.v:12080.46-12080.68" */
wire _038_;
/* src = "generated/sv2v_out.v:12080.73-12080.95" */
wire _039_;
/* src = "generated/sv2v_out.v:12081.46-12081.68" */
wire _040_;
/* src = "generated/sv2v_out.v:12081.73-12081.95" */
wire _041_;
/* src = "generated/sv2v_out.v:12080.45-12080.96" */
wire _042_;
/* src = "generated/sv2v_out.v:12081.45-12081.96" */
wire _043_;
/* src = "generated/sv2v_out.v:12094.52-12094.70" */
wire _044_;
/* src = "generated/sv2v_out.v:12094.51-12094.87" */
wire _045_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12094.51-12094.87" */
wire _046_;
wire [31:0] _047_;
/* cellift = 32'd1 */
wire [31:0] _048_;
wire [31:0] _049_;
/* cellift = 32'd1 */
wire [31:0] _050_;
wire [31:0] _051_;
/* cellift = 32'd1 */
wire [31:0] _052_;
/* src = "generated/sv2v_out.v:12066.13-12066.23" */
wire [31:0] branch_imm;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12066.13-12066.23" */
wire [31:0] branch_imm_t0;
/* src = "generated/sv2v_out.v:12055.13-12055.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:12058.20-12058.30" */
input [31:0] fetch_pc_i;
wire [31:0] fetch_pc_i;
/* cellift = 32'd1 */
input [31:0] fetch_pc_i_t0;
wire [31:0] fetch_pc_i_t0;
/* src = "generated/sv2v_out.v:12057.20-12057.33" */
input [31:0] fetch_rdata_i;
wire [31:0] fetch_rdata_i;
/* cellift = 32'd1 */
input [31:0] fetch_rdata_i_t0;
wire [31:0] fetch_rdata_i_t0;
/* src = "generated/sv2v_out.v:12059.13-12059.26" */
input fetch_valid_i;
wire fetch_valid_i;
/* cellift = 32'd1 */
input fetch_valid_i_t0;
wire fetch_valid_i_t0;
/* src = "generated/sv2v_out.v:12069.7-12069.14" */
wire instr_b;
/* src = "generated/sv2v_out.v:12072.7-12072.20" */
wire instr_b_taken;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12072.7-12072.20" */
wire instr_b_taken_t0;
/* src = "generated/sv2v_out.v:12071.7-12071.15" */
wire instr_cb;
/* src = "generated/sv2v_out.v:12070.7-12070.15" */
wire instr_cj;
/* src = "generated/sv2v_out.v:12068.7-12068.14" */
wire instr_j;
/* src = "generated/sv2v_out.v:12061.21-12061.40" */
output [31:0] predict_branch_pc_o;
wire [31:0] predict_branch_pc_o;
/* cellift = 32'd1 */
output [31:0] predict_branch_pc_o_t0;
wire [31:0] predict_branch_pc_o_t0;
/* src = "generated/sv2v_out.v:12060.14-12060.36" */
output predict_branch_taken_o;
wire predict_branch_taken_o;
/* cellift = 32'd1 */
output predict_branch_taken_o_t0;
wire predict_branch_taken_o_t0;
/* src = "generated/sv2v_out.v:12056.13-12056.19" */
input rst_ni;
wire rst_ni;
assign predict_branch_pc_o = fetch_pc_i + /* src = "generated/sv2v_out.v:12095.31-12095.54" */ branch_imm;
assign instr_cb = _037_ & /* src = "generated/sv2v_out.v:12080.20-12080.97" */ _042_;
assign instr_cj = _037_ & /* src = "generated/sv2v_out.v:12081.20-12081.97" */ _043_;
assign _000_ = instr_b & /* src = "generated/sv2v_out.v:12093.26-12093.50" */ fetch_rdata_i[31];
assign _002_ = instr_cb & /* src = "generated/sv2v_out.v:12093.55-12093.81" */ fetch_rdata_i[12];
assign predict_branch_taken_o = fetch_valid_i & /* src = "generated/sv2v_out.v:12094.34-12094.88" */ _045_;
assign _004_ = ~ fetch_pc_i_t0;
assign _005_ = ~ branch_imm_t0;
assign _013_ = fetch_pc_i & _004_;
assign _014_ = branch_imm & _005_;
assign _035_ = _013_ + _014_;
assign _029_ = fetch_pc_i | fetch_pc_i_t0;
assign _030_ = branch_imm | branch_imm_t0;
assign _036_ = _029_ + _030_;
assign _034_ = _035_ ^ _036_;
assign _031_ = _034_ | fetch_pc_i_t0;
assign predict_branch_pc_o_t0 = _031_ | branch_imm_t0;
assign _015_ = fetch_valid_i_t0 & _045_;
assign _001_ = fetch_rdata_i_t0[31] & instr_b;
assign _003_ = fetch_rdata_i_t0[12] & instr_cb;
assign _016_ = _046_ & fetch_valid_i;
assign _017_ = fetch_valid_i_t0 & _046_;
assign _032_ = _015_ | _016_;
assign predict_branch_taken_o_t0 = _032_ | _017_;
assign _006_ = ~ { instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb };
assign _007_ = ~ { instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj };
assign _008_ = ~ { instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b };
assign _009_ = ~ { instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j };
assign _021_ = _006_ & { fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[7], fetch_rdata_i_t0[30:25], fetch_rdata_i_t0[11:8], 1'h0 };
assign _023_ = _007_ & _048_;
assign _025_ = _008_ & _050_;
assign _027_ = _009_ & _052_;
assign _022_ = { instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb, instr_cb } & { fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[6:5], fetch_rdata_i_t0[2], fetch_rdata_i_t0[11:10], fetch_rdata_i_t0[4:3], 1'h0 };
assign _024_ = { instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj, instr_cj } & { fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[12], fetch_rdata_i_t0[8], fetch_rdata_i_t0[10:9], fetch_rdata_i_t0[6], fetch_rdata_i_t0[7], fetch_rdata_i_t0[2], fetch_rdata_i_t0[11], fetch_rdata_i_t0[5:3], 1'h0 };
assign _026_ = { instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b, instr_b } & { fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[7], fetch_rdata_i_t0[30:25], fetch_rdata_i_t0[11:8], 1'h0 };
assign _028_ = { instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j, instr_j } & { fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[31], fetch_rdata_i_t0[19:12], fetch_rdata_i_t0[20], fetch_rdata_i_t0[30:21], 1'h0 };
assign _048_ = _021_ | _022_;
assign _050_ = _023_ | _024_;
assign _052_ = _025_ | _026_;
assign branch_imm_t0 = _027_ | _028_;
assign _010_ = ~ _000_;
assign _011_ = ~ _044_;
assign _012_ = ~ _002_;
assign _018_ = _001_ & _012_;
assign _019_ = _003_ & _010_;
assign _046_ = instr_b_taken_t0 & _011_;
assign _020_ = _001_ & _003_;
assign _033_ = _018_ | _019_;
assign instr_b_taken_t0 = _033_ | _020_;
assign instr_b = fetch_rdata_i[6:0] == /* src = "generated/sv2v_out.v:12078.19-12078.38" */ 7'h63;
assign instr_j = fetch_rdata_i[6:0] == /* src = "generated/sv2v_out.v:12079.19-12079.38" */ 7'h6f;
assign _038_ = fetch_rdata_i[15:13] == /* src = "generated/sv2v_out.v:12080.46-12080.68" */ 3'h6;
assign _039_ = fetch_rdata_i[15:13] == /* src = "generated/sv2v_out.v:12080.73-12080.95" */ 3'h7;
assign _037_ = fetch_rdata_i[1:0] == /* src = "generated/sv2v_out.v:12081.21-12081.40" */ 2'h1;
assign _040_ = fetch_rdata_i[15:13] == /* src = "generated/sv2v_out.v:12081.46-12081.68" */ 3'h5;
assign _041_ = fetch_rdata_i[15:13] == /* src = "generated/sv2v_out.v:12081.73-12081.95" */ 3'h1;
assign _042_ = _038_ | /* src = "generated/sv2v_out.v:12080.45-12080.96" */ _039_;
assign _043_ = _040_ | /* src = "generated/sv2v_out.v:12081.45-12081.96" */ _041_;
assign instr_b_taken = _000_ | /* src = "generated/sv2v_out.v:12093.25-12093.82" */ _002_;
assign _044_ = instr_j | /* src = "generated/sv2v_out.v:12094.52-12094.70" */ instr_cj;
assign _045_ = _044_ | /* src = "generated/sv2v_out.v:12094.51-12094.87" */ instr_b_taken;
assign _047_ = instr_cb ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12084.3-12091.10" */ { fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[6:5], fetch_rdata_i[2], fetch_rdata_i[11:10], fetch_rdata_i[4:3], 1'h0 } : { fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[7], fetch_rdata_i[30:25], fetch_rdata_i[11:8], 1'h0 };
assign _049_ = instr_cj ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12084.3-12091.10" */ { fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[12], fetch_rdata_i[8], fetch_rdata_i[10:9], fetch_rdata_i[6], fetch_rdata_i[7], fetch_rdata_i[2], fetch_rdata_i[11], fetch_rdata_i[5:3], 1'h0 } : _047_;
assign _051_ = instr_b ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12084.3-12091.10" */ { fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[7], fetch_rdata_i[30:25], fetch_rdata_i[11:8], 1'h0 } : _049_;
assign branch_imm = instr_j ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12084.3-12091.10" */ { fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[31], fetch_rdata_i[19:12], fetch_rdata_i[20], fetch_rdata_i[30:21], 1'h0 } : _051_;
endmodule

module ibex_compressed_decoder(clk_i, rst_ni, valid_i, instr_i, instr_o, is_compressed_o, illegal_instr_o, valid_i_t0, instr_o_t0, instr_i_t0, illegal_instr_o_t0, is_compressed_o_t0);
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire _000_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _001_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _002_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire _003_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _005_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire _006_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire _007_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire _008_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _009_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _010_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire _011_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _013_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire _014_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _015_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _016_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire _017_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _018_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _019_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire _020_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _021_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _022_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _023_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _024_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire _025_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _026_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _027_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire _028_;
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _029_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12115.2-12201.5" */
wire [31:0] _030_;
wire [31:0] _031_;
wire [31:0] _032_;
wire [31:0] _033_;
wire [31:0] _034_;
wire [31:0] _035_;
wire [31:0] _036_;
wire [31:0] _037_;
wire [31:0] _038_;
wire [31:0] _039_;
wire [31:0] _040_;
wire [31:0] _041_;
wire [31:0] _042_;
wire [31:0] _043_;
wire [31:0] _044_;
wire [31:0] _045_;
wire [31:0] _046_;
wire [31:0] _047_;
wire [31:0] _048_;
wire [31:0] _049_;
wire [31:0] _050_;
wire [31:0] _051_;
wire [31:0] _052_;
wire _053_;
wire _054_;
wire _055_;
wire [31:0] _056_;
wire [31:0] _057_;
wire [31:0] _058_;
wire [31:0] _059_;
wire [31:0] _060_;
wire [31:0] _061_;
wire [31:0] _062_;
wire [31:0] _063_;
wire [31:0] _064_;
wire [31:0] _065_;
wire [31:0] _066_;
wire [31:0] _067_;
wire [31:0] _068_;
wire [31:0] _069_;
wire [31:0] _070_;
wire [31:0] _071_;
wire [31:0] _072_;
wire [31:0] _073_;
wire [31:0] _074_;
wire [31:0] _075_;
wire [31:0] _076_;
wire [31:0] _077_;
wire [31:0] _078_;
wire [31:0] _079_;
wire [31:0] _080_;
wire [31:0] _081_;
wire [31:0] _082_;
wire [31:0] _083_;
wire [31:0] _084_;
wire [31:0] _085_;
wire [31:0] _086_;
wire [31:0] _087_;
wire [31:0] _088_;
wire [31:0] _089_;
wire [31:0] _090_;
wire [31:0] _091_;
wire [31:0] _092_;
wire [31:0] _093_;
wire [31:0] _094_;
wire [31:0] _095_;
wire [31:0] _096_;
wire [31:0] _097_;
wire [31:0] _098_;
wire [31:0] _099_;
wire [31:0] _100_;
wire [31:0] _101_;
wire [31:0] _102_;
wire [31:0] _103_;
wire [31:0] _104_;
wire [31:0] _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire [31:0] _113_;
/* cellift = 32'd1 */
wire [31:0] _114_;
wire [31:0] _115_;
/* cellift = 32'd1 */
wire [31:0] _116_;
wire [31:0] _117_;
/* cellift = 32'd1 */
wire [31:0] _118_;
wire [31:0] _119_;
/* cellift = 32'd1 */
wire [31:0] _120_;
wire [31:0] _121_;
/* cellift = 32'd1 */
wire [31:0] _122_;
wire [31:0] _123_;
/* cellift = 32'd1 */
wire [31:0] _124_;
wire _125_;
wire [31:0] _126_;
/* cellift = 32'd1 */
wire [31:0] _127_;
wire [31:0] _128_;
/* cellift = 32'd1 */
wire [31:0] _129_;
wire [31:0] _130_;
/* cellift = 32'd1 */
wire [31:0] _131_;
wire [31:0] _132_;
/* cellift = 32'd1 */
wire [31:0] _133_;
wire [31:0] _134_;
/* cellift = 32'd1 */
wire [31:0] _135_;
wire _136_;
wire _137_;
wire [31:0] _138_;
/* cellift = 32'd1 */
wire [31:0] _139_;
wire [31:0] _140_;
/* cellift = 32'd1 */
wire [31:0] _141_;
wire _142_;
wire _143_;
wire [31:0] _144_;
/* cellift = 32'd1 */
wire [31:0] _145_;
wire [31:0] _146_;
/* cellift = 32'd1 */
wire [31:0] _147_;
/* src = "generated/sv2v_out.v:12123.11-12123.39" */
wire _148_;
/* src = "generated/sv2v_out.v:12138.11-12138.33" */
wire _149_;
/* src = "generated/sv2v_out.v:12140.11-12140.51" */
wire _150_;
/* src = "generated/sv2v_out.v:12174.11-12174.36" */
wire _151_;
/* src = "generated/sv2v_out.v:12179.12-12179.36" */
wire _152_;
/* src = "generated/sv2v_out.v:12134.164-12134.176" */
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire [3:0] _158_;
wire _159_;
wire _160_;
wire [3:0] _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
/* src = "generated/sv2v_out.v:12106.13-12106.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:12112.13-12112.28" */
output illegal_instr_o;
wire illegal_instr_o;
/* cellift = 32'd1 */
output illegal_instr_o_t0;
wire illegal_instr_o_t0;
/* src = "generated/sv2v_out.v:12109.20-12109.27" */
input [31:0] instr_i;
wire [31:0] instr_i;
/* cellift = 32'd1 */
input [31:0] instr_i_t0;
wire [31:0] instr_i_t0;
/* src = "generated/sv2v_out.v:12110.20-12110.27" */
output [31:0] instr_o;
wire [31:0] instr_o;
/* cellift = 32'd1 */
output [31:0] instr_o_t0;
wire [31:0] instr_o_t0;
/* src = "generated/sv2v_out.v:12111.14-12111.29" */
output is_compressed_o;
wire is_compressed_o;
/* cellift = 32'd1 */
output is_compressed_o_t0;
wire is_compressed_o_t0;
/* src = "generated/sv2v_out.v:12107.13-12107.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:12108.13-12108.20" */
input valid_i;
wire valid_i;
/* cellift = 32'd1 */
input valid_i_t0;
wire valid_i_t0;
assign _031_ = ~ { _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_ };
assign _033_ = ~ { _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_ };
assign _034_ = ~ { _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_ };
assign _035_ = ~ { _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_ };
assign _036_ = ~ { _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_ };
assign _037_ = ~ { _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_ };
assign _038_ = ~ { _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_ };
assign _039_ = ~ { _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_ };
assign _040_ = ~ { _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_ };
assign _041_ = ~ { _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_ };
assign _042_ = ~ { _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_ };
assign _043_ = ~ { _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_ };
assign _044_ = ~ { _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_ };
assign _032_ = ~ { _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_ };
assign _045_ = ~ { _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_ };
assign _046_ = ~ { _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_ };
assign _047_ = ~ { _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_ };
assign _048_ = ~ { _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_ };
assign _049_ = ~ { _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_, _151_ };
assign _050_ = ~ { _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_ };
assign _051_ = ~ { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12] };
assign _052_ = ~ { _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_ };
assign _056_ = _031_ & { 4'h0, instr_i_t0[8:7], instr_i_t0[12], instr_i_t0[6:2], 8'h00, instr_i_t0[11:9], 9'h000 };
assign _058_ = _032_ & { 7'h00, instr_i_t0[6:2], instr_i_t0[11:7], 3'h0, instr_i_t0[11:7], 7'h00 };
assign _060_ = _033_ & _116_;
assign _062_ = _034_ & _118_;
assign _064_ = _035_ & { 9'h000, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 };
assign _066_ = _036_ & { 9'h000, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 };
assign _068_ = _037_ & _122_;
assign _070_ = _038_ & _124_;
assign _072_ = _039_ & { 1'h0, instr_i_t0[10], 5'h00, instr_i_t0[6:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 };
assign _074_ = _040_ & _127_;
assign _076_ = _033_ & _016_;
assign _078_ = _041_ & _129_;
assign _080_ = _042_ & { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:2], instr_i_t0[11:7], 3'h0, instr_i_t0[11:7], 7'h00 };
assign _082_ = _032_ & _133_;
assign _084_ = _043_ & _135_;
assign _086_ = _044_ & { 5'h00, instr_i_t0[5], instr_i_t0[12], 2'h0, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 3'h0, instr_i_t0[11:10], instr_i_t0[6], 9'h000 };
assign _088_ = _032_ & { 2'h0, instr_i_t0[10:7], instr_i_t0[12:11], instr_i_t0[5], instr_i_t0[6], 12'h000, instr_i_t0[4:2], 7'h00 };
assign _090_ = _045_ & _141_;
assign _092_ = _046_ & _024_;
assign _094_ = _047_ & _010_;
assign _096_ = _048_ & _147_;
assign _005_ = _049_ & { 12'h000, instr_i_t0[11:7], 15'h0000 };
assign _098_ = _050_ & _005_;
assign _100_ = _050_ & { 12'h000, instr_i_t0[11:7], 15'h0000 };
assign _102_ = _051_ & _030_;
assign _104_ = _052_ & { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:2], instr_i_t0[11:7], 7'h00 };
assign _057_ = { _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_, _159_ } & instr_i_t0;
assign _059_ = { _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_ } & { 4'h0, instr_i_t0[3:2], instr_i_t0[12], instr_i_t0[6:4], 10'h000, instr_i_t0[11:7], 7'h00 };
assign _061_ = { _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_ } & _027_;
assign _063_ = { _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_, _106_ } & _114_;
assign _065_ = { _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_, _162_ } & instr_i_t0;
assign _067_ = { _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_, _165_ } & { 9'h000, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 };
assign _069_ = { _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_, _164_ } & { 9'h000, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 };
assign _071_ = { _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_, _107_ } & _120_;
assign _073_ = { _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_, _168_ } & { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 };
assign _075_ = { _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_, _166_ } & _022_;
assign _077_ = { _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_, _154_ } & _019_;
assign _079_ = { _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_, _169_ } & { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:5], instr_i_t0[2], 7'h00, instr_i_t0[9:7], 2'h0, instr_i_t0[13], instr_i_t0[11:10], instr_i_t0[4:3], instr_i_t0[12], 7'h00 };
assign _081_ = { _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_, _170_ } & { instr_i_t0[12], instr_i_t0[8], instr_i_t0[10:9], instr_i_t0[6], instr_i_t0[7], instr_i_t0[2], instr_i_t0[11], instr_i_t0[5:3], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], 4'h0, instr_i_t0[15], 7'h00 };
assign _083_ = { _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_ } & { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:2], 8'h00, instr_i_t0[11:7], 7'h00 };
assign _085_ = { _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_, _053_ } & _131_;
assign _087_ = { _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_, _171_ } & instr_i_t0;
assign _089_ = { _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_, _156_ } & { 5'h00, instr_i_t0[5], instr_i_t0[12:10], instr_i_t0[6], 4'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[4:2], 7'h00 };
assign _091_ = { _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_, _108_ } & _139_;
assign _093_ = { _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_, _172_ } & instr_i_t0;
assign _095_ = { _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_, _167_ } & _013_;
assign _097_ = { _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_, _109_ } & _145_;
assign _099_ = { _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_ } & { 7'h00, instr_i_t0[6:2], instr_i_t0[11:7], 3'h0, instr_i_t0[11:7], 7'h00 };
assign _101_ = { _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_, _152_ } & { 7'h00, instr_i_t0[6:2], 8'h00, instr_i_t0[11:7], 7'h00 };
assign _103_ = { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12] } & _002_;
assign _105_ = { _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_, _149_ } & { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[4:3], instr_i_t0[5], instr_i_t0[2], instr_i_t0[6], 24'h000000 };
assign _114_ = _056_ | _057_;
assign _116_ = _058_ | _059_;
assign _118_ = _060_ | _061_;
assign _024_ = _062_ | _063_;
assign _120_ = _064_ | _065_;
assign _122_ = _066_ | _067_;
assign _124_ = _068_ | _069_;
assign _022_ = _070_ | _071_;
assign _127_ = _072_ | _073_;
assign _019_ = _074_ | _075_;
assign _129_ = _076_ | _077_;
assign _131_ = _078_ | _079_;
assign _133_ = _080_ | _081_;
assign _135_ = _082_ | _083_;
assign _013_ = _084_ | _085_;
assign _139_ = _086_ | _087_;
assign _141_ = _088_ | _089_;
assign _010_ = _090_ | _091_;
assign _145_ = _092_ | _093_;
assign _147_ = _094_ | _095_;
assign instr_o_t0 = _096_ | _097_;
assign _002_ = _098_ | _099_;
assign _030_ = _100_ | _101_;
assign _027_ = _102_ | _103_;
assign _016_ = _104_ | _105_;
assign _054_ = | { _160_, _156_ };
assign _055_ = | { _160_, _158_[3:2], _158_[0], _157_, _156_ };
assign _106_ = _160_ | _159_;
assign _107_ = _163_ | _162_;
assign _108_ = _160_ | _171_;
assign _109_ = _155_ | _172_;
assign _053_ = | { _160_, _158_[3], _158_[1], _154_ };
assign _110_ = _159_ ? 1'h1 : 1'h0;
assign _111_ = _156_ ? _003_ : _000_;
assign _112_ = _154_ ? _006_ : _111_;
assign _028_ = _106_ ? _110_ : _112_;
assign _113_ = _159_ ? instr_i : { 4'h0, instr_i[8:7], instr_i[12], instr_i[6:2], 8'h12, instr_i[11:9], 9'h023 };
assign _115_ = _156_ ? { 4'h0, instr_i[3:2], instr_i[12], instr_i[6:4], 10'h012, instr_i[11:7], 7'h03 } : { 7'h00, instr_i[6:2], instr_i[11:7], 3'h1, instr_i[11:7], 7'h13 };
assign _117_ = _154_ ? _026_ : _115_;
assign _023_ = _106_ ? _113_ : _117_;
assign _119_ = _162_ ? instr_i : { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h1d, instr_i[9:7], 7'h33 };
assign _121_ = _165_ ? { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h11, instr_i[9:7], 7'h33 } : { 9'h081, instr_i[4:2], 2'h1, instr_i[9:7], 5'h01, instr_i[9:7], 7'h33 };
assign _123_ = _164_ ? { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h19, instr_i[9:7], 7'h33 } : _121_;
assign _021_ = _107_ ? _119_ : _123_;
assign _025_ = _162_ ? 1'h1 : 1'h0;
assign _125_ = _168_ ? 1'h0 : _000_;
assign _020_ = _166_ ? _025_ : _125_;
assign _126_ = _168_ ? { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], 2'h1, instr_i[9:7], 5'h1d, instr_i[9:7], 7'h13 } : { 1'h0, instr_i[10], 5'h00, instr_i[6:2], 2'h1, instr_i[9:7], 5'h15, instr_i[9:7], 7'h13 };
assign _018_ = _166_ ? _021_ : _126_;
assign _128_ = _154_ ? _018_ : _015_;
assign _130_ = _169_ ? { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:5], instr_i[2], 7'h01, instr_i[9:7], 2'h0, instr_i[13], instr_i[11:10], instr_i[4:3], instr_i[12], 7'h63 } : _128_;
assign _132_ = _170_ ? { instr_i[12], instr_i[8], instr_i[10:9], instr_i[6], instr_i[7], instr_i[2], instr_i[11], instr_i[5:3], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], 4'h0, _153_, 7'h6f } : { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], instr_i[11:7], 3'h0, instr_i[11:7], 7'h13 };
assign _134_ = _156_ ? { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], 8'h00, instr_i[11:7], 7'h13 } : _132_;
assign _012_ = _053_ ? _130_ : _134_;
assign _136_ = _154_ ? _020_ : _017_;
assign _014_ = _055_ ? 1'h0 : _136_;
assign _137_ = _054_ ? 1'h0 : _011_;
assign _008_ = _171_ ? 1'h1 : _137_;
assign _138_ = _171_ ? instr_i : { 5'h00, instr_i[5], instr_i[12], 2'h1, instr_i[4:2], 2'h1, instr_i[9:7], 3'h2, instr_i[11:10], instr_i[6], 9'h023 };
assign _140_ = _156_ ? { 5'h00, instr_i[5], instr_i[12:10], instr_i[6], 4'h1, instr_i[9:7], 5'h09, instr_i[4:2], 7'h03 } : { 2'h0, instr_i[10:7], instr_i[12:11], instr_i[5], instr_i[6], 12'h041, instr_i[4:2], 7'h13 };
assign _009_ = _108_ ? _138_ : _140_;
assign _142_ = _172_ ? 1'h0 : _028_;
assign _143_ = _167_ ? _014_ : _008_;
assign illegal_instr_o = _109_ ? _142_ : _143_;
assign _144_ = _172_ ? instr_i : _023_;
assign _146_ = _167_ ? _012_ : _009_;
assign instr_o = _109_ ? _144_ : _146_;
assign _148_ = ! /* src = "generated/sv2v_out.v:12123.11-12123.39" */ instr_i[12:5];
assign _149_ = instr_i[11:7] == /* src = "generated/sv2v_out.v:12138.11-12138.33" */ 5'h02;
assign _150_ = ! /* src = "generated/sv2v_out.v:12140.11-12140.51" */ { instr_i[12], instr_i[6:2] };
assign _151_ = ! /* src = "generated/sv2v_out.v:12189.16-12189.41" */ instr_i[11:7];
assign _152_ = | /* src = "generated/sv2v_out.v:12187.16-12187.40" */ instr_i[6:2];
assign is_compressed_o = instr_i[1:0] != /* src = "generated/sv2v_out.v:12202.27-12202.48" */ 2'h3;
assign _153_ = ~ /* src = "generated/sv2v_out.v:12134.164-12134.176" */ instr_i[15];
assign _004_ = _151_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12189.16-12189.41|generated/sv2v_out.v:12189.12-12192.77" */ 32'd1048691 : { 12'h000, instr_i[11:7], 15'h00e7 };
assign _001_ = _152_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12187.16-12187.40|generated/sv2v_out.v:12187.12-12192.77" */ { 7'h00, instr_i[6:2], instr_i[11:7], 3'h0, instr_i[11:7], 7'h33 } : _004_;
assign _029_ = _152_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12179.12-12179.36|generated/sv2v_out.v:12179.8-12185.11" */ { 7'h00, instr_i[6:2], 8'h00, instr_i[11:7], 7'h33 } : { 12'h000, instr_i[11:7], 15'h0067 };
assign _007_ = _152_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12179.12-12179.36|generated/sv2v_out.v:12179.8-12185.11" */ 1'h0 : _003_;
assign _006_ = instr_i[12] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12178.11-12178.30|generated/sv2v_out.v:12178.7-12192.77" */ 1'h0 : _007_;
assign _026_ = instr_i[12] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12178.11-12178.30|generated/sv2v_out.v:12178.7-12192.77" */ _001_ : _029_;
assign _003_ = _151_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12174.11-12174.36|generated/sv2v_out.v:12174.7-12175.31" */ 1'h1 : 1'h0;
assign _000_ = instr_i[12] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12169.11-12169.30|generated/sv2v_out.v:12169.7-12170.31" */ 1'h1 : 1'h0;
assign _159_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12166.5-12196.12" */ _158_;
assign _162_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12152.9-12159.16" */ _161_;
assign _161_[0] = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12152.9-12159.16" */ 3'h4;
assign _161_[1] = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12152.9-12159.16" */ 3'h5;
assign _161_[2] = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12152.9-12159.16" */ 3'h6;
assign _161_[3] = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12152.9-12159.16" */ 3'h7;
assign _163_ = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12152.9-12159.16" */ 3'h3;
assign _164_ = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12152.9-12159.16" */ 3'h2;
assign _165_ = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12152.9-12159.16" */ 3'h1;
assign _166_ = instr_i[11:10] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12144.7-12161.14" */ 2'h3;
assign _168_ = instr_i[11:10] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12144.7-12161.14" */ 2'h2;
assign _017_ = _150_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12140.11-12140.51|generated/sv2v_out.v:12140.7-12141.31" */ 1'h1 : 1'h0;
assign _015_ = _149_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12138.11-12138.33|generated/sv2v_out.v:12138.7-12139.126" */ { instr_i[12], instr_i[12], instr_i[12], instr_i[4:3], instr_i[5], instr_i[2], instr_i[6], 24'h010113 } : { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], instr_i[11:7], 7'h37 };
assign _169_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12132.5-12164.12" */ { _160_, _158_[3] };
assign _170_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12132.5-12164.12" */ { _158_[2], _158_[0] };
assign _011_ = _148_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12123.11-12123.39|generated/sv2v_out.v:12123.7-12124.31" */ 1'h1 : 1'h0;
assign _171_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12120.5-12130.12" */ { _158_, _154_ };
assign _158_[0] = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12120.5-12130.12" */ 3'h1;
assign _158_[1] = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12120.5-12130.12" */ 3'h3;
assign _154_ = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12120.5-12130.12" */ 3'h4;
assign _158_[2] = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12120.5-12130.12" */ 3'h5;
assign _158_[3] = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12120.5-12130.12" */ 3'h7;
assign _160_ = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12120.5-12130.12" */ 3'h6;
assign _156_ = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12120.5-12130.12" */ 3'h2;
assign _157_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12120.5-12130.12" */ instr_i[15:13];
assign _167_ = instr_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12118.3-12200.10" */ 2'h1;
assign _172_ = instr_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12118.3-12200.10" */ 2'h3;
assign _155_ = instr_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12118.3-12200.10" */ 2'h2;
assign illegal_instr_o_t0 = 1'h0;
assign is_compressed_o_t0 = 1'h0;
endmodule

module ibex_multdiv_slow(clk_i, rst_ni, mult_en_i, div_en_i, mult_sel_i, div_sel_i, operator_i, signed_mode_i, op_a_i, op_b_i, alu_adder_ext_i, alu_adder_i, equal_to_zero_i, data_ind_timing_i, alu_operand_a_o, alu_operand_b_o, imd_val_q_i, imd_val_d_o, imd_val_we_o, multdiv_ready_id_i, multdiv_result_o
, valid_o, data_ind_timing_i_t0, alu_adder_ext_i_t0, alu_adder_i_t0, alu_operand_a_o_t0, alu_operand_b_o_t0, div_en_i_t0, div_sel_i_t0, equal_to_zero_i_t0, imd_val_d_o_t0, imd_val_q_i_t0, imd_val_we_o_t0, mult_en_i_t0, mult_sel_i_t0, multdiv_ready_id_i_t0, multdiv_result_o_t0, op_a_i_t0, op_b_i_t0, operator_i_t0, signed_mode_i_t0, valid_o_t0
);
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _001_;
/* src = "generated/sv2v_out.v:19607.2-19640.5" */
wire [32:0] _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19607.2-19640.5" */
wire [32:0] _003_;
/* src = "generated/sv2v_out.v:19607.2-19640.5" */
wire [32:0] _004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19607.2-19640.5" */
wire [32:0] _005_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [2:0] _006_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [4:0] _007_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire _008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire _009_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _011_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _013_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [31:0] _014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [31:0] _015_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _016_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _017_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire _018_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [2:0] _019_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire _020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire _021_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _022_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _023_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _024_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _025_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _026_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _027_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [2:0] _028_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _029_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _030_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _031_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _032_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _033_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _034_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [2:0] _035_;
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _036_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19654.2-19766.5" */
wire [32:0] _037_;
/* src = "generated/sv2v_out.v:19669.55-19669.88" */
wire [31:0] _038_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19669.55-19669.88" */
wire [31:0] _039_;
/* src = "generated/sv2v_out.v:19669.28-19669.52" */
wire _040_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19669.28-19669.52" */
wire _041_;
/* src = "generated/sv2v_out.v:19675.61-19675.94" */
wire [30:0] _042_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19675.61-19675.94" */
wire [30:0] _043_;
/* src = "generated/sv2v_out.v:19783.43-19783.111" */
wire _044_;
wire _045_;
wire _046_;
wire [32:0] _047_;
wire [32:0] _048_;
wire _049_;
wire [32:0] _050_;
wire [32:0] _051_;
wire [32:0] _052_;
wire [32:0] _053_;
wire [32:0] _054_;
wire [32:0] _055_;
wire [32:0] _056_;
wire [32:0] _057_;
wire [32:0] _058_;
wire [32:0] _059_;
wire _060_;
wire [32:0] _061_;
wire [31:0] _062_;
wire [31:0] _063_;
wire [32:0] _064_;
wire [32:0] _065_;
wire [31:0] _066_;
wire [32:0] _067_;
wire [31:0] _068_;
wire [32:0] _069_;
wire [32:0] _070_;
wire [32:0] _071_;
wire [31:0] _072_;
wire [32:0] _073_;
wire _074_;
wire [32:0] _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire [31:0] _096_;
wire [31:0] _097_;
wire [31:0] _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire [31:0] _108_;
wire [31:0] _109_;
wire [31:0] _110_;
wire [30:0] _111_;
wire [30:0] _112_;
wire [30:0] _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire [32:0] _120_;
wire [32:0] _121_;
wire [32:0] _122_;
wire [32:0] _123_;
wire [32:0] _124_;
wire [32:0] _125_;
wire [32:0] _126_;
wire [32:0] _127_;
wire [32:0] _128_;
wire [32:0] _129_;
wire [32:0] _130_;
wire [32:0] _131_;
wire [32:0] _132_;
wire [32:0] _133_;
wire [32:0] _134_;
wire [32:0] _135_;
wire [32:0] _136_;
wire [32:0] _137_;
wire [32:0] _138_;
wire [32:0] _139_;
wire [32:0] _140_;
wire [32:0] _141_;
wire [32:0] _142_;
wire [32:0] _143_;
wire [32:0] _144_;
wire [32:0] _145_;
wire [32:0] _146_;
wire [32:0] _147_;
wire [32:0] _148_;
wire [32:0] _149_;
wire [32:0] _150_;
wire [32:0] _151_;
wire [32:0] _152_;
wire [32:0] _153_;
wire [32:0] _154_;
wire [32:0] _155_;
wire [32:0] _156_;
wire [32:0] _157_;
wire [32:0] _158_;
wire [32:0] _159_;
wire _160_;
wire _161_;
wire [32:0] _162_;
wire [32:0] _163_;
wire [32:0] _164_;
wire [32:0] _165_;
wire [32:0] _166_;
wire [32:0] _167_;
wire [32:0] _168_;
wire [32:0] _169_;
wire [32:0] _170_;
wire [32:0] _171_;
wire [32:0] _172_;
wire [32:0] _173_;
wire [32:0] _174_;
wire [32:0] _175_;
wire [32:0] _176_;
wire _177_;
wire _178_;
wire _179_;
wire [31:0] _180_;
wire [31:0] _181_;
wire [31:0] _182_;
wire [31:0] _183_;
wire [32:0] _184_;
wire [32:0] _185_;
wire [32:0] _186_;
wire [32:0] _187_;
wire [31:0] _188_;
wire [31:0] _189_;
wire [32:0] _190_;
wire [32:0] _191_;
wire [31:0] _192_;
wire [31:0] _193_;
wire [32:0] _194_;
wire [32:0] _195_;
wire [32:0] _196_;
wire [32:0] _197_;
wire [32:0] _198_;
wire [32:0] _199_;
wire [31:0] _200_;
wire [31:0] _201_;
wire _202_;
wire _203_;
wire _204_;
wire [31:0] _205_;
wire _206_;
wire _207_;
wire _208_;
wire [31:0] _209_;
wire [30:0] _210_;
wire _211_;
wire _212_;
wire [32:0] _213_;
wire [32:0] _214_;
wire [32:0] _215_;
wire _216_;
wire [32:0] _217_;
/* cellift = 32'd1 */
wire [32:0] _218_;
wire [32:0] _219_;
/* cellift = 32'd1 */
wire [32:0] _220_;
wire [32:0] _221_;
/* cellift = 32'd1 */
wire [32:0] _222_;
wire [2:0] _223_;
wire [32:0] _224_;
/* cellift = 32'd1 */
wire [32:0] _225_;
wire [32:0] _226_;
/* cellift = 32'd1 */
wire [32:0] _227_;
wire [32:0] _228_;
/* cellift = 32'd1 */
wire [32:0] _229_;
wire [32:0] _230_;
/* cellift = 32'd1 */
wire [32:0] _231_;
wire [32:0] _232_;
/* cellift = 32'd1 */
wire [32:0] _233_;
wire [32:0] _234_;
/* cellift = 32'd1 */
wire [32:0] _235_;
wire [32:0] _236_;
/* cellift = 32'd1 */
wire [32:0] _237_;
wire [32:0] _238_;
/* cellift = 32'd1 */
wire [32:0] _239_;
wire [2:0] _240_;
wire [2:0] _241_;
wire [2:0] _242_;
wire [2:0] _243_;
wire [2:0] _244_;
wire _245_;
/* cellift = 32'd1 */
wire _246_;
wire [32:0] _247_;
/* cellift = 32'd1 */
wire [32:0] _248_;
wire [32:0] _249_;
/* cellift = 32'd1 */
wire [32:0] _250_;
wire [32:0] _251_;
/* cellift = 32'd1 */
wire [32:0] _252_;
/* src = "generated/sv2v_out.v:19611.29-19611.47" */
wire _253_;
/* src = "generated/sv2v_out.v:19648.29-19648.67" */
wire _254_;
/* src = "generated/sv2v_out.v:19671.45-19671.65" */
wire _255_;
/* src = "generated/sv2v_out.v:19710.46-19710.63" */
wire _256_;
/* src = "generated/sv2v_out.v:19710.70-19710.93" */
wire _257_;
/* src = "generated/sv2v_out.v:19783.20-19783.38" */
wire _258_;
/* src = "generated/sv2v_out.v:19783.68-19783.86" */
wire _259_;
/* src = "generated/sv2v_out.v:19783.91-19783.109" */
wire _260_;
/* src = "generated/sv2v_out.v:19671.22-19671.66" */
wire _261_;
/* src = "generated/sv2v_out.v:19681.22-19681.59" */
wire _262_;
/* src = "generated/sv2v_out.v:19710.23-19710.64" */
wire _263_;
/* src = "generated/sv2v_out.v:19671.22-19671.40" */
wire _264_;
/* src = "generated/sv2v_out.v:19663.7-19663.30" */
wire _265_;
/* src = "generated/sv2v_out.v:19710.22-19710.94" */
wire _266_;
/* src = "generated/sv2v_out.v:19616.26-19616.33" */
wire [31:0] _267_;
/* src = "generated/sv2v_out.v:19620.26-19620.33" */
wire [31:0] _268_;
/* src = "generated/sv2v_out.v:19628.26-19628.47" */
wire [31:0] _269_;
/* src = "generated/sv2v_out.v:19632.26-19632.45" */
wire [31:0] _270_;
/* src = "generated/sv2v_out.v:19648.70-19648.86" */
wire _271_;
/* src = "generated/sv2v_out.v:19652.47-19652.61" */
wire _272_;
/* src = "generated/sv2v_out.v:19669.26-19669.53" */
wire _273_;
/* src = "generated/sv2v_out.v:19732.23-19732.42" */
wire _274_;
/* src = "generated/sv2v_out.v:19651.45-19651.69" */
wire [32:0] _275_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19651.45-19651.69" */
wire [32:0] _276_;
/* src = "generated/sv2v_out.v:19767.23-19767.43" */
wire _277_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19767.23-19767.43" */
wire _278_;
/* src = "generated/sv2v_out.v:19783.67-19783.110" */
wire _279_;
wire _280_;
wire _281_;
wire _282_;
wire _283_;
wire _284_;
wire _285_;
wire _286_;
/* src = "generated/sv2v_out.v:0.0-0.0" */
wire _287_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:0.0-0.0" */
wire _288_;
/* src = "generated/sv2v_out.v:19704.24-19704.47" */
wire [4:0] _289_;
/* src = "generated/sv2v_out.v:19611.29-19611.78" */
wire [32:0] _290_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19611.29-19611.78" */
wire [32:0] _291_;
/* src = "generated/sv2v_out.v:19671.22-19671.80" */
wire [2:0] _292_;
/* src = "generated/sv2v_out.v:19681.22-19681.73" */
wire [2:0] _293_;
/* src = "generated/sv2v_out.v:19695.24-19695.53" */
wire [31:0] _294_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19695.24-19695.53" */
wire [31:0] _295_;
/* src = "generated/sv2v_out.v:19700.22-19700.67" */
wire [32:0] _296_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19700.22-19700.67" */
wire [32:0] _297_;
/* src = "generated/sv2v_out.v:19710.22-19710.108" */
wire [2:0] _298_;
/* src = "generated/sv2v_out.v:19716.22-19716.59" */
wire [2:0] _299_;
/* src = "generated/sv2v_out.v:19754.31-19754.85" */
wire [32:0] _300_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19754.31-19754.85" */
wire [32:0] _301_;
/* src = "generated/sv2v_out.v:19755.31-19755.85" */
wire [32:0] _302_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19755.31-19755.85" */
wire [32:0] _303_;
/* src = "generated/sv2v_out.v:19652.28-19652.43" */
wire _304_;
/* src = "generated/sv2v_out.v:19567.13-19567.27" */
wire [32:0] accum_window_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19567.13-19567.27" */
wire [32:0] accum_window_d_t0;
/* src = "generated/sv2v_out.v:19552.20-19552.35" */
input [33:0] alu_adder_ext_i;
wire [33:0] alu_adder_ext_i;
/* cellift = 32'd1 */
input [33:0] alu_adder_ext_i_t0;
wire [33:0] alu_adder_ext_i_t0;
/* src = "generated/sv2v_out.v:19553.20-19553.31" */
input [31:0] alu_adder_i;
wire [31:0] alu_adder_i;
/* cellift = 32'd1 */
input [31:0] alu_adder_i_t0;
wire [31:0] alu_adder_i_t0;
/* src = "generated/sv2v_out.v:19556.20-19556.35" */
output [32:0] alu_operand_a_o;
wire [32:0] alu_operand_a_o;
/* cellift = 32'd1 */
output [32:0] alu_operand_a_o_t0;
wire [32:0] alu_operand_a_o_t0;
/* src = "generated/sv2v_out.v:19557.20-19557.35" */
output [32:0] alu_operand_b_o;
wire [32:0] alu_operand_b_o;
/* cellift = 32'd1 */
output [32:0] alu_operand_b_o_t0;
wire [32:0] alu_operand_b_o_t0;
/* src = "generated/sv2v_out.v:19542.13-19542.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:19555.13-19555.30" */
input data_ind_timing_i;
wire data_ind_timing_i;
/* cellift = 32'd1 */
input data_ind_timing_i_t0;
wire data_ind_timing_i_t0;
/* src = "generated/sv2v_out.v:19594.6-19594.19" */
reg div_by_zero_q;
/* src = "generated/sv2v_out.v:19591.7-19591.22" */
wire div_change_sign;
/* src = "generated/sv2v_out.v:19545.13-19545.21" */
input div_en_i;
wire div_en_i;
/* cellift = 32'd1 */
input div_en_i_t0;
wire div_en_i_t0;
/* src = "generated/sv2v_out.v:19547.13-19547.22" */
input div_sel_i;
wire div_sel_i;
/* cellift = 32'd1 */
input div_sel_i_t0;
wire div_sel_i_t0;
/* src = "generated/sv2v_out.v:19554.13-19554.28" */
input equal_to_zero_i;
wire equal_to_zero_i;
/* cellift = 32'd1 */
input equal_to_zero_i_t0;
wire equal_to_zero_i_t0;
/* src = "generated/sv2v_out.v:19559.21-19559.32" */
output [67:0] imd_val_d_o;
wire [67:0] imd_val_d_o;
/* cellift = 32'd1 */
output [67:0] imd_val_d_o_t0;
wire [67:0] imd_val_d_o_t0;
/* src = "generated/sv2v_out.v:19558.20-19558.31" */
input [67:0] imd_val_q_i;
wire [67:0] imd_val_q_i;
/* cellift = 32'd1 */
input [67:0] imd_val_q_i_t0;
wire [67:0] imd_val_q_i_t0;
/* src = "generated/sv2v_out.v:19560.20-19560.32" */
output [1:0] imd_val_we_o;
wire [1:0] imd_val_we_o;
/* cellift = 32'd1 */
output [1:0] imd_val_we_o_t0;
wire [1:0] imd_val_we_o_t0;
/* src = "generated/sv2v_out.v:19590.7-19590.23" */
wire is_greater_equal;
/* src = "generated/sv2v_out.v:19564.12-19564.22" */
reg [2:0] md_state_q;
/* src = "generated/sv2v_out.v:19544.13-19544.22" */
input mult_en_i;
wire mult_en_i;
/* cellift = 32'd1 */
input mult_en_i_t0;
wire mult_en_i_t0;
/* src = "generated/sv2v_out.v:19546.13-19546.23" */
input mult_sel_i;
wire mult_sel_i;
/* cellift = 32'd1 */
input mult_sel_i_t0;
wire mult_sel_i_t0;
/* src = "generated/sv2v_out.v:19572.12-19572.27" */
reg [4:0] multdiv_count_q;
/* src = "generated/sv2v_out.v:19596.7-19596.17" */
wire multdiv_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19596.7-19596.17" */
wire multdiv_en_t0;
/* src = "generated/sv2v_out.v:19595.6-19595.18" */
wire multdiv_hold;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19595.6-19595.18" */
wire multdiv_hold_t0;
/* src = "generated/sv2v_out.v:19561.13-19561.31" */
input multdiv_ready_id_i;
wire multdiv_ready_id_i;
/* cellift = 32'd1 */
input multdiv_ready_id_i_t0;
wire multdiv_ready_id_i_t0;
/* src = "generated/sv2v_out.v:19562.21-19562.37" */
output [31:0] multdiv_result_o;
wire [31:0] multdiv_result_o;
/* cellift = 32'd1 */
output [31:0] multdiv_result_o_t0;
wire [31:0] multdiv_result_o_t0;
/* src = "generated/sv2v_out.v:19586.14-19586.27" */
wire [32:0] next_quotient;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19586.14-19586.27" */
wire [32:0] next_quotient_t0;
/* src = "generated/sv2v_out.v:19587.14-19587.28" */
wire [31:0] next_remainder;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19587.14-19587.28" */
wire [31:0] next_remainder_t0;
/* src = "generated/sv2v_out.v:19580.14-19580.23" */
wire [32:0] one_shift;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19580.14-19580.23" */
wire [32:0] one_shift_t0;
/* src = "generated/sv2v_out.v:19582.14-19582.29" */
wire [32:0] op_a_bw_last_pp;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19582.14-19582.29" */
wire [32:0] op_a_bw_last_pp_t0;
/* src = "generated/sv2v_out.v:19581.14-19581.24" */
wire [32:0] op_a_bw_pp;
/* src = "generated/sv2v_out.v:19550.20-19550.26" */
input [31:0] op_a_i;
wire [31:0] op_a_i;
/* cellift = 32'd1 */
input [31:0] op_a_i_t0;
wire [31:0] op_a_i_t0;
/* src = "generated/sv2v_out.v:19576.13-19576.25" */
reg [32:0] op_a_shift_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19576.13-19576.25" */
reg [32:0] op_a_shift_q_t0;
/* src = "generated/sv2v_out.v:19551.20-19551.26" */
input [31:0] op_b_i;
wire [31:0] op_b_i;
/* cellift = 32'd1 */
input [31:0] op_b_i_t0;
wire [31:0] op_b_i_t0;
/* src = "generated/sv2v_out.v:19574.13-19574.25" */
reg [32:0] op_b_shift_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19574.13-19574.25" */
reg [32:0] op_b_shift_q_t0;
/* src = "generated/sv2v_out.v:19589.13-19589.27" */
wire [31:0] op_numerator_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.13-19589.27" */
wire [31:0] op_numerator_d_t0;
/* src = "generated/sv2v_out.v:19548.19-19548.29" */
input [1:0] operator_i;
wire [1:0] operator_i;
/* cellift = 32'd1 */
input [1:0] operator_i_t0;
wire [1:0] operator_i_t0;
/* src = "generated/sv2v_out.v:19592.7-19592.22" */
wire rem_change_sign;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19592.7-19592.22" */
wire rem_change_sign_t0;
/* src = "generated/sv2v_out.v:19543.13-19543.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:19585.7-19585.13" */
wire sign_b;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19585.7-19585.13" */
wire sign_b_t0;
/* src = "generated/sv2v_out.v:19549.19-19549.32" */
input [1:0] signed_mode_i;
wire [1:0] signed_mode_i;
/* cellift = 32'd1 */
input [1:0] signed_mode_i_t0;
wire [1:0] signed_mode_i_t0;
/* src = "generated/sv2v_out.v:19563.14-19563.21" */
output valid_o;
wire valid_o;
/* cellift = 32'd1 */
output valid_o_t0;
wire valid_o_t0;
assign op_a_bw_pp[31:0] = op_a_shift_q[31:0] & /* src = "generated/sv2v_out.v:19643.66-19643.90" */ { op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0] };
assign op_a_bw_last_pp[32] = op_a_shift_q[32] & /* src = "generated/sv2v_out.v:19643.28-19643.62" */ op_b_shift_q[0];
assign rem_change_sign = op_a_i[31] & /* src = "generated/sv2v_out.v:19644.18-19644.47" */ signed_mode_i[0];
assign sign_b = op_b_i[31] & /* src = "generated/sv2v_out.v:19645.18-19645.47" */ signed_mode_i[1];
assign div_change_sign = _304_ & /* src = "generated/sv2v_out.v:19652.27-19652.61" */ _272_;
assign _038_ = op_a_i & /* src = "generated/sv2v_out.v:19669.55-19669.88" */ { op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0] };
assign _042_ = op_a_i[31:1] & /* src = "generated/sv2v_out.v:19675.61-19675.94" */ { op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0] };
assign _040_ = rem_change_sign & /* src = "generated/sv2v_out.v:19675.34-19675.58" */ op_b_i[0];
assign multdiv_en = _277_ & /* src = "generated/sv2v_out.v:19767.22-19767.60" */ imd_val_we_o[0];
assign _044_ = _253_ & /* src = "generated/sv2v_out.v:19783.43-19783.111" */ _279_;
assign _045_ = ~ _089_;
assign _046_ = ~ _090_;
assign _120_ = { _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_, _089_ } & _013_;
assign _122_ = { _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_, _090_ } & _011_;
assign _121_ = { _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_, _045_ } & op_b_shift_q_t0;
assign _123_ = { _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_, _046_ } & op_a_shift_q_t0;
assign _213_ = _120_ | _121_;
assign _214_ = _122_ | _123_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME op_b_shift_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) op_b_shift_q_t0 <= 33'h000000000;
else op_b_shift_q_t0 <= _213_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME op_a_shift_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) op_a_shift_q_t0 <= 33'h000000000;
else op_a_shift_q_t0 <= _214_;
assign _096_ = op_a_shift_q_t0[31:0] & { op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0] };
assign _099_ = op_a_shift_q_t0[32] & op_b_shift_q[0];
assign _102_ = op_a_i_t0[31] & signed_mode_i[0];
assign _105_ = op_b_i_t0[31] & signed_mode_i[1];
assign _108_ = op_a_i_t0 & { op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0] };
assign _111_ = op_a_i_t0[31:1] & { op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0] };
assign _114_ = rem_change_sign_t0 & op_b_i[0];
assign _117_ = _278_ & imd_val_we_o[0];
assign _097_ = { op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0] } & op_a_shift_q[31:0];
assign _100_ = op_b_shift_q_t0[0] & op_a_shift_q[32];
assign _103_ = signed_mode_i_t0[0] & op_a_i[31];
assign _106_ = signed_mode_i_t0[1] & op_b_i[31];
assign _109_ = { op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0] } & op_a_i;
assign _112_ = { op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0] } & op_a_i[31:1];
assign _115_ = op_b_i_t0[0] & rem_change_sign;
assign _118_ = multdiv_hold_t0 & _277_;
assign _098_ = op_a_shift_q_t0[31:0] & { op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0] };
assign _101_ = op_a_shift_q_t0[32] & op_b_shift_q_t0[0];
assign _104_ = op_a_i_t0[31] & signed_mode_i_t0[0];
assign _107_ = op_b_i_t0[31] & signed_mode_i_t0[1];
assign _110_ = op_a_i_t0 & { op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0] };
assign _113_ = op_a_i_t0[31:1] & { op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0] };
assign _116_ = rem_change_sign_t0 & op_b_i_t0[0];
assign _119_ = _278_ & multdiv_hold_t0;
assign _205_ = _096_ | _097_;
assign _206_ = _099_ | _100_;
assign _207_ = _102_ | _103_;
assign _208_ = _105_ | _106_;
assign _209_ = _108_ | _109_;
assign _210_ = _111_ | _112_;
assign _211_ = _114_ | _115_;
assign _212_ = _117_ | _118_;
assign op_a_bw_last_pp_t0[31:0] = _205_ | _098_;
assign op_a_bw_last_pp_t0[32] = _206_ | _101_;
assign rem_change_sign_t0 = _207_ | _104_;
assign sign_b_t0 = _208_ | _107_;
assign _039_ = _209_ | _110_;
assign _043_ = _210_ | _113_;
assign _041_ = _211_ | _116_;
assign multdiv_en_t0 = _212_ | _119_;
/* src = "generated/sv2v_out.v:19768.2-19782.6" */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME md_state_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) md_state_q <= 3'h0;
else if (_087_) md_state_q <= _006_;
/* src = "generated/sv2v_out.v:19768.2-19782.6" */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME multdiv_count_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) multdiv_count_q <= 5'h00;
else if (_088_) multdiv_count_q <= _007_;
/* src = "generated/sv2v_out.v:19768.2-19782.6" */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME op_b_shift_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) op_b_shift_q <= 33'h000000000;
else if (_089_) op_b_shift_q <= _012_;
/* src = "generated/sv2v_out.v:19768.2-19782.6" */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME op_a_shift_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) op_a_shift_q <= 33'h000000000;
else if (_090_) op_a_shift_q <= _010_;
/* src = "generated/sv2v_out.v:19768.2-19782.6" */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME div_by_zero_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) div_by_zero_q <= 1'h0;
else if (_091_) div_by_zero_q <= _018_;
assign _047_ = ~ { _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_ };
assign _048_ = ~ { _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_ };
assign _049_ = ~ _077_;
assign _050_ = ~ { _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_ };
assign _051_ = ~ { _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_ };
assign _052_ = ~ { _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_ };
assign _053_ = ~ { _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_ };
assign _054_ = ~ { _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_ };
assign _055_ = ~ { _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_ };
assign _056_ = ~ { _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_ };
assign _057_ = ~ { _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_ };
assign _058_ = ~ { _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_ };
assign _059_ = ~ { _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_ };
assign _060_ = ~ _258_;
assign _061_ = ~ { _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_ };
assign _062_ = ~ { _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_ };
assign _063_ = ~ { _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_ };
assign _064_ = ~ { _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_ };
assign _065_ = ~ { _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_, _078_ };
assign _066_ = ~ { is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal };
assign _067_ = ~ { is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal };
assign _068_ = ~ { rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign };
assign _069_ = ~ { sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b };
assign _070_ = ~ { div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign };
assign _071_ = ~ { rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign };
assign _072_ = ~ { div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i };
assign _124_ = _047_ & imd_val_q_i_t0[66:34];
assign _126_ = _048_ & _218_;
assign _021_ = _049_ & multdiv_ready_id_i_t0;
assign _128_ = _047_ & alu_adder_ext_i_t0[32:0];
assign _130_ = _048_ & _220_;
assign _132_ = _050_ & { op_a_shift_q_t0[31:0], 1'h0 };
assign _134_ = _051_ & alu_adder_ext_i_t0[32:0];
assign _136_ = _050_ & _222_;
assign _138_ = _051_ & { _041_, _039_ };
assign _140_ = _052_ & _227_;
assign _142_ = _051_ & { op_a_i_t0, 1'h0 };
assign _229_ = _053_ & _023_;
assign _144_ = _054_ & _229_;
assign _146_ = _055_ & _025_;
assign _148_ = _054_ & _231_;
assign _150_ = _056_ & _027_;
assign _152_ = _057_ & _233_;
assign _154_ = _058_ & imd_val_q_i_t0[66:34];
assign _156_ = _055_ & _237_;
assign _158_ = _059_ & _239_;
assign _160_ = _060_ & _246_;
assign _162_ = _057_ & { op_b_i_t0, 1'h0 };
assign _164_ = _053_ & { op_b_shift_q_t0[31:0], 1'h0 };
assign _166_ = _061_ & _250_;
assign _168_ = _051_ & op_a_bw_last_pp_t0;
assign _170_ = _050_ & _252_;
assign _172_ = _050_ & imd_val_q_i_t0[66:34];
assign _180_ = _062_ & imd_val_q_i_t0[31:0];
assign _182_ = _063_ & imd_val_q_i_t0[31:0];
assign _184_ = _064_ & imd_val_q_i_t0[66:34];
assign _003_ = _065_ & { imd_val_q_i_t0[65:34], 1'h0 };
assign _186_ = _056_ & op_a_bw_last_pp_t0;
assign _188_ = _066_ & imd_val_q_i_t0[65:34];
assign _190_ = _067_ & op_a_shift_q_t0;
assign _192_ = _068_ & op_a_i_t0;
assign _194_ = _069_ & { 1'h0, op_b_i_t0 };
assign _196_ = _070_ & imd_val_q_i_t0[66:34];
assign _198_ = _071_ & imd_val_q_i_t0[66:34];
assign _200_ = _072_ & alu_adder_ext_i_t0[31:0];
assign _125_ = { _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_ } & _301_;
assign _127_ = { _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_ } & _303_;
assign _129_ = { _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_, _281_ } & next_quotient_t0;
assign _131_ = { _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_ } & { 1'h0, next_remainder_t0 };
assign _133_ = { _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_ } & next_quotient_t0;
assign _135_ = { _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_ } & alu_adder_ext_i_t0[33:1];
assign _137_ = { _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_ } & { next_remainder_t0, _288_ };
assign _225_ = { _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_, _280_ } & { rem_change_sign_t0, op_a_i_t0 };
assign _139_ = { _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_ } & { 1'h0, _041_, _043_ };
assign _141_ = { _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_, _202_ } & _225_;
assign _143_ = { _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_ } & { rem_change_sign_t0, op_a_i_t0 };
assign _145_ = { _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_ } & _030_;
assign _147_ = { _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_ } & _297_;
assign _149_ = { _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_, _283_ } & _032_;
assign _151_ = { _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_ } & _034_;
assign _153_ = { _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_ } & _037_;
assign _155_ = { _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_, _284_ } & _017_;
assign _157_ = { _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_, _286_ } & { 32'h00000000, imd_val_q_i_t0[31] };
assign _159_ = { _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_, _079_ } & _235_;
assign _246_ = _253_ & _021_;
assign _161_ = _258_ & multdiv_ready_id_i_t0;
assign _163_ = { _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_, _282_ } & { imd_val_q_i_t0[65:34], 1'h0 };
assign _165_ = { _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_ } & { op_a_i_t0, 1'h0 };
assign _167_ = { _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_, _204_ } & _248_;
assign _169_ = { _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_, _260_ } & _291_;
assign _171_ = { _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_ } & _005_;
assign _173_ = { _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_, _077_ } & _003_;
assign _032_ = { _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_ } & { 1'h0, op_b_shift_q_t0[32:1] };
assign _025_ = { _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_, _093_ } & { 1'h0, sign_b_t0, op_b_i_t0[31:1] };
assign _181_ = { _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_, _285_ } & _295_;
assign multdiv_hold_t0 = _265_ & _009_;
assign _183_ = { _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_ } & _015_;
assign _185_ = { _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_, _265_ } & _001_;
assign _187_ = { _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_, _253_ } & op_a_bw_last_pp_t0;
assign _189_ = { is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal } & alu_adder_ext_i_t0[32:1];
assign _191_ = { is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal } & _276_;
assign _193_ = { rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign } & alu_adder_i_t0;
assign _195_ = { sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b } & { 1'h0, alu_adder_i_t0 };
assign _197_ = { div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign } & { 1'h0, alu_adder_i_t0 };
assign _199_ = { rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign } & { 1'h0, alu_adder_i_t0 };
assign _201_ = { div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i } & imd_val_q_i_t0[65:34];
assign _218_ = _124_ | _125_;
assign _037_ = _126_ | _127_;
assign _220_ = _128_ | _129_;
assign _034_ = _130_ | _131_;
assign _030_ = _132_ | _133_;
assign _222_ = _134_ | _135_;
assign _027_ = _136_ | _137_;
assign _227_ = _138_ | _139_;
assign _017_ = _140_ | _141_;
assign _023_ = _142_ | _143_;
assign _011_ = _144_ | _145_;
assign _231_ = _146_ | _147_;
assign _013_ = _148_ | _149_;
assign _233_ = _150_ | _151_;
assign _235_ = _152_ | _153_;
assign _237_ = _154_ | _155_;
assign _239_ = _156_ | _157_;
assign _001_ = _158_ | _159_;
assign _009_ = _160_ | _161_;
assign _248_ = _162_ | _163_;
assign _250_ = _164_ | _165_;
assign _005_ = _166_ | _167_;
assign _252_ = _168_ | _169_;
assign alu_operand_b_o_t0 = _170_ | _171_;
assign alu_operand_a_o_t0 = _172_ | _173_;
assign _015_ = _180_ | _181_;
assign op_numerator_d_t0 = _182_ | _183_;
assign accum_window_d_t0 = _184_ | _185_;
assign _291_ = _186_ | _187_;
assign next_remainder_t0 = _188_ | _189_;
assign next_quotient_t0 = _190_ | _191_;
assign _295_ = _192_ | _193_;
assign _297_ = _194_ | _195_;
assign _301_ = _196_ | _197_;
assign _303_ = _198_ | _199_;
assign multdiv_result_o_t0 = _200_ | _201_;
assign _080_ = | { _284_, _283_ };
assign _081_ = { _283_, _077_ } != 2'h3;
assign _082_ = { _284_, _077_ } != 2'h3;
assign _083_ = | { _286_, _284_, _283_ };
assign _084_ = { _283_, _260_ } != 2'h3;
assign _085_ = | { _285_, _284_, _283_ };
assign _086_ = ~ _092_;
assign _087_ = & { _265_, multdiv_en };
assign _088_ = & { _080_, _265_, multdiv_en };
assign _089_ = & { _265_, multdiv_en, _081_, _082_, _083_ };
assign _090_ = & { _265_, multdiv_en, _084_, _085_, _082_ };
assign _091_ = & { _284_, _265_, multdiv_en, _086_ };
assign _092_ = | { _280_, _260_, _259_ };
assign _094_ = | { _286_, _284_ };
assign _093_ = | { _260_, _259_ };
assign _095_ = | { _281_, _280_, _260_ };
assign _073_ = ~ op_a_shift_q;
assign _074_ = ~ mult_en_i;
assign _075_ = ~ one_shift;
assign _076_ = ~ div_en_i;
assign _174_ = op_a_shift_q_t0 & _075_;
assign _177_ = mult_en_i_t0 & _076_;
assign _175_ = one_shift_t0 & _073_;
assign _178_ = div_en_i_t0 & _074_;
assign _176_ = op_a_shift_q_t0 & one_shift_t0;
assign _179_ = mult_en_i_t0 & div_en_i_t0;
assign _215_ = _174_ | _175_;
assign _216_ = _177_ | _178_;
assign _276_ = _215_ | _176_;
assign _278_ = _216_ | _179_;
assign _077_ = | { _281_, _280_ };
assign _078_ = | { _286_, _285_, _284_, _282_ };
assign _202_ = _281_ | _280_;
assign _203_ = _285_ | _286_;
assign _204_ = _094_ | _282_;
assign _079_ = | { _283_, _282_, _253_ };
assign _217_ = _281_ ? _300_ : imd_val_q_i[66:34];
assign _036_ = _280_ ? _302_ : _217_;
assign _020_ = _077_ ? 1'h0 : _274_;
assign _035_ = _077_ ? 3'h5 : 3'h0;
assign _219_ = _281_ ? next_quotient : alu_adder_ext_i[32:0];
assign _033_ = _280_ ? { 1'h0, next_remainder } : _219_;
assign _028_ = _095_ ? _299_ : _298_;
assign _029_ = _077_ ? next_quotient : { op_a_shift_q[31:0], 1'h0 };
assign _221_ = _260_ ? alu_adder_ext_i[33:1] : alu_adder_ext_i[32:0];
assign _026_ = _077_ ? { next_remainder, _287_ } : _221_;
assign _223_ = _260_ ? 3'h3 : _292_;
assign _019_ = _077_ ? _293_ : _223_;
assign _224_ = _280_ ? { rem_change_sign, op_a_i } : 33'h1ffffffff;
assign _226_ = _260_ ? { 1'h1, _273_, _042_ } : { _273_, _038_ };
assign _016_ = _202_ ? _224_ : _226_;
assign _022_ = _260_ ? { rem_change_sign, op_a_i } : { op_a_i, 1'h0 };
assign _007_ = _283_ ? _289_ : 5'h1f;
assign _228_ = _285_ ? 33'h000000000 : _022_;
assign _010_ = _283_ ? _029_ : _228_;
assign _230_ = _286_ ? _296_ : _024_;
assign _012_ = _283_ ? _031_ : _230_;
assign _232_ = _253_ ? _033_ : _026_;
assign _234_ = _282_ ? _036_ : _232_;
assign _236_ = _284_ ? _016_ : imd_val_q_i[66:34];
assign _238_ = _286_ ? { 32'h00000000, imd_val_q_i[31] } : _236_;
assign _000_ = _079_ ? _234_ : _238_;
assign _240_ = _253_ ? _035_ : _028_;
assign _241_ = _282_ ? 3'h6 : _240_;
assign _242_ = _286_ ? 3'h3 : 3'h2;
assign _243_ = _284_ ? _019_ : 3'h0;
assign _244_ = _203_ ? _242_ : _243_;
assign _006_ = _079_ ? _241_ : _244_;
assign _245_ = _253_ ? _020_ : 1'h0;
assign _008_ = _258_ ? _274_ : _245_;
assign _247_ = _282_ ? { _269_, 1'h1 } : { _267_, 1'h1 };
assign _249_ = _285_ ? { _268_, 1'h1 } : { _270_, 1'h1 };
assign _004_ = _204_ ? _247_ : _249_;
assign _251_ = _260_ ? _290_ : op_a_bw_pp;
assign alu_operand_b_o = _077_ ? _004_ : _251_;
assign alu_operand_a_o = _077_ ? _002_ : imd_val_q_i[66:34];
assign _288_ = imd_val_q_i_t0[31:0] >> _289_;
assign one_shift_t0 = 33'h000000000 << multdiv_count_q;
assign _254_ = imd_val_q_i[65] == /* src = "generated/sv2v_out.v:19648.29-19648.67" */ op_b_shift_q[31];
assign _255_ = ! /* src = "generated/sv2v_out.v:19671.45-19671.65" */ { 1'h0, sign_b, op_b_i[31:1] };
assign _256_ = ! /* src = "generated/sv2v_out.v:19710.46-19710.63" */ { 1'h0, op_b_shift_q[32:1] };
assign _257_ = multdiv_count_q == /* src = "generated/sv2v_out.v:19721.22-19721.45" */ 5'h01;
assign _261_ = _264_ && /* src = "generated/sv2v_out.v:19671.22-19671.66" */ _255_;
assign _262_ = _264_ && /* src = "generated/sv2v_out.v:19686.22-19686.59" */ equal_to_zero_i;
assign _263_ = _264_ && /* src = "generated/sv2v_out.v:19710.23-19710.64" */ _256_;
assign _264_ = ! /* src = "generated/sv2v_out.v:19710.23-19710.41" */ data_ind_timing_i;
assign _265_ = mult_sel_i || /* src = "generated/sv2v_out.v:19663.7-19663.30" */ div_sel_i;
assign _266_ = _263_ || /* src = "generated/sv2v_out.v:19710.22-19710.94" */ _257_;
assign _268_ = ~ /* src = "generated/sv2v_out.v:19620.26-19620.33" */ op_a_i;
assign _267_ = ~ /* src = "generated/sv2v_out.v:19624.26-19624.33" */ op_b_i;
assign _269_ = ~ /* src = "generated/sv2v_out.v:19628.26-19628.47" */ imd_val_q_i[65:34];
assign _270_ = ~ /* src = "generated/sv2v_out.v:19637.24-19637.43" */ op_b_shift_q[31:0];
assign op_a_bw_pp[32] = ~ /* src = "generated/sv2v_out.v:19642.23-19642.60" */ op_a_bw_last_pp[32];
assign op_a_bw_last_pp[31:0] = ~ /* src = "generated/sv2v_out.v:19643.64-19643.91" */ op_a_bw_pp[31:0];
assign _271_ = ~ /* src = "generated/sv2v_out.v:19648.70-19648.86" */ alu_adder_ext_i[32];
assign _272_ = ~ /* src = "generated/sv2v_out.v:19652.47-19652.61" */ div_by_zero_q;
assign _273_ = ~ /* src = "generated/sv2v_out.v:19675.32-19675.59" */ _040_;
assign _274_ = ~ /* src = "generated/sv2v_out.v:19762.21-19762.40" */ multdiv_ready_id_i;
assign imd_val_we_o[0] = ~ /* src = "generated/sv2v_out.v:19767.47-19767.60" */ multdiv_hold;
assign _275_ = op_a_shift_q | /* src = "generated/sv2v_out.v:19651.45-19651.69" */ one_shift;
assign _277_ = mult_en_i | /* src = "generated/sv2v_out.v:19767.23-19767.43" */ div_en_i;
assign _279_ = _259_ | /* src = "generated/sv2v_out.v:19783.67-19783.110" */ _260_;
assign valid_o = _258_ | /* src = "generated/sv2v_out.v:19783.19-19783.112" */ _044_;
assign _031_ = _093_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19705.6-19725.13" */ { 1'h0, op_b_shift_q[32:1] } : 33'hxxxxxxxxx;
assign _024_ = _093_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19666.6-19690.13" */ { 1'h0, sign_b, op_b_i[31:1] } : 33'hxxxxxxxxx;
assign _018_ = _281_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19666.6-19690.13" */ equal_to_zero_i : 1'hx;
assign _283_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19664.4-19765.11" */ 3'h3;
assign _258_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19664.4-19765.11" */ 3'h6;
assign _253_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19664.4-19765.11" */ 3'h4;
assign _014_ = _285_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19664.4-19765.11" */ _294_ : imd_val_q_i[31:0];
assign multdiv_hold = _265_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:19663.7-19663.30|generated/sv2v_out.v:19663.3-19765.11" */ _008_ : 1'h0;
assign op_numerator_d = _265_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:19663.7-19663.30|generated/sv2v_out.v:19663.3-19765.11" */ _014_ : imd_val_q_i[31:0];
assign accum_window_d = _265_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:19663.7-19663.30|generated/sv2v_out.v:19663.3-19765.11" */ _000_ : imd_val_q_i[66:34];
assign _002_ = _078_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19613.5-19634.12" */ 33'h000000001 : { imd_val_q_i[65:34], 1'h1 };
assign _282_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19613.5-19634.12" */ 3'h5;
assign _286_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19613.5-19634.12" */ 3'h2;
assign _285_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19613.5-19634.12" */ 3'h1;
assign _284_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19613.5-19634.12" */ md_state_q;
assign _260_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19609.3-19639.10" */ 2'h1;
assign _259_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19609.3-19639.10" */ operator_i;
assign _281_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19609.3-19639.10" */ 2'h2;
assign _280_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19609.3-19639.10" */ 2'h3;
wire [31:0] _651_ = imd_val_q_i[31:0];
assign _287_ = _651_[_289_ +: 1];
assign one_shift = 33'h000000001 << /* src = "generated/sv2v_out.v:19649.21-19649.77" */ multdiv_count_q;
assign _289_ = multdiv_count_q - /* src = "generated/sv2v_out.v:19704.24-19704.47" */ 5'h01;
assign _290_ = _253_ ? /* src = "generated/sv2v_out.v:19611.29-19611.78" */ op_a_bw_last_pp : op_a_bw_pp;
assign is_greater_equal = _254_ ? /* src = "generated/sv2v_out.v:19648.29-19648.107" */ _271_ : imd_val_q_i[65];
assign next_remainder = is_greater_equal ? /* src = "generated/sv2v_out.v:19650.27-19650.86" */ alu_adder_ext_i[32:1] : imd_val_q_i[65:34];
assign next_quotient = is_greater_equal ? /* src = "generated/sv2v_out.v:19651.26-19651.84" */ _275_ : op_a_shift_q;
assign _292_ = _261_ ? /* src = "generated/sv2v_out.v:19671.22-19671.80" */ 3'h4 : 3'h3;
assign _293_ = _262_ ? /* src = "generated/sv2v_out.v:19686.22-19686.73" */ 3'h6 : 3'h1;
assign _294_ = rem_change_sign ? /* src = "generated/sv2v_out.v:19695.24-19695.53" */ alu_adder_i : op_a_i;
assign _296_ = sign_b ? /* src = "generated/sv2v_out.v:19700.22-19700.67" */ { 1'h0, alu_adder_i } : { 1'h0, op_b_i };
assign _298_ = _266_ ? /* src = "generated/sv2v_out.v:19710.22-19710.108" */ 3'h4 : 3'h3;
assign _299_ = _257_ ? /* src = "generated/sv2v_out.v:19721.22-19721.59" */ 3'h4 : 3'h3;
assign _300_ = div_change_sign ? /* src = "generated/sv2v_out.v:19754.31-19754.85" */ { 1'h0, alu_adder_i } : imd_val_q_i[66:34];
assign _302_ = rem_change_sign ? /* src = "generated/sv2v_out.v:19755.31-19755.85" */ { 1'h0, alu_adder_i } : imd_val_q_i[66:34];
assign multdiv_result_o = div_en_i ? /* src = "generated/sv2v_out.v:19784.29-19784.80" */ imd_val_q_i[65:34] : alu_adder_ext_i[31:0];
assign _304_ = rem_change_sign ^ /* src = "generated/sv2v_out.v:19652.28-19652.43" */ sign_b;
assign imd_val_d_o = { 1'h0, accum_window_d, 2'h0, op_numerator_d };
assign imd_val_d_o_t0 = { 1'h0, accum_window_d_t0, 2'h0, op_numerator_d_t0 };
assign imd_val_we_o[1] = multdiv_en;
assign imd_val_we_o_t0 = { multdiv_en_t0, multdiv_hold_t0 };
assign valid_o_t0 = 1'h0;
endmodule

module ibex_top(clk_i, rst_ni, test_en_i, ram_cfg_i, hart_id_i, boot_addr_i, instr_req_o, instr_gnt_i, instr_rvalid_i, instr_addr_o, instr_rdata_i, instr_rdata_intg_i, instr_err_i, data_req_o, data_gnt_i, data_rvalid_i, data_we_o, data_be_o, data_addr_o, data_wdata_o, data_wdata_intg_o
, data_rdata_i, data_rdata_intg_i, data_err_i, irq_software_i, irq_timer_i, irq_external_i, irq_fast_i, irq_nm_i, scramble_key_valid_i, scramble_key_i, scramble_nonce_i, scramble_req_o, debug_req_i, crash_dump_o, double_fault_seen_o, fetch_enable_i, alert_minor_o, alert_major_internal_o, alert_major_bus_o, core_sleep_o, scan_rst_ni
, debug_req_i_t0, boot_addr_i_t0, irq_nm_i_t0, data_we_o_t0, data_req_o_t0, instr_rvalid_i_t0, instr_req_o_t0, instr_rdata_i_t0, instr_gnt_i_t0, instr_err_i_t0, instr_addr_o_t0, test_en_i_t0, data_addr_o_t0, data_be_o_t0, data_gnt_i_t0, data_rdata_i_t0, data_rvalid_i_t0, data_wdata_o_t0, double_fault_seen_o_t0, hart_id_i_t0, irq_external_i_t0
, irq_fast_i_t0, irq_software_i_t0, irq_timer_i_t0, alert_major_bus_o_t0, alert_major_internal_o_t0, alert_minor_o_t0, crash_dump_o_t0, data_err_i_t0, fetch_enable_i_t0, core_sleep_o_t0, data_rdata_intg_i_t0, data_wdata_intg_o_t0, instr_rdata_intg_i_t0, ram_cfg_i_t0, scan_rst_ni_t0, scramble_key_i_t0, scramble_key_valid_i_t0, scramble_nonce_i_t0, scramble_req_o_t0);
wire _00_;
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
/* src = "generated/sv2v_out.v:20400.25-20400.60" */
wire _19_;
/* src = "generated/sv2v_out.v:20400.24-20400.75" */
wire _20_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20400.24-20400.75" */
wire _21_;
/* src = "generated/sv2v_out.v:20400.23-20400.90" */
wire _22_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20400.23-20400.90" */
wire _23_;
/* src = "generated/sv2v_out.v:20315.14-20315.31" */
output alert_major_bus_o;
wire alert_major_bus_o;
/* cellift = 32'd1 */
output alert_major_bus_o_t0;
wire alert_major_bus_o_t0;
/* src = "generated/sv2v_out.v:20314.14-20314.36" */
output alert_major_internal_o;
wire alert_major_internal_o;
/* cellift = 32'd1 */
output alert_major_internal_o_t0;
wire alert_major_internal_o_t0;
/* src = "generated/sv2v_out.v:20313.14-20313.27" */
output alert_minor_o;
wire alert_minor_o;
/* cellift = 32'd1 */
output alert_minor_o_t0;
wire alert_minor_o_t0;
/* src = "generated/sv2v_out.v:20281.20-20281.31" */
input [31:0] boot_addr_i;
wire [31:0] boot_addr_i;
/* cellift = 32'd1 */
input [31:0] boot_addr_i_t0;
wire [31:0] boot_addr_i_t0;
/* src = "generated/sv2v_out.v:20343.7-20343.10" */
wire clk;
/* src = "generated/sv2v_out.v:20276.13-20276.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:20346.7-20346.15" */
wire clock_en;
/* src = "generated/sv2v_out.v:20373.7-20373.32" */
wire core_alert_major_internal;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20373.7-20373.32" */
wire core_alert_major_internal_t0;
/* src = "generated/sv2v_out.v:20344.13-20344.24" */
wire [3:0] core_busy_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20344.13-20344.24" */
wire [3:0] core_busy_d_t0;
/* src = "generated/sv2v_out.v:20345.12-20345.23" */
wire [3:0] core_busy_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20345.12-20345.23" */
/* unused_bits = "0 1 2 3" */
wire [3:0] core_busy_q_t0;
/* src = "generated/sv2v_out.v:20316.14-20316.26" */
output core_sleep_o;
wire core_sleep_o;
/* cellift = 32'd1 */
output core_sleep_o_t0;
wire core_sleep_o_t0;
/* src = "generated/sv2v_out.v:20310.22-20310.34" */
output [159:0] crash_dump_o;
wire [159:0] crash_dump_o;
/* cellift = 32'd1 */
output [159:0] crash_dump_o_t0;
wire [159:0] crash_dump_o_t0;
/* src = "generated/sv2v_out.v:20294.21-20294.32" */
output [31:0] data_addr_o;
wire [31:0] data_addr_o;
/* cellift = 32'd1 */
output [31:0] data_addr_o_t0;
wire [31:0] data_addr_o_t0;
/* src = "generated/sv2v_out.v:20293.20-20293.29" */
output [3:0] data_be_o;
wire [3:0] data_be_o;
/* cellift = 32'd1 */
output [3:0] data_be_o_t0;
wire [3:0] data_be_o_t0;
/* src = "generated/sv2v_out.v:20299.13-20299.23" */
input data_err_i;
wire data_err_i;
/* cellift = 32'd1 */
input data_err_i_t0;
wire data_err_i_t0;
/* src = "generated/sv2v_out.v:20290.13-20290.23" */
input data_gnt_i;
wire data_gnt_i;
/* cellift = 32'd1 */
input data_gnt_i_t0;
wire data_gnt_i_t0;
/* src = "generated/sv2v_out.v:20297.20-20297.32" */
input [31:0] data_rdata_i;
wire [31:0] data_rdata_i;
/* cellift = 32'd1 */
input [31:0] data_rdata_i_t0;
wire [31:0] data_rdata_i_t0;
/* src = "generated/sv2v_out.v:20298.19-20298.36" */
input [6:0] data_rdata_intg_i;
wire [6:0] data_rdata_intg_i;
/* cellift = 32'd1 */
input [6:0] data_rdata_intg_i_t0;
wire [6:0] data_rdata_intg_i_t0;
/* src = "generated/sv2v_out.v:20289.14-20289.24" */
output data_req_o;
wire data_req_o;
/* cellift = 32'd1 */
output data_req_o_t0;
wire data_req_o_t0;
/* src = "generated/sv2v_out.v:20291.13-20291.26" */
input data_rvalid_i;
wire data_rvalid_i;
/* cellift = 32'd1 */
input data_rvalid_i_t0;
wire data_rvalid_i_t0;
/* src = "generated/sv2v_out.v:20359.28-20359.43" */
wire [38:0] data_wdata_core;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20359.28-20359.43" */
wire [38:0] data_wdata_core_t0;
/* src = "generated/sv2v_out.v:20296.20-20296.37" */
output [6:0] data_wdata_intg_o;
wire [6:0] data_wdata_intg_o;
/* cellift = 32'd1 */
output [6:0] data_wdata_intg_o_t0;
wire [6:0] data_wdata_intg_o_t0;
/* src = "generated/sv2v_out.v:20295.21-20295.33" */
output [31:0] data_wdata_o;
wire [31:0] data_wdata_o;
/* cellift = 32'd1 */
output [31:0] data_wdata_o_t0;
wire [31:0] data_wdata_o_t0;
/* src = "generated/sv2v_out.v:20292.14-20292.23" */
output data_we_o;
wire data_we_o;
/* cellift = 32'd1 */
output data_we_o_t0;
wire data_we_o_t0;
/* src = "generated/sv2v_out.v:20309.13-20309.24" */
input debug_req_i;
wire debug_req_i;
/* cellift = 32'd1 */
input debug_req_i_t0;
wire debug_req_i_t0;
/* src = "generated/sv2v_out.v:20311.14-20311.33" */
output double_fault_seen_o;
wire double_fault_seen_o;
/* cellift = 32'd1 */
output double_fault_seen_o_t0;
wire double_fault_seen_o_t0;
/* src = "generated/sv2v_out.v:20348.7-20348.21" */
wire dummy_instr_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20348.7-20348.21" */
wire dummy_instr_id_t0;
/* src = "generated/sv2v_out.v:20349.7-20349.21" */
wire dummy_instr_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20349.7-20349.21" */
wire dummy_instr_wb_t0;
/* src = "generated/sv2v_out.v:20385.13-20385.29" */
wire [3:0] fetch_enable_buf;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20385.13-20385.29" */
wire [3:0] fetch_enable_buf_t0;
/* src = "generated/sv2v_out.v:20312.19-20312.33" */
input [3:0] fetch_enable_i;
wire [3:0] fetch_enable_i;
/* cellift = 32'd1 */
input [3:0] fetch_enable_i_t0;
wire [3:0] fetch_enable_i_t0;
/* src = "generated/sv2v_out.v:20280.20-20280.29" */
input [31:0] hart_id_i;
wire [31:0] hart_id_i;
/* cellift = 32'd1 */
input [31:0] hart_id_i_t0;
wire [31:0] hart_id_i_t0;
/* src = "generated/sv2v_out.v:20369.35-20369.47" */
/* unused_bits = "0 1 2 3 4 5 6 7" */
wire [7:0] ic_data_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20369.35-20369.47" */
/* unused_bits = "0 1 2 3 4 5 6 7" */
wire [7:0] ic_data_addr_t0;
/* src = "generated/sv2v_out.v:20367.13-20367.24" */
/* unused_bits = "0 1" */
wire [1:0] ic_data_req;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20367.13-20367.24" */
/* unused_bits = "0 1" */
wire [1:0] ic_data_req_t0;
/* src = "generated/sv2v_out.v:20370.27-20370.40" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63" */
wire [63:0] ic_data_wdata;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20370.27-20370.40" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63" */
wire [63:0] ic_data_wdata_t0;
/* src = "generated/sv2v_out.v:20368.7-20368.20" */
/* unused_bits = "0" */
wire ic_data_write;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20368.7-20368.20" */
/* unused_bits = "0" */
wire ic_data_write_t0;
/* src = "generated/sv2v_out.v:20372.7-20372.21" */
/* unused_bits = "0" */
wire ic_scr_key_req;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20372.7-20372.21" */
/* unused_bits = "0" */
wire ic_scr_key_req_t0;
/* src = "generated/sv2v_out.v:20364.35-20364.46" */
/* unused_bits = "0 1 2 3 4 5 6 7" */
wire [7:0] ic_tag_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20364.35-20364.46" */
/* unused_bits = "0 1 2 3 4 5 6 7" */
wire [7:0] ic_tag_addr_t0;
/* src = "generated/sv2v_out.v:20362.13-20362.23" */
/* unused_bits = "0 1" */
wire [1:0] ic_tag_req;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20362.13-20362.23" */
/* unused_bits = "0 1" */
wire [1:0] ic_tag_req_t0;
/* src = "generated/sv2v_out.v:20365.26-20365.38" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21" */
wire [21:0] ic_tag_wdata;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20365.26-20365.38" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21" */
wire [21:0] ic_tag_wdata_t0;
/* src = "generated/sv2v_out.v:20363.7-20363.19" */
/* unused_bits = "0" */
wire ic_tag_write;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20363.7-20363.19" */
/* unused_bits = "0" */
wire ic_tag_write_t0;
/* src = "generated/sv2v_out.v:20285.21-20285.33" */
output [31:0] instr_addr_o;
wire [31:0] instr_addr_o;
/* cellift = 32'd1 */
output [31:0] instr_addr_o_t0;
wire [31:0] instr_addr_o_t0;
/* src = "generated/sv2v_out.v:20288.13-20288.24" */
input instr_err_i;
wire instr_err_i;
/* cellift = 32'd1 */
input instr_err_i_t0;
wire instr_err_i_t0;
/* src = "generated/sv2v_out.v:20283.13-20283.24" */
input instr_gnt_i;
wire instr_gnt_i;
/* cellift = 32'd1 */
input instr_gnt_i_t0;
wire instr_gnt_i_t0;
/* src = "generated/sv2v_out.v:20286.20-20286.33" */
input [31:0] instr_rdata_i;
wire [31:0] instr_rdata_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_i_t0;
wire [31:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:20287.19-20287.37" */
input [6:0] instr_rdata_intg_i;
wire [6:0] instr_rdata_intg_i;
/* cellift = 32'd1 */
input [6:0] instr_rdata_intg_i_t0;
wire [6:0] instr_rdata_intg_i_t0;
/* src = "generated/sv2v_out.v:20282.14-20282.25" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:20284.13-20284.27" */
input instr_rvalid_i;
wire instr_rvalid_i;
/* cellift = 32'd1 */
input instr_rvalid_i_t0;
wire instr_rvalid_i_t0;
/* src = "generated/sv2v_out.v:20302.13-20302.27" */
input irq_external_i;
wire irq_external_i;
/* cellift = 32'd1 */
input irq_external_i_t0;
wire irq_external_i_t0;
/* src = "generated/sv2v_out.v:20303.20-20303.30" */
input [14:0] irq_fast_i;
wire [14:0] irq_fast_i;
/* cellift = 32'd1 */
input [14:0] irq_fast_i_t0;
wire [14:0] irq_fast_i_t0;
/* src = "generated/sv2v_out.v:20304.13-20304.21" */
input irq_nm_i;
wire irq_nm_i;
/* cellift = 32'd1 */
input irq_nm_i_t0;
wire irq_nm_i_t0;
/* src = "generated/sv2v_out.v:20347.7-20347.18" */
wire irq_pending;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20347.7-20347.18" */
wire irq_pending_t0;
/* src = "generated/sv2v_out.v:20300.13-20300.27" */
input irq_software_i;
wire irq_software_i;
/* cellift = 32'd1 */
input irq_software_i_t0;
wire irq_software_i_t0;
/* src = "generated/sv2v_out.v:20301.13-20301.24" */
input irq_timer_i;
wire irq_timer_i;
/* cellift = 32'd1 */
input irq_timer_i_t0;
wire irq_timer_i_t0;
/* src = "generated/sv2v_out.v:20279.19-20279.28" */
input [9:0] ram_cfg_i;
wire [9:0] ram_cfg_i;
/* cellift = 32'd1 */
input [9:0] ram_cfg_i_t0;
wire [9:0] ram_cfg_i_t0;
/* src = "generated/sv2v_out.v:20530.7-20530.30" */
wire rf_alert_major_internal;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20530.7-20530.30" */
wire rf_alert_major_internal_t0;
/* src = "generated/sv2v_out.v:20350.13-20350.23" */
wire [4:0] rf_raddr_a;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20350.13-20350.23" */
wire [4:0] rf_raddr_a_t0;
/* src = "generated/sv2v_out.v:20351.13-20351.23" */
wire [4:0] rf_raddr_b;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20351.13-20351.23" */
wire [4:0] rf_raddr_b_t0;
/* src = "generated/sv2v_out.v:20355.32-20355.46" */
wire [38:0] rf_rdata_a_ecc;
/* src = "generated/sv2v_out.v:20356.32-20356.50" */
wire [38:0] rf_rdata_a_ecc_buf;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20356.32-20356.50" */
wire [38:0] rf_rdata_a_ecc_buf_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20355.32-20355.46" */
wire [38:0] rf_rdata_a_ecc_t0;
/* src = "generated/sv2v_out.v:20357.32-20357.46" */
wire [38:0] rf_rdata_b_ecc;
/* src = "generated/sv2v_out.v:20358.32-20358.50" */
wire [38:0] rf_rdata_b_ecc_buf;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20358.32-20358.50" */
wire [38:0] rf_rdata_b_ecc_buf_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20357.32-20357.46" */
wire [38:0] rf_rdata_b_ecc_t0;
/* src = "generated/sv2v_out.v:20352.13-20352.24" */
wire [4:0] rf_waddr_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20352.13-20352.24" */
wire [4:0] rf_waddr_wb_t0;
/* src = "generated/sv2v_out.v:20354.32-20354.47" */
wire [38:0] rf_wdata_wb_ecc;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20354.32-20354.47" */
wire [38:0] rf_wdata_wb_ecc_t0;
/* src = "generated/sv2v_out.v:20353.7-20353.15" */
wire rf_we_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20353.7-20353.15" */
wire rf_we_wb_t0;
/* src = "generated/sv2v_out.v:20277.13-20277.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:20317.13-20317.24" */
input scan_rst_ni;
wire scan_rst_ni;
/* cellift = 32'd1 */
input scan_rst_ni_t0;
wire scan_rst_ni_t0;
/* src = "generated/sv2v_out.v:20306.21-20306.35" */
input [127:0] scramble_key_i;
wire [127:0] scramble_key_i;
/* cellift = 32'd1 */
input [127:0] scramble_key_i_t0;
wire [127:0] scramble_key_i_t0;
/* src = "generated/sv2v_out.v:20305.13-20305.33" */
input scramble_key_valid_i;
wire scramble_key_valid_i;
/* cellift = 32'd1 */
input scramble_key_valid_i_t0;
wire scramble_key_valid_i_t0;
/* src = "generated/sv2v_out.v:20307.20-20307.36" */
input [63:0] scramble_nonce_i;
wire [63:0] scramble_nonce_i;
/* cellift = 32'd1 */
input [63:0] scramble_nonce_i_t0;
wire [63:0] scramble_nonce_i_t0;
/* src = "generated/sv2v_out.v:20308.14-20308.28" */
output scramble_req_o;
wire scramble_req_o;
/* cellift = 32'd1 */
output scramble_req_o_t0;
wire scramble_req_o_t0;
/* src = "generated/sv2v_out.v:20278.13-20278.22" */
input test_en_i;
wire test_en_i;
/* cellift = 32'd1 */
input test_en_i_t0;
wire test_en_i_t0;
assign _00_ = ~ _19_;
assign _01_ = ~ _20_;
assign _02_ = ~ _22_;
assign _03_ = ~ core_alert_major_internal;
assign _04_ = ~ irq_pending;
assign _05_ = ~ irq_nm_i;
assign _06_ = ~ rf_alert_major_internal;
assign _07_ = _21_ & _04_;
assign _10_ = _23_ & _05_;
assign _13_ = core_alert_major_internal_t0 & _06_;
assign _21_ = debug_req_i_t0 & _00_;
assign _08_ = irq_pending_t0 & _01_;
assign _11_ = irq_nm_i_t0 & _02_;
assign _14_ = rf_alert_major_internal_t0 & _03_;
assign _09_ = _21_ & irq_pending_t0;
assign _12_ = _23_ & irq_nm_i_t0;
assign _15_ = core_alert_major_internal_t0 & rf_alert_major_internal_t0;
assign _16_ = _07_ | _08_;
assign _17_ = _10_ | _11_;
assign _18_ = _13_ | _14_;
assign _23_ = _16_ | _09_;
assign core_sleep_o_t0 = _17_ | _12_;
assign alert_major_internal_o_t0 = _18_ | _15_;
assign _19_ = core_busy_q != /* src = "generated/sv2v_out.v:20400.25-20400.60" */ 4'ha;
assign core_sleep_o = ~ /* src = "generated/sv2v_out.v:20413.24-20413.33" */ clock_en;
assign _20_ = _19_ | /* src = "generated/sv2v_out.v:20400.24-20400.75" */ debug_req_i;
assign _22_ = _20_ | /* src = "generated/sv2v_out.v:20400.23-20400.90" */ irq_pending;
assign clock_en = _22_ | /* src = "generated/sv2v_out.v:20400.22-20400.102" */ irq_nm_i;
assign alert_major_internal_o = core_alert_major_internal | /* src = "generated/sv2v_out.v:20942.34-20942.119" */ rf_alert_major_internal;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20414.20-20419.3" */
prim_clock_gating core_clock_gate_i (
.clk_i(clk_i),
.clk_o(clk),
.en_i(clock_en),
.en_i_t0(core_sleep_o_t0),
.test_en_i(test_en_i),
.test_en_i_t0(test_en_i_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20394.6-20399.5" */
\$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_flop  \g_clock_en_secure.u_prim_core_busy_flop  (
.clk_i(clk_i),
.d_i(core_busy_d),
.d_i_t0(core_busy_d_t0),
.q_o(core_busy_q),
.q_o_t0(core_busy_q_t0),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20753.26-20756.5" */
\$paramod\prim_buf\Width=s32'00000000000000000000000000000111  \gen_mem_wdata_ecc.u_prim_buf_data_wdata_intg  (
.in_i(data_wdata_core[38:32]),
.in_i_t0(data_wdata_core_t0[38:32]),
.out_o(data_wdata_intg_o),
.out_o_t0(data_wdata_intg_o_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20544.6-20558.5" */
\$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  \gen_regfile_ff.register_file_i  (
.clk_i(clk),
.dummy_instr_id_i(dummy_instr_id),
.dummy_instr_id_i_t0(dummy_instr_id_t0),
.dummy_instr_wb_i(dummy_instr_wb),
.dummy_instr_wb_i_t0(dummy_instr_wb_t0),
.err_o(rf_alert_major_internal),
.err_o_t0(rf_alert_major_internal_t0),
.raddr_a_i(rf_raddr_a),
.raddr_a_i_t0(rf_raddr_a_t0),
.raddr_b_i(rf_raddr_b),
.raddr_b_i_t0(rf_raddr_b_t0),
.rdata_a_o(rf_rdata_a_ecc),
.rdata_a_o_t0(rf_rdata_a_ecc_t0),
.rdata_b_o(rf_rdata_b_ecc),
.rdata_b_o_t0(rf_rdata_b_ecc_t0),
.rst_ni(rst_ni),
.test_en_i(test_en_i),
.test_en_i_t0(test_en_i_t0),
.waddr_a_i(rf_waddr_wb),
.waddr_a_i_t0(rf_waddr_wb_t0),
.wdata_a_i(rf_wdata_wb_ecc),
.wdata_a_i_t0(rf_wdata_wb_ecc_t0),
.we_a_i(rf_we_wb),
.we_a_i_t0(rf_we_wb_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20420.24-20423.3" */
\$paramod\prim_buf\Width=s32'00000000000000000000000000000100  u_fetch_enable_buf (
.in_i(fetch_enable_i),
.in_i_t0(fetch_enable_i_t0),
.out_o(fetch_enable_buf),
.out_o_t0(fetch_enable_buf_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20474.4-20529.3" */
\$paramod$8d906854a94bfc59042b9faf57c7a7f19e3f03e7\ibex_core  u_ibex_core (
.alert_major_bus_o(alert_major_bus_o),
.alert_major_bus_o_t0(alert_major_bus_o_t0),
.alert_major_internal_o(core_alert_major_internal),
.alert_major_internal_o_t0(core_alert_major_internal_t0),
.alert_minor_o(alert_minor_o),
.alert_minor_o_t0(alert_minor_o_t0),
.boot_addr_i(boot_addr_i),
.boot_addr_i_t0(boot_addr_i_t0),
.clk_i(clk),
.core_busy_o(core_busy_d),
.core_busy_o_t0(core_busy_d_t0),
.crash_dump_o(crash_dump_o),
.crash_dump_o_t0(crash_dump_o_t0),
.data_addr_o(data_addr_o),
.data_addr_o_t0(data_addr_o_t0),
.data_be_o(data_be_o),
.data_be_o_t0(data_be_o_t0),
.data_err_i(data_err_i),
.data_err_i_t0(data_err_i_t0),
.data_gnt_i(data_gnt_i),
.data_gnt_i_t0(data_gnt_i_t0),
.data_rdata_i({ data_rdata_intg_i, data_rdata_i }),
.data_rdata_i_t0({ data_rdata_intg_i_t0, data_rdata_i_t0 }),
.data_req_o(data_req_o),
.data_req_o_t0(data_req_o_t0),
.data_rvalid_i(data_rvalid_i),
.data_rvalid_i_t0(data_rvalid_i_t0),
.data_wdata_o(data_wdata_core),
.data_wdata_o_t0(data_wdata_core_t0),
.data_we_o(data_we_o),
.data_we_o_t0(data_we_o_t0),
.debug_req_i(debug_req_i),
.debug_req_i_t0(debug_req_i_t0),
.double_fault_seen_o(double_fault_seen_o),
.double_fault_seen_o_t0(double_fault_seen_o_t0),
.dummy_instr_id_o(dummy_instr_id),
.dummy_instr_id_o_t0(dummy_instr_id_t0),
.dummy_instr_wb_o(dummy_instr_wb),
.dummy_instr_wb_o_t0(dummy_instr_wb_t0),
.fetch_enable_i(fetch_enable_buf),
.fetch_enable_i_t0(fetch_enable_buf_t0),
.hart_id_i(hart_id_i),
.hart_id_i_t0(hart_id_i_t0),
.ic_data_addr_o(ic_data_addr),
.ic_data_addr_o_t0(ic_data_addr_t0),
.ic_data_rdata_i(128'h00000000000000000000000000000000),
.ic_data_rdata_i_t0(128'h00000000000000000000000000000000),
.ic_data_req_o(ic_data_req),
.ic_data_req_o_t0(ic_data_req_t0),
.ic_data_wdata_o(ic_data_wdata),
.ic_data_wdata_o_t0(ic_data_wdata_t0),
.ic_data_write_o(ic_data_write),
.ic_data_write_o_t0(ic_data_write_t0),
.ic_scr_key_req_o(ic_scr_key_req),
.ic_scr_key_req_o_t0(ic_scr_key_req_t0),
.ic_scr_key_valid_i(1'h1),
.ic_scr_key_valid_i_t0(1'h0),
.ic_tag_addr_o(ic_tag_addr),
.ic_tag_addr_o_t0(ic_tag_addr_t0),
.ic_tag_rdata_i(44'h00000000000),
.ic_tag_rdata_i_t0(44'h00000000000),
.ic_tag_req_o(ic_tag_req),
.ic_tag_req_o_t0(ic_tag_req_t0),
.ic_tag_wdata_o(ic_tag_wdata),
.ic_tag_wdata_o_t0(ic_tag_wdata_t0),
.ic_tag_write_o(ic_tag_write),
.ic_tag_write_o_t0(ic_tag_write_t0),
.instr_addr_o(instr_addr_o),
.instr_addr_o_t0(instr_addr_o_t0),
.instr_err_i(instr_err_i),
.instr_err_i_t0(instr_err_i_t0),
.instr_gnt_i(instr_gnt_i),
.instr_gnt_i_t0(instr_gnt_i_t0),
.instr_rdata_i({ instr_rdata_intg_i, instr_rdata_i }),
.instr_rdata_i_t0({ instr_rdata_intg_i_t0, instr_rdata_i_t0 }),
.instr_req_o(instr_req_o),
.instr_req_o_t0(instr_req_o_t0),
.instr_rvalid_i(instr_rvalid_i),
.instr_rvalid_i_t0(instr_rvalid_i_t0),
.irq_external_i(irq_external_i),
.irq_external_i_t0(irq_external_i_t0),
.irq_fast_i(irq_fast_i),
.irq_fast_i_t0(irq_fast_i_t0),
.irq_nm_i(irq_nm_i),
.irq_nm_i_t0(irq_nm_i_t0),
.irq_pending_o(irq_pending),
.irq_pending_o_t0(irq_pending_t0),
.irq_software_i(irq_software_i),
.irq_software_i_t0(irq_software_i_t0),
.irq_timer_i(irq_timer_i),
.irq_timer_i_t0(irq_timer_i_t0),
.rf_raddr_a_o(rf_raddr_a),
.rf_raddr_a_o_t0(rf_raddr_a_t0),
.rf_raddr_b_o(rf_raddr_b),
.rf_raddr_b_o_t0(rf_raddr_b_t0),
.rf_rdata_a_ecc_i(rf_rdata_a_ecc_buf),
.rf_rdata_a_ecc_i_t0(rf_rdata_a_ecc_buf_t0),
.rf_rdata_b_ecc_i(rf_rdata_b_ecc_buf),
.rf_rdata_b_ecc_i_t0(rf_rdata_b_ecc_buf_t0),
.rf_waddr_wb_o(rf_waddr_wb),
.rf_waddr_wb_o_t0(rf_waddr_wb_t0),
.rf_wdata_wb_ecc_o(rf_wdata_wb_ecc),
.rf_wdata_wb_ecc_o_t0(rf_wdata_wb_ecc_t0),
.rf_we_wb_o(rf_we_wb),
.rf_we_wb_o_t0(rf_we_wb_t0),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20424.39-20427.3" */
\$paramod\prim_buf\Width=32'00000000000000000000000000100111  u_rf_rdata_a_ecc_buf (
.in_i(rf_rdata_a_ecc),
.in_i_t0(rf_rdata_a_ecc_t0),
.out_o(rf_rdata_a_ecc_buf),
.out_o_t0(rf_rdata_a_ecc_buf_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20428.39-20431.3" */
\$paramod\prim_buf\Width=32'00000000000000000000000000100111  u_rf_rdata_b_ecc_buf (
.in_i(rf_rdata_b_ecc),
.in_i_t0(rf_rdata_b_ecc_t0),
.out_o(rf_rdata_b_ecc_buf),
.out_o_t0(rf_rdata_b_ecc_buf_t0)
);
assign data_wdata_o = data_wdata_core[31:0];
assign data_wdata_o_t0 = data_wdata_core_t0[31:0];
assign scramble_req_o = 1'h0;
assign scramble_req_o_t0 = 1'h0;
endmodule

module prim_clock_gating(clk_i, en_i, test_en_i, clk_o, clk_o_t0, en_i_t0, test_en_i_t0);
/* src = "generated/sv2v_out.v:23125.2-23127.32" */
wire _00_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:23125.2-23127.32" */
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
/* src = "generated/sv2v_out.v:23120.8-23120.13" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:23123.14-23123.19" */
output clk_o;
wire clk_o;
/* cellift = 32'd1 */
output clk_o_t0;
wire clk_o_t0;
/* src = "generated/sv2v_out.v:23121.8-23121.12" */
input en_i;
wire en_i;
/* cellift = 32'd1 */
input en_i_t0;
wire en_i_t0;
/* src = "generated/sv2v_out.v:23124.6-23124.14" */
reg en_latch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:23124.6-23124.14" */
reg en_latch_t0;
/* src = "generated/sv2v_out.v:23122.8-23122.17" */
input test_en_i;
wire test_en_i;
/* cellift = 32'd1 */
input test_en_i_t0;
wire test_en_i_t0;
assign clk_o = en_latch & /* src = "generated/sv2v_out.v:23128.17-23128.33" */ clk_i;
assign clk_o_t0 = en_latch_t0 & clk_i;
/* taint_latch = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME prim_clock_gating */
/* PC_TAINT_INFO STATE_NAME en_latch_t0 */
always_latch
if (!clk_i) en_latch_t0 = _01_;
assign _02_ = ~ en_i;
assign _03_ = ~ test_en_i;
assign _04_ = en_i_t0 & _03_;
assign _05_ = test_en_i_t0 & _02_;
assign _06_ = en_i_t0 & test_en_i_t0;
assign _07_ = _04_ | _05_;
assign _01_ = _07_ | _06_;
/* src = "generated/sv2v_out.v:23125.2-23127.32" */
/* PC_TAINT_INFO MODULE_NAME prim_clock_gating */
/* PC_TAINT_INFO STATE_NAME en_latch */
always_latch
if (!clk_i) en_latch = _00_;
assign _00_ = en_i | /* src = "generated/sv2v_out.v:23127.15-23127.31" */ test_en_i;
endmodule

module prim_secded_inv_39_32_dec(data_i, data_o, syndrome_o, err_o, syndrome_o_t0, err_o_t0, data_o_t0, data_i_t0);
/* src = "generated/sv2v_out.v:29338.21-29338.63" */
wire [38:0] _000_;
/* src = "generated/sv2v_out.v:29340.21-29340.63" */
wire [38:0] _001_;
/* src = "generated/sv2v_out.v:29342.21-29342.63" */
wire [38:0] _002_;
/* src = "generated/sv2v_out.v:29344.16-29344.35" */
wire _003_;
/* src = "generated/sv2v_out.v:29345.16-29345.35" */
wire _004_;
/* src = "generated/sv2v_out.v:29346.16-29346.35" */
wire _005_;
/* src = "generated/sv2v_out.v:29347.16-29347.35" */
wire _006_;
/* src = "generated/sv2v_out.v:29348.16-29348.35" */
wire _007_;
/* src = "generated/sv2v_out.v:29349.16-29349.35" */
wire _008_;
/* src = "generated/sv2v_out.v:29350.16-29350.35" */
wire _009_;
/* src = "generated/sv2v_out.v:29351.16-29351.35" */
wire _010_;
/* src = "generated/sv2v_out.v:29352.16-29352.35" */
wire _011_;
/* src = "generated/sv2v_out.v:29353.16-29353.35" */
wire _012_;
/* src = "generated/sv2v_out.v:29354.17-29354.36" */
wire _013_;
/* src = "generated/sv2v_out.v:29355.17-29355.36" */
wire _014_;
/* src = "generated/sv2v_out.v:29356.17-29356.36" */
wire _015_;
/* src = "generated/sv2v_out.v:29357.17-29357.36" */
wire _016_;
/* src = "generated/sv2v_out.v:29358.17-29358.36" */
wire _017_;
/* src = "generated/sv2v_out.v:29359.17-29359.36" */
wire _018_;
/* src = "generated/sv2v_out.v:29360.17-29360.36" */
wire _019_;
/* src = "generated/sv2v_out.v:29361.17-29361.36" */
wire _020_;
/* src = "generated/sv2v_out.v:29362.17-29362.36" */
wire _021_;
/* src = "generated/sv2v_out.v:29363.17-29363.36" */
wire _022_;
/* src = "generated/sv2v_out.v:29364.17-29364.36" */
wire _023_;
/* src = "generated/sv2v_out.v:29365.17-29365.36" */
wire _024_;
/* src = "generated/sv2v_out.v:29366.17-29366.36" */
wire _025_;
/* src = "generated/sv2v_out.v:29367.17-29367.36" */
wire _026_;
/* src = "generated/sv2v_out.v:29368.17-29368.36" */
wire _027_;
/* src = "generated/sv2v_out.v:29369.17-29369.36" */
wire _028_;
/* src = "generated/sv2v_out.v:29370.17-29370.36" */
wire _029_;
/* src = "generated/sv2v_out.v:29371.17-29371.36" */
wire _030_;
/* src = "generated/sv2v_out.v:29372.17-29372.36" */
wire _031_;
/* src = "generated/sv2v_out.v:29373.17-29373.36" */
wire _032_;
/* src = "generated/sv2v_out.v:29374.17-29374.36" */
wire _033_;
/* src = "generated/sv2v_out.v:29375.17-29375.36" */
wire _034_;
/* src = "generated/sv2v_out.v:29377.14-29377.23" */
wire _035_;
/* src = "generated/sv2v_out.v:29377.26-29377.37" */
wire _036_;
/* src = "generated/sv2v_out.v:29332.15-29332.21" */
input [38:0] data_i;
wire [38:0] data_i;
/* cellift = 32'd1 */
input [38:0] data_i_t0;
wire [38:0] data_i_t0;
/* src = "generated/sv2v_out.v:29333.20-29333.26" */
output [31:0] data_o;
wire [31:0] data_o;
/* cellift = 32'd1 */
output [31:0] data_o_t0;
wire [31:0] data_o_t0;
/* src = "generated/sv2v_out.v:29335.19-29335.24" */
output [1:0] err_o;
wire [1:0] err_o;
/* cellift = 32'd1 */
output [1:0] err_o_t0;
wire [1:0] err_o_t0;
/* src = "generated/sv2v_out.v:29334.19-29334.29" */
output [6:0] syndrome_o;
wire [6:0] syndrome_o;
/* cellift = 32'd1 */
output [6:0] syndrome_o_t0;
wire [6:0] syndrome_o_t0;
assign err_o[1] = _035_ & /* src = "generated/sv2v_out.v:29377.14-29377.37" */ _036_;
assign { _002_[37], _001_[35], _000_[33] } = ~ { data_i[37], data_i[35], data_i[33] };
assign _003_ = syndrome_o == /* src = "generated/sv2v_out.v:29344.16-29344.35" */ 7'h19;
assign _004_ = syndrome_o == /* src = "generated/sv2v_out.v:29345.16-29345.35" */ 7'h54;
assign _005_ = syndrome_o == /* src = "generated/sv2v_out.v:29346.16-29346.35" */ 7'h61;
assign _006_ = syndrome_o == /* src = "generated/sv2v_out.v:29347.16-29347.35" */ 7'h34;
assign _007_ = syndrome_o == /* src = "generated/sv2v_out.v:29348.16-29348.35" */ 7'h1a;
assign _008_ = syndrome_o == /* src = "generated/sv2v_out.v:29349.16-29349.35" */ 7'h15;
assign _009_ = syndrome_o == /* src = "generated/sv2v_out.v:29350.16-29350.35" */ 7'h2a;
assign _010_ = syndrome_o == /* src = "generated/sv2v_out.v:29351.16-29351.35" */ 7'h4c;
assign _011_ = syndrome_o == /* src = "generated/sv2v_out.v:29352.16-29352.35" */ 7'h45;
assign _012_ = syndrome_o == /* src = "generated/sv2v_out.v:29353.16-29353.35" */ 7'h38;
assign _013_ = syndrome_o == /* src = "generated/sv2v_out.v:29354.17-29354.36" */ 7'h49;
assign _014_ = syndrome_o == /* src = "generated/sv2v_out.v:29355.17-29355.36" */ 7'h0d;
assign _015_ = syndrome_o == /* src = "generated/sv2v_out.v:29356.17-29356.36" */ 7'h51;
assign _016_ = syndrome_o == /* src = "generated/sv2v_out.v:29357.17-29357.36" */ 7'h31;
assign _017_ = syndrome_o == /* src = "generated/sv2v_out.v:29358.17-29358.36" */ 7'h68;
assign _018_ = syndrome_o == /* src = "generated/sv2v_out.v:29359.17-29359.36" */ 7'h07;
assign _019_ = syndrome_o == /* src = "generated/sv2v_out.v:29360.17-29360.36" */ 7'h1c;
assign _020_ = syndrome_o == /* src = "generated/sv2v_out.v:29361.17-29361.36" */ 7'h0b;
assign _021_ = syndrome_o == /* src = "generated/sv2v_out.v:29362.17-29362.36" */ 7'h25;
assign _022_ = syndrome_o == /* src = "generated/sv2v_out.v:29363.17-29363.36" */ 7'h26;
assign _023_ = syndrome_o == /* src = "generated/sv2v_out.v:29364.17-29364.36" */ 7'h46;
assign _024_ = syndrome_o == /* src = "generated/sv2v_out.v:29365.17-29365.36" */ 7'h0e;
assign _025_ = syndrome_o == /* src = "generated/sv2v_out.v:29366.17-29366.36" */ 7'h70;
assign _026_ = syndrome_o == /* src = "generated/sv2v_out.v:29367.17-29367.36" */ 7'h32;
assign _027_ = syndrome_o == /* src = "generated/sv2v_out.v:29368.17-29368.36" */ 7'h2c;
assign _028_ = syndrome_o == /* src = "generated/sv2v_out.v:29369.17-29369.36" */ 7'h13;
assign _029_ = syndrome_o == /* src = "generated/sv2v_out.v:29370.17-29370.36" */ 7'h23;
assign _030_ = syndrome_o == /* src = "generated/sv2v_out.v:29371.17-29371.36" */ 7'h62;
assign _031_ = syndrome_o == /* src = "generated/sv2v_out.v:29372.17-29372.36" */ 7'h4a;
assign _032_ = syndrome_o == /* src = "generated/sv2v_out.v:29373.17-29373.36" */ 7'h29;
assign _033_ = syndrome_o == /* src = "generated/sv2v_out.v:29374.17-29374.36" */ 7'h16;
assign _034_ = syndrome_o == /* src = "generated/sv2v_out.v:29375.17-29375.36" */ 7'h52;
assign _035_ = ~ /* src = "generated/sv2v_out.v:29377.14-29377.23" */ err_o[0];
assign _036_ = | /* src = "generated/sv2v_out.v:29377.26-29377.37" */ syndrome_o;
assign syndrome_o[0] = ^ /* src = "generated/sv2v_out.v:29337.19-29337.64" */ { 6'h00, data_i[32], 2'h0, data_i[29], 2'h0, data_i[26:25], 6'h00, data_i[18:17], 1'h0, data_i[15], 1'h0, data_i[13:10], 1'h0, data_i[8], 2'h0, data_i[5], 2'h0, data_i[2], 1'h0, data_i[0] };
assign syndrome_o[1] = ^ /* src = "generated/sv2v_out.v:29338.19-29338.64" */ { 5'h00, _000_[33], 1'h0, data_i[31:30], 1'h0, data_i[28:25], 1'h0, data_i[23], 1'h0, data_i[21:19], 1'h0, data_i[17], 1'h0, data_i[15], 8'h00, data_i[6], 1'h0, data_i[4], 4'h0 };
assign syndrome_o[2] = ^ /* src = "generated/sv2v_out.v:29339.19-29339.64" */ { 4'h0, data_i[34], 3'h0, data_i[30], 5'h00, data_i[24], 2'h0, data_i[21:18], 1'h0, data_i[16:15], 3'h0, data_i[11], 2'h0, data_i[8:7], 1'h0, data_i[5], 1'h0, data_i[3], 1'h0, data_i[1], 1'h0 };
assign syndrome_o[3] = ^ /* src = "generated/sv2v_out.v:29340.19-29340.64" */ { 3'h0, _001_[35], 5'h00, data_i[29:28], 3'h0, data_i[24], 2'h0, data_i[21], 3'h0, data_i[17:16], 1'h0, data_i[14], 2'h0, data_i[11:9], 1'h0, data_i[7:6], 1'h0, data_i[4], 3'h0, data_i[0] };
assign syndrome_o[4] = ^ /* src = "generated/sv2v_out.v:29341.19-29341.64" */ { 2'h0, data_i[36], 4'h0, data_i[31:30], 4'h0, data_i[25], 1'h0, data_i[23:22], 5'h00, data_i[16], 2'h0, data_i[13:12], 2'h0, data_i[9], 3'h0, data_i[5:3], 1'h0, data_i[1:0] };
assign syndrome_o[5] = ^ /* src = "generated/sv2v_out.v:29342.19-29342.64" */ { 1'h0, _002_[37], 7'h00, data_i[29], 1'h0, data_i[27:26], 1'h0, data_i[24:22], 2'h0, data_i[19:18], 3'h0, data_i[14:13], 3'h0, data_i[9], 2'h0, data_i[6], 2'h0, data_i[3:2], 2'h0 };
assign syndrome_o[6] = ^ /* src = "generated/sv2v_out.v:29343.19-29343.64" */ { data_i[38], 6'h00, data_i[31], 2'h0, data_i[28:27], 4'h0, data_i[22], 1'h0, data_i[20], 5'h00, data_i[14], 1'h0, data_i[12], 1'h0, data_i[10], 1'h0, data_i[8:7], 4'h0, data_i[2:1], 1'h0 };
assign err_o[0] = ^ /* src = "generated/sv2v_out.v:29376.14-29376.25" */ syndrome_o;
assign data_o[0] = _003_ ^ /* src = "generated/sv2v_out.v:29344.15-29344.48" */ data_i[0];
assign data_o[1] = _004_ ^ /* src = "generated/sv2v_out.v:29345.15-29345.48" */ data_i[1];
assign data_o[2] = _005_ ^ /* src = "generated/sv2v_out.v:29346.15-29346.48" */ data_i[2];
assign data_o[3] = _006_ ^ /* src = "generated/sv2v_out.v:29347.15-29347.48" */ data_i[3];
assign data_o[4] = _007_ ^ /* src = "generated/sv2v_out.v:29348.15-29348.48" */ data_i[4];
assign data_o[5] = _008_ ^ /* src = "generated/sv2v_out.v:29349.15-29349.48" */ data_i[5];
assign data_o[6] = _009_ ^ /* src = "generated/sv2v_out.v:29350.15-29350.48" */ data_i[6];
assign data_o[7] = _010_ ^ /* src = "generated/sv2v_out.v:29351.15-29351.48" */ data_i[7];
assign data_o[8] = _011_ ^ /* src = "generated/sv2v_out.v:29352.15-29352.48" */ data_i[8];
assign data_o[9] = _012_ ^ /* src = "generated/sv2v_out.v:29353.15-29353.48" */ data_i[9];
assign data_o[10] = _013_ ^ /* src = "generated/sv2v_out.v:29354.16-29354.50" */ data_i[10];
assign data_o[11] = _014_ ^ /* src = "generated/sv2v_out.v:29355.16-29355.50" */ data_i[11];
assign data_o[12] = _015_ ^ /* src = "generated/sv2v_out.v:29356.16-29356.50" */ data_i[12];
assign data_o[13] = _016_ ^ /* src = "generated/sv2v_out.v:29357.16-29357.50" */ data_i[13];
assign data_o[14] = _017_ ^ /* src = "generated/sv2v_out.v:29358.16-29358.50" */ data_i[14];
assign data_o[15] = _018_ ^ /* src = "generated/sv2v_out.v:29359.16-29359.50" */ data_i[15];
assign data_o[16] = _019_ ^ /* src = "generated/sv2v_out.v:29360.16-29360.50" */ data_i[16];
assign data_o[17] = _020_ ^ /* src = "generated/sv2v_out.v:29361.16-29361.50" */ data_i[17];
assign data_o[18] = _021_ ^ /* src = "generated/sv2v_out.v:29362.16-29362.50" */ data_i[18];
assign data_o[19] = _022_ ^ /* src = "generated/sv2v_out.v:29363.16-29363.50" */ data_i[19];
assign data_o[20] = _023_ ^ /* src = "generated/sv2v_out.v:29364.16-29364.50" */ data_i[20];
assign data_o[21] = _024_ ^ /* src = "generated/sv2v_out.v:29365.16-29365.50" */ data_i[21];
assign data_o[22] = _025_ ^ /* src = "generated/sv2v_out.v:29366.16-29366.50" */ data_i[22];
assign data_o[23] = _026_ ^ /* src = "generated/sv2v_out.v:29367.16-29367.50" */ data_i[23];
assign data_o[24] = _027_ ^ /* src = "generated/sv2v_out.v:29368.16-29368.50" */ data_i[24];
assign data_o[25] = _028_ ^ /* src = "generated/sv2v_out.v:29369.16-29369.50" */ data_i[25];
assign data_o[26] = _029_ ^ /* src = "generated/sv2v_out.v:29370.16-29370.50" */ data_i[26];
assign data_o[27] = _030_ ^ /* src = "generated/sv2v_out.v:29371.16-29371.50" */ data_i[27];
assign data_o[28] = _031_ ^ /* src = "generated/sv2v_out.v:29372.16-29372.50" */ data_i[28];
assign data_o[29] = _032_ ^ /* src = "generated/sv2v_out.v:29373.16-29373.50" */ data_i[29];
assign data_o[30] = _033_ ^ /* src = "generated/sv2v_out.v:29374.16-29374.50" */ data_i[30];
assign data_o[31] = _034_ ^ /* src = "generated/sv2v_out.v:29375.16-29375.50" */ data_i[31];
assign { _000_[38:34], _000_[32:0] } = { 6'h00, data_i[31:30], 1'h0, data_i[28:25], 1'h0, data_i[23], 1'h0, data_i[21:19], 1'h0, data_i[17], 1'h0, data_i[15], 8'h00, data_i[6], 1'h0, data_i[4], 4'h0 };
assign { _001_[38:36], _001_[34:0] } = { 8'h00, data_i[29:28], 3'h0, data_i[24], 2'h0, data_i[21], 3'h0, data_i[17:16], 1'h0, data_i[14], 2'h0, data_i[11:9], 1'h0, data_i[7:6], 1'h0, data_i[4], 3'h0, data_i[0] };
assign { _002_[38], _002_[36:0] } = { 8'h00, data_i[29], 1'h0, data_i[27:26], 1'h0, data_i[24:22], 2'h0, data_i[19:18], 3'h0, data_i[14:13], 3'h0, data_i[9], 2'h0, data_i[6], 2'h0, data_i[3:2], 2'h0 };
assign data_o_t0 = data_i_t0[31:0];
assign err_o_t0 = 2'h0;
assign syndrome_o_t0 = 7'h00;
endmodule

module prim_secded_inv_39_32_enc(data_i, data_o, data_o_t0, data_i_t0);
/* src = "generated/sv2v_out.v:29393.16-29393.42" */
wire _00_;
/* src = "generated/sv2v_out.v:29395.16-29395.42" */
wire _01_;
/* src = "generated/sv2v_out.v:29397.16-29397.42" */
wire _02_;
/* src = "generated/sv2v_out.v:29384.15-29384.21" */
input [31:0] data_i;
wire [31:0] data_i;
/* cellift = 32'd1 */
input [31:0] data_i_t0;
wire [31:0] data_i_t0;
/* src = "generated/sv2v_out.v:29385.20-29385.26" */
output [38:0] data_o;
wire [38:0] data_o;
/* cellift = 32'd1 */
output [38:0] data_o_t0;
wire [38:0] data_o_t0;
assign { data_o[37], data_o[35], data_o[33] } = ~ { _02_, _01_, _00_ };
assign data_o[32] = ^ /* src = "generated/sv2v_out.v:29392.16-29392.42" */ { 9'h000, data_i[29], 2'h0, data_i[26:25], 6'h00, data_i[18:17], 1'h0, data_i[15], 1'h0, data_i[13:10], 1'h0, data_i[8], 2'h0, data_i[5], 2'h0, data_i[2], 1'h0, data_i[0] };
assign _00_ = ^ /* src = "generated/sv2v_out.v:29393.16-29393.42" */ { 7'h00, data_i[31:30], 1'h0, data_i[28:25], 1'h0, data_i[23], 1'h0, data_i[21:19], 1'h0, data_i[17], 1'h0, data_i[15], 8'h00, data_i[6], 1'h0, data_i[4], 4'h0 };
assign data_o[34] = ^ /* src = "generated/sv2v_out.v:29394.16-29394.42" */ { 8'h00, data_i[30], 5'h00, data_i[24], 2'h0, data_i[21:18], 1'h0, data_i[16:15], 3'h0, data_i[11], 2'h0, data_i[8:7], 1'h0, data_i[5], 1'h0, data_i[3], 1'h0, data_i[1], 1'h0 };
assign _01_ = ^ /* src = "generated/sv2v_out.v:29395.16-29395.42" */ { 9'h000, data_i[29:28], 3'h0, data_i[24], 2'h0, data_i[21], 3'h0, data_i[17:16], 1'h0, data_i[14], 2'h0, data_i[11:9], 1'h0, data_i[7:6], 1'h0, data_i[4], 3'h0, data_i[0] };
assign data_o[36] = ^ /* src = "generated/sv2v_out.v:29396.16-29396.42" */ { 7'h00, data_i[31:30], 4'h0, data_i[25], 1'h0, data_i[23:22], 5'h00, data_i[16], 2'h0, data_i[13:12], 2'h0, data_i[9], 3'h0, data_i[5:3], 1'h0, data_i[1:0] };
assign _02_ = ^ /* src = "generated/sv2v_out.v:29397.16-29397.42" */ { 9'h000, data_i[29], 1'h0, data_i[27:26], 1'h0, data_i[24:22], 2'h0, data_i[19:18], 3'h0, data_i[14:13], 3'h0, data_i[9], 2'h0, data_i[6], 2'h0, data_i[3:2], 2'h0 };
assign data_o[38] = ^ /* src = "generated/sv2v_out.v:29398.16-29398.42" */ { 7'h00, data_i[31], 2'h0, data_i[28:27], 4'h0, data_i[22], 1'h0, data_i[20], 5'h00, data_i[14], 1'h0, data_i[12], 1'h0, data_i[10], 1'h0, data_i[8:7], 4'h0, data_i[2:1], 1'h0 };
assign data_o[31:0] = data_i;
assign data_o_t0 = { 7'h00, data_i_t0 };
endmodule