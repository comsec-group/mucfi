bit gen_uc_rs1;
assign gen_uc_rs1 = ((1'h1));
