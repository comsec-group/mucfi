module cellift_scarv_fpv 
(
g_clk,
g_resetn,
trs_pc,
trs_instr,
trs_valid,
leak_prng,
leak_fence_unc0,
leak_fence_unc1,
leak_fence_unc2,
rng_req_valid,
rng_req_op,
rng_req_data,
rng_req_ready,
rng_rsp_valid,
rng_rsp_status,
rng_rsp_data,
rng_rsp_ready,
int_nmi,
int_external,
int_extern_cause,
int_software,
int_mtime,
imem_req,
imem_wen,
imem_strb,
imem_wdata,
imem_addr,
imem_gnt,
imem_recv,
imem_ack,
imem_error,
imem_rdata,
dmem_req,
dmem_wen,
dmem_strb,
dmem_wdata,
dmem_addr,
dmem_gnt,
dmem_recv,
dmem_ack,
dmem_error,
dmem_rdata,
leak_prng_t0,
imem_wen_t0,
imem_wdata_t0,
imem_strb_t0,
imem_req_t0,
imem_recv_t0,
imem_rdata_t0,
imem_gnt_t0,
imem_error_t0,
imem_addr_t0,
imem_ack_t0,
rng_req_data_t0,
rng_req_op_t0,
rng_req_ready_t0,
rng_req_valid_t0,
rng_rsp_data_t0,
rng_rsp_ready_t0,
rng_rsp_status_t0,
rng_rsp_valid_t0,
dmem_addr_t0,
dmem_gnt_t0,
dmem_req_t0,
dmem_strb_t0,
dmem_wdata_t0,
dmem_wen_t0,
leak_fence_unc0_t0,
leak_fence_unc1_t0,
leak_fence_unc2_t0,
dmem_ack_t0,
dmem_error_t0,
dmem_rdata_t0,
dmem_recv_t0,
trs_instr_t0,
trs_pc_t0,
trs_valid_t0,
int_extern_cause_t0,
int_external_t0,
int_mtime_t0,
int_nmi_t0,
int_software_t0,
ctr_cycle_t0,
ctr_cycle,
ctr_instret_t0,
ctr_instret,
ctr_time_t0,
ctr_time,
inhibit_cy_t0,
inhibit_cy,
inhibit_ir_t0,
inhibit_ir,
inhibit_tm_t0,
inhibit_tm,
instr_ret_t0,
instr_ret,
int_trap_ack_t0,
int_trap_ack,
int_trap_cause_t0,
int_trap_cause,
int_trap_req_t0,
int_trap_req,
mie_meie_t0,
mie_meie,
mie_msie_t0,
mie_msie,
mie_mtie_t0,
mie_mtie,
mip_meip_t0,
mip_meip,
mip_msip_t0,
mip_msip,
mmio_addr_t0,
mmio_addr,
mmio_en_t0,
mmio_en,
mmio_error_t0,
mmio_error,
mmio_rdata_t0,
mmio_rdata,
mmio_wdata_t0,
mmio_wdata,
mmio_wen_t0,
mmio_wen,
mstatus_mie_t0,
mstatus_mie,
ti_pending_t0,
ti_pending,
i_counters__g_clk,
i_counters__g_resetn,
i_counters__instr_ret,
i_counters__timer_interrupt,
i_counters__ctr_time,
i_counters__ctr_cycle,
i_counters__ctr_instret,
i_counters__inhibit_cy,
i_counters__inhibit_tm,
i_counters__inhibit_ir,
i_counters__mmio_en,
i_counters__mmio_wen,
i_counters__mmio_addr,
i_counters__mmio_wdata,
i_counters__mmio_rdata,
i_counters__mmio_error,
i_counters__timer_interrupt_t0,
i_counters__mmio_wen_t0,
i_counters__mmio_wdata_t0,
i_counters__mmio_rdata_t0,
i_counters__mmio_error_t0,
i_counters__mmio_en_t0,
i_counters__mmio_addr_t0,
i_counters__instr_ret_t0,
i_counters__inhibit_tm_t0,
i_counters__inhibit_ir_t0,
i_counters__inhibit_cy_t0,
i_counters__ctr_time_t0,
i_counters__ctr_instret_t0,
i_counters__ctr_cycle_t0,
i_counters__addr_mtime_hi_t0,
i_counters__addr_mtime_hi,
i_counters__addr_mtime_lo_t0,
i_counters__addr_mtime_lo,
i_counters__addr_mtimecmp_hi_t0,
i_counters__addr_mtimecmp_hi,
i_counters__addr_mtimecmp_lo_t0,
i_counters__addr_mtimecmp_lo,
i_counters__mapped_mtimecmp_t0,
i_counters__mapped_mtimecmp,
i_counters__n_ctr_cycle_t0,
i_counters__n_ctr_cycle,
i_counters__n_ctr_instret_t0,
i_counters__n_ctr_instret,
i_counters__n_mapped_mtime_t0,
i_counters__n_mapped_mtime,
i_counters__n_mmio_error_t0,
i_counters__n_mmio_error,
i_counters__n_mmio_rdata_t0,
i_counters__n_mmio_rdata,
i_counters__n_timer_interrupt_t0,
i_counters__n_timer_interrupt,
i_counters__wr_mtime_hi_t0,
i_counters__wr_mtime_hi,
i_counters__wr_mtime_lo_t0,
i_counters__wr_mtime_lo,
i_counters__wr_mtimecmp_hi_t0,
i_counters__wr_mtimecmp_hi,
i_counters__wr_mtimecmp_lo_t0,
i_counters__wr_mtimecmp_lo,
i_interrupts__g_clk,
i_interrupts__g_resetn,
i_interrupts__mstatus_mie,
i_interrupts__mie_meie,
i_interrupts__mie_mtie,
i_interrupts__mie_msie,
i_interrupts__nmi_pending,
i_interrupts__ex_pending,
i_interrupts__ex_cause,
i_interrupts__ti_pending,
i_interrupts__sw_pending,
i_interrupts__mip_meip,
i_interrupts__mip_mtip,
i_interrupts__mip_msip,
i_interrupts__int_trap_req,
i_interrupts__int_trap_cause,
i_interrupts__int_trap_ack,
i_interrupts__nmi_pending_t0,
i_interrupts__mstatus_mie_t0,
i_interrupts__mip_mtip_t0,
i_interrupts__mie_mtie_t0,
i_interrupts__mie_msie_t0,
i_interrupts__sw_pending_t0,
i_interrupts__ti_pending_t0,
i_interrupts__int_trap_req_t0,
i_interrupts__ex_cause_t0,
i_interrupts__ex_pending_t0,
i_interrupts__int_trap_cause_t0,
i_interrupts__int_trap_ack_t0,
i_interrupts__mie_meie_t0,
i_interrupts__mip_msip_t0,
i_interrupts__mip_meip_t0,
i_interrupts__extern_cause_t0,
i_interrupts__extern_cause,
i_interrupts__mip_nmi_t0,
i_interrupts__mip_nmi,
i_interrupts__n_int_trap_cause_t0,
i_interrupts__n_int_trap_cause,
i_interrupts__raise_mei_t0,
i_interrupts__raise_mei,
i_interrupts__raise_msi_t0,
i_interrupts__raise_msi,
i_interrupts__raise_mti_t0,
i_interrupts__raise_mti,
i_interrupts__raise_nmi_t0,
i_interrupts__raise_nmi,
i_interrupts__use_extern_cause_t0,
i_interrupts__use_extern_cause,
i_pipeline__g_clk,
i_pipeline__g_resetn,
i_pipeline__trs_pc,
i_pipeline__trs_instr,
i_pipeline__trs_valid,
i_pipeline__leak_prng,
i_pipeline__leak_fence_unc0,
i_pipeline__leak_fence_unc1,
i_pipeline__leak_fence_unc2,
i_pipeline__rng_req_valid,
i_pipeline__rng_req_op,
i_pipeline__rng_req_data,
i_pipeline__rng_req_ready,
i_pipeline__rng_rsp_valid,
i_pipeline__rng_rsp_status,
i_pipeline__rng_rsp_data,
i_pipeline__rng_rsp_ready,
i_pipeline__instr_ret,
i_pipeline__mstatus_mie,
i_pipeline__mie_meie,
i_pipeline__mie_mtie,
i_pipeline__mie_msie,
i_pipeline__mip_meip,
i_pipeline__mip_mtip,
i_pipeline__mip_msip,
i_pipeline__ctr_time,
i_pipeline__ctr_cycle,
i_pipeline__ctr_instret,
i_pipeline__int_trap_req,
i_pipeline__int_trap_cause,
i_pipeline__int_trap_ack,
i_pipeline__inhibit_cy,
i_pipeline__inhibit_tm,
i_pipeline__inhibit_ir,
i_pipeline__mmio_en,
i_pipeline__mmio_wen,
i_pipeline__mmio_addr,
i_pipeline__mmio_wdata,
i_pipeline__mmio_rdata,
i_pipeline__mmio_error,
i_pipeline__imem_req,
i_pipeline__imem_wen,
i_pipeline__imem_strb,
i_pipeline__imem_wdata,
i_pipeline__imem_addr,
i_pipeline__imem_gnt,
i_pipeline__imem_recv,
i_pipeline__imem_ack,
i_pipeline__imem_error,
i_pipeline__imem_rdata,
i_pipeline__dmem_req,
i_pipeline__dmem_wen,
i_pipeline__dmem_strb,
i_pipeline__dmem_wdata,
i_pipeline__dmem_addr,
i_pipeline__dmem_gnt,
i_pipeline__dmem_recv,
i_pipeline__dmem_ack,
i_pipeline__dmem_error,
i_pipeline__dmem_rdata,
i_pipeline__mstatus_mie_t0,
i_pipeline__mip_mtip_t0,
i_pipeline__mie_mtie_t0,
i_pipeline__mie_msie_t0,
i_pipeline__leak_prng_t0,
i_pipeline__imem_wen_t0,
i_pipeline__imem_wdata_t0,
i_pipeline__imem_strb_t0,
i_pipeline__imem_req_t0,
i_pipeline__imem_recv_t0,
i_pipeline__imem_rdata_t0,
i_pipeline__imem_gnt_t0,
i_pipeline__imem_error_t0,
i_pipeline__imem_addr_t0,
i_pipeline__imem_ack_t0,
i_pipeline__int_trap_req_t0,
i_pipeline__mmio_wen_t0,
i_pipeline__mmio_wdata_t0,
i_pipeline__mmio_rdata_t0,
i_pipeline__mmio_error_t0,
i_pipeline__mmio_en_t0,
i_pipeline__mmio_addr_t0,
i_pipeline__instr_ret_t0,
i_pipeline__inhibit_tm_t0,
i_pipeline__inhibit_ir_t0,
i_pipeline__inhibit_cy_t0,
i_pipeline__ctr_time_t0,
i_pipeline__ctr_instret_t0,
i_pipeline__ctr_cycle_t0,
i_pipeline__int_trap_cause_t0,
i_pipeline__int_trap_ack_t0,
i_pipeline__mie_meie_t0,
i_pipeline__mip_msip_t0,
i_pipeline__mip_meip_t0,
i_pipeline__rng_req_data_t0,
i_pipeline__rng_req_op_t0,
i_pipeline__rng_req_ready_t0,
i_pipeline__rng_req_valid_t0,
i_pipeline__rng_rsp_data_t0,
i_pipeline__rng_rsp_ready_t0,
i_pipeline__rng_rsp_status_t0,
i_pipeline__rng_rsp_valid_t0,
i_pipeline__dmem_addr_t0,
i_pipeline__dmem_gnt_t0,
i_pipeline__dmem_req_t0,
i_pipeline__dmem_strb_t0,
i_pipeline__dmem_wdata_t0,
i_pipeline__dmem_wen_t0,
i_pipeline__leak_fence_unc0_t0,
i_pipeline__leak_fence_unc1_t0,
i_pipeline__leak_fence_unc2_t0,
i_pipeline__dmem_ack_t0,
i_pipeline__dmem_error_t0,
i_pipeline__dmem_rdata_t0,
i_pipeline__dmem_recv_t0,
i_pipeline__trs_instr_t0,
i_pipeline__trs_pc_t0,
i_pipeline__trs_valid_t0,
i_pipeline__cf_ack_t0,
i_pipeline__cf_ack,
i_pipeline__cf_req_t0,
i_pipeline__cf_req,
i_pipeline__cf_target_t0,
i_pipeline__cf_target,
i_pipeline__csr_addr_t0,
i_pipeline__csr_addr,
i_pipeline__csr_en_t0,
i_pipeline__csr_en,
i_pipeline__csr_error_t0,
i_pipeline__csr_error,
i_pipeline__csr_mepc_t0,
i_pipeline__csr_mepc,
i_pipeline__csr_mtvec_t0,
i_pipeline__csr_mtvec,
i_pipeline__csr_rdata_t0,
i_pipeline__csr_rdata,
i_pipeline__csr_wdata_t0,
i_pipeline__csr_wdata,
i_pipeline__csr_wr_clr_t0,
i_pipeline__csr_wr_clr,
i_pipeline__csr_wr_set_t0,
i_pipeline__csr_wr_set,
i_pipeline__csr_wr_t0,
i_pipeline__csr_wr,
i_pipeline__exec_mret_t0,
i_pipeline__exec_mret,
i_pipeline__fwd_rs1_rdata_t0,
i_pipeline__fwd_rs1_rdata,
i_pipeline__fwd_rs2_rdata_t0,
i_pipeline__fwd_rs2_rdata,
i_pipeline__fwd_rs3_rdata_t0,
i_pipeline__fwd_rs3_rdata,
i_pipeline__fwd_s2_csr_t0,
i_pipeline__fwd_s2_csr,
i_pipeline__fwd_s2_load_t0,
i_pipeline__fwd_s2_load,
i_pipeline__fwd_s2_rd_t0,
i_pipeline__fwd_s2_rd,
i_pipeline__fwd_s2_rs1_hi_t0,
i_pipeline__fwd_s2_rs1_hi,
i_pipeline__fwd_s2_rs2_hi_t0,
i_pipeline__fwd_s2_rs2_hi,
i_pipeline__fwd_s2_rs3_hi_t0,
i_pipeline__fwd_s2_rs3_hi,
i_pipeline__fwd_s2_wdata_hi_t0,
i_pipeline__fwd_s2_wdata_hi,
i_pipeline__fwd_s2_wdata_t0,
i_pipeline__fwd_s2_wdata,
i_pipeline__fwd_s2_wide_t0,
i_pipeline__fwd_s2_wide,
i_pipeline__fwd_s3_csr_t0,
i_pipeline__fwd_s3_csr,
i_pipeline__fwd_s3_load_t0,
i_pipeline__fwd_s3_load,
i_pipeline__fwd_s3_rd_t0,
i_pipeline__fwd_s3_rd,
i_pipeline__fwd_s3_rs1_hi_t0,
i_pipeline__fwd_s3_rs1_hi,
i_pipeline__fwd_s3_rs2_hi_t0,
i_pipeline__fwd_s3_rs2_hi,
i_pipeline__fwd_s3_rs3_hi_t0,
i_pipeline__fwd_s3_rs3_hi,
i_pipeline__fwd_s3_wdata_hi_t0,
i_pipeline__fwd_s3_wdata_hi,
i_pipeline__fwd_s3_wdata_t0,
i_pipeline__fwd_s3_wdata,
i_pipeline__fwd_s3_wide_t0,
i_pipeline__fwd_s3_wide,
i_pipeline__fwd_s4_csr_t0,
i_pipeline__fwd_s4_csr,
i_pipeline__fwd_s4_load_t0,
i_pipeline__fwd_s4_load,
i_pipeline__fwd_s4_rd_t0,
i_pipeline__fwd_s4_rd,
i_pipeline__fwd_s4_rs1_hi_t0,
i_pipeline__fwd_s4_rs1_hi,
i_pipeline__fwd_s4_rs2_hi_t0,
i_pipeline__fwd_s4_rs2_hi,
i_pipeline__fwd_s4_rs3_hi_t0,
i_pipeline__fwd_s4_rs3_hi,
i_pipeline__fwd_s4_wdata_t0,
i_pipeline__fwd_s4_wdata,
i_pipeline__gpr_rd_t0,
i_pipeline__gpr_rd,
i_pipeline__gpr_wdata_hi_t0,
i_pipeline__gpr_wdata_hi,
i_pipeline__gpr_wdata_t0,
i_pipeline__gpr_wdata,
i_pipeline__gpr_wen_t0,
i_pipeline__gpr_wen,
i_pipeline__gpr_wide_t0,
i_pipeline__gpr_wide,
i_pipeline__hold_lsu_req_t0,
i_pipeline__hold_lsu_req,
i_pipeline__hzd_rs1_s2_t0,
i_pipeline__hzd_rs1_s2,
i_pipeline__hzd_rs1_s3_t0,
i_pipeline__hzd_rs1_s3,
i_pipeline__hzd_rs1_s4_t0,
i_pipeline__hzd_rs1_s4,
i_pipeline__hzd_rs2_s2_t0,
i_pipeline__hzd_rs2_s2,
i_pipeline__hzd_rs2_s3_t0,
i_pipeline__hzd_rs2_s3,
i_pipeline__hzd_rs2_s4_t0,
i_pipeline__hzd_rs2_s4,
i_pipeline__hzd_rs3_s2_t0,
i_pipeline__hzd_rs3_s2,
i_pipeline__hzd_rs3_s3_t0,
i_pipeline__hzd_rs3_s3,
i_pipeline__hzd_rs3_s4_t0,
i_pipeline__hzd_rs3_s4,
i_pipeline__leak_lkgcfg_t0,
i_pipeline__leak_lkgcfg,
i_pipeline__nz_s1_rs1_t0,
i_pipeline__nz_s1_rs1,
i_pipeline__nz_s1_rs2_t0,
i_pipeline__nz_s1_rs2,
i_pipeline__nz_s1_rs3_t0,
i_pipeline__nz_s1_rs3,
i_pipeline__s0_flush_t0,
i_pipeline__s0_flush,
i_pipeline__s1_bubble_from_s2_t0,
i_pipeline__s1_bubble_from_s2,
i_pipeline__s1_bubble_from_s3_t0,
i_pipeline__s1_bubble_from_s3,
i_pipeline__s1_bubble_from_s4_t0,
i_pipeline__s1_bubble_from_s4,
i_pipeline__s1_bubble_no_instr_t0,
i_pipeline__s1_bubble_no_instr,
i_pipeline__s1_bubble_t0,
i_pipeline__s1_bubble,
i_pipeline__s1_busy_t0,
i_pipeline__s1_busy,
i_pipeline__s1_data_t0,
i_pipeline__s1_data,
i_pipeline__s1_error_t0,
i_pipeline__s1_error,
i_pipeline__s1_leak_fence_t0,
i_pipeline__s1_leak_fence,
i_pipeline__s1_rs1_addr_t0,
i_pipeline__s1_rs1_addr,
i_pipeline__s1_rs1_rdata_t0,
i_pipeline__s1_rs1_rdata,
i_pipeline__s1_rs2_addr_t0,
i_pipeline__s1_rs2_addr,
i_pipeline__s1_rs2_rdata_t0,
i_pipeline__s1_rs2_rdata,
i_pipeline__s1_rs3_addr_t0,
i_pipeline__s1_rs3_addr,
i_pipeline__s1_rs3_rdata_t0,
i_pipeline__s1_rs3_rdata,
i_pipeline__s1_valid_t0,
i_pipeline__s1_valid,
i_pipeline__s2_busy_t0,
i_pipeline__s2_busy,
i_pipeline__s2_fu_t0,
i_pipeline__s2_fu,
i_pipeline__s2_instr_t0,
i_pipeline__s2_instr,
i_pipeline__s2_opr_a_t0,
i_pipeline__s2_opr_a,
i_pipeline__s2_opr_b_t0,
i_pipeline__s2_opr_b,
i_pipeline__s2_opr_c_t0,
i_pipeline__s2_opr_c,
i_pipeline__s2_pw_t0,
i_pipeline__s2_pw,
i_pipeline__s2_rd_t0,
i_pipeline__s2_rd,
i_pipeline__s2_size_t0,
i_pipeline__s2_size,
i_pipeline__s2_trap_t0,
i_pipeline__s2_trap,
i_pipeline__s2_uop_t0,
i_pipeline__s2_uop,
i_pipeline__s2_valid_t0,
i_pipeline__s2_valid,
i_pipeline__s3_busy_t0,
i_pipeline__s3_busy,
i_pipeline__s3_fu_t0,
i_pipeline__s3_fu,
i_pipeline__s3_instr_t0,
i_pipeline__s3_instr,
i_pipeline__s3_opr_a_t0,
i_pipeline__s3_opr_a,
i_pipeline__s3_opr_b_t0,
i_pipeline__s3_opr_b,
i_pipeline__s3_rd_t0,
i_pipeline__s3_rd,
i_pipeline__s3_size_t0,
i_pipeline__s3_size,
i_pipeline__s3_trap_t0,
i_pipeline__s3_trap,
i_pipeline__s3_uop_t0,
i_pipeline__s3_uop,
i_pipeline__s3_valid_t0,
i_pipeline__s3_valid,
i_pipeline__s4_busy_t0,
i_pipeline__s4_busy,
i_pipeline__s4_fu_t0,
i_pipeline__s4_fu,
i_pipeline__s4_instr_t0,
i_pipeline__s4_instr,
i_pipeline__s4_opr_a_t0,
i_pipeline__s4_opr_a,
i_pipeline__s4_opr_b_t0,
i_pipeline__s4_opr_b,
i_pipeline__s4_rd_t0,
i_pipeline__s4_rd,
i_pipeline__s4_size_t0,
i_pipeline__s4_size,
i_pipeline__s4_trap_t0,
i_pipeline__s4_trap,
i_pipeline__s4_uop_t0,
i_pipeline__s4_uop,
i_pipeline__s4_valid_t0,
i_pipeline__s4_valid,
i_pipeline__trap_cause_t0,
i_pipeline__trap_cause,
i_pipeline__trap_cpu_t0,
i_pipeline__trap_cpu,
i_pipeline__trap_int_t0,
i_pipeline__trap_int,
i_pipeline__trap_mtval_t0,
i_pipeline__trap_mtval,
i_pipeline__trap_pc_t0,
i_pipeline__trap_pc,
i_pipeline__uxcrypto_b0_t0,
i_pipeline__uxcrypto_b0,
i_pipeline__uxcrypto_b1_t0,
i_pipeline__uxcrypto_b1,
i_pipeline__uxcrypto_ct_t0,
i_pipeline__uxcrypto_ct,
i_pipeline__vector_intrs_t0,
i_pipeline__vector_intrs,
i_pipeline__i_csrs__g_clk,
i_pipeline__i_csrs__g_resetn,
i_pipeline__i_csrs__csr_en,
i_pipeline__i_csrs__csr_wr,
i_pipeline__i_csrs__csr_wr_set,
i_pipeline__i_csrs__csr_wr_clr,
i_pipeline__i_csrs__csr_addr,
i_pipeline__i_csrs__csr_wdata,
i_pipeline__i_csrs__csr_rdata,
i_pipeline__i_csrs__csr_error,
i_pipeline__i_csrs__csr_mepc,
i_pipeline__i_csrs__csr_mtvec,
i_pipeline__i_csrs__vector_intrs,
i_pipeline__i_csrs__exec_mret,
i_pipeline__i_csrs__mstatus_mie,
i_pipeline__i_csrs__mie_meie,
i_pipeline__i_csrs__mie_mtie,
i_pipeline__i_csrs__mie_msie,
i_pipeline__i_csrs__mip_meip,
i_pipeline__i_csrs__mip_mtip,
i_pipeline__i_csrs__mip_msip,
i_pipeline__i_csrs__ctr_time,
i_pipeline__i_csrs__ctr_cycle,
i_pipeline__i_csrs__ctr_instret,
i_pipeline__i_csrs__inhibit_cy,
i_pipeline__i_csrs__inhibit_tm,
i_pipeline__i_csrs__inhibit_ir,
i_pipeline__i_csrs__uxcrypto_ct,
i_pipeline__i_csrs__uxcrypto_b0,
i_pipeline__i_csrs__uxcrypto_b1,
i_pipeline__i_csrs__leak_lkgcfg,
i_pipeline__i_csrs__trap_cpu,
i_pipeline__i_csrs__trap_int,
i_pipeline__i_csrs__trap_cause,
i_pipeline__i_csrs__trap_mtval,
i_pipeline__i_csrs__trap_pc,
i_pipeline__i_csrs__mstatus_mie_t0,
i_pipeline__i_csrs__mip_mtip_t0,
i_pipeline__i_csrs__mie_mtie_t0,
i_pipeline__i_csrs__mie_msie_t0,
i_pipeline__i_csrs__leak_lkgcfg_t0,
i_pipeline__i_csrs__inhibit_tm_t0,
i_pipeline__i_csrs__inhibit_ir_t0,
i_pipeline__i_csrs__inhibit_cy_t0,
i_pipeline__i_csrs__ctr_time_t0,
i_pipeline__i_csrs__ctr_instret_t0,
i_pipeline__i_csrs__ctr_cycle_t0,
i_pipeline__i_csrs__mie_meie_t0,
i_pipeline__i_csrs__mip_msip_t0,
i_pipeline__i_csrs__mip_meip_t0,
i_pipeline__i_csrs__trap_cause_t0,
i_pipeline__i_csrs__uxcrypto_b0_t0,
i_pipeline__i_csrs__uxcrypto_b1_t0,
i_pipeline__i_csrs__uxcrypto_ct_t0,
i_pipeline__i_csrs__csr_addr_t0,
i_pipeline__i_csrs__csr_en_t0,
i_pipeline__i_csrs__csr_error_t0,
i_pipeline__i_csrs__csr_mepc_t0,
i_pipeline__i_csrs__csr_mtvec_t0,
i_pipeline__i_csrs__csr_rdata_t0,
i_pipeline__i_csrs__csr_wdata_t0,
i_pipeline__i_csrs__csr_wr_t0,
i_pipeline__i_csrs__csr_wr_clr_t0,
i_pipeline__i_csrs__csr_wr_set_t0,
i_pipeline__i_csrs__exec_mret_t0,
i_pipeline__i_csrs__trap_cpu_t0,
i_pipeline__i_csrs__trap_int_t0,
i_pipeline__i_csrs__trap_mtval_t0,
i_pipeline__i_csrs__trap_pc_t0,
i_pipeline__i_csrs__vector_intrs_t0,
i_pipeline__i_csrs__int_pulse_t0,
i_pipeline__i_csrs__int_pulse,
i_pipeline__i_csrs__invalid_addr_t0,
i_pipeline__i_csrs__invalid_addr,
i_pipeline__i_csrs__mtvec_bad_write_t0,
i_pipeline__i_csrs__mtvec_bad_write,
i_pipeline__i_csrs__n_mcause_cause_t0,
i_pipeline__i_csrs__n_mcause_cause,
i_pipeline__i_csrs__n_mepc_t0,
i_pipeline__i_csrs__n_mepc,
i_pipeline__i_csrs__n_mstatus_mie_t0,
i_pipeline__i_csrs__n_mstatus_mie,
i_pipeline__i_csrs__n_mstatus_mpie_t0,
i_pipeline__i_csrs__n_mstatus_mpie,
i_pipeline__i_csrs__n_mtvec_base_t0,
i_pipeline__i_csrs__n_mtvec_base,
i_pipeline__i_csrs__n_mtvec_mode_t0,
i_pipeline__i_csrs__n_mtvec_mode,
i_pipeline__i_csrs__n_reg_lkgcfg_t0,
i_pipeline__i_csrs__n_reg_lkgcfg,
i_pipeline__i_csrs__n_reg_mie_t0,
i_pipeline__i_csrs__n_reg_mie,
i_pipeline__i_csrs__n_reg_mscratch_t0,
i_pipeline__i_csrs__n_reg_mscratch,
i_pipeline__i_csrs__n_reg_mtval_t0,
i_pipeline__i_csrs__n_reg_mtval,
i_pipeline__i_csrs__n_uxcrypto_b0_t0,
i_pipeline__i_csrs__n_uxcrypto_b0,
i_pipeline__i_csrs__n_uxcrypto_b1_t0,
i_pipeline__i_csrs__n_uxcrypto_b1,
i_pipeline__i_csrs__n_uxcrypto_ct_t0,
i_pipeline__i_csrs__n_uxcrypto_ct,
i_pipeline__i_csrs__p_trap_int_t0,
i_pipeline__i_csrs__p_trap_int,
i_pipeline__i_csrs__read_cycle_t0,
i_pipeline__i_csrs__read_cycle,
i_pipeline__i_csrs__read_cycleh_t0,
i_pipeline__i_csrs__read_cycleh,
i_pipeline__i_csrs__read_instret_t0,
i_pipeline__i_csrs__read_instret,
i_pipeline__i_csrs__read_instreth_t0,
i_pipeline__i_csrs__read_instreth,
i_pipeline__i_csrs__read_lkgcfg_t0,
i_pipeline__i_csrs__read_lkgcfg,
i_pipeline__i_csrs__read_marchid_t0,
i_pipeline__i_csrs__read_marchid,
i_pipeline__i_csrs__read_mcause_t0,
i_pipeline__i_csrs__read_mcause,
i_pipeline__i_csrs__read_mcountin_t0,
i_pipeline__i_csrs__read_mcountin,
i_pipeline__i_csrs__read_mcycle_t0,
i_pipeline__i_csrs__read_mcycle,
i_pipeline__i_csrs__read_mcycleh_t0,
i_pipeline__i_csrs__read_mcycleh,
i_pipeline__i_csrs__read_medeleg_t0,
i_pipeline__i_csrs__read_medeleg,
i_pipeline__i_csrs__read_mepc_t0,
i_pipeline__i_csrs__read_mepc,
i_pipeline__i_csrs__read_mhartid_t0,
i_pipeline__i_csrs__read_mhartid,
i_pipeline__i_csrs__read_mideleg_t0,
i_pipeline__i_csrs__read_mideleg,
i_pipeline__i_csrs__read_mie_t0,
i_pipeline__i_csrs__read_mie,
i_pipeline__i_csrs__read_mimpid_t0,
i_pipeline__i_csrs__read_mimpid,
i_pipeline__i_csrs__read_minstret_t0,
i_pipeline__i_csrs__read_minstret,
i_pipeline__i_csrs__read_minstreth_t0,
i_pipeline__i_csrs__read_minstreth,
i_pipeline__i_csrs__read_mip_t0,
i_pipeline__i_csrs__read_mip,
i_pipeline__i_csrs__read_misa_t0,
i_pipeline__i_csrs__read_misa,
i_pipeline__i_csrs__read_mscratch_t0,
i_pipeline__i_csrs__read_mscratch,
i_pipeline__i_csrs__read_mstatus_t0,
i_pipeline__i_csrs__read_mstatus,
i_pipeline__i_csrs__read_mtval_t0,
i_pipeline__i_csrs__read_mtval,
i_pipeline__i_csrs__read_mtvec_t0,
i_pipeline__i_csrs__read_mtvec,
i_pipeline__i_csrs__read_mvendorid_t0,
i_pipeline__i_csrs__read_mvendorid,
i_pipeline__i_csrs__read_time_t0,
i_pipeline__i_csrs__read_time,
i_pipeline__i_csrs__read_timeh_t0,
i_pipeline__i_csrs__read_timeh,
i_pipeline__i_csrs__read_uxcrypto_t0,
i_pipeline__i_csrs__read_uxcrypto,
i_pipeline__i_csrs__reg_mcause_cause_t0,
i_pipeline__i_csrs__reg_mcause_cause,
i_pipeline__i_csrs__reg_mcause_interrupt_t0,
i_pipeline__i_csrs__reg_mcause_interrupt,
i_pipeline__i_csrs__reg_mepc_mepc_t0,
i_pipeline__i_csrs__reg_mepc_mepc,
i_pipeline__i_csrs__reg_mscratch_t0,
i_pipeline__i_csrs__reg_mscratch,
i_pipeline__i_csrs__reg_mstatus_mpie_t0,
i_pipeline__i_csrs__reg_mstatus_mpie,
i_pipeline__i_csrs__reg_mstatus_wpri1_t0,
i_pipeline__i_csrs__reg_mstatus_wpri1,
i_pipeline__i_csrs__reg_mstatus_wpri2_t0,
i_pipeline__i_csrs__reg_mstatus_wpri2,
i_pipeline__i_csrs__reg_mstatus_wpri3_t0,
i_pipeline__i_csrs__reg_mstatus_wpri3,
i_pipeline__i_csrs__reg_mstatus_wpri4_t0,
i_pipeline__i_csrs__reg_mstatus_wpri4,
i_pipeline__i_csrs__reg_mtval_t0,
i_pipeline__i_csrs__reg_mtval,
i_pipeline__i_csrs__reg_mtvec_base_t0,
i_pipeline__i_csrs__reg_mtvec_base,
i_pipeline__i_csrs__reg_mtvec_mode_t0,
i_pipeline__i_csrs__reg_mtvec_mode,
i_pipeline__i_csrs__wen_lkgcfg_t0,
i_pipeline__i_csrs__wen_lkgcfg,
i_pipeline__i_csrs__wen_mcause_t0,
i_pipeline__i_csrs__wen_mcause,
i_pipeline__i_csrs__wen_mcountin_t0,
i_pipeline__i_csrs__wen_mcountin,
i_pipeline__i_csrs__wen_mepc_t0,
i_pipeline__i_csrs__wen_mepc,
i_pipeline__i_csrs__wen_mie_t0,
i_pipeline__i_csrs__wen_mie,
i_pipeline__i_csrs__wen_mscratch_t0,
i_pipeline__i_csrs__wen_mscratch,
i_pipeline__i_csrs__wen_mstatus_mie_t0,
i_pipeline__i_csrs__wen_mstatus_mie,
i_pipeline__i_csrs__wen_mstatus_t0,
i_pipeline__i_csrs__wen_mstatus,
i_pipeline__i_csrs__wen_mtval_t0,
i_pipeline__i_csrs__wen_mtval,
i_pipeline__i_csrs__wen_mtvec_t0,
i_pipeline__i_csrs__wen_mtvec,
i_pipeline__i_csrs__wen_uxcrypto_t0,
i_pipeline__i_csrs__wen_uxcrypto,
i_pipeline__i_csrs__wen_valid_mcause_t0,
i_pipeline__i_csrs__wen_valid_mcause,
i_pipeline__i_gprs__g_clk,
i_pipeline__i_gprs__g_resetn,
i_pipeline__i_gprs__rs1_addr,
i_pipeline__i_gprs__rs1_data,
i_pipeline__i_gprs__rs2_addr,
i_pipeline__i_gprs__rs2_data,
i_pipeline__i_gprs__rs3_addr,
i_pipeline__i_gprs__rs3_data,
i_pipeline__i_gprs__rd_wen,
i_pipeline__i_gprs__rd_wide,
i_pipeline__i_gprs__rd_addr,
i_pipeline__i_gprs__rd_wdata,
i_pipeline__i_gprs__rd_wdata_hi,
i_pipeline__i_gprs__rs3_data_t0,
i_pipeline__i_gprs__rs3_addr_t0,
i_pipeline__i_gprs__rs2_data_t0,
i_pipeline__i_gprs__rs2_addr_t0,
i_pipeline__i_gprs__rs1_data_t0,
i_pipeline__i_gprs__rs1_addr_t0,
i_pipeline__i_gprs__rd_wide_t0,
i_pipeline__i_gprs__rd_wen_t0,
i_pipeline__i_gprs__rd_wdata_hi_t0,
i_pipeline__i_gprs__rd_wdata_t0,
i_pipeline__i_gprs__rd_addr_t0,
i_pipeline__i_gprs__gprs_10__t0,
i_pipeline__i_gprs__gprs_10_,
i_pipeline__i_gprs__gprs_11__t0,
i_pipeline__i_gprs__gprs_11_,
i_pipeline__i_gprs__gprs_12__t0,
i_pipeline__i_gprs__gprs_12_,
i_pipeline__i_gprs__gprs_13__t0,
i_pipeline__i_gprs__gprs_13_,
i_pipeline__i_gprs__gprs_14__t0,
i_pipeline__i_gprs__gprs_14_,
i_pipeline__i_gprs__gprs_15__t0,
i_pipeline__i_gprs__gprs_15_,
i_pipeline__i_gprs__gprs_16__t0,
i_pipeline__i_gprs__gprs_16_,
i_pipeline__i_gprs__gprs_17__t0,
i_pipeline__i_gprs__gprs_17_,
i_pipeline__i_gprs__gprs_18__t0,
i_pipeline__i_gprs__gprs_18_,
i_pipeline__i_gprs__gprs_19__t0,
i_pipeline__i_gprs__gprs_19_,
i_pipeline__i_gprs__gprs_1__t0,
i_pipeline__i_gprs__gprs_1_,
i_pipeline__i_gprs__gprs_20__t0,
i_pipeline__i_gprs__gprs_20_,
i_pipeline__i_gprs__gprs_21__t0,
i_pipeline__i_gprs__gprs_21_,
i_pipeline__i_gprs__gprs_22__t0,
i_pipeline__i_gprs__gprs_22_,
i_pipeline__i_gprs__gprs_23__t0,
i_pipeline__i_gprs__gprs_23_,
i_pipeline__i_gprs__gprs_24__t0,
i_pipeline__i_gprs__gprs_24_,
i_pipeline__i_gprs__gprs_25__t0,
i_pipeline__i_gprs__gprs_25_,
i_pipeline__i_gprs__gprs_26__t0,
i_pipeline__i_gprs__gprs_26_,
i_pipeline__i_gprs__gprs_27__t0,
i_pipeline__i_gprs__gprs_27_,
i_pipeline__i_gprs__gprs_28__t0,
i_pipeline__i_gprs__gprs_28_,
i_pipeline__i_gprs__gprs_29__t0,
i_pipeline__i_gprs__gprs_29_,
i_pipeline__i_gprs__gprs_2__t0,
i_pipeline__i_gprs__gprs_2_,
i_pipeline__i_gprs__gprs_30__t0,
i_pipeline__i_gprs__gprs_30_,
i_pipeline__i_gprs__gprs_31__t0,
i_pipeline__i_gprs__gprs_31_,
i_pipeline__i_gprs__gprs_3__t0,
i_pipeline__i_gprs__gprs_3_,
i_pipeline__i_gprs__gprs_4__t0,
i_pipeline__i_gprs__gprs_4_,
i_pipeline__i_gprs__gprs_5__t0,
i_pipeline__i_gprs__gprs_5_,
i_pipeline__i_gprs__gprs_6__t0,
i_pipeline__i_gprs__gprs_6_,
i_pipeline__i_gprs__gprs_7__t0,
i_pipeline__i_gprs__gprs_7_,
i_pipeline__i_gprs__gprs_8__t0,
i_pipeline__i_gprs__gprs_8_,
i_pipeline__i_gprs__gprs_9__t0,
i_pipeline__i_gprs__gprs_9_,
i_pipeline__i_gprs__rd_wdata_odd_t0,
i_pipeline__i_gprs__rd_wdata_odd,
i_pipeline__i_gprs__rd_wen_even_t0,
i_pipeline__i_gprs__rd_wen_even,
i_pipeline__i_gprs__rd_wen_odd_t0,
i_pipeline__i_gprs__rd_wen_odd,
i_pipeline__i_pipeline_s0_fetch__g_clk,
i_pipeline__i_pipeline_s0_fetch__g_resetn,
i_pipeline__i_pipeline_s0_fetch__cf_req,
i_pipeline__i_pipeline_s0_fetch__cf_target,
i_pipeline__i_pipeline_s0_fetch__cf_ack,
i_pipeline__i_pipeline_s0_fetch__imem_req,
i_pipeline__i_pipeline_s0_fetch__imem_wen,
i_pipeline__i_pipeline_s0_fetch__imem_strb,
i_pipeline__i_pipeline_s0_fetch__imem_wdata,
i_pipeline__i_pipeline_s0_fetch__imem_addr,
i_pipeline__i_pipeline_s0_fetch__imem_gnt,
i_pipeline__i_pipeline_s0_fetch__imem_ack,
i_pipeline__i_pipeline_s0_fetch__imem_recv,
i_pipeline__i_pipeline_s0_fetch__imem_error,
i_pipeline__i_pipeline_s0_fetch__imem_rdata,
i_pipeline__i_pipeline_s0_fetch__s0_flush,
i_pipeline__i_pipeline_s0_fetch__s1_busy,
i_pipeline__i_pipeline_s0_fetch__s1_valid,
i_pipeline__i_pipeline_s0_fetch__s1_data,
i_pipeline__i_pipeline_s0_fetch__s1_error,
i_pipeline__i_pipeline_s0_fetch__s1_valid_t0,
i_pipeline__i_pipeline_s0_fetch__s1_error_t0,
i_pipeline__i_pipeline_s0_fetch__s1_data_t0,
i_pipeline__i_pipeline_s0_fetch__s1_busy_t0,
i_pipeline__i_pipeline_s0_fetch__s0_flush_t0,
i_pipeline__i_pipeline_s0_fetch__imem_wen_t0,
i_pipeline__i_pipeline_s0_fetch__imem_wdata_t0,
i_pipeline__i_pipeline_s0_fetch__imem_strb_t0,
i_pipeline__i_pipeline_s0_fetch__imem_req_t0,
i_pipeline__i_pipeline_s0_fetch__imem_recv_t0,
i_pipeline__i_pipeline_s0_fetch__imem_rdata_t0,
i_pipeline__i_pipeline_s0_fetch__imem_gnt_t0,
i_pipeline__i_pipeline_s0_fetch__imem_error_t0,
i_pipeline__i_pipeline_s0_fetch__imem_addr_t0,
i_pipeline__i_pipeline_s0_fetch__imem_ack_t0,
i_pipeline__i_pipeline_s0_fetch__cf_target_t0,
i_pipeline__i_pipeline_s0_fetch__cf_req_t0,
i_pipeline__i_pipeline_s0_fetch__cf_ack_t0,
i_pipeline__i_pipeline_s0_fetch__allow_new_mem_req_t0,
i_pipeline__i_pipeline_s0_fetch__allow_new_mem_req,
i_pipeline__i_pipeline_s0_fetch__buf_16_t0,
i_pipeline__i_pipeline_s0_fetch__buf_16,
i_pipeline__i_pipeline_s0_fetch__buf_32_t0,
i_pipeline__i_pipeline_s0_fetch__buf_32,
i_pipeline__i_pipeline_s0_fetch__buf_depth_t0,
i_pipeline__i_pipeline_s0_fetch__buf_depth,
i_pipeline__i_pipeline_s0_fetch__buf_out_2_t0,
i_pipeline__i_pipeline_s0_fetch__buf_out_2,
i_pipeline__i_pipeline_s0_fetch__buf_out_4_t0,
i_pipeline__i_pipeline_s0_fetch__buf_out_4,
i_pipeline__i_pipeline_s0_fetch__buf_ready_t0,
i_pipeline__i_pipeline_s0_fetch__buf_ready,
i_pipeline__i_pipeline_s0_fetch__cf_change_t0,
i_pipeline__i_pipeline_s0_fetch__cf_change,
i_pipeline__i_pipeline_s0_fetch__drop_response_t0,
i_pipeline__i_pipeline_s0_fetch__drop_response,
i_pipeline__i_pipeline_s0_fetch__f_2byte_t0,
i_pipeline__i_pipeline_s0_fetch__f_2byte,
i_pipeline__i_pipeline_s0_fetch__f_4byte_t0,
i_pipeline__i_pipeline_s0_fetch__f_4byte,
i_pipeline__i_pipeline_s0_fetch__fetch_misaligned_t0,
i_pipeline__i_pipeline_s0_fetch__fetch_misaligned,
i_pipeline__i_pipeline_s0_fetch__ignore_rsps_t0,
i_pipeline__i_pipeline_s0_fetch__ignore_rsps,
i_pipeline__i_pipeline_s0_fetch__incomplete_instr_t0,
i_pipeline__i_pipeline_s0_fetch__incomplete_instr,
i_pipeline__i_pipeline_s0_fetch__n_fetch_misaligned_t0,
i_pipeline__i_pipeline_s0_fetch__n_fetch_misaligned,
i_pipeline__i_pipeline_s0_fetch__n_ignore_rsps_t0,
i_pipeline__i_pipeline_s0_fetch__n_ignore_rsps,
i_pipeline__i_pipeline_s0_fetch__n_imem_addr_t0,
i_pipeline__i_pipeline_s0_fetch__n_imem_addr,
i_pipeline__i_pipeline_s0_fetch__n_imem_req_t0,
i_pipeline__i_pipeline_s0_fetch__n_imem_req,
i_pipeline__i_pipeline_s0_fetch__n_reqs_outstanding_t0,
i_pipeline__i_pipeline_s0_fetch__n_reqs_outstanding,
i_pipeline__i_pipeline_s0_fetch__new_mem_req_t0,
i_pipeline__i_pipeline_s0_fetch__new_mem_req,
i_pipeline__i_pipeline_s0_fetch__progress_imem_addr_t0,
i_pipeline__i_pipeline_s0_fetch__progress_imem_addr,
i_pipeline__i_pipeline_s0_fetch__reqs_outstanding_t0,
i_pipeline__i_pipeline_s0_fetch__reqs_outstanding,
i_pipeline__i_pipeline_s0_fetch__rsp_recv_t0,
i_pipeline__i_pipeline_s0_fetch__rsp_recv,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__g_clk,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__g_resetn,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__flush,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_4byte,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_2byte,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_err,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_in,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_ready,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_depth,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_16,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_32,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out_2,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out_4,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_err,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_valid,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_ready,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_16_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_32_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_depth_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_err_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out_2_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out_4_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_ready_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_valid_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_2byte_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_4byte_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_err_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_in_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_ready_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__flush_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buffer_err_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buffer_err,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buffer_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buffer,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__eat_2_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__eat_2,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__eat_4_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__eat_4,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__insert_at_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__insert_at,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_bdepth_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_bdepth,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_d_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_d,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_err_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_err,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_or_in_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_or_in,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_shf_out_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_shf_out,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_err_in_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_err_in,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_err_or_in_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_err_or_in,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_err_shf_out_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_err_shf_out,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__update_buffer_t0,
i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__update_buffer,
i_pipeline__i_pipeline_s1_decode__g_clk,
i_pipeline__i_pipeline_s1_decode__g_resetn,
i_pipeline__i_pipeline_s1_decode__s1_valid,
i_pipeline__i_pipeline_s1_decode__s1_busy,
i_pipeline__i_pipeline_s1_decode__s1_data,
i_pipeline__i_pipeline_s1_decode__s1_error,
i_pipeline__i_pipeline_s1_decode__s1_flush,
i_pipeline__i_pipeline_s1_decode__s1_bubble,
i_pipeline__i_pipeline_s1_decode__s1_rs1_addr,
i_pipeline__i_pipeline_s1_decode__s1_rs2_addr,
i_pipeline__i_pipeline_s1_decode__s1_rs3_addr,
i_pipeline__i_pipeline_s1_decode__s1_rs1_rdata,
i_pipeline__i_pipeline_s1_decode__s1_rs2_rdata,
i_pipeline__i_pipeline_s1_decode__s1_rs3_rdata,
i_pipeline__i_pipeline_s1_decode__leak_prng,
i_pipeline__i_pipeline_s1_decode__leak_lkgcfg,
i_pipeline__i_pipeline_s1_decode__s1_leak_fence,
i_pipeline__i_pipeline_s1_decode__cf_req,
i_pipeline__i_pipeline_s1_decode__cf_target,
i_pipeline__i_pipeline_s1_decode__cf_ack,
i_pipeline__i_pipeline_s1_decode__s2_valid,
i_pipeline__i_pipeline_s1_decode__s2_busy,
i_pipeline__i_pipeline_s1_decode__s2_rd,
i_pipeline__i_pipeline_s1_decode__s2_opr_a,
i_pipeline__i_pipeline_s1_decode__s2_opr_b,
i_pipeline__i_pipeline_s1_decode__s2_opr_c,
i_pipeline__i_pipeline_s1_decode__s2_uop,
i_pipeline__i_pipeline_s1_decode__s2_fu,
i_pipeline__i_pipeline_s1_decode__s2_pw,
i_pipeline__i_pipeline_s1_decode__s2_trap,
i_pipeline__i_pipeline_s1_decode__s2_size,
i_pipeline__i_pipeline_s1_decode__s2_instr,
i_pipeline__i_pipeline_s1_decode__s2_valid_t0,
i_pipeline__i_pipeline_s1_decode__s2_uop_t0,
i_pipeline__i_pipeline_s1_decode__s2_trap_t0,
i_pipeline__i_pipeline_s1_decode__s2_size_t0,
i_pipeline__i_pipeline_s1_decode__s2_rd_t0,
i_pipeline__i_pipeline_s1_decode__s2_pw_t0,
i_pipeline__i_pipeline_s1_decode__s2_opr_c_t0,
i_pipeline__i_pipeline_s1_decode__s2_opr_b_t0,
i_pipeline__i_pipeline_s1_decode__s2_opr_a_t0,
i_pipeline__i_pipeline_s1_decode__s2_instr_t0,
i_pipeline__i_pipeline_s1_decode__s2_fu_t0,
i_pipeline__i_pipeline_s1_decode__s2_busy_t0,
i_pipeline__i_pipeline_s1_decode__s1_rs3_rdata_t0,
i_pipeline__i_pipeline_s1_decode__s1_rs3_addr_t0,
i_pipeline__i_pipeline_s1_decode__s1_rs2_rdata_t0,
i_pipeline__i_pipeline_s1_decode__s1_rs2_addr_t0,
i_pipeline__i_pipeline_s1_decode__s1_rs1_rdata_t0,
i_pipeline__i_pipeline_s1_decode__s1_rs1_addr_t0,
i_pipeline__i_pipeline_s1_decode__s1_leak_fence_t0,
i_pipeline__i_pipeline_s1_decode__s1_flush_t0,
i_pipeline__i_pipeline_s1_decode__s1_bubble_t0,
i_pipeline__i_pipeline_s1_decode__leak_lkgcfg_t0,
i_pipeline__i_pipeline_s1_decode__leak_prng_t0,
i_pipeline__i_pipeline_s1_decode__s1_valid_t0,
i_pipeline__i_pipeline_s1_decode__s1_error_t0,
i_pipeline__i_pipeline_s1_decode__s1_data_t0,
i_pipeline__i_pipeline_s1_decode__s1_busy_t0,
i_pipeline__i_pipeline_s1_decode__cf_target_t0,
i_pipeline__i_pipeline_s1_decode__cf_req_t0,
i_pipeline__i_pipeline_s1_decode__cf_ack_t0,
i_pipeline__i_pipeline_s1_decode__cfu_no_rd_t0,
i_pipeline__i_pipeline_s1_decode__cfu_no_rd,
i_pipeline__i_pipeline_s1_decode__clr_rd_lsb_t0,
i_pipeline__i_pipeline_s1_decode__clr_rd_lsb,
i_pipeline__i_pipeline_s1_decode__csr_no_read_t0,
i_pipeline__i_pipeline_s1_decode__csr_no_read,
i_pipeline__i_pipeline_s1_decode__csr_no_write_t0,
i_pipeline__i_pipeline_s1_decode__csr_no_write,
i_pipeline__i_pipeline_s1_decode__csr_op_t0,
i_pipeline__i_pipeline_s1_decode__csr_op,
i_pipeline__i_pipeline_s1_decode__dec_add_t0,
i_pipeline__i_pipeline_s1_decode__dec_add,
i_pipeline__i_pipeline_s1_decode__dec_addi_t0,
i_pipeline__i_pipeline_s1_decode__dec_addi,
i_pipeline__i_pipeline_s1_decode__dec_and_t0,
i_pipeline__i_pipeline_s1_decode__dec_and,
i_pipeline__i_pipeline_s1_decode__dec_andi_t0,
i_pipeline__i_pipeline_s1_decode__dec_andi,
i_pipeline__i_pipeline_s1_decode__dec_auipc_t0,
i_pipeline__i_pipeline_s1_decode__dec_auipc,
i_pipeline__i_pipeline_s1_decode__dec_b_bdep_t0,
i_pipeline__i_pipeline_s1_decode__dec_b_bdep,
i_pipeline__i_pipeline_s1_decode__dec_b_bext_t0,
i_pipeline__i_pipeline_s1_decode__dec_b_bext,
i_pipeline__i_pipeline_s1_decode__dec_b_clmul_t0,
i_pipeline__i_pipeline_s1_decode__dec_b_clmul,
i_pipeline__i_pipeline_s1_decode__dec_b_clmulh_t0,
i_pipeline__i_pipeline_s1_decode__dec_b_clmulh,
i_pipeline__i_pipeline_s1_decode__dec_b_clmulr_t0,
i_pipeline__i_pipeline_s1_decode__dec_b_clmulr,
i_pipeline__i_pipeline_s1_decode__dec_b_cmov_t0,
i_pipeline__i_pipeline_s1_decode__dec_b_cmov,
i_pipeline__i_pipeline_s1_decode__dec_b_fsl_t0,
i_pipeline__i_pipeline_s1_decode__dec_b_fsl,
i_pipeline__i_pipeline_s1_decode__dec_b_fsr_t0,
i_pipeline__i_pipeline_s1_decode__dec_b_fsr,
i_pipeline__i_pipeline_s1_decode__dec_b_fsri_t0,
i_pipeline__i_pipeline_s1_decode__dec_b_fsri,
i_pipeline__i_pipeline_s1_decode__dec_b_grev_t0,
i_pipeline__i_pipeline_s1_decode__dec_b_grev,
i_pipeline__i_pipeline_s1_decode__dec_b_grevi_t0,
i_pipeline__i_pipeline_s1_decode__dec_b_grevi,
i_pipeline__i_pipeline_s1_decode__dec_b_ror_t0,
i_pipeline__i_pipeline_s1_decode__dec_b_ror,
i_pipeline__i_pipeline_s1_decode__dec_b_rori_t0,
i_pipeline__i_pipeline_s1_decode__dec_b_rori,
i_pipeline__i_pipeline_s1_decode__dec_beq_t0,
i_pipeline__i_pipeline_s1_decode__dec_beq,
i_pipeline__i_pipeline_s1_decode__dec_bge_t0,
i_pipeline__i_pipeline_s1_decode__dec_bge,
i_pipeline__i_pipeline_s1_decode__dec_bgeu_t0,
i_pipeline__i_pipeline_s1_decode__dec_bgeu,
i_pipeline__i_pipeline_s1_decode__dec_blt_t0,
i_pipeline__i_pipeline_s1_decode__dec_blt,
i_pipeline__i_pipeline_s1_decode__dec_bltu_t0,
i_pipeline__i_pipeline_s1_decode__dec_bltu,
i_pipeline__i_pipeline_s1_decode__dec_bne_t0,
i_pipeline__i_pipeline_s1_decode__dec_bne,
i_pipeline__i_pipeline_s1_decode__dec_c_add_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_add,
i_pipeline__i_pipeline_s1_decode__dec_c_addi16sp_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_addi16sp,
i_pipeline__i_pipeline_s1_decode__dec_c_addi4spn_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_addi4spn,
i_pipeline__i_pipeline_s1_decode__dec_c_addi_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_addi,
i_pipeline__i_pipeline_s1_decode__dec_c_and_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_and,
i_pipeline__i_pipeline_s1_decode__dec_c_andi_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_andi,
i_pipeline__i_pipeline_s1_decode__dec_c_beqz_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_beqz,
i_pipeline__i_pipeline_s1_decode__dec_c_bnez_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_bnez,
i_pipeline__i_pipeline_s1_decode__dec_c_ebreak_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_ebreak,
i_pipeline__i_pipeline_s1_decode__dec_c_j_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_j,
i_pipeline__i_pipeline_s1_decode__dec_c_jal_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_jal,
i_pipeline__i_pipeline_s1_decode__dec_c_jalr_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_jalr,
i_pipeline__i_pipeline_s1_decode__dec_c_jr_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_jr,
i_pipeline__i_pipeline_s1_decode__dec_c_li_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_li,
i_pipeline__i_pipeline_s1_decode__dec_c_lui_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_lui,
i_pipeline__i_pipeline_s1_decode__dec_c_lw_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_lw,
i_pipeline__i_pipeline_s1_decode__dec_c_lwsp_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_lwsp,
i_pipeline__i_pipeline_s1_decode__dec_c_mv_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_mv,
i_pipeline__i_pipeline_s1_decode__dec_c_nop_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_nop,
i_pipeline__i_pipeline_s1_decode__dec_c_or_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_or,
i_pipeline__i_pipeline_s1_decode__dec_c_slli_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_slli,
i_pipeline__i_pipeline_s1_decode__dec_c_srai_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_srai,
i_pipeline__i_pipeline_s1_decode__dec_c_srli_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_srli,
i_pipeline__i_pipeline_s1_decode__dec_c_sub_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_sub,
i_pipeline__i_pipeline_s1_decode__dec_c_sw_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_sw,
i_pipeline__i_pipeline_s1_decode__dec_c_swsp_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_swsp,
i_pipeline__i_pipeline_s1_decode__dec_c_xor_t0,
i_pipeline__i_pipeline_s1_decode__dec_c_xor,
i_pipeline__i_pipeline_s1_decode__dec_csrrc_t0,
i_pipeline__i_pipeline_s1_decode__dec_csrrc,
i_pipeline__i_pipeline_s1_decode__dec_csrrci_t0,
i_pipeline__i_pipeline_s1_decode__dec_csrrci,
i_pipeline__i_pipeline_s1_decode__dec_csrrs_t0,
i_pipeline__i_pipeline_s1_decode__dec_csrrs,
i_pipeline__i_pipeline_s1_decode__dec_csrrsi_t0,
i_pipeline__i_pipeline_s1_decode__dec_csrrsi,
i_pipeline__i_pipeline_s1_decode__dec_csrrw_t0,
i_pipeline__i_pipeline_s1_decode__dec_csrrw,
i_pipeline__i_pipeline_s1_decode__dec_csrrwi_t0,
i_pipeline__i_pipeline_s1_decode__dec_csrrwi,
i_pipeline__i_pipeline_s1_decode__dec_div_t0,
i_pipeline__i_pipeline_s1_decode__dec_div,
i_pipeline__i_pipeline_s1_decode__dec_divu_t0,
i_pipeline__i_pipeline_s1_decode__dec_divu,
i_pipeline__i_pipeline_s1_decode__dec_ebreak_t0,
i_pipeline__i_pipeline_s1_decode__dec_ebreak,
i_pipeline__i_pipeline_s1_decode__dec_ecall_t0,
i_pipeline__i_pipeline_s1_decode__dec_ecall,
i_pipeline__i_pipeline_s1_decode__dec_fence_i_t0,
i_pipeline__i_pipeline_s1_decode__dec_fence_i,
i_pipeline__i_pipeline_s1_decode__dec_fence_t0,
i_pipeline__i_pipeline_s1_decode__dec_fence,
i_pipeline__i_pipeline_s1_decode__dec_jal_t0,
i_pipeline__i_pipeline_s1_decode__dec_jal,
i_pipeline__i_pipeline_s1_decode__dec_jalr_t0,
i_pipeline__i_pipeline_s1_decode__dec_jalr,
i_pipeline__i_pipeline_s1_decode__dec_lb_t0,
i_pipeline__i_pipeline_s1_decode__dec_lb,
i_pipeline__i_pipeline_s1_decode__dec_lbu_t0,
i_pipeline__i_pipeline_s1_decode__dec_lbu,
i_pipeline__i_pipeline_s1_decode__dec_lh_t0,
i_pipeline__i_pipeline_s1_decode__dec_lh,
i_pipeline__i_pipeline_s1_decode__dec_lhu_t0,
i_pipeline__i_pipeline_s1_decode__dec_lhu,
i_pipeline__i_pipeline_s1_decode__dec_lui_t0,
i_pipeline__i_pipeline_s1_decode__dec_lui,
i_pipeline__i_pipeline_s1_decode__dec_lw_t0,
i_pipeline__i_pipeline_s1_decode__dec_lw,
i_pipeline__i_pipeline_s1_decode__dec_mret_t0,
i_pipeline__i_pipeline_s1_decode__dec_mret,
i_pipeline__i_pipeline_s1_decode__dec_mul_t0,
i_pipeline__i_pipeline_s1_decode__dec_mul,
i_pipeline__i_pipeline_s1_decode__dec_mulh_t0,
i_pipeline__i_pipeline_s1_decode__dec_mulh,
i_pipeline__i_pipeline_s1_decode__dec_mulhsu_t0,
i_pipeline__i_pipeline_s1_decode__dec_mulhsu,
i_pipeline__i_pipeline_s1_decode__dec_mulhu_t0,
i_pipeline__i_pipeline_s1_decode__dec_mulhu,
i_pipeline__i_pipeline_s1_decode__dec_or_t0,
i_pipeline__i_pipeline_s1_decode__dec_or,
i_pipeline__i_pipeline_s1_decode__dec_ori_t0,
i_pipeline__i_pipeline_s1_decode__dec_ori,
i_pipeline__i_pipeline_s1_decode__dec_rd_16_t0,
i_pipeline__i_pipeline_s1_decode__dec_rd_16,
i_pipeline__i_pipeline_s1_decode__dec_rd_32_t0,
i_pipeline__i_pipeline_s1_decode__dec_rd_32,
i_pipeline__i_pipeline_s1_decode__dec_rem_t0,
i_pipeline__i_pipeline_s1_decode__dec_rem,
i_pipeline__i_pipeline_s1_decode__dec_remu_t0,
i_pipeline__i_pipeline_s1_decode__dec_remu,
i_pipeline__i_pipeline_s1_decode__dec_rs1_16_t0,
i_pipeline__i_pipeline_s1_decode__dec_rs1_16,
i_pipeline__i_pipeline_s1_decode__dec_rs2_16_t0,
i_pipeline__i_pipeline_s1_decode__dec_rs2_16,
i_pipeline__i_pipeline_s1_decode__dec_sb_t0,
i_pipeline__i_pipeline_s1_decode__dec_sb,
i_pipeline__i_pipeline_s1_decode__dec_sh_t0,
i_pipeline__i_pipeline_s1_decode__dec_sh,
i_pipeline__i_pipeline_s1_decode__dec_sll_t0,
i_pipeline__i_pipeline_s1_decode__dec_sll,
i_pipeline__i_pipeline_s1_decode__dec_slli_t0,
i_pipeline__i_pipeline_s1_decode__dec_slli,
i_pipeline__i_pipeline_s1_decode__dec_slt_t0,
i_pipeline__i_pipeline_s1_decode__dec_slt,
i_pipeline__i_pipeline_s1_decode__dec_slti_t0,
i_pipeline__i_pipeline_s1_decode__dec_slti,
i_pipeline__i_pipeline_s1_decode__dec_sltiu_t0,
i_pipeline__i_pipeline_s1_decode__dec_sltiu,
i_pipeline__i_pipeline_s1_decode__dec_sltu_t0,
i_pipeline__i_pipeline_s1_decode__dec_sltu,
i_pipeline__i_pipeline_s1_decode__dec_sra_t0,
i_pipeline__i_pipeline_s1_decode__dec_sra,
i_pipeline__i_pipeline_s1_decode__dec_srai_t0,
i_pipeline__i_pipeline_s1_decode__dec_srai,
i_pipeline__i_pipeline_s1_decode__dec_srl_t0,
i_pipeline__i_pipeline_s1_decode__dec_srl,
i_pipeline__i_pipeline_s1_decode__dec_srli_t0,
i_pipeline__i_pipeline_s1_decode__dec_srli,
i_pipeline__i_pipeline_s1_decode__dec_sub_t0,
i_pipeline__i_pipeline_s1_decode__dec_sub,
i_pipeline__i_pipeline_s1_decode__dec_sw_t0,
i_pipeline__i_pipeline_s1_decode__dec_sw,
i_pipeline__i_pipeline_s1_decode__dec_wfi_t0,
i_pipeline__i_pipeline_s1_decode__dec_wfi,
i_pipeline__i_pipeline_s1_decode__dec_xc_aesmix_dec_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_aesmix_dec,
i_pipeline__i_pipeline_s1_decode__dec_xc_aesmix_enc_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_aesmix_enc,
i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_dec_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_dec,
i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_decrot_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_decrot,
i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_enc_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_enc,
i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_encrot_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_encrot,
i_pipeline__i_pipeline_s1_decode__dec_xc_bop_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_bop,
i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_b_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_b,
i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_bu_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_bu,
i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_h_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_h,
i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_hu_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_hu,
i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_w_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_w,
i_pipeline__i_pipeline_s1_decode__dec_xc_lkgfence_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_lkgfence,
i_pipeline__i_pipeline_s1_decode__dec_xc_lut_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_lut,
i_pipeline__i_pipeline_s1_decode__dec_xc_macc_1_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_macc_1,
i_pipeline__i_pipeline_s1_decode__dec_xc_madd_3_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_madd_3,
i_pipeline__i_pipeline_s1_decode__dec_xc_mmul_3_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_mmul_3,
i_pipeline__i_pipeline_s1_decode__dec_xc_mror_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_mror,
i_pipeline__i_pipeline_s1_decode__dec_xc_msub_3_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_msub_3,
i_pipeline__i_pipeline_s1_decode__dec_xc_padd_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_padd,
i_pipeline__i_pipeline_s1_decode__dec_xc_pclmul_h_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_pclmul_h,
i_pipeline__i_pipeline_s1_decode__dec_xc_pclmul_l_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_pclmul_l,
i_pipeline__i_pipeline_s1_decode__dec_xc_pmul_h_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_pmul_h,
i_pipeline__i_pipeline_s1_decode__dec_xc_pmul_l_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_pmul_l,
i_pipeline__i_pipeline_s1_decode__dec_xc_pror_i_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_pror_i,
i_pipeline__i_pipeline_s1_decode__dec_xc_pror_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_pror,
i_pipeline__i_pipeline_s1_decode__dec_xc_psll_i_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_psll_i,
i_pipeline__i_pipeline_s1_decode__dec_xc_psll_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_psll,
i_pipeline__i_pipeline_s1_decode__dec_xc_psrl_i_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_psrl_i,
i_pipeline__i_pipeline_s1_decode__dec_xc_psrl_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_psrl,
i_pipeline__i_pipeline_s1_decode__dec_xc_psub_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_psub,
i_pipeline__i_pipeline_s1_decode__dec_xc_rngsamp_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_rngsamp,
i_pipeline__i_pipeline_s1_decode__dec_xc_rngseed_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_rngseed,
i_pipeline__i_pipeline_s1_decode__dec_xc_rngtest_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_rngtest,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s0_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s0,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s1_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s1,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s2_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s2,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s3_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s3,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_x1_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_x1,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_x2_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_x2,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_x4_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_x4,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_xy_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_xy,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_yx_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_yx,
i_pipeline__i_pipeline_s1_decode__dec_xc_str_b_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_str_b,
i_pipeline__i_pipeline_s1_decode__dec_xc_str_h_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_str_h,
i_pipeline__i_pipeline_s1_decode__dec_xc_str_w_t0,
i_pipeline__i_pipeline_s1_decode__dec_xc_str_w,
i_pipeline__i_pipeline_s1_decode__dec_xor_t0,
i_pipeline__i_pipeline_s1_decode__dec_xor,
i_pipeline__i_pipeline_s1_decode__dec_xori_t0,
i_pipeline__i_pipeline_s1_decode__dec_xori,
i_pipeline__i_pipeline_s1_decode__instr_16bit_t0,
i_pipeline__i_pipeline_s1_decode__instr_16bit,
i_pipeline__i_pipeline_s1_decode__invalid_instr_t0,
i_pipeline__i_pipeline_s1_decode__invalid_instr,
i_pipeline__i_pipeline_s1_decode__leak_stall_t0,
i_pipeline__i_pipeline_s1_decode__leak_stall,
i_pipeline__i_pipeline_s1_decode__lf_count_ld_t0,
i_pipeline__i_pipeline_s1_decode__lf_count_ld,
i_pipeline__i_pipeline_s1_decode__lf_count_t0,
i_pipeline__i_pipeline_s1_decode__lf_count,
i_pipeline__i_pipeline_s1_decode__lsu_no_rd_t0,
i_pipeline__i_pipeline_s1_decode__lsu_no_rd,
i_pipeline__i_pipeline_s1_decode__lsu_width_t0,
i_pipeline__i_pipeline_s1_decode__lsu_width,
i_pipeline__i_pipeline_s1_decode__n_lf_count_t0,
i_pipeline__i_pipeline_s1_decode__n_lf_count,
i_pipeline__i_pipeline_s1_decode__n_program_counter_t0,
i_pipeline__i_pipeline_s1_decode__n_program_counter,
i_pipeline__i_pipeline_s1_decode__n_s2_fu_t0,
i_pipeline__i_pipeline_s1_decode__n_s2_fu,
i_pipeline__i_pipeline_s1_decode__n_s2_imm_pc_t0,
i_pipeline__i_pipeline_s1_decode__n_s2_imm_pc,
i_pipeline__i_pipeline_s1_decode__n_s2_imm_t0,
i_pipeline__i_pipeline_s1_decode__n_s2_imm,
i_pipeline__i_pipeline_s1_decode__n_s2_instr_t0,
i_pipeline__i_pipeline_s1_decode__n_s2_instr,
i_pipeline__i_pipeline_s1_decode__n_s2_opr_a_t0,
i_pipeline__i_pipeline_s1_decode__n_s2_opr_a,
i_pipeline__i_pipeline_s1_decode__n_s2_opr_b_t0,
i_pipeline__i_pipeline_s1_decode__n_s2_opr_b,
i_pipeline__i_pipeline_s1_decode__n_s2_opr_c_t0,
i_pipeline__i_pipeline_s1_decode__n_s2_opr_c,
i_pipeline__i_pipeline_s1_decode__n_s2_pw_t0,
i_pipeline__i_pipeline_s1_decode__n_s2_pw,
i_pipeline__i_pipeline_s1_decode__n_s2_rd_t0,
i_pipeline__i_pipeline_s1_decode__n_s2_rd,
i_pipeline__i_pipeline_s1_decode__n_s2_trap_t0,
i_pipeline__i_pipeline_s1_decode__n_s2_trap,
i_pipeline__i_pipeline_s1_decode__n_s2_uop_t0,
i_pipeline__i_pipeline_s1_decode__n_s2_uop,
i_pipeline__i_pipeline_s1_decode__n_s2_valid_t0,
i_pipeline__i_pipeline_s1_decode__n_s2_valid,
i_pipeline__i_pipeline_s1_decode__opra_flush_t0,
i_pipeline__i_pipeline_s1_decode__opra_flush,
i_pipeline__i_pipeline_s1_decode__opra_ld_en_t0,
i_pipeline__i_pipeline_s1_decode__opra_ld_en,
i_pipeline__i_pipeline_s1_decode__opra_src_csri_t0,
i_pipeline__i_pipeline_s1_decode__opra_src_csri,
i_pipeline__i_pipeline_s1_decode__opra_src_rs1_t0,
i_pipeline__i_pipeline_s1_decode__opra_src_rs1,
i_pipeline__i_pipeline_s1_decode__opra_src_zero_t0,
i_pipeline__i_pipeline_s1_decode__opra_src_zero,
i_pipeline__i_pipeline_s1_decode__oprb_flush_t0,
i_pipeline__i_pipeline_s1_decode__oprb_flush,
i_pipeline__i_pipeline_s1_decode__oprb_ld_en_t0,
i_pipeline__i_pipeline_s1_decode__oprb_ld_en,
i_pipeline__i_pipeline_s1_decode__oprb_rs2_shf_1_t0,
i_pipeline__i_pipeline_s1_decode__oprb_rs2_shf_1,
i_pipeline__i_pipeline_s1_decode__oprb_rs2_shf_2_t0,
i_pipeline__i_pipeline_s1_decode__oprb_rs2_shf_2,
i_pipeline__i_pipeline_s1_decode__oprb_src_imm_t0,
i_pipeline__i_pipeline_s1_decode__oprb_src_imm,
i_pipeline__i_pipeline_s1_decode__oprb_src_rs2_t0,
i_pipeline__i_pipeline_s1_decode__oprb_src_rs2,
i_pipeline__i_pipeline_s1_decode__oprb_src_zero_t0,
i_pipeline__i_pipeline_s1_decode__oprb_src_zero,
i_pipeline__i_pipeline_s1_decode__oprc_flush_t0,
i_pipeline__i_pipeline_s1_decode__oprc_flush,
i_pipeline__i_pipeline_s1_decode__oprc_ld_en_t0,
i_pipeline__i_pipeline_s1_decode__oprc_ld_en,
i_pipeline__i_pipeline_s1_decode__oprc_src_pcim_t0,
i_pipeline__i_pipeline_s1_decode__oprc_src_pcim,
i_pipeline__i_pipeline_s1_decode__oprc_src_rs2_t0,
i_pipeline__i_pipeline_s1_decode__oprc_src_rs2,
i_pipeline__i_pipeline_s1_decode__oprc_src_rs3_t0,
i_pipeline__i_pipeline_s1_decode__oprc_src_rs3,
i_pipeline__i_pipeline_s1_decode__p_in_t0,
i_pipeline__i_pipeline_s1_decode__p_in,
i_pipeline__i_pipeline_s1_decode__p_mr_t0,
i_pipeline__i_pipeline_s1_decode__p_mr,
i_pipeline__i_pipeline_s1_decode__p_out_t0,
i_pipeline__i_pipeline_s1_decode__p_out,
i_pipeline__i_pipeline_s1_decode__p_s2_busy_t0,
i_pipeline__i_pipeline_s1_decode__p_s2_busy,
i_pipeline__i_pipeline_s1_decode__packed_instruction_t0,
i_pipeline__i_pipeline_s1_decode__packed_instruction,
i_pipeline__i_pipeline_s1_decode__pc_plus_imm_t0,
i_pipeline__i_pipeline_s1_decode__pc_plus_imm,
i_pipeline__i_pipeline_s1_decode__pipe_progress_t0,
i_pipeline__i_pipeline_s1_decode__pipe_progress,
i_pipeline__i_pipeline_s1_decode__program_counter_t0,
i_pipeline__i_pipeline_s1_decode__program_counter,
i_pipeline__i_pipeline_s1_decode__s1_rs2_shf_t0,
i_pipeline__i_pipeline_s1_decode__s1_rs2_shf,
i_pipeline__i_pipeline_s1_decode__trap_cause_t0,
i_pipeline__i_pipeline_s1_decode__trap_cause,
i_pipeline__i_pipeline_s1_decode__uop_alu_t0,
i_pipeline__i_pipeline_s1_decode__uop_alu,
i_pipeline__i_pipeline_s1_decode__uop_asi_t0,
i_pipeline__i_pipeline_s1_decode__uop_asi,
i_pipeline__i_pipeline_s1_decode__uop_bit_t0,
i_pipeline__i_pipeline_s1_decode__uop_bit,
i_pipeline__i_pipeline_s1_decode__uop_cfu_t0,
i_pipeline__i_pipeline_s1_decode__uop_cfu,
i_pipeline__i_pipeline_s1_decode__uop_csr_t0,
i_pipeline__i_pipeline_s1_decode__uop_csr,
i_pipeline__i_pipeline_s1_decode__uop_lsu_t0,
i_pipeline__i_pipeline_s1_decode__uop_lsu,
i_pipeline__i_pipeline_s1_decode__uop_mul_t0,
i_pipeline__i_pipeline_s1_decode__uop_mul,
i_pipeline__i_pipeline_s1_decode__uop_rng_t0,
i_pipeline__i_pipeline_s1_decode__uop_rng,
i_pipeline__i_pipeline_s1_decode__use_imm32_b_t0,
i_pipeline__i_pipeline_s1_decode__use_imm32_b,
i_pipeline__i_pipeline_s1_decode__use_imm32_i_t0,
i_pipeline__i_pipeline_s1_decode__use_imm32_i,
i_pipeline__i_pipeline_s1_decode__use_imm32_s_t0,
i_pipeline__i_pipeline_s1_decode__use_imm32_s,
i_pipeline__i_pipeline_s1_decode__use_imm32_u_t0,
i_pipeline__i_pipeline_s1_decode__use_imm32_u,
i_pipeline__i_pipeline_s1_decode__use_imm_csr_t0,
i_pipeline__i_pipeline_s1_decode__use_imm_csr,
i_pipeline__i_pipeline_s1_decode__use_imm_sha3_t0,
i_pipeline__i_pipeline_s1_decode__use_imm_sha3,
i_pipeline__i_pipeline_s1_decode__use_imm_shfi_t0,
i_pipeline__i_pipeline_s1_decode__use_imm_shfi,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__g_clk,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__g_resetn,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_data,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_valid,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_busy,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__mr_data,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__flush,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__flush_dat,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_data,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_valid,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_busy,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__flush_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_valid_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_data_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_busy_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__mr_data_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_valid_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_data_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_busy_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__flush_dat_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__genblk1__progress_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__genblk1__progress,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__g_clk,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__g_resetn,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_data,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_valid,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_busy,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__mr_data,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__flush,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__flush_dat,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_data,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_valid,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_busy,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__flush_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_valid_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_data_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_busy_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__mr_data_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_valid_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_data_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_busy_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__flush_dat_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__genblk1__progress_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__genblk1__progress,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__g_clk,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__g_resetn,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_data,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_valid,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_busy,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__mr_data,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__flush,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__flush_dat,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_data,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_valid,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_busy,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__flush_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_valid_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_data_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_busy_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__mr_data_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_valid_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_data_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_busy_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__flush_dat_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__genblk1__progress_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__genblk1__progress,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__g_clk,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__g_resetn,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_data,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_valid,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_busy,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__mr_data,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__flush,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__flush_dat,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_data,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_valid,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_busy,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__flush_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_valid_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_data_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_busy_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__mr_data_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_valid_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_data_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_busy_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__flush_dat_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__genblk1__progress_t0,
i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__genblk1__progress,
i_pipeline__i_pipeline_s1_decode__i_frv_leak__g_clk,
i_pipeline__i_pipeline_s1_decode__i_frv_leak__g_resetn,
i_pipeline__i_pipeline_s1_decode__i_frv_leak__leak_prng,
i_pipeline__i_pipeline_s1_decode__i_frv_leak__leak_fence,
i_pipeline__i_pipeline_s1_decode__i_frv_leak__leak_prng_t0,
i_pipeline__i_pipeline_s1_decode__i_frv_leak__leak_fence_t0,
i_pipeline__i_pipeline_s1_decode__i_frv_leak__genblk1__genblk1__n_prng_lsb_t0,
i_pipeline__i_pipeline_s1_decode__i_frv_leak__genblk1__genblk1__n_prng_lsb,
i_pipeline__i_pipeline_s2_execute__g_clk,
i_pipeline__i_pipeline_s2_execute__g_resetn,
i_pipeline__i_pipeline_s2_execute__s2_rd,
i_pipeline__i_pipeline_s2_execute__s2_opr_a,
i_pipeline__i_pipeline_s2_execute__s2_opr_b,
i_pipeline__i_pipeline_s2_execute__s2_opr_c,
i_pipeline__i_pipeline_s2_execute__s2_uop,
i_pipeline__i_pipeline_s2_execute__s2_fu,
i_pipeline__i_pipeline_s2_execute__s2_pw,
i_pipeline__i_pipeline_s2_execute__s2_trap,
i_pipeline__i_pipeline_s2_execute__s2_size,
i_pipeline__i_pipeline_s2_execute__s2_instr,
i_pipeline__i_pipeline_s2_execute__s2_busy,
i_pipeline__i_pipeline_s2_execute__s2_valid,
i_pipeline__i_pipeline_s2_execute__leak_prng,
i_pipeline__i_pipeline_s2_execute__leak_lkgcfg,
i_pipeline__i_pipeline_s2_execute__rng_req_valid,
i_pipeline__i_pipeline_s2_execute__rng_req_op,
i_pipeline__i_pipeline_s2_execute__rng_req_data,
i_pipeline__i_pipeline_s2_execute__rng_req_ready,
i_pipeline__i_pipeline_s2_execute__rng_rsp_valid,
i_pipeline__i_pipeline_s2_execute__rng_rsp_status,
i_pipeline__i_pipeline_s2_execute__rng_rsp_data,
i_pipeline__i_pipeline_s2_execute__rng_rsp_ready,
i_pipeline__i_pipeline_s2_execute__uxcrypto_ct,
i_pipeline__i_pipeline_s2_execute__uxcrypto_b0,
i_pipeline__i_pipeline_s2_execute__uxcrypto_b1,
i_pipeline__i_pipeline_s2_execute__flush,
i_pipeline__i_pipeline_s2_execute__fwd_s2_rd,
i_pipeline__i_pipeline_s2_execute__fwd_s2_wide,
i_pipeline__i_pipeline_s2_execute__fwd_s2_wdata,
i_pipeline__i_pipeline_s2_execute__fwd_s2_wdata_hi,
i_pipeline__i_pipeline_s2_execute__fwd_s2_load,
i_pipeline__i_pipeline_s2_execute__fwd_s2_csr,
i_pipeline__i_pipeline_s2_execute__s3_rd,
i_pipeline__i_pipeline_s2_execute__s3_opr_a,
i_pipeline__i_pipeline_s2_execute__s3_opr_b,
i_pipeline__i_pipeline_s2_execute__s3_uop,
i_pipeline__i_pipeline_s2_execute__s3_fu,
i_pipeline__i_pipeline_s2_execute__s3_trap,
i_pipeline__i_pipeline_s2_execute__s3_size,
i_pipeline__i_pipeline_s2_execute__s3_instr,
i_pipeline__i_pipeline_s2_execute__s3_busy,
i_pipeline__i_pipeline_s2_execute__s3_valid,
i_pipeline__i_pipeline_s2_execute__flush_t0,
i_pipeline__i_pipeline_s2_execute__s2_valid_t0,
i_pipeline__i_pipeline_s2_execute__s2_uop_t0,
i_pipeline__i_pipeline_s2_execute__s2_trap_t0,
i_pipeline__i_pipeline_s2_execute__s2_size_t0,
i_pipeline__i_pipeline_s2_execute__s2_rd_t0,
i_pipeline__i_pipeline_s2_execute__s2_pw_t0,
i_pipeline__i_pipeline_s2_execute__s2_opr_c_t0,
i_pipeline__i_pipeline_s2_execute__s2_opr_b_t0,
i_pipeline__i_pipeline_s2_execute__s2_opr_a_t0,
i_pipeline__i_pipeline_s2_execute__s2_instr_t0,
i_pipeline__i_pipeline_s2_execute__s2_fu_t0,
i_pipeline__i_pipeline_s2_execute__s2_busy_t0,
i_pipeline__i_pipeline_s2_execute__leak_lkgcfg_t0,
i_pipeline__i_pipeline_s2_execute__leak_prng_t0,
i_pipeline__i_pipeline_s2_execute__rng_req_data_t0,
i_pipeline__i_pipeline_s2_execute__rng_req_op_t0,
i_pipeline__i_pipeline_s2_execute__rng_req_ready_t0,
i_pipeline__i_pipeline_s2_execute__rng_req_valid_t0,
i_pipeline__i_pipeline_s2_execute__rng_rsp_data_t0,
i_pipeline__i_pipeline_s2_execute__rng_rsp_ready_t0,
i_pipeline__i_pipeline_s2_execute__rng_rsp_status_t0,
i_pipeline__i_pipeline_s2_execute__rng_rsp_valid_t0,
i_pipeline__i_pipeline_s2_execute__fwd_s2_csr_t0,
i_pipeline__i_pipeline_s2_execute__fwd_s2_load_t0,
i_pipeline__i_pipeline_s2_execute__fwd_s2_rd_t0,
i_pipeline__i_pipeline_s2_execute__fwd_s2_wdata_t0,
i_pipeline__i_pipeline_s2_execute__fwd_s2_wdata_hi_t0,
i_pipeline__i_pipeline_s2_execute__fwd_s2_wide_t0,
i_pipeline__i_pipeline_s2_execute__s3_busy_t0,
i_pipeline__i_pipeline_s2_execute__s3_fu_t0,
i_pipeline__i_pipeline_s2_execute__s3_instr_t0,
i_pipeline__i_pipeline_s2_execute__s3_opr_a_t0,
i_pipeline__i_pipeline_s2_execute__s3_opr_b_t0,
i_pipeline__i_pipeline_s2_execute__s3_rd_t0,
i_pipeline__i_pipeline_s2_execute__s3_size_t0,
i_pipeline__i_pipeline_s2_execute__s3_trap_t0,
i_pipeline__i_pipeline_s2_execute__s3_uop_t0,
i_pipeline__i_pipeline_s2_execute__s3_valid_t0,
i_pipeline__i_pipeline_s2_execute__uxcrypto_b0_t0,
i_pipeline__i_pipeline_s2_execute__uxcrypto_b1_t0,
i_pipeline__i_pipeline_s2_execute__uxcrypto_ct_t0,
i_pipeline__i_pipeline_s2_execute__alu_add_result_t0,
i_pipeline__i_pipeline_s2_execute__alu_add_result,
i_pipeline__i_pipeline_s2_execute__alu_eq_t0,
i_pipeline__i_pipeline_s2_execute__alu_eq,
i_pipeline__i_pipeline_s2_execute__alu_lt_t0,
i_pipeline__i_pipeline_s2_execute__alu_lt,
i_pipeline__i_pipeline_s2_execute__alu_op_add_t0,
i_pipeline__i_pipeline_s2_execute__alu_op_add,
i_pipeline__i_pipeline_s2_execute__alu_op_and_t0,
i_pipeline__i_pipeline_s2_execute__alu_op_and,
i_pipeline__i_pipeline_s2_execute__alu_op_cmp_t0,
i_pipeline__i_pipeline_s2_execute__alu_op_cmp,
i_pipeline__i_pipeline_s2_execute__alu_op_or_t0,
i_pipeline__i_pipeline_s2_execute__alu_op_or,
i_pipeline__i_pipeline_s2_execute__alu_op_rot_t0,
i_pipeline__i_pipeline_s2_execute__alu_op_rot,
i_pipeline__i_pipeline_s2_execute__alu_op_shf_arith_t0,
i_pipeline__i_pipeline_s2_execute__alu_op_shf_arith,
i_pipeline__i_pipeline_s2_execute__alu_op_shf_left_t0,
i_pipeline__i_pipeline_s2_execute__alu_op_shf_left,
i_pipeline__i_pipeline_s2_execute__alu_op_shf_t0,
i_pipeline__i_pipeline_s2_execute__alu_op_shf,
i_pipeline__i_pipeline_s2_execute__alu_op_sub_t0,
i_pipeline__i_pipeline_s2_execute__alu_op_sub,
i_pipeline__i_pipeline_s2_execute__alu_op_unsigned_t0,
i_pipeline__i_pipeline_s2_execute__alu_op_unsigned,
i_pipeline__i_pipeline_s2_execute__alu_op_xor_t0,
i_pipeline__i_pipeline_s2_execute__alu_op_xor,
i_pipeline__i_pipeline_s2_execute__alu_ready_t0,
i_pipeline__i_pipeline_s2_execute__alu_ready,
i_pipeline__i_pipeline_s2_execute__alu_result_t0,
i_pipeline__i_pipeline_s2_execute__alu_result,
i_pipeline__i_pipeline_s2_execute__asi_done_t0,
i_pipeline__i_pipeline_s2_execute__asi_done,
i_pipeline__i_pipeline_s2_execute__asi_finished_t0,
i_pipeline__i_pipeline_s2_execute__asi_finished,
i_pipeline__i_pipeline_s2_execute__asi_flush_aesmix_t0,
i_pipeline__i_pipeline_s2_execute__asi_flush_aesmix,
i_pipeline__i_pipeline_s2_execute__asi_flush_aessub_t0,
i_pipeline__i_pipeline_s2_execute__asi_flush_aessub,
i_pipeline__i_pipeline_s2_execute__asi_ready_t0,
i_pipeline__i_pipeline_s2_execute__asi_ready,
i_pipeline__i_pipeline_s2_execute__asi_result_t0,
i_pipeline__i_pipeline_s2_execute__asi_result,
i_pipeline__i_pipeline_s2_execute__bitw_bop_lut_t0,
i_pipeline__i_pipeline_s2_execute__bitw_bop_lut,
i_pipeline__i_pipeline_s2_execute__bitw_bop_t0,
i_pipeline__i_pipeline_s2_execute__bitw_bop,
i_pipeline__i_pipeline_s2_execute__bitw_cmov_t0,
i_pipeline__i_pipeline_s2_execute__bitw_cmov,
i_pipeline__i_pipeline_s2_execute__bitw_flush_t0,
i_pipeline__i_pipeline_s2_execute__bitw_flush,
i_pipeline__i_pipeline_s2_execute__bitw_fsl_t0,
i_pipeline__i_pipeline_s2_execute__bitw_fsl,
i_pipeline__i_pipeline_s2_execute__bitw_fsr_t0,
i_pipeline__i_pipeline_s2_execute__bitw_fsr,
i_pipeline__i_pipeline_s2_execute__bitw_gpr_wide_t0,
i_pipeline__i_pipeline_s2_execute__bitw_gpr_wide,
i_pipeline__i_pipeline_s2_execute__bitw_lut_t0,
i_pipeline__i_pipeline_s2_execute__bitw_lut,
i_pipeline__i_pipeline_s2_execute__bitw_ready_t0,
i_pipeline__i_pipeline_s2_execute__bitw_ready,
i_pipeline__i_pipeline_s2_execute__bitw_result_wide_t0,
i_pipeline__i_pipeline_s2_execute__bitw_result_wide,
i_pipeline__i_pipeline_s2_execute__cfu_cond_t0,
i_pipeline__i_pipeline_s2_execute__cfu_cond,
i_pipeline__i_pipeline_s2_execute__cfu_cond_taken_t0,
i_pipeline__i_pipeline_s2_execute__cfu_cond_taken,
i_pipeline__i_pipeline_s2_execute__cfu_jalr_t0,
i_pipeline__i_pipeline_s2_execute__cfu_jalr,
i_pipeline__i_pipeline_s2_execute__cond_beq_t0,
i_pipeline__i_pipeline_s2_execute__cond_beq,
i_pipeline__i_pipeline_s2_execute__cond_bge_t0,
i_pipeline__i_pipeline_s2_execute__cond_bge,
i_pipeline__i_pipeline_s2_execute__cond_bgeu_t0,
i_pipeline__i_pipeline_s2_execute__cond_bgeu,
i_pipeline__i_pipeline_s2_execute__cond_blt_t0,
i_pipeline__i_pipeline_s2_execute__cond_blt,
i_pipeline__i_pipeline_s2_execute__cond_bltu_t0,
i_pipeline__i_pipeline_s2_execute__cond_bltu,
i_pipeline__i_pipeline_s2_execute__cond_bne_t0,
i_pipeline__i_pipeline_s2_execute__cond_bne,
i_pipeline__i_pipeline_s2_execute__imul_clmul_r_t0,
i_pipeline__i_pipeline_s2_execute__imul_clmul_r,
i_pipeline__i_pipeline_s2_execute__imul_clmul_t0,
i_pipeline__i_pipeline_s2_execute__imul_clmul,
i_pipeline__i_pipeline_s2_execute__imul_div_t0,
i_pipeline__i_pipeline_s2_execute__imul_div,
i_pipeline__i_pipeline_s2_execute__imul_divu_t0,
i_pipeline__i_pipeline_s2_execute__imul_divu,
i_pipeline__i_pipeline_s2_execute__imul_flush_t0,
i_pipeline__i_pipeline_s2_execute__imul_flush,
i_pipeline__i_pipeline_s2_execute__imul_gpr_wide_t0,
i_pipeline__i_pipeline_s2_execute__imul_gpr_wide,
i_pipeline__i_pipeline_s2_execute__imul_macc_t0,
i_pipeline__i_pipeline_s2_execute__imul_macc,
i_pipeline__i_pipeline_s2_execute__imul_madd_t0,
i_pipeline__i_pipeline_s2_execute__imul_madd,
i_pipeline__i_pipeline_s2_execute__imul_mmul_t0,
i_pipeline__i_pipeline_s2_execute__imul_mmul,
i_pipeline__i_pipeline_s2_execute__imul_msub_t0,
i_pipeline__i_pipeline_s2_execute__imul_msub,
i_pipeline__i_pipeline_s2_execute__imul_mul_t0,
i_pipeline__i_pipeline_s2_execute__imul_mul,
i_pipeline__i_pipeline_s2_execute__imul_mulhsu_t0,
i_pipeline__i_pipeline_s2_execute__imul_mulhsu,
i_pipeline__i_pipeline_s2_execute__imul_mulhu_t0,
i_pipeline__i_pipeline_s2_execute__imul_mulhu,
i_pipeline__i_pipeline_s2_execute__imul_pclmul_t0,
i_pipeline__i_pipeline_s2_execute__imul_pclmul,
i_pipeline__i_pipeline_s2_execute__imul_pmul_t0,
i_pipeline__i_pipeline_s2_execute__imul_pmul,
i_pipeline__i_pipeline_s2_execute__imul_pw_16_t0,
i_pipeline__i_pipeline_s2_execute__imul_pw_16,
i_pipeline__i_pipeline_s2_execute__imul_pw_2_t0,
i_pipeline__i_pipeline_s2_execute__imul_pw_2,
i_pipeline__i_pipeline_s2_execute__imul_pw_32_t0,
i_pipeline__i_pipeline_s2_execute__imul_pw_32,
i_pipeline__i_pipeline_s2_execute__imul_pw_4_t0,
i_pipeline__i_pipeline_s2_execute__imul_pw_4,
i_pipeline__i_pipeline_s2_execute__imul_pw_8_t0,
i_pipeline__i_pipeline_s2_execute__imul_pw_8,
i_pipeline__i_pipeline_s2_execute__imul_ready_t0,
i_pipeline__i_pipeline_s2_execute__imul_ready,
i_pipeline__i_pipeline_s2_execute__imul_rem_t0,
i_pipeline__i_pipeline_s2_execute__imul_rem,
i_pipeline__i_pipeline_s2_execute__imul_remu_t0,
i_pipeline__i_pipeline_s2_execute__imul_remu,
i_pipeline__i_pipeline_s2_execute__imul_result_hi_t0,
i_pipeline__i_pipeline_s2_execute__imul_result_hi,
i_pipeline__i_pipeline_s2_execute__imul_result_t0,
i_pipeline__i_pipeline_s2_execute__imul_result,
i_pipeline__i_pipeline_s2_execute__imul_result_wide_t0,
i_pipeline__i_pipeline_s2_execute__imul_result_wide,
i_pipeline__i_pipeline_s2_execute__leak_fence_t0,
i_pipeline__i_pipeline_s2_execute__leak_fence,
i_pipeline__i_pipeline_s2_execute__lsu_load_t0,
i_pipeline__i_pipeline_s2_execute__lsu_load,
i_pipeline__i_pipeline_s2_execute__lsu_store_t0,
i_pipeline__i_pipeline_s2_execute__lsu_store,
i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_cfu_t0,
i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_cfu,
i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_mul_t0,
i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_mul,
i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_rng_t0,
i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_rng,
i_pipeline__i_pipeline_s2_execute__n_s3_opr_b_t0,
i_pipeline__i_pipeline_s2_execute__n_s3_opr_b,
i_pipeline__i_pipeline_s2_execute__n_s3_uop_cfu_t0,
i_pipeline__i_pipeline_s2_execute__n_s3_uop_cfu,
i_pipeline__i_pipeline_s2_execute__n_s3_uop_t0,
i_pipeline__i_pipeline_s2_execute__n_s3_uop,
i_pipeline__i_pipeline_s2_execute__opra_flush_t0,
i_pipeline__i_pipeline_s2_execute__opra_flush,
i_pipeline__i_pipeline_s2_execute__opra_ld_en_t0,
i_pipeline__i_pipeline_s2_execute__opra_ld_en,
i_pipeline__i_pipeline_s2_execute__oprb_flush_t0,
i_pipeline__i_pipeline_s2_execute__oprb_flush,
i_pipeline__i_pipeline_s2_execute__oprb_ld_en_t0,
i_pipeline__i_pipeline_s2_execute__oprb_ld_en,
i_pipeline__i_pipeline_s2_execute__p_busy_t0,
i_pipeline__i_pipeline_s2_execute__p_busy,
i_pipeline__i_pipeline_s2_execute__p_valid_t0,
i_pipeline__i_pipeline_s2_execute__p_valid,
i_pipeline__i_pipeline_s2_execute__pipe_reg_out_t0,
i_pipeline__i_pipeline_s2_execute__pipe_reg_out,
i_pipeline__i_pipeline_s2_execute__rng_if_ready_t0,
i_pipeline__i_pipeline_s2_execute__rng_if_ready,
i_pipeline__i_pipeline_s2_execute__rng_ready_t0,
i_pipeline__i_pipeline_s2_execute__rng_ready,
i_pipeline__i_pipeline_s2_execute__rng_uop_samp_t0,
i_pipeline__i_pipeline_s2_execute__rng_uop_samp,
i_pipeline__i_pipeline_s2_execute__rng_uop_seed_t0,
i_pipeline__i_pipeline_s2_execute__rng_uop_seed,
i_pipeline__i_pipeline_s2_execute__rng_uop_test_t0,
i_pipeline__i_pipeline_s2_execute__rng_uop_test,
i_pipeline__i_pipeline_s2_execute__rng_valid_t0,
i_pipeline__i_pipeline_s2_execute__rng_valid,
i_pipeline__i_pipeline_s2_execute__i_alu__g_clk,
i_pipeline__i_pipeline_s2_execute__i_alu__g_resetn,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_valid,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_flush,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_ready,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_pw,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_add,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_sub,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_xor,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_or,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_and,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_rot,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf_left,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf_arith,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_cmp,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_unsigned,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_lt,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_eq,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_add_result,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_lhs,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_rhs,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_result,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_add_result_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_eq_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_flush_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_lt_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_add_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_and_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_cmp_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_or_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_rot_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf_arith_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf_left_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_sub_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_unsigned_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_xor_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_pw_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_ready_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_result_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_valid_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_lt_signed_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_lt_signed,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_lt_unsigned_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__alu_lt_unsigned,
i_pipeline__i_pipeline_s2_execute__i_alu__bw_result_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__bw_result,
i_pipeline__i_pipeline_s2_execute__i_alu__out_adder_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__out_adder,
i_pipeline__i_pipeline_s2_execute__i_alu__out_bw_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__out_bw,
i_pipeline__i_pipeline_s2_execute__i_alu__out_shift_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__out_shift,
i_pipeline__i_pipeline_s2_execute__i_alu__pw_d_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__pw_d,
i_pipeline__i_pipeline_s2_execute__i_alu__shift_arith_mask_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__shift_arith_mask,
i_pipeline__i_pipeline_s2_execute__i_alu__shift_arith_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__shift_arith,
i_pipeline__i_pipeline_s2_execute__i_alu__shift_out_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__shift_out,
i_pipeline__i_pipeline_s2_execute__i_alu__shift_result_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__shift_result,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__lhs,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__rhs,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__pw,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__cin,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__sub,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__c_en,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__c_out,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__result,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__c_en_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__c_out_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__cin_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__pw_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__result_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__sub_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__carry_mask_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__carry_mask,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_0___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_0___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_0___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_0___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_10___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_10___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_10___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_10___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_11___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_11___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_11___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_11___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_11___force_carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_11___force_carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_12___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_12___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_12___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_12___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_13___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_13___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_13___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_13___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_13___force_carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_13___force_carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_14___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_14___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_14___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_14___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_15___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_15___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_15___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_15___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_15___force_carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_15___force_carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_16___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_16___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_16___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_16___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_17___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_17___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_17___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_17___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_18___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_18___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_18___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_18___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_19___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_19___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_19___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_19___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_1___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_1___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_1___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_1___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_20___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_20___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_20___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_20___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_21___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_21___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_21___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_21___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_22___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_22___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_22___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_22___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_23___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_23___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_23___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_23___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_23___force_carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_23___force_carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_24___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_24___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_24___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_24___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_25___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_25___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_25___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_25___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_26___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_26___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_26___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_26___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_27___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_27___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_27___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_27___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_28___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_28___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_28___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_28___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_29___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_29___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_29___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_29___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_2___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_2___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_2___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_2___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_30___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_30___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_30___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_30___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_31___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_31___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_31___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_31___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_3___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_3___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_3___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_3___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_4___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_4___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_4___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_4___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_5___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_5___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_5___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_5___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_6___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_6___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_6___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_6___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_7___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_7___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_7___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_7___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_8___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_8___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_8___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_8___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_9___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_9___c_in,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_9___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_9___carry,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__rhs_m_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__rhs_m,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__crs1,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__shamt,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__pw,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__shift,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__rotate,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__left,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__right,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__result,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__pw_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__result_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__crs1_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__left_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__right_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__rotate_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__shamt_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__shift_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_16_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_16,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_32_left_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_32_left,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_32_right_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_32_right,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_16_left_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_16_left,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_16_right_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_16_right,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_2_left_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_2_left,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_2_right_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_2_right,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_16_left_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_16_left,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_16_right_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_16_right,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_2_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_2,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_4_left_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_4_left,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_4_right_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_4_right,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_16_left_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_16_left,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_16_right_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_16_right,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_2_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_2,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_8_left_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_8_left,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_8_right_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_8_right,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_16_left_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_16_left,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_16_right_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_16_right,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_2_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_2,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_16_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_16,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_2_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_2,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_32_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_32,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_4_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_4,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_8_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_8,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_16_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_16,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_2_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_2,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_32_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_32,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_4_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_4,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_8_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_8,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_16_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_16,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_2_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_2,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_32_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_32,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_4_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_4,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_8_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_8,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_16_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_16,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_2_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_2,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_32_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_32,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_4_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_4,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_8_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_8,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_2_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_2,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_16_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_16,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_32_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_32,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_4_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_4,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_8_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_8,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_16_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_16,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_32_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_32,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_4_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_4,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_8_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_8,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_16_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_16,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_2_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_2,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_32_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_32,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_4_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_4,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_8_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_8,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_16_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_16,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_2_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_2,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_32_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_32,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_4_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_4,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_8_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_8,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_16_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_16,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_2_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_2,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_32_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_32,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_4_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_4,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_8_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_8,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_16_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_16,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_2_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_2,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_32_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_32,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_4_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_4,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_8_t0,
i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_8,
i_pipeline__i_pipeline_s2_execute__i_asi__g_clk,
i_pipeline__i_pipeline_s2_execute__i_asi__g_resetn,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_valid,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_ready,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_aessub,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_aesmix,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_data,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_uop,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_rs1,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_rs2,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_shamt,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_result,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_aesmix_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_aessub_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_data_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_ready_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_result_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_rs2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_shamt_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_uop_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__asi_valid_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_ready_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_ready,
i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_rs1,
i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_rs2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_rs2,
i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_ready_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_ready,
i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_rs1,
i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_rs2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_rs2,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_aes_mix_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_aes_mix,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_aes_sub_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_aes_sub,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_aes_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_aes,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha2,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_x1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_x1,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_x2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_x2,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_x4_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_x4,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_xy_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_xy,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_yx_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_yx,
i_pipeline__i_pipeline_s2_execute__i_asi__result_aesmix_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__result_aesmix,
i_pipeline__i_pipeline_s2_execute__i_asi__result_aessub_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__result_aessub,
i_pipeline__i_pipeline_s2_execute__i_asi__result_sha2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__result_sha2,
i_pipeline__i_pipeline_s2_execute__i_asi__result_sha3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__result_sha3,
i_pipeline__i_pipeline_s2_execute__i_asi__sha2_rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__sha2_rs1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__clock,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__reset,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__flush,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__flush_data,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__valid,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__rs1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__rs2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__enc,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__ready,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__result,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__flush_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__result_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__ready_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__rs2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__valid_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__flush_data_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__enc_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__b_0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__b_0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__b_1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__b_1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__b_2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__b_2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__b_3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__b_3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_0_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_0_lhs,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_0_out_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_0_out,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_1_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_1_lhs,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_1_out_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_1_out,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_2_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_2_lhs,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_2_out_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_2_out,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_3_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_3_lhs,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_3_out_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_3_out,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_byte_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_byte,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_byte_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_byte,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x0_in_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x0_in,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x1_in_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x1_in,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x2_in_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x2_in,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x2_out_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x2_out,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x3_in_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x3_in,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x3_out_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x3_out,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__fsm_0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__fsm_0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__fsm_1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__fsm_1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__fsm_2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__fsm_2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__fsm_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__fsm,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__n_fsm_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__n_fsm,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__clock,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__reset,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__flush,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__flush_data,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__valid,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rs1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rs2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__enc,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rot,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__ready,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__result,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__flush_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__result_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__ready_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rs2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__valid_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__flush_data_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__enc_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rot_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__b_0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__b_0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__b_1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__b_1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__b_2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__b_2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__fsm_0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__fsm_0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__fsm_1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__fsm_1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__fsm_2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__fsm_2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__fsm_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__fsm,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__n_fsm_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__n_fsm,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_in_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_in,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_out_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_out,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__in,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__inv,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__in_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__inv_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out_fwd_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out_fwd,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out_inv_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out_inv,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__in,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__out,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__in_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__out_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s4_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s4,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s5_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s5,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s6_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s6,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s7_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s7,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t10_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t10,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t11_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t11,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t12_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t12,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t13_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t13,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t14_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t14,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t15_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t15,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t16_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t16,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t17_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t17,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t18_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t18,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t19_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t19,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t20_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t20,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t21_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t21,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t22_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t22,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t23_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t23,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t24_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t24,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t25_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t25,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t26_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t26,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t27_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t27,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t28_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t28,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t29_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t29,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t30_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t30,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t31_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t31,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t32_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t32,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t33_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t33,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t34_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t34,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t35_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t35,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t36_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t36,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t37_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t37,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t38_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t38,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t39_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t39,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t40_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t40,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t41_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t41,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t42_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t42,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t43_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t43,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t44_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t44,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t45_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t45,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t4_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t4,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t5_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t5,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t6_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t6,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t7_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t7,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t8_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t8,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t9_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t9,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc10_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc10,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc11_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc11,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc12_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc12,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc13_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc13,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc14_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc14,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc16_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc16,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc17_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc17,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc18_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc18,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc20_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc20,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc21_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc21,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc26_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc26,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc4_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc4,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc5_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc5,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc6_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc6,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc7_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc7,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc8_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc8,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc9_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc9,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y10_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y10,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y11_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y11,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y12_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y12,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y13_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y13,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y14_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y14,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y15_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y15,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y16_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y16,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y17_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y17,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y18_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y18,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y19_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y19,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y20_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y20,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y21_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y21,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y4_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y4,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y5_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y5,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y6_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y6,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y7_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y7,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y8_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y8,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y9_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y9,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z10_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z10,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z11_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z11,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z12_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z12,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z13_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z13,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z14_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z14,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z15_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z15,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z16_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z16,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z17_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z17,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z4_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z4,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z5_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z5,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z6_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z6,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z7_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z7,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z8_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z8,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z9_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z9,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__in,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__out,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__in_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__out_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__aa_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__aa,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab20_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab20,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab21_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab21,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab22_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab22,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab23_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab23,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd4_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd4,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd5_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd5,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd6_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd6,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ah_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ah,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__al_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__al,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__bb_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__bb,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__bh_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__bh,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__bl_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__bl,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp4_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp4,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__dd_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__dd,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__dh_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__dh,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__dl_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__dl,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p4_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p4,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p6_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p6,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p7_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p7,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph01_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph01,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph02_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph02,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph03_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph03,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph11_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph11,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph12_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph12,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph13_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph13,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl01_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl01,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl02_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl02,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl03_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl03,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl11_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl11,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl12_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl12,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl13_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl13,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pr1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pr1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pr2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pr2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pr3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pr3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__qr1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__qr1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__qr2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__qr2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__qr3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__qr3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r10_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r10,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r11_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r11,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r4_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r4,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r5_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r5,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r6_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r6,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r7_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r7,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r8_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r8,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r9_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r9,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rr1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rr1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rr2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rr2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rtl0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rtl0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rtl1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rtl1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rtl2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rtl2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s4_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s4,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s5_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s5,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s6_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s6,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s7_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s7,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sa0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sa0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sa1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sa1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sb0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sb0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sb1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sb1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sd0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sd0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sd1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sd1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__t01_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__t01,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__t02_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__t02,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv10_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv10,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv11_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv11,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv12_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv12,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv13_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv13,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv4_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv4,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv5_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv5,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv6_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv6,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv7_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv7,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv8_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv8,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv9_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv9,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__vr1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__vr1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__vr2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__vr2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__vr3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__vr3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__wr1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__wr1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__wr2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__wr2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__wr3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__wr3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x11_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x11,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x13_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x13,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x14_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x14,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x16_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x16,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x18_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x18,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x19_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x19,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y4_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y4,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y5_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y5,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y6_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y6,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y7_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y7,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__rs1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__ss,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__result,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__result_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__ss_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s0_result_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s0_result,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s0_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s1_result_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s1_result,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s2_result_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s2_result,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s3_result_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s3_result,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s3_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s3,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__rs1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__rs2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shamt,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_xy,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x4,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_yx,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__result,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__result_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shamt_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__rs2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x4_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_xy_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_yx_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__in_x_plus_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__in_x_plus,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__in_y_plus_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__in_y_plus,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_in_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_in_lhs,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_in_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_in_rhs,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_out_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_out_lhs,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_out_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_out_rhs,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__result_sum_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__result_sum,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shf_1_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shf_1,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shf_2_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shf_2,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__sum_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__sum_rhs,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__g_clk,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__g_resetn,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_data,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_valid,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_busy,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__mr_data,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__flush,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__flush_dat,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_data,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_valid,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_busy,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__flush_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_valid_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_data_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_busy_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__mr_data_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_valid_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_data_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_busy_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__flush_dat_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__genblk1__progress_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__genblk1__progress,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__g_clk,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__g_resetn,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_data,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_valid,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_busy,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__mr_data,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__flush,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__flush_dat,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_data,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_valid,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_busy,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__flush_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_valid_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_data_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_busy_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__mr_data_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_valid_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_data_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_busy_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__flush_dat_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__genblk1__progress_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__genblk1__progress,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__g_clk,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__g_resetn,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_data,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_valid,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_busy,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__mr_data,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__flush,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__flush_dat,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_data,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_valid,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_busy,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__flush_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_valid_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_data_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_busy_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__mr_data_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_valid_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_data_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_busy_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__flush_dat_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__genblk1__progress_t0,
i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__genblk1__progress,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs1,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs2,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs3,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__bop_lut,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__flush,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__valid,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_fsl,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_fsr,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_mror,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_cmov,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_lut,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_bop,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__ready,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__flush_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__ready_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs2_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__valid_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs3_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__bop_lut_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_bop_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_cmov_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_fsl_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_fsr_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_lut_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_mror_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__r_in_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__r_in,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__r_out_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__r_out,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__ramt_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__ramt,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_bop_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_bop,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_cmov_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_cmov,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_fsl_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_fsl,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_lut_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_lut,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_0_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_1_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_1,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_2_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_2,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_3_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_3,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_4_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_4,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_5_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_5,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rword_l_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rword_l,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs1,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs2,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs3,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__result,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__result_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs1_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs2_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs3_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rd,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rs1,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rs2,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__lut,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__result,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__result_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rs2_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__lut_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rd_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__g_clk,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__g_resetn,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__flush,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__pipeline_progress,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__valid,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rs1,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_valid,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_op,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_data,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_ready,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_valid,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_status,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_data,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_ready,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_test,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_seed,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_samp,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__result,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__ready,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__flush_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__result_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__ready_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__valid_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__pipeline_progress_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_data_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_op_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_ready_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_valid_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_data_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_ready_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_status_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_valid_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_samp_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_seed_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_test_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__n_req_done_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__n_req_done,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__req_done_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__req_done,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__status_healthy_t0,
i_pipeline__i_pipeline_s2_execute__i_frv_rngif__status_healthy,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__clock,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__resetn,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs1,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs2,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs3,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__flush,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__flush_data,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__valid,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_div,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_divu,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_rem,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_remu,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mul,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mulu,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mulsu,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_clmul,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_pmul,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_pclmul,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_madd,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_msub,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_macc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mmul,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_32,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_16,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_8,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_4,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_2,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__result,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__ready,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__flush_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mul_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__result_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_16_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_2_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_32_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_4_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_8_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__ready_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs2_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__valid_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs3_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_macc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_madd_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mmul_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_msub_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__flush_data_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_clmul_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_div_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_divu_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mulsu_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mulu_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_pclmul_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_pmul_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_rem_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_remu_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__arg_0_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__arg_0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__arg_1_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__arg_1,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__count_en_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__count_en,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__count_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__count,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__do_mulu_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__do_mulu,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__fsm_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__fsm,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__insn_divrem_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__insn_divrem,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__insn_long_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__insn_long,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__insn_mdr_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__insn_mdr,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__ld_long_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__ld_long,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__ld_mdr_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__ld_mdr,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__ld_on_init_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__ld_on_init,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_n_acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_n_acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_n_carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_n_carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_cin_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_cin,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_lhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_rhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_sub_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_sub,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_ready_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_ready,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_result_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_result,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_arg_0_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_arg_0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_arg_1_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_arg_1,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_cen_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_cen,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_cin_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_cin,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_lhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_rhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_sub_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_sub,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_ready_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_ready,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_result_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_result,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_arg_0_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_arg_0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_count_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_count,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_fsm_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_fsm,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_cen_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_cen,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_cin_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_cin,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_cout_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_cout,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_lhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_result_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_result,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_rhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_sub_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_sub,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__reg_ld_en_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__reg_ld_en,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__clock,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__resetn,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs1,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs2,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs3,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__flush,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__valid,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_div,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_divu,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_rem,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_remu,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mul,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mulu,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mulsu,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_clmul,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_pmul,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_pclmul,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_32,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_16,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_8,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_4,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_2,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__count,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_1,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_arg_0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_arg_1,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_lhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_rhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_sub,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cin,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cen,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cout,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_result,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__result,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__ready,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__flush_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__result_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_0_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__count_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_arg_0_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cen_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cin_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cout_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_result_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_sub_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_16_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_2_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_32_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_4_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_8_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__ready_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs2_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_1_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_arg_1_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__valid_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_clmul_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_div_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_divu_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mul_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mulsu_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mulu_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_pclmul_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_pmul_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_rem_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_remu_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs3_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_sel_neg_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_sel_neg,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_sel_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_sel,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_n_acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_n_acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_n_arg_0_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_n_arg_0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_outsign_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_outsign,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_ready_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_ready,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_signed_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_signed,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__divrem_result_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__divrem_result,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_carryless_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_carryless,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_lhs_sign_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_lhs_sign,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_n_acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_n_acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_n_arg_0_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_n_arg_0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_cen_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_cen,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_cin_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_cin,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_lhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_rhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_sub_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_sub,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_ready_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_ready,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_n_acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_n_acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_n_arg_0_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_n_arg_0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_cen_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_cen,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_lhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_rhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_sub_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_sub,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_ready_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_ready,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_result_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_result,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rem_outsign_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rem_outsign,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__result_div_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__result_div,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__result_rem_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__result_rem,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__route_div_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__route_div,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__route_mul_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__route_mul,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__route_pmul_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__route_pmul,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__rs1,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__rs2,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__count,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__arg_0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__carryless,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_16,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_8,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_4,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_2,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_lhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_rhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_sub,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_cen,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_cout,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_result,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__n_acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__n_arg_0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__result,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__ready,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__result_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__arg_0_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__carryless_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__count_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__n_acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__n_arg_0_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_cen_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_cout_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_result_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_sub_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_16_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_2_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_4_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_8_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__ready_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__rs2_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_mask_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_mask,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pmul_result_0_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pmul_result_0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__clock,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__resetn,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__rs1,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__rs2,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__valid,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__op_signed,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__flush,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__count,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__arg_0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__arg_1,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_arg_0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_arg_1,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__ready,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__flush_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__arg_0_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__count_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_arg_0_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__ready_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__rs2_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__arg_1_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_arg_1_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__op_signed_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__valid_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__div_less_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__div_less,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__div_run_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__div_run,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__div_start_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__div_start,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__divisor_start_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__divisor_start,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__qmask_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__qmask,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__signed_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__signed_lhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__signed_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__signed_rhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__sub_result_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__sub_result,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rs1,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rs2,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__count,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__arg_0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__carryless,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_32,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_16,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_8,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_4,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_2,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__lhs_sign,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rhs_sign,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_lhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_rhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_sub,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cin,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cen,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cout,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_result,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__n_acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__n_arg_0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__ready,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__arg_0_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__carryless_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__count_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__lhs_sign_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__n_acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__n_arg_0_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cen_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cin_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cout_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_result_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_sub_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_16_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_2_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_32_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_4_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_8_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__ready_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rhs_sign_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rs2_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_32_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_32,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_lhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_rhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__lhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__rhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__pw,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__cin,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__sub,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__c_en,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__c_out,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__result,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__c_en_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__c_out_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__cin_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__pw_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__result_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__sub_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__carry_mask_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__carry_mask,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_0___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_0___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_0___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_0___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_10___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_10___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_10___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_10___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_11___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_11___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_11___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_11___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_11___force_carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_11___force_carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_12___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_12___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_12___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_12___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_13___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_13___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_13___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_13___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_13___force_carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_13___force_carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_14___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_14___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_14___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_14___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_15___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_15___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_15___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_15___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_15___force_carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_15___force_carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_16___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_16___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_16___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_16___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_17___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_17___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_17___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_17___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_18___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_18___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_18___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_18___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_19___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_19___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_19___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_19___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_1___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_1___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_1___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_1___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_20___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_20___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_20___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_20___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_21___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_21___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_21___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_21___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_22___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_22___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_22___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_22___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_23___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_23___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_23___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_23___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_23___force_carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_23___force_carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_24___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_24___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_24___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_24___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_25___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_25___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_25___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_25___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_26___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_26___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_26___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_26___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_27___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_27___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_27___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_27___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_28___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_28___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_28___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_28___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_29___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_29___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_29___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_29___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_2___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_2___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_2___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_2___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_30___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_30___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_30___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_30___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_31___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_31___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_31___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_31___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_3___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_3___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_3___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_3___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_4___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_4___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_4___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_4___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_5___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_5___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_5___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_5___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_6___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_6___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_6___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_6___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_7___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_7___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_7___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_7___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_8___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_8___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_8___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_8___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_9___c_in_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_9___c_in,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_9___carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_9___carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__rhs_m_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__rhs_m,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs1,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs2,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs3,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_init,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mdr,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_msub_1,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_macc_1,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mmul_1,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mmul_2,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_done,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__count,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_lhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_rhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_cin,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_sub,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_cout,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_result,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_madd,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_msub,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_macc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_mmul,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__n_carry,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__n_acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__result,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__ready,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__result_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__count_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__n_acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_cin_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_cout_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_result_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_sub_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__ready_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs1_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs2_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs3_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_done_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_init_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_macc_1_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mdr_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mmul_1_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mmul_2_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_msub_1_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__n_carry_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_macc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_madd_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_mmul_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_msub_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_lhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_n_acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_n_acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_rhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_lhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_n_acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_n_acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_rhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__msub_lhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__msub_lhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__msub_rhs_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__msub_rhs,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__result_acc_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__result_acc,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__sub_result_t0,
i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__sub_result,
i_pipeline__i_pipeline_s3_memory__g_clk,
i_pipeline__i_pipeline_s3_memory__g_resetn,
i_pipeline__i_pipeline_s3_memory__flush,
i_pipeline__i_pipeline_s3_memory__s3_rd,
i_pipeline__i_pipeline_s3_memory__s3_opr_a,
i_pipeline__i_pipeline_s3_memory__s3_opr_b,
i_pipeline__i_pipeline_s3_memory__s3_uop,
i_pipeline__i_pipeline_s3_memory__s3_fu,
i_pipeline__i_pipeline_s3_memory__s3_trap,
i_pipeline__i_pipeline_s3_memory__s3_size,
i_pipeline__i_pipeline_s3_memory__s3_instr,
i_pipeline__i_pipeline_s3_memory__s3_busy,
i_pipeline__i_pipeline_s3_memory__s3_valid,
i_pipeline__i_pipeline_s3_memory__leak_prng,
i_pipeline__i_pipeline_s3_memory__leak_lkgcfg,
i_pipeline__i_pipeline_s3_memory__leak_fence_unc0,
i_pipeline__i_pipeline_s3_memory__leak_fence_unc1,
i_pipeline__i_pipeline_s3_memory__leak_fence_unc2,
i_pipeline__i_pipeline_s3_memory__fwd_s3_rd,
i_pipeline__i_pipeline_s3_memory__fwd_s3_wide,
i_pipeline__i_pipeline_s3_memory__fwd_s3_wdata,
i_pipeline__i_pipeline_s3_memory__fwd_s3_wdata_hi,
i_pipeline__i_pipeline_s3_memory__fwd_s3_load,
i_pipeline__i_pipeline_s3_memory__fwd_s3_csr,
i_pipeline__i_pipeline_s3_memory__hold_lsu_req,
i_pipeline__i_pipeline_s3_memory__mmio_en,
i_pipeline__i_pipeline_s3_memory__mmio_wen,
i_pipeline__i_pipeline_s3_memory__mmio_addr,
i_pipeline__i_pipeline_s3_memory__mmio_wdata,
i_pipeline__i_pipeline_s3_memory__dmem_req,
i_pipeline__i_pipeline_s3_memory__dmem_wen,
i_pipeline__i_pipeline_s3_memory__dmem_strb,
i_pipeline__i_pipeline_s3_memory__dmem_wdata,
i_pipeline__i_pipeline_s3_memory__dmem_addr,
i_pipeline__i_pipeline_s3_memory__dmem_gnt,
i_pipeline__i_pipeline_s3_memory__s4_rd,
i_pipeline__i_pipeline_s3_memory__s4_opr_a,
i_pipeline__i_pipeline_s3_memory__s4_opr_b,
i_pipeline__i_pipeline_s3_memory__s4_uop,
i_pipeline__i_pipeline_s3_memory__s4_fu,
i_pipeline__i_pipeline_s3_memory__s4_trap,
i_pipeline__i_pipeline_s3_memory__s4_size,
i_pipeline__i_pipeline_s3_memory__s4_instr,
i_pipeline__i_pipeline_s3_memory__s4_busy,
i_pipeline__i_pipeline_s3_memory__s4_valid,
i_pipeline__i_pipeline_s3_memory__flush_t0,
i_pipeline__i_pipeline_s3_memory__leak_lkgcfg_t0,
i_pipeline__i_pipeline_s3_memory__leak_prng_t0,
i_pipeline__i_pipeline_s3_memory__mmio_wen_t0,
i_pipeline__i_pipeline_s3_memory__mmio_wdata_t0,
i_pipeline__i_pipeline_s3_memory__mmio_en_t0,
i_pipeline__i_pipeline_s3_memory__mmio_addr_t0,
i_pipeline__i_pipeline_s3_memory__s3_busy_t0,
i_pipeline__i_pipeline_s3_memory__s3_fu_t0,
i_pipeline__i_pipeline_s3_memory__s3_instr_t0,
i_pipeline__i_pipeline_s3_memory__s3_opr_a_t0,
i_pipeline__i_pipeline_s3_memory__s3_opr_b_t0,
i_pipeline__i_pipeline_s3_memory__s3_rd_t0,
i_pipeline__i_pipeline_s3_memory__s3_size_t0,
i_pipeline__i_pipeline_s3_memory__s3_trap_t0,
i_pipeline__i_pipeline_s3_memory__s3_uop_t0,
i_pipeline__i_pipeline_s3_memory__s3_valid_t0,
i_pipeline__i_pipeline_s3_memory__dmem_addr_t0,
i_pipeline__i_pipeline_s3_memory__dmem_gnt_t0,
i_pipeline__i_pipeline_s3_memory__dmem_req_t0,
i_pipeline__i_pipeline_s3_memory__dmem_strb_t0,
i_pipeline__i_pipeline_s3_memory__dmem_wdata_t0,
i_pipeline__i_pipeline_s3_memory__dmem_wen_t0,
i_pipeline__i_pipeline_s3_memory__hold_lsu_req_t0,
i_pipeline__i_pipeline_s3_memory__fwd_s3_csr_t0,
i_pipeline__i_pipeline_s3_memory__fwd_s3_load_t0,
i_pipeline__i_pipeline_s3_memory__fwd_s3_rd_t0,
i_pipeline__i_pipeline_s3_memory__fwd_s3_wdata_t0,
i_pipeline__i_pipeline_s3_memory__fwd_s3_wdata_hi_t0,
i_pipeline__i_pipeline_s3_memory__fwd_s3_wide_t0,
i_pipeline__i_pipeline_s3_memory__leak_fence_unc0_t0,
i_pipeline__i_pipeline_s3_memory__leak_fence_unc1_t0,
i_pipeline__i_pipeline_s3_memory__leak_fence_unc2_t0,
i_pipeline__i_pipeline_s3_memory__s4_busy_t0,
i_pipeline__i_pipeline_s3_memory__s4_fu_t0,
i_pipeline__i_pipeline_s3_memory__s4_instr_t0,
i_pipeline__i_pipeline_s3_memory__s4_opr_a_t0,
i_pipeline__i_pipeline_s3_memory__s4_opr_b_t0,
i_pipeline__i_pipeline_s3_memory__s4_rd_t0,
i_pipeline__i_pipeline_s3_memory__s4_size_t0,
i_pipeline__i_pipeline_s3_memory__s4_trap_t0,
i_pipeline__i_pipeline_s3_memory__s4_uop_t0,
i_pipeline__i_pipeline_s3_memory__s4_valid_t0,
i_pipeline__i_pipeline_s3_memory__bitw_gpr_wide_t0,
i_pipeline__i_pipeline_s3_memory__bitw_gpr_wide,
i_pipeline__i_pipeline_s3_memory__imul_gpr_wide_t0,
i_pipeline__i_pipeline_s3_memory__imul_gpr_wide,
i_pipeline__i_pipeline_s3_memory__leak_fence_t0,
i_pipeline__i_pipeline_s3_memory__leak_fence,
i_pipeline__i_pipeline_s3_memory__lsu_a_error_t0,
i_pipeline__i_pipeline_s3_memory__lsu_a_error,
i_pipeline__i_pipeline_s3_memory__lsu_byte_t0,
i_pipeline__i_pipeline_s3_memory__lsu_byte,
i_pipeline__i_pipeline_s3_memory__lsu_cause_t0,
i_pipeline__i_pipeline_s3_memory__lsu_cause,
i_pipeline__i_pipeline_s3_memory__lsu_half_t0,
i_pipeline__i_pipeline_s3_memory__lsu_half,
i_pipeline__i_pipeline_s3_memory__lsu_mmio_t0,
i_pipeline__i_pipeline_s3_memory__lsu_mmio,
i_pipeline__i_pipeline_s3_memory__lsu_ready_t0,
i_pipeline__i_pipeline_s3_memory__lsu_ready,
i_pipeline__i_pipeline_s3_memory__lsu_word_t0,
i_pipeline__i_pipeline_s3_memory__lsu_word,
i_pipeline__i_pipeline_s3_memory__n_s4_opr_a_t0,
i_pipeline__i_pipeline_s3_memory__n_s4_opr_a,
i_pipeline__i_pipeline_s3_memory__n_s4_opr_b_t0,
i_pipeline__i_pipeline_s3_memory__n_s4_opr_b,
i_pipeline__i_pipeline_s3_memory__n_s4_rd_t0,
i_pipeline__i_pipeline_s3_memory__n_s4_rd,
i_pipeline__i_pipeline_s3_memory__n_s4_trap_t0,
i_pipeline__i_pipeline_s3_memory__n_s4_trap,
i_pipeline__i_pipeline_s3_memory__opra_flush_t0,
i_pipeline__i_pipeline_s3_memory__opra_flush,
i_pipeline__i_pipeline_s3_memory__opra_ld_en_t0,
i_pipeline__i_pipeline_s3_memory__opra_ld_en,
i_pipeline__i_pipeline_s3_memory__oprb_flush_t0,
i_pipeline__i_pipeline_s3_memory__oprb_flush,
i_pipeline__i_pipeline_s3_memory__oprb_ld_en_t0,
i_pipeline__i_pipeline_s3_memory__oprb_ld_en,
i_pipeline__i_pipeline_s3_memory__p_busy_t0,
i_pipeline__i_pipeline_s3_memory__p_busy,
i_pipeline__i_pipeline_s3_memory__p_valid_t0,
i_pipeline__i_pipeline_s3_memory__p_valid,
i_pipeline__i_pipeline_s3_memory__pipe_reg_out_t0,
i_pipeline__i_pipeline_s3_memory__pipe_reg_out,
i_pipeline__i_pipeline_s3_memory__i_lsu__g_clk,
i_pipeline__i_pipeline_s3_memory__i_lsu__g_resetn,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_valid,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_a_error,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_ready,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_mmio,
i_pipeline__i_pipeline_s3_memory__i_lsu__pipe_prog,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_addr,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_wdata,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_load,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_store,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_byte,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_half,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_word,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_signed,
i_pipeline__i_pipeline_s3_memory__i_lsu__hold_lsu_req,
i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_en,
i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_wen,
i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_addr,
i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_wdata,
i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_req,
i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_wen,
i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_strb,
i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_wdata,
i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_addr,
i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_gnt,
i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_wen_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_wdata_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_en_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_addr_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_load_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_store_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_addr_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_gnt_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_req_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_strb_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_wdata_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_wen_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__hold_lsu_req_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_a_error_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_addr_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_byte_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_half_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_mmio_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_ready_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_signed_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_valid_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_wdata_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_word_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__pipe_prog_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_txn_done_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_txn_done,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_finished_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_finished,
i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_done_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_done,
i_pipeline__i_pipeline_s3_memory__i_lsu__n_lsu_finished_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__n_lsu_finished,
i_pipeline__i_pipeline_s3_memory__i_lsu__n_mmio_done_t0,
i_pipeline__i_pipeline_s3_memory__i_lsu__n_mmio_done,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__g_clk,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__g_resetn,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_data,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_valid,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_busy,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__mr_data,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__flush,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__flush_dat,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_data,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_valid,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_busy,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__flush_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_valid_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_data_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_busy_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__mr_data_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_valid_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_data_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_busy_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__flush_dat_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__genblk1__progress_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__genblk1__progress,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__g_clk,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__g_resetn,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_data,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_valid,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_busy,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__mr_data,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__flush,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__flush_dat,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_data,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_valid,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_busy,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__flush_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_valid_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_data_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_busy_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__mr_data_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_valid_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_data_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_busy_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__flush_dat_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__genblk1__progress_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__genblk1__progress,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__g_clk,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__g_resetn,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_data,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_valid,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_busy,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__mr_data,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__flush,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__flush_dat,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_data,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_valid,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_busy,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__flush_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_valid_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_data_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_busy_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__mr_data_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_valid_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_data_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_busy_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__flush_dat_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__genblk1__progress_t0,
i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__genblk1__progress,
i_pipeline__i_pipeline_s4_writeback__g_clk,
i_pipeline__i_pipeline_s4_writeback__g_resetn,
i_pipeline__i_pipeline_s4_writeback__s4_rd,
i_pipeline__i_pipeline_s4_writeback__s4_opr_a,
i_pipeline__i_pipeline_s4_writeback__s4_opr_b,
i_pipeline__i_pipeline_s4_writeback__s4_uop,
i_pipeline__i_pipeline_s4_writeback__s4_fu,
i_pipeline__i_pipeline_s4_writeback__s4_trap,
i_pipeline__i_pipeline_s4_writeback__s4_size,
i_pipeline__i_pipeline_s4_writeback__s4_instr,
i_pipeline__i_pipeline_s4_writeback__s4_busy,
i_pipeline__i_pipeline_s4_writeback__s4_valid,
i_pipeline__i_pipeline_s4_writeback__fwd_s4_rd,
i_pipeline__i_pipeline_s4_writeback__fwd_s4_wdata,
i_pipeline__i_pipeline_s4_writeback__fwd_s4_load,
i_pipeline__i_pipeline_s4_writeback__fwd_s4_csr,
i_pipeline__i_pipeline_s4_writeback__gpr_wen,
i_pipeline__i_pipeline_s4_writeback__gpr_wide,
i_pipeline__i_pipeline_s4_writeback__gpr_rd,
i_pipeline__i_pipeline_s4_writeback__gpr_wdata,
i_pipeline__i_pipeline_s4_writeback__gpr_wdata_hi,
i_pipeline__i_pipeline_s4_writeback__int_trap_req,
i_pipeline__i_pipeline_s4_writeback__int_trap_cause,
i_pipeline__i_pipeline_s4_writeback__int_trap_ack,
i_pipeline__i_pipeline_s4_writeback__trap_cpu,
i_pipeline__i_pipeline_s4_writeback__trap_int,
i_pipeline__i_pipeline_s4_writeback__trap_cause,
i_pipeline__i_pipeline_s4_writeback__trap_mtval,
i_pipeline__i_pipeline_s4_writeback__trap_pc,
i_pipeline__i_pipeline_s4_writeback__exec_mret,
i_pipeline__i_pipeline_s4_writeback__csr_mepc,
i_pipeline__i_pipeline_s4_writeback__csr_mtvec,
i_pipeline__i_pipeline_s4_writeback__vector_intrs,
i_pipeline__i_pipeline_s4_writeback__trs_pc,
i_pipeline__i_pipeline_s4_writeback__trs_instr,
i_pipeline__i_pipeline_s4_writeback__trs_valid,
i_pipeline__i_pipeline_s4_writeback__csr_en,
i_pipeline__i_pipeline_s4_writeback__csr_wr,
i_pipeline__i_pipeline_s4_writeback__csr_wr_set,
i_pipeline__i_pipeline_s4_writeback__csr_wr_clr,
i_pipeline__i_pipeline_s4_writeback__csr_addr,
i_pipeline__i_pipeline_s4_writeback__csr_wdata,
i_pipeline__i_pipeline_s4_writeback__csr_rdata,
i_pipeline__i_pipeline_s4_writeback__csr_error,
i_pipeline__i_pipeline_s4_writeback__cf_req,
i_pipeline__i_pipeline_s4_writeback__cf_target,
i_pipeline__i_pipeline_s4_writeback__cf_ack,
i_pipeline__i_pipeline_s4_writeback__hold_lsu_req,
i_pipeline__i_pipeline_s4_writeback__mmio_rdata,
i_pipeline__i_pipeline_s4_writeback__mmio_error,
i_pipeline__i_pipeline_s4_writeback__dmem_recv,
i_pipeline__i_pipeline_s4_writeback__dmem_ack,
i_pipeline__i_pipeline_s4_writeback__dmem_error,
i_pipeline__i_pipeline_s4_writeback__dmem_rdata,
i_pipeline__i_pipeline_s4_writeback__cf_target_t0,
i_pipeline__i_pipeline_s4_writeback__cf_req_t0,
i_pipeline__i_pipeline_s4_writeback__cf_ack_t0,
i_pipeline__i_pipeline_s4_writeback__int_trap_req_t0,
i_pipeline__i_pipeline_s4_writeback__mmio_rdata_t0,
i_pipeline__i_pipeline_s4_writeback__mmio_error_t0,
i_pipeline__i_pipeline_s4_writeback__int_trap_cause_t0,
i_pipeline__i_pipeline_s4_writeback__int_trap_ack_t0,
i_pipeline__i_pipeline_s4_writeback__trap_cause_t0,
i_pipeline__i_pipeline_s4_writeback__hold_lsu_req_t0,
i_pipeline__i_pipeline_s4_writeback__s4_busy_t0,
i_pipeline__i_pipeline_s4_writeback__s4_fu_t0,
i_pipeline__i_pipeline_s4_writeback__s4_instr_t0,
i_pipeline__i_pipeline_s4_writeback__s4_opr_a_t0,
i_pipeline__i_pipeline_s4_writeback__s4_opr_b_t0,
i_pipeline__i_pipeline_s4_writeback__s4_rd_t0,
i_pipeline__i_pipeline_s4_writeback__s4_size_t0,
i_pipeline__i_pipeline_s4_writeback__s4_trap_t0,
i_pipeline__i_pipeline_s4_writeback__s4_uop_t0,
i_pipeline__i_pipeline_s4_writeback__s4_valid_t0,
i_pipeline__i_pipeline_s4_writeback__csr_addr_t0,
i_pipeline__i_pipeline_s4_writeback__csr_en_t0,
i_pipeline__i_pipeline_s4_writeback__csr_error_t0,
i_pipeline__i_pipeline_s4_writeback__csr_mepc_t0,
i_pipeline__i_pipeline_s4_writeback__csr_mtvec_t0,
i_pipeline__i_pipeline_s4_writeback__csr_rdata_t0,
i_pipeline__i_pipeline_s4_writeback__csr_wdata_t0,
i_pipeline__i_pipeline_s4_writeback__csr_wr_t0,
i_pipeline__i_pipeline_s4_writeback__csr_wr_clr_t0,
i_pipeline__i_pipeline_s4_writeback__csr_wr_set_t0,
i_pipeline__i_pipeline_s4_writeback__dmem_ack_t0,
i_pipeline__i_pipeline_s4_writeback__dmem_error_t0,
i_pipeline__i_pipeline_s4_writeback__dmem_rdata_t0,
i_pipeline__i_pipeline_s4_writeback__dmem_recv_t0,
i_pipeline__i_pipeline_s4_writeback__exec_mret_t0,
i_pipeline__i_pipeline_s4_writeback__fwd_s4_csr_t0,
i_pipeline__i_pipeline_s4_writeback__fwd_s4_load_t0,
i_pipeline__i_pipeline_s4_writeback__fwd_s4_rd_t0,
i_pipeline__i_pipeline_s4_writeback__fwd_s4_wdata_t0,
i_pipeline__i_pipeline_s4_writeback__gpr_rd_t0,
i_pipeline__i_pipeline_s4_writeback__gpr_wdata_t0,
i_pipeline__i_pipeline_s4_writeback__gpr_wdata_hi_t0,
i_pipeline__i_pipeline_s4_writeback__gpr_wen_t0,
i_pipeline__i_pipeline_s4_writeback__gpr_wide_t0,
i_pipeline__i_pipeline_s4_writeback__trap_cpu_t0,
i_pipeline__i_pipeline_s4_writeback__trap_int_t0,
i_pipeline__i_pipeline_s4_writeback__trap_mtval_t0,
i_pipeline__i_pipeline_s4_writeback__trap_pc_t0,
i_pipeline__i_pipeline_s4_writeback__trs_instr_t0,
i_pipeline__i_pipeline_s4_writeback__trs_pc_t0,
i_pipeline__i_pipeline_s4_writeback__trs_valid_t0,
i_pipeline__i_pipeline_s4_writeback__vector_intrs_t0,
i_pipeline__i_pipeline_s4_writeback__cf_req_noint_t0,
i_pipeline__i_pipeline_s4_writeback__cf_req_noint,
i_pipeline__i_pipeline_s4_writeback__cf_target_noint_t0,
i_pipeline__i_pipeline_s4_writeback__cf_target_noint,
i_pipeline__i_pipeline_s4_writeback__cfu_busy_t0,
i_pipeline__i_pipeline_s4_writeback__cfu_busy,
i_pipeline__i_pipeline_s4_writeback__cfu_cf_taken_t0,
i_pipeline__i_pipeline_s4_writeback__cfu_cf_taken,
i_pipeline__i_pipeline_s4_writeback__cfu_done_t0,
i_pipeline__i_pipeline_s4_writeback__cfu_done,
i_pipeline__i_pipeline_s4_writeback__cfu_ebreak_t0,
i_pipeline__i_pipeline_s4_writeback__cfu_ebreak,
i_pipeline__i_pipeline_s4_writeback__cfu_ecall_t0,
i_pipeline__i_pipeline_s4_writeback__cfu_ecall,
i_pipeline__i_pipeline_s4_writeback__cfu_finish_now_t0,
i_pipeline__i_pipeline_s4_writeback__cfu_finish_now,
i_pipeline__i_pipeline_s4_writeback__cfu_gpr_wdata_t0,
i_pipeline__i_pipeline_s4_writeback__cfu_gpr_wdata,
i_pipeline__i_pipeline_s4_writeback__cfu_gpr_wen_t0,
i_pipeline__i_pipeline_s4_writeback__cfu_gpr_wen,
i_pipeline__i_pipeline_s4_writeback__cfu_mret_t0,
i_pipeline__i_pipeline_s4_writeback__cfu_mret,
i_pipeline__i_pipeline_s4_writeback__cfu_tgt_trap_t0,
i_pipeline__i_pipeline_s4_writeback__cfu_tgt_trap,
i_pipeline__i_pipeline_s4_writeback__cfu_trap_t0,
i_pipeline__i_pipeline_s4_writeback__cfu_trap,
i_pipeline__i_pipeline_s4_writeback__csr_done_t0,
i_pipeline__i_pipeline_s4_writeback__csr_done,
i_pipeline__i_pipeline_s4_writeback__csr_gpr_wen_t0,
i_pipeline__i_pipeline_s4_writeback__csr_gpr_wen,
i_pipeline__i_pipeline_s4_writeback__csr_read_t0,
i_pipeline__i_pipeline_s4_writeback__csr_read,
i_pipeline__i_pipeline_s4_writeback__dmem_error_seen_t0,
i_pipeline__i_pipeline_s4_writeback__dmem_error_seen,
i_pipeline__i_pipeline_s4_writeback__lsu_b_error_t0,
i_pipeline__i_pipeline_s4_writeback__lsu_b_error,
i_pipeline__i_pipeline_s4_writeback__lsu_busy_t0,
i_pipeline__i_pipeline_s4_writeback__lsu_busy,
i_pipeline__i_pipeline_s4_writeback__lsu_byte_t0,
i_pipeline__i_pipeline_s4_writeback__lsu_byte,
i_pipeline__i_pipeline_s4_writeback__lsu_gpr_wen_t0,
i_pipeline__i_pipeline_s4_writeback__lsu_gpr_wen,
i_pipeline__i_pipeline_s4_writeback__lsu_half_t0,
i_pipeline__i_pipeline_s4_writeback__lsu_half,
i_pipeline__i_pipeline_s4_writeback__lsu_load_t0,
i_pipeline__i_pipeline_s4_writeback__lsu_load,
i_pipeline__i_pipeline_s4_writeback__lsu_mmio_t0,
i_pipeline__i_pipeline_s4_writeback__lsu_mmio,
i_pipeline__i_pipeline_s4_writeback__lsu_rsp_seen_t0,
i_pipeline__i_pipeline_s4_writeback__lsu_rsp_seen,
i_pipeline__i_pipeline_s4_writeback__lsu_store_t0,
i_pipeline__i_pipeline_s4_writeback__lsu_store,
i_pipeline__i_pipeline_s4_writeback__lsu_txn_recv_t0,
i_pipeline__i_pipeline_s4_writeback__lsu_txn_recv,
i_pipeline__i_pipeline_s4_writeback__lsu_word_t0,
i_pipeline__i_pipeline_s4_writeback__lsu_word,
i_pipeline__i_pipeline_s4_writeback__mem_rdata_t0,
i_pipeline__i_pipeline_s4_writeback__mem_rdata,
i_pipeline__i_pipeline_s4_writeback__n_cfu_done_t0,
i_pipeline__i_pipeline_s4_writeback__n_cfu_done,
i_pipeline__i_pipeline_s4_writeback__n_csr_done_t0,
i_pipeline__i_pipeline_s4_writeback__n_csr_done,
i_pipeline__i_pipeline_s4_writeback__n_dmem_error_seen_t0,
i_pipeline__i_pipeline_s4_writeback__n_dmem_error_seen,
i_pipeline__i_pipeline_s4_writeback__n_lsu_rsp_seen_t0,
i_pipeline__i_pipeline_s4_writeback__n_lsu_rsp_seen,
i_pipeline__i_pipeline_s4_writeback__pipe_progress_t0,
i_pipeline__i_pipeline_s4_writeback__pipe_progress,
i_pipeline__i_pipeline_s4_writeback__rdata_b0_t0,
i_pipeline__i_pipeline_s4_writeback__rdata_b0,
i_pipeline__i_pipeline_s4_writeback__rdata_b1_t0,
i_pipeline__i_pipeline_s4_writeback__rdata_b1,
i_pipeline__i_pipeline_s4_writeback__rdata_h1_t0,
i_pipeline__i_pipeline_s4_writeback__rdata_h1,
i_pipeline__i_pipeline_s4_writeback__rng_gpr_wen_t0,
i_pipeline__i_pipeline_s4_writeback__rng_gpr_wen,
i_pipeline__i_pipeline_s4_writeback__trap_int_pending_t0,
i_pipeline__i_pipeline_s4_writeback__trap_int_pending,
i_pipeline__i_pipeline_s4_writeback__trap_target_addr_t0,
i_pipeline__i_pipeline_s4_writeback__trap_target_addr,
i_pipeline__i_pipeline_s4_writeback__trap_vector_offset_t0,
i_pipeline__i_pipeline_s4_writeback__trap_vector_offset);


input logic g_clk;
input logic g_resetn;
input logic [31:0] trs_pc;
input logic [31:0] trs_instr;
input logic trs_valid;
input logic [31:0] leak_prng;
input logic leak_fence_unc0;
input logic leak_fence_unc1;
input logic leak_fence_unc2;
input logic rng_req_valid;
input logic [2:0] rng_req_op;
input logic [31:0] rng_req_data;
input logic rng_req_ready;
input logic rng_rsp_valid;
input logic [2:0] rng_rsp_status;
input logic [31:0] rng_rsp_data;
input logic rng_rsp_ready;
input logic int_nmi;
input logic int_external;
input logic [3:0] int_extern_cause;
input logic int_software;
input logic int_mtime;
input logic imem_req;
input logic imem_wen;
input logic [3:0] imem_strb;
input logic [31:0] imem_wdata;
input logic [31:0] imem_addr;
input logic imem_gnt;
input logic imem_recv;
input logic imem_ack;
input logic imem_error;
input logic [31:0] imem_rdata;
input logic dmem_req;
input logic dmem_wen;
input logic [3:0] dmem_strb;
input logic [31:0] dmem_wdata;
input logic [31:0] dmem_addr;
input logic dmem_gnt;
input logic dmem_recv;
input logic dmem_ack;
input logic dmem_error;
input logic [31:0] dmem_rdata;
input logic [31:0] leak_prng_t0;
input logic imem_wen_t0;
input logic [31:0] imem_wdata_t0;
input logic [3:0] imem_strb_t0;
input logic imem_req_t0;
input logic imem_recv_t0;
input logic [31:0] imem_rdata_t0;
input logic imem_gnt_t0;
input logic imem_error_t0;
input logic [31:0] imem_addr_t0;
input logic imem_ack_t0;
input logic [31:0] rng_req_data_t0;
input logic [2:0] rng_req_op_t0;
input logic rng_req_ready_t0;
input logic rng_req_valid_t0;
input logic [31:0] rng_rsp_data_t0;
input logic rng_rsp_ready_t0;
input logic [2:0] rng_rsp_status_t0;
input logic rng_rsp_valid_t0;
input logic [31:0] dmem_addr_t0;
input logic dmem_gnt_t0;
input logic dmem_req_t0;
input logic [3:0] dmem_strb_t0;
input logic [31:0] dmem_wdata_t0;
input logic dmem_wen_t0;
input logic leak_fence_unc0_t0;
input logic leak_fence_unc1_t0;
input logic leak_fence_unc2_t0;
input logic dmem_ack_t0;
input logic dmem_error_t0;
input logic [31:0] dmem_rdata_t0;
input logic dmem_recv_t0;
input logic [31:0] trs_instr_t0;
input logic [31:0] trs_pc_t0;
input logic trs_valid_t0;
input logic [3:0] int_extern_cause_t0;
input logic int_external_t0;
input logic int_mtime_t0;
input logic int_nmi_t0;
input logic int_software_t0;
input logic [63:0] ctr_cycle_t0;
input logic [63:0] ctr_cycle;
input logic [63:0] ctr_instret_t0;
input logic [63:0] ctr_instret;
input logic [63:0] ctr_time_t0;
input logic [63:0] ctr_time;
input logic inhibit_cy_t0;
input logic inhibit_cy;
input logic inhibit_ir_t0;
input logic inhibit_ir;
input logic inhibit_tm_t0;
input logic inhibit_tm;
input logic instr_ret_t0;
input logic instr_ret;
input logic int_trap_ack_t0;
input logic int_trap_ack;
input logic [5:0] int_trap_cause_t0;
input logic [5:0] int_trap_cause;
input logic int_trap_req_t0;
input logic int_trap_req;
input logic mie_meie_t0;
input logic mie_meie;
input logic mie_msie_t0;
input logic mie_msie;
input logic mie_mtie_t0;
input logic mie_mtie;
input logic mip_meip_t0;
input logic mip_meip;
input logic mip_msip_t0;
input logic mip_msip;
input logic [31:0] mmio_addr_t0;
input logic [31:0] mmio_addr;
input logic mmio_en_t0;
input logic mmio_en;
input logic mmio_error_t0;
input logic mmio_error;
input logic [31:0] mmio_rdata_t0;
input logic [31:0] mmio_rdata;
input logic [31:0] mmio_wdata_t0;
input logic [31:0] mmio_wdata;
input logic mmio_wen_t0;
input logic mmio_wen;
input logic mstatus_mie_t0;
input logic mstatus_mie;
input logic ti_pending_t0;
input logic ti_pending;
input logic i_counters__g_clk;
input logic i_counters__g_resetn;
input logic i_counters__instr_ret;
input logic i_counters__timer_interrupt;
input logic [63:0] i_counters__ctr_time;
input logic [63:0] i_counters__ctr_cycle;
input logic [63:0] i_counters__ctr_instret;
input logic i_counters__inhibit_cy;
input logic i_counters__inhibit_tm;
input logic i_counters__inhibit_ir;
input logic i_counters__mmio_en;
input logic i_counters__mmio_wen;
input logic [31:0] i_counters__mmio_addr;
input logic [31:0] i_counters__mmio_wdata;
input logic [31:0] i_counters__mmio_rdata;
input logic i_counters__mmio_error;
input logic i_counters__timer_interrupt_t0;
input logic i_counters__mmio_wen_t0;
input logic [31:0] i_counters__mmio_wdata_t0;
input logic [31:0] i_counters__mmio_rdata_t0;
input logic i_counters__mmio_error_t0;
input logic i_counters__mmio_en_t0;
input logic [31:0] i_counters__mmio_addr_t0;
input logic i_counters__instr_ret_t0;
input logic i_counters__inhibit_tm_t0;
input logic i_counters__inhibit_ir_t0;
input logic i_counters__inhibit_cy_t0;
input logic [63:0] i_counters__ctr_time_t0;
input logic [63:0] i_counters__ctr_instret_t0;
input logic [63:0] i_counters__ctr_cycle_t0;
input logic i_counters__addr_mtime_hi_t0;
input logic i_counters__addr_mtime_hi;
input logic i_counters__addr_mtime_lo_t0;
input logic i_counters__addr_mtime_lo;
input logic i_counters__addr_mtimecmp_hi_t0;
input logic i_counters__addr_mtimecmp_hi;
input logic i_counters__addr_mtimecmp_lo_t0;
input logic i_counters__addr_mtimecmp_lo;
input logic [63:0] i_counters__mapped_mtimecmp_t0;
input logic [63:0] i_counters__mapped_mtimecmp;
input logic [63:0] i_counters__n_ctr_cycle_t0;
input logic [63:0] i_counters__n_ctr_cycle;
input logic [63:0] i_counters__n_ctr_instret_t0;
input logic [63:0] i_counters__n_ctr_instret;
input logic [63:0] i_counters__n_mapped_mtime_t0;
input logic [63:0] i_counters__n_mapped_mtime;
input logic i_counters__n_mmio_error_t0;
input logic i_counters__n_mmio_error;
input logic [31:0] i_counters__n_mmio_rdata_t0;
input logic [31:0] i_counters__n_mmio_rdata;
input logic i_counters__n_timer_interrupt_t0;
input logic i_counters__n_timer_interrupt;
input logic i_counters__wr_mtime_hi_t0;
input logic i_counters__wr_mtime_hi;
input logic i_counters__wr_mtime_lo_t0;
input logic i_counters__wr_mtime_lo;
input logic i_counters__wr_mtimecmp_hi_t0;
input logic i_counters__wr_mtimecmp_hi;
input logic i_counters__wr_mtimecmp_lo_t0;
input logic i_counters__wr_mtimecmp_lo;
input logic i_interrupts__g_clk;
input logic i_interrupts__g_resetn;
input logic i_interrupts__mstatus_mie;
input logic i_interrupts__mie_meie;
input logic i_interrupts__mie_mtie;
input logic i_interrupts__mie_msie;
input logic i_interrupts__nmi_pending;
input logic i_interrupts__ex_pending;
input logic [3:0] i_interrupts__ex_cause;
input logic i_interrupts__ti_pending;
input logic i_interrupts__sw_pending;
input logic i_interrupts__mip_meip;
input logic i_interrupts__mip_mtip;
input logic i_interrupts__mip_msip;
input logic i_interrupts__int_trap_req;
input logic [5:0] i_interrupts__int_trap_cause;
input logic i_interrupts__int_trap_ack;
input logic i_interrupts__nmi_pending_t0;
input logic i_interrupts__mstatus_mie_t0;
input logic i_interrupts__mip_mtip_t0;
input logic i_interrupts__mie_mtie_t0;
input logic i_interrupts__mie_msie_t0;
input logic i_interrupts__sw_pending_t0;
input logic i_interrupts__ti_pending_t0;
input logic i_interrupts__int_trap_req_t0;
input logic [3:0] i_interrupts__ex_cause_t0;
input logic i_interrupts__ex_pending_t0;
input logic [5:0] i_interrupts__int_trap_cause_t0;
input logic i_interrupts__int_trap_ack_t0;
input logic i_interrupts__mie_meie_t0;
input logic i_interrupts__mip_msip_t0;
input logic i_interrupts__mip_meip_t0;
input logic [5:0] i_interrupts__extern_cause_t0;
input logic [5:0] i_interrupts__extern_cause;
input logic i_interrupts__mip_nmi_t0;
input logic i_interrupts__mip_nmi;
input logic [5:0] i_interrupts__n_int_trap_cause_t0;
input logic [5:0] i_interrupts__n_int_trap_cause;
input logic i_interrupts__raise_mei_t0;
input logic i_interrupts__raise_mei;
input logic i_interrupts__raise_msi_t0;
input logic i_interrupts__raise_msi;
input logic i_interrupts__raise_mti_t0;
input logic i_interrupts__raise_mti;
input logic i_interrupts__raise_nmi_t0;
input logic i_interrupts__raise_nmi;
input logic i_interrupts__use_extern_cause_t0;
input logic i_interrupts__use_extern_cause;
input logic i_pipeline__g_clk;
input logic i_pipeline__g_resetn;
input logic [31:0] i_pipeline__trs_pc;
input logic [31:0] i_pipeline__trs_instr;
input logic i_pipeline__trs_valid;
input logic [31:0] i_pipeline__leak_prng;
input logic i_pipeline__leak_fence_unc0;
input logic i_pipeline__leak_fence_unc1;
input logic i_pipeline__leak_fence_unc2;
input logic i_pipeline__rng_req_valid;
input logic [2:0] i_pipeline__rng_req_op;
input logic [31:0] i_pipeline__rng_req_data;
input logic i_pipeline__rng_req_ready;
input logic i_pipeline__rng_rsp_valid;
input logic [2:0] i_pipeline__rng_rsp_status;
input logic [31:0] i_pipeline__rng_rsp_data;
input logic i_pipeline__rng_rsp_ready;
input logic i_pipeline__instr_ret;
input logic i_pipeline__mstatus_mie;
input logic i_pipeline__mie_meie;
input logic i_pipeline__mie_mtie;
input logic i_pipeline__mie_msie;
input logic i_pipeline__mip_meip;
input logic i_pipeline__mip_mtip;
input logic i_pipeline__mip_msip;
input logic [63:0] i_pipeline__ctr_time;
input logic [63:0] i_pipeline__ctr_cycle;
input logic [63:0] i_pipeline__ctr_instret;
input logic i_pipeline__int_trap_req;
input logic [5:0] i_pipeline__int_trap_cause;
input logic i_pipeline__int_trap_ack;
input logic i_pipeline__inhibit_cy;
input logic i_pipeline__inhibit_tm;
input logic i_pipeline__inhibit_ir;
input logic i_pipeline__mmio_en;
input logic i_pipeline__mmio_wen;
input logic [31:0] i_pipeline__mmio_addr;
input logic [31:0] i_pipeline__mmio_wdata;
input logic [31:0] i_pipeline__mmio_rdata;
input logic i_pipeline__mmio_error;
input logic i_pipeline__imem_req;
input logic i_pipeline__imem_wen;
input logic [3:0] i_pipeline__imem_strb;
input logic [31:0] i_pipeline__imem_wdata;
input logic [31:0] i_pipeline__imem_addr;
input logic i_pipeline__imem_gnt;
input logic i_pipeline__imem_recv;
input logic i_pipeline__imem_ack;
input logic i_pipeline__imem_error;
input logic [31:0] i_pipeline__imem_rdata;
input logic i_pipeline__dmem_req;
input logic i_pipeline__dmem_wen;
input logic [3:0] i_pipeline__dmem_strb;
input logic [31:0] i_pipeline__dmem_wdata;
input logic [31:0] i_pipeline__dmem_addr;
input logic i_pipeline__dmem_gnt;
input logic i_pipeline__dmem_recv;
input logic i_pipeline__dmem_ack;
input logic i_pipeline__dmem_error;
input logic [31:0] i_pipeline__dmem_rdata;
input logic i_pipeline__mstatus_mie_t0;
input logic i_pipeline__mip_mtip_t0;
input logic i_pipeline__mie_mtie_t0;
input logic i_pipeline__mie_msie_t0;
input logic [31:0] i_pipeline__leak_prng_t0;
input logic i_pipeline__imem_wen_t0;
input logic [31:0] i_pipeline__imem_wdata_t0;
input logic [3:0] i_pipeline__imem_strb_t0;
input logic i_pipeline__imem_req_t0;
input logic i_pipeline__imem_recv_t0;
input logic [31:0] i_pipeline__imem_rdata_t0;
input logic i_pipeline__imem_gnt_t0;
input logic i_pipeline__imem_error_t0;
input logic [31:0] i_pipeline__imem_addr_t0;
input logic i_pipeline__imem_ack_t0;
input logic i_pipeline__int_trap_req_t0;
input logic i_pipeline__mmio_wen_t0;
input logic [31:0] i_pipeline__mmio_wdata_t0;
input logic [31:0] i_pipeline__mmio_rdata_t0;
input logic i_pipeline__mmio_error_t0;
input logic i_pipeline__mmio_en_t0;
input logic [31:0] i_pipeline__mmio_addr_t0;
input logic i_pipeline__instr_ret_t0;
input logic i_pipeline__inhibit_tm_t0;
input logic i_pipeline__inhibit_ir_t0;
input logic i_pipeline__inhibit_cy_t0;
input logic [63:0] i_pipeline__ctr_time_t0;
input logic [63:0] i_pipeline__ctr_instret_t0;
input logic [63:0] i_pipeline__ctr_cycle_t0;
input logic [5:0] i_pipeline__int_trap_cause_t0;
input logic i_pipeline__int_trap_ack_t0;
input logic i_pipeline__mie_meie_t0;
input logic i_pipeline__mip_msip_t0;
input logic i_pipeline__mip_meip_t0;
input logic [31:0] i_pipeline__rng_req_data_t0;
input logic [2:0] i_pipeline__rng_req_op_t0;
input logic i_pipeline__rng_req_ready_t0;
input logic i_pipeline__rng_req_valid_t0;
input logic [31:0] i_pipeline__rng_rsp_data_t0;
input logic i_pipeline__rng_rsp_ready_t0;
input logic [2:0] i_pipeline__rng_rsp_status_t0;
input logic i_pipeline__rng_rsp_valid_t0;
input logic [31:0] i_pipeline__dmem_addr_t0;
input logic i_pipeline__dmem_gnt_t0;
input logic i_pipeline__dmem_req_t0;
input logic [3:0] i_pipeline__dmem_strb_t0;
input logic [31:0] i_pipeline__dmem_wdata_t0;
input logic i_pipeline__dmem_wen_t0;
input logic i_pipeline__leak_fence_unc0_t0;
input logic i_pipeline__leak_fence_unc1_t0;
input logic i_pipeline__leak_fence_unc2_t0;
input logic i_pipeline__dmem_ack_t0;
input logic i_pipeline__dmem_error_t0;
input logic [31:0] i_pipeline__dmem_rdata_t0;
input logic i_pipeline__dmem_recv_t0;
input logic [31:0] i_pipeline__trs_instr_t0;
input logic [31:0] i_pipeline__trs_pc_t0;
input logic i_pipeline__trs_valid_t0;
input logic i_pipeline__cf_ack_t0;
input logic i_pipeline__cf_ack;
input logic i_pipeline__cf_req_t0;
input logic i_pipeline__cf_req;
input logic [31:0] i_pipeline__cf_target_t0;
input logic [31:0] i_pipeline__cf_target;
input logic [11:0] i_pipeline__csr_addr_t0;
input logic [11:0] i_pipeline__csr_addr;
input logic i_pipeline__csr_en_t0;
input logic i_pipeline__csr_en;
input logic i_pipeline__csr_error_t0;
input logic i_pipeline__csr_error;
input logic [31:0] i_pipeline__csr_mepc_t0;
input logic [31:0] i_pipeline__csr_mepc;
input logic [31:0] i_pipeline__csr_mtvec_t0;
input logic [31:0] i_pipeline__csr_mtvec;
input logic [31:0] i_pipeline__csr_rdata_t0;
input logic [31:0] i_pipeline__csr_rdata;
input logic [31:0] i_pipeline__csr_wdata_t0;
input logic [31:0] i_pipeline__csr_wdata;
input logic i_pipeline__csr_wr_clr_t0;
input logic i_pipeline__csr_wr_clr;
input logic i_pipeline__csr_wr_set_t0;
input logic i_pipeline__csr_wr_set;
input logic i_pipeline__csr_wr_t0;
input logic i_pipeline__csr_wr;
input logic i_pipeline__exec_mret_t0;
input logic i_pipeline__exec_mret;
input logic [31:0] i_pipeline__fwd_rs1_rdata_t0;
input logic [31:0] i_pipeline__fwd_rs1_rdata;
input logic [31:0] i_pipeline__fwd_rs2_rdata_t0;
input logic [31:0] i_pipeline__fwd_rs2_rdata;
input logic [31:0] i_pipeline__fwd_rs3_rdata_t0;
input logic [31:0] i_pipeline__fwd_rs3_rdata;
input logic i_pipeline__fwd_s2_csr_t0;
input logic i_pipeline__fwd_s2_csr;
input logic i_pipeline__fwd_s2_load_t0;
input logic i_pipeline__fwd_s2_load;
input logic [4:0] i_pipeline__fwd_s2_rd_t0;
input logic [4:0] i_pipeline__fwd_s2_rd;
input logic i_pipeline__fwd_s2_rs1_hi_t0;
input logic i_pipeline__fwd_s2_rs1_hi;
input logic i_pipeline__fwd_s2_rs2_hi_t0;
input logic i_pipeline__fwd_s2_rs2_hi;
input logic i_pipeline__fwd_s2_rs3_hi_t0;
input logic i_pipeline__fwd_s2_rs3_hi;
input logic [31:0] i_pipeline__fwd_s2_wdata_hi_t0;
input logic [31:0] i_pipeline__fwd_s2_wdata_hi;
input logic [31:0] i_pipeline__fwd_s2_wdata_t0;
input logic [31:0] i_pipeline__fwd_s2_wdata;
input logic i_pipeline__fwd_s2_wide_t0;
input logic i_pipeline__fwd_s2_wide;
input logic i_pipeline__fwd_s3_csr_t0;
input logic i_pipeline__fwd_s3_csr;
input logic i_pipeline__fwd_s3_load_t0;
input logic i_pipeline__fwd_s3_load;
input logic [4:0] i_pipeline__fwd_s3_rd_t0;
input logic [4:0] i_pipeline__fwd_s3_rd;
input logic i_pipeline__fwd_s3_rs1_hi_t0;
input logic i_pipeline__fwd_s3_rs1_hi;
input logic i_pipeline__fwd_s3_rs2_hi_t0;
input logic i_pipeline__fwd_s3_rs2_hi;
input logic i_pipeline__fwd_s3_rs3_hi_t0;
input logic i_pipeline__fwd_s3_rs3_hi;
input logic [31:0] i_pipeline__fwd_s3_wdata_hi_t0;
input logic [31:0] i_pipeline__fwd_s3_wdata_hi;
input logic [31:0] i_pipeline__fwd_s3_wdata_t0;
input logic [31:0] i_pipeline__fwd_s3_wdata;
input logic i_pipeline__fwd_s3_wide_t0;
input logic i_pipeline__fwd_s3_wide;
input logic i_pipeline__fwd_s4_csr_t0;
input logic i_pipeline__fwd_s4_csr;
input logic i_pipeline__fwd_s4_load_t0;
input logic i_pipeline__fwd_s4_load;
input logic [4:0] i_pipeline__fwd_s4_rd_t0;
input logic [4:0] i_pipeline__fwd_s4_rd;
input logic i_pipeline__fwd_s4_rs1_hi_t0;
input logic i_pipeline__fwd_s4_rs1_hi;
input logic i_pipeline__fwd_s4_rs2_hi_t0;
input logic i_pipeline__fwd_s4_rs2_hi;
input logic i_pipeline__fwd_s4_rs3_hi_t0;
input logic i_pipeline__fwd_s4_rs3_hi;
input logic [31:0] i_pipeline__fwd_s4_wdata_t0;
input logic [31:0] i_pipeline__fwd_s4_wdata;
input logic [4:0] i_pipeline__gpr_rd_t0;
input logic [4:0] i_pipeline__gpr_rd;
input logic [31:0] i_pipeline__gpr_wdata_hi_t0;
input logic [31:0] i_pipeline__gpr_wdata_hi;
input logic [31:0] i_pipeline__gpr_wdata_t0;
input logic [31:0] i_pipeline__gpr_wdata;
input logic i_pipeline__gpr_wen_t0;
input logic i_pipeline__gpr_wen;
input logic i_pipeline__gpr_wide_t0;
input logic i_pipeline__gpr_wide;
input logic i_pipeline__hold_lsu_req_t0;
input logic i_pipeline__hold_lsu_req;
input logic i_pipeline__hzd_rs1_s2_t0;
input logic i_pipeline__hzd_rs1_s2;
input logic i_pipeline__hzd_rs1_s3_t0;
input logic i_pipeline__hzd_rs1_s3;
input logic i_pipeline__hzd_rs1_s4_t0;
input logic i_pipeline__hzd_rs1_s4;
input logic i_pipeline__hzd_rs2_s2_t0;
input logic i_pipeline__hzd_rs2_s2;
input logic i_pipeline__hzd_rs2_s3_t0;
input logic i_pipeline__hzd_rs2_s3;
input logic i_pipeline__hzd_rs2_s4_t0;
input logic i_pipeline__hzd_rs2_s4;
input logic i_pipeline__hzd_rs3_s2_t0;
input logic i_pipeline__hzd_rs3_s2;
input logic i_pipeline__hzd_rs3_s3_t0;
input logic i_pipeline__hzd_rs3_s3;
input logic i_pipeline__hzd_rs3_s4_t0;
input logic i_pipeline__hzd_rs3_s4;
input logic [12:0] i_pipeline__leak_lkgcfg_t0;
input logic [12:0] i_pipeline__leak_lkgcfg;
input logic i_pipeline__nz_s1_rs1_t0;
input logic i_pipeline__nz_s1_rs1;
input logic i_pipeline__nz_s1_rs2_t0;
input logic i_pipeline__nz_s1_rs2;
input logic i_pipeline__nz_s1_rs3_t0;
input logic i_pipeline__nz_s1_rs3;
input logic i_pipeline__s0_flush_t0;
input logic i_pipeline__s0_flush;
input logic i_pipeline__s1_bubble_from_s2_t0;
input logic i_pipeline__s1_bubble_from_s2;
input logic i_pipeline__s1_bubble_from_s3_t0;
input logic i_pipeline__s1_bubble_from_s3;
input logic i_pipeline__s1_bubble_from_s4_t0;
input logic i_pipeline__s1_bubble_from_s4;
input logic i_pipeline__s1_bubble_no_instr_t0;
input logic i_pipeline__s1_bubble_no_instr;
input logic i_pipeline__s1_bubble_t0;
input logic i_pipeline__s1_bubble;
input logic i_pipeline__s1_busy_t0;
input logic i_pipeline__s1_busy;
input logic [31:0] i_pipeline__s1_data_t0;
input logic [31:0] i_pipeline__s1_data;
input logic i_pipeline__s1_error_t0;
input logic i_pipeline__s1_error;
input logic i_pipeline__s1_leak_fence_t0;
input logic i_pipeline__s1_leak_fence;
input logic [4:0] i_pipeline__s1_rs1_addr_t0;
input logic [4:0] i_pipeline__s1_rs1_addr;
input logic [31:0] i_pipeline__s1_rs1_rdata_t0;
input logic [31:0] i_pipeline__s1_rs1_rdata;
input logic [4:0] i_pipeline__s1_rs2_addr_t0;
input logic [4:0] i_pipeline__s1_rs2_addr;
input logic [31:0] i_pipeline__s1_rs2_rdata_t0;
input logic [31:0] i_pipeline__s1_rs2_rdata;
input logic [4:0] i_pipeline__s1_rs3_addr_t0;
input logic [4:0] i_pipeline__s1_rs3_addr;
input logic [31:0] i_pipeline__s1_rs3_rdata_t0;
input logic [31:0] i_pipeline__s1_rs3_rdata;
input logic i_pipeline__s1_valid_t0;
input logic i_pipeline__s1_valid;
input logic i_pipeline__s2_busy_t0;
input logic i_pipeline__s2_busy;
input logic [7:0] i_pipeline__s2_fu_t0;
input logic [7:0] i_pipeline__s2_fu;
input logic [31:0] i_pipeline__s2_instr_t0;
input logic [31:0] i_pipeline__s2_instr;
input logic [31:0] i_pipeline__s2_opr_a_t0;
input logic [31:0] i_pipeline__s2_opr_a;
input logic [31:0] i_pipeline__s2_opr_b_t0;
input logic [31:0] i_pipeline__s2_opr_b;
input logic [31:0] i_pipeline__s2_opr_c_t0;
input logic [31:0] i_pipeline__s2_opr_c;
input logic [2:0] i_pipeline__s2_pw_t0;
input logic [2:0] i_pipeline__s2_pw;
input logic [4:0] i_pipeline__s2_rd_t0;
input logic [4:0] i_pipeline__s2_rd;
input logic [1:0] i_pipeline__s2_size_t0;
input logic [1:0] i_pipeline__s2_size;
input logic i_pipeline__s2_trap_t0;
input logic i_pipeline__s2_trap;
input logic [4:0] i_pipeline__s2_uop_t0;
input logic [4:0] i_pipeline__s2_uop;
input logic i_pipeline__s2_valid_t0;
input logic i_pipeline__s2_valid;
input logic i_pipeline__s3_busy_t0;
input logic i_pipeline__s3_busy;
input logic [7:0] i_pipeline__s3_fu_t0;
input logic [7:0] i_pipeline__s3_fu;
input logic [31:0] i_pipeline__s3_instr_t0;
input logic [31:0] i_pipeline__s3_instr;
input logic [31:0] i_pipeline__s3_opr_a_t0;
input logic [31:0] i_pipeline__s3_opr_a;
input logic [31:0] i_pipeline__s3_opr_b_t0;
input logic [31:0] i_pipeline__s3_opr_b;
input logic [4:0] i_pipeline__s3_rd_t0;
input logic [4:0] i_pipeline__s3_rd;
input logic [1:0] i_pipeline__s3_size_t0;
input logic [1:0] i_pipeline__s3_size;
input logic i_pipeline__s3_trap_t0;
input logic i_pipeline__s3_trap;
input logic [4:0] i_pipeline__s3_uop_t0;
input logic [4:0] i_pipeline__s3_uop;
input logic i_pipeline__s3_valid_t0;
input logic i_pipeline__s3_valid;
input logic i_pipeline__s4_busy_t0;
input logic i_pipeline__s4_busy;
input logic [7:0] i_pipeline__s4_fu_t0;
input logic [7:0] i_pipeline__s4_fu;
input logic [31:0] i_pipeline__s4_instr_t0;
input logic [31:0] i_pipeline__s4_instr;
input logic [31:0] i_pipeline__s4_opr_a_t0;
input logic [31:0] i_pipeline__s4_opr_a;
input logic [31:0] i_pipeline__s4_opr_b_t0;
input logic [31:0] i_pipeline__s4_opr_b;
input logic [4:0] i_pipeline__s4_rd_t0;
input logic [4:0] i_pipeline__s4_rd;
input logic [1:0] i_pipeline__s4_size_t0;
input logic [1:0] i_pipeline__s4_size;
input logic i_pipeline__s4_trap_t0;
input logic i_pipeline__s4_trap;
input logic [4:0] i_pipeline__s4_uop_t0;
input logic [4:0] i_pipeline__s4_uop;
input logic i_pipeline__s4_valid_t0;
input logic i_pipeline__s4_valid;
input logic [5:0] i_pipeline__trap_cause_t0;
input logic [5:0] i_pipeline__trap_cause;
input logic i_pipeline__trap_cpu_t0;
input logic i_pipeline__trap_cpu;
input logic i_pipeline__trap_int_t0;
input logic i_pipeline__trap_int;
input logic [31:0] i_pipeline__trap_mtval_t0;
input logic [31:0] i_pipeline__trap_mtval;
input logic [31:0] i_pipeline__trap_pc_t0;
input logic [31:0] i_pipeline__trap_pc;
input logic [7:0] i_pipeline__uxcrypto_b0_t0;
input logic [7:0] i_pipeline__uxcrypto_b0;
input logic [7:0] i_pipeline__uxcrypto_b1_t0;
input logic [7:0] i_pipeline__uxcrypto_b1;
input logic i_pipeline__uxcrypto_ct_t0;
input logic i_pipeline__uxcrypto_ct;
input logic i_pipeline__vector_intrs_t0;
input logic i_pipeline__vector_intrs;
input logic i_pipeline__i_csrs__g_clk;
input logic i_pipeline__i_csrs__g_resetn;
input logic i_pipeline__i_csrs__csr_en;
input logic i_pipeline__i_csrs__csr_wr;
input logic i_pipeline__i_csrs__csr_wr_set;
input logic i_pipeline__i_csrs__csr_wr_clr;
input logic [11:0] i_pipeline__i_csrs__csr_addr;
input logic [31:0] i_pipeline__i_csrs__csr_wdata;
input logic [31:0] i_pipeline__i_csrs__csr_rdata;
input logic i_pipeline__i_csrs__csr_error;
input logic [31:0] i_pipeline__i_csrs__csr_mepc;
input logic [31:0] i_pipeline__i_csrs__csr_mtvec;
input logic i_pipeline__i_csrs__vector_intrs;
input logic i_pipeline__i_csrs__exec_mret;
input logic i_pipeline__i_csrs__mstatus_mie;
input logic i_pipeline__i_csrs__mie_meie;
input logic i_pipeline__i_csrs__mie_mtie;
input logic i_pipeline__i_csrs__mie_msie;
input logic i_pipeline__i_csrs__mip_meip;
input logic i_pipeline__i_csrs__mip_mtip;
input logic i_pipeline__i_csrs__mip_msip;
input logic [63:0] i_pipeline__i_csrs__ctr_time;
input logic [63:0] i_pipeline__i_csrs__ctr_cycle;
input logic [63:0] i_pipeline__i_csrs__ctr_instret;
input logic i_pipeline__i_csrs__inhibit_cy;
input logic i_pipeline__i_csrs__inhibit_tm;
input logic i_pipeline__i_csrs__inhibit_ir;
input logic i_pipeline__i_csrs__uxcrypto_ct;
input logic [7:0] i_pipeline__i_csrs__uxcrypto_b0;
input logic [7:0] i_pipeline__i_csrs__uxcrypto_b1;
input logic [12:0] i_pipeline__i_csrs__leak_lkgcfg;
input logic i_pipeline__i_csrs__trap_cpu;
input logic i_pipeline__i_csrs__trap_int;
input logic [5:0] i_pipeline__i_csrs__trap_cause;
input logic [31:0] i_pipeline__i_csrs__trap_mtval;
input logic [31:0] i_pipeline__i_csrs__trap_pc;
input logic i_pipeline__i_csrs__mstatus_mie_t0;
input logic i_pipeline__i_csrs__mip_mtip_t0;
input logic i_pipeline__i_csrs__mie_mtie_t0;
input logic i_pipeline__i_csrs__mie_msie_t0;
input logic [12:0] i_pipeline__i_csrs__leak_lkgcfg_t0;
input logic i_pipeline__i_csrs__inhibit_tm_t0;
input logic i_pipeline__i_csrs__inhibit_ir_t0;
input logic i_pipeline__i_csrs__inhibit_cy_t0;
input logic [63:0] i_pipeline__i_csrs__ctr_time_t0;
input logic [63:0] i_pipeline__i_csrs__ctr_instret_t0;
input logic [63:0] i_pipeline__i_csrs__ctr_cycle_t0;
input logic i_pipeline__i_csrs__mie_meie_t0;
input logic i_pipeline__i_csrs__mip_msip_t0;
input logic i_pipeline__i_csrs__mip_meip_t0;
input logic [5:0] i_pipeline__i_csrs__trap_cause_t0;
input logic [7:0] i_pipeline__i_csrs__uxcrypto_b0_t0;
input logic [7:0] i_pipeline__i_csrs__uxcrypto_b1_t0;
input logic i_pipeline__i_csrs__uxcrypto_ct_t0;
input logic [11:0] i_pipeline__i_csrs__csr_addr_t0;
input logic i_pipeline__i_csrs__csr_en_t0;
input logic i_pipeline__i_csrs__csr_error_t0;
input logic [31:0] i_pipeline__i_csrs__csr_mepc_t0;
input logic [31:0] i_pipeline__i_csrs__csr_mtvec_t0;
input logic [31:0] i_pipeline__i_csrs__csr_rdata_t0;
input logic [31:0] i_pipeline__i_csrs__csr_wdata_t0;
input logic i_pipeline__i_csrs__csr_wr_t0;
input logic i_pipeline__i_csrs__csr_wr_clr_t0;
input logic i_pipeline__i_csrs__csr_wr_set_t0;
input logic i_pipeline__i_csrs__exec_mret_t0;
input logic i_pipeline__i_csrs__trap_cpu_t0;
input logic i_pipeline__i_csrs__trap_int_t0;
input logic [31:0] i_pipeline__i_csrs__trap_mtval_t0;
input logic [31:0] i_pipeline__i_csrs__trap_pc_t0;
input logic i_pipeline__i_csrs__vector_intrs_t0;
input logic i_pipeline__i_csrs__int_pulse_t0;
input logic i_pipeline__i_csrs__int_pulse;
input logic i_pipeline__i_csrs__invalid_addr_t0;
input logic i_pipeline__i_csrs__invalid_addr;
input logic i_pipeline__i_csrs__mtvec_bad_write_t0;
input logic i_pipeline__i_csrs__mtvec_bad_write;
input logic [30:0] i_pipeline__i_csrs__n_mcause_cause_t0;
input logic [30:0] i_pipeline__i_csrs__n_mcause_cause;
input logic [30:0] i_pipeline__i_csrs__n_mepc_t0;
input logic [30:0] i_pipeline__i_csrs__n_mepc;
input logic i_pipeline__i_csrs__n_mstatus_mie_t0;
input logic i_pipeline__i_csrs__n_mstatus_mie;
input logic i_pipeline__i_csrs__n_mstatus_mpie_t0;
input logic i_pipeline__i_csrs__n_mstatus_mpie;
input logic [29:0] i_pipeline__i_csrs__n_mtvec_base_t0;
input logic [29:0] i_pipeline__i_csrs__n_mtvec_base;
input logic [1:0] i_pipeline__i_csrs__n_mtvec_mode_t0;
input logic [1:0] i_pipeline__i_csrs__n_mtvec_mode;
input logic [12:0] i_pipeline__i_csrs__n_reg_lkgcfg_t0;
input logic [12:0] i_pipeline__i_csrs__n_reg_lkgcfg;
input logic [31:0] i_pipeline__i_csrs__n_reg_mie_t0;
input logic [31:0] i_pipeline__i_csrs__n_reg_mie;
input logic [31:0] i_pipeline__i_csrs__n_reg_mscratch_t0;
input logic [31:0] i_pipeline__i_csrs__n_reg_mscratch;
input logic [31:0] i_pipeline__i_csrs__n_reg_mtval_t0;
input logic [31:0] i_pipeline__i_csrs__n_reg_mtval;
input logic [7:0] i_pipeline__i_csrs__n_uxcrypto_b0_t0;
input logic [7:0] i_pipeline__i_csrs__n_uxcrypto_b0;
input logic [7:0] i_pipeline__i_csrs__n_uxcrypto_b1_t0;
input logic [7:0] i_pipeline__i_csrs__n_uxcrypto_b1;
input logic i_pipeline__i_csrs__n_uxcrypto_ct_t0;
input logic i_pipeline__i_csrs__n_uxcrypto_ct;
input logic i_pipeline__i_csrs__p_trap_int_t0;
input logic i_pipeline__i_csrs__p_trap_int;
input logic i_pipeline__i_csrs__read_cycle_t0;
input logic i_pipeline__i_csrs__read_cycle;
input logic i_pipeline__i_csrs__read_cycleh_t0;
input logic i_pipeline__i_csrs__read_cycleh;
input logic i_pipeline__i_csrs__read_instret_t0;
input logic i_pipeline__i_csrs__read_instret;
input logic i_pipeline__i_csrs__read_instreth_t0;
input logic i_pipeline__i_csrs__read_instreth;
input logic i_pipeline__i_csrs__read_lkgcfg_t0;
input logic i_pipeline__i_csrs__read_lkgcfg;
input logic i_pipeline__i_csrs__read_marchid_t0;
input logic i_pipeline__i_csrs__read_marchid;
input logic i_pipeline__i_csrs__read_mcause_t0;
input logic i_pipeline__i_csrs__read_mcause;
input logic i_pipeline__i_csrs__read_mcountin_t0;
input logic i_pipeline__i_csrs__read_mcountin;
input logic i_pipeline__i_csrs__read_mcycle_t0;
input logic i_pipeline__i_csrs__read_mcycle;
input logic i_pipeline__i_csrs__read_mcycleh_t0;
input logic i_pipeline__i_csrs__read_mcycleh;
input logic i_pipeline__i_csrs__read_medeleg_t0;
input logic i_pipeline__i_csrs__read_medeleg;
input logic i_pipeline__i_csrs__read_mepc_t0;
input logic i_pipeline__i_csrs__read_mepc;
input logic i_pipeline__i_csrs__read_mhartid_t0;
input logic i_pipeline__i_csrs__read_mhartid;
input logic i_pipeline__i_csrs__read_mideleg_t0;
input logic i_pipeline__i_csrs__read_mideleg;
input logic i_pipeline__i_csrs__read_mie_t0;
input logic i_pipeline__i_csrs__read_mie;
input logic i_pipeline__i_csrs__read_mimpid_t0;
input logic i_pipeline__i_csrs__read_mimpid;
input logic i_pipeline__i_csrs__read_minstret_t0;
input logic i_pipeline__i_csrs__read_minstret;
input logic i_pipeline__i_csrs__read_minstreth_t0;
input logic i_pipeline__i_csrs__read_minstreth;
input logic i_pipeline__i_csrs__read_mip_t0;
input logic i_pipeline__i_csrs__read_mip;
input logic i_pipeline__i_csrs__read_misa_t0;
input logic i_pipeline__i_csrs__read_misa;
input logic i_pipeline__i_csrs__read_mscratch_t0;
input logic i_pipeline__i_csrs__read_mscratch;
input logic i_pipeline__i_csrs__read_mstatus_t0;
input logic i_pipeline__i_csrs__read_mstatus;
input logic i_pipeline__i_csrs__read_mtval_t0;
input logic i_pipeline__i_csrs__read_mtval;
input logic i_pipeline__i_csrs__read_mtvec_t0;
input logic i_pipeline__i_csrs__read_mtvec;
input logic i_pipeline__i_csrs__read_mvendorid_t0;
input logic i_pipeline__i_csrs__read_mvendorid;
input logic i_pipeline__i_csrs__read_time_t0;
input logic i_pipeline__i_csrs__read_time;
input logic i_pipeline__i_csrs__read_timeh_t0;
input logic i_pipeline__i_csrs__read_timeh;
input logic i_pipeline__i_csrs__read_uxcrypto_t0;
input logic i_pipeline__i_csrs__read_uxcrypto;
input logic [30:0] i_pipeline__i_csrs__reg_mcause_cause_t0;
input logic [30:0] i_pipeline__i_csrs__reg_mcause_cause;
input logic i_pipeline__i_csrs__reg_mcause_interrupt_t0;
input logic i_pipeline__i_csrs__reg_mcause_interrupt;
input logic [30:0] i_pipeline__i_csrs__reg_mepc_mepc_t0;
input logic [30:0] i_pipeline__i_csrs__reg_mepc_mepc;
input logic [31:0] i_pipeline__i_csrs__reg_mscratch_t0;
input logic [31:0] i_pipeline__i_csrs__reg_mscratch;
input logic i_pipeline__i_csrs__reg_mstatus_mpie_t0;
input logic i_pipeline__i_csrs__reg_mstatus_mpie;
input logic [7:0] i_pipeline__i_csrs__reg_mstatus_wpri1_t0;
input logic [7:0] i_pipeline__i_csrs__reg_mstatus_wpri1;
input logic [1:0] i_pipeline__i_csrs__reg_mstatus_wpri2_t0;
input logic [1:0] i_pipeline__i_csrs__reg_mstatus_wpri2;
input logic i_pipeline__i_csrs__reg_mstatus_wpri3_t0;
input logic i_pipeline__i_csrs__reg_mstatus_wpri3;
input logic i_pipeline__i_csrs__reg_mstatus_wpri4_t0;
input logic i_pipeline__i_csrs__reg_mstatus_wpri4;
input logic [31:0] i_pipeline__i_csrs__reg_mtval_t0;
input logic [31:0] i_pipeline__i_csrs__reg_mtval;
input logic [29:0] i_pipeline__i_csrs__reg_mtvec_base_t0;
input logic [29:0] i_pipeline__i_csrs__reg_mtvec_base;
input logic [1:0] i_pipeline__i_csrs__reg_mtvec_mode_t0;
input logic [1:0] i_pipeline__i_csrs__reg_mtvec_mode;
input logic i_pipeline__i_csrs__wen_lkgcfg_t0;
input logic i_pipeline__i_csrs__wen_lkgcfg;
input logic i_pipeline__i_csrs__wen_mcause_t0;
input logic i_pipeline__i_csrs__wen_mcause;
input logic i_pipeline__i_csrs__wen_mcountin_t0;
input logic i_pipeline__i_csrs__wen_mcountin;
input logic i_pipeline__i_csrs__wen_mepc_t0;
input logic i_pipeline__i_csrs__wen_mepc;
input logic i_pipeline__i_csrs__wen_mie_t0;
input logic i_pipeline__i_csrs__wen_mie;
input logic i_pipeline__i_csrs__wen_mscratch_t0;
input logic i_pipeline__i_csrs__wen_mscratch;
input logic i_pipeline__i_csrs__wen_mstatus_mie_t0;
input logic i_pipeline__i_csrs__wen_mstatus_mie;
input logic i_pipeline__i_csrs__wen_mstatus_t0;
input logic i_pipeline__i_csrs__wen_mstatus;
input logic i_pipeline__i_csrs__wen_mtval_t0;
input logic i_pipeline__i_csrs__wen_mtval;
input logic i_pipeline__i_csrs__wen_mtvec_t0;
input logic i_pipeline__i_csrs__wen_mtvec;
input logic i_pipeline__i_csrs__wen_uxcrypto_t0;
input logic i_pipeline__i_csrs__wen_uxcrypto;
input logic i_pipeline__i_csrs__wen_valid_mcause_t0;
input logic i_pipeline__i_csrs__wen_valid_mcause;
input logic i_pipeline__i_gprs__g_clk;
input logic i_pipeline__i_gprs__g_resetn;
input logic [4:0] i_pipeline__i_gprs__rs1_addr;
input logic [31:0] i_pipeline__i_gprs__rs1_data;
input logic [4:0] i_pipeline__i_gprs__rs2_addr;
input logic [31:0] i_pipeline__i_gprs__rs2_data;
input logic [4:0] i_pipeline__i_gprs__rs3_addr;
input logic [31:0] i_pipeline__i_gprs__rs3_data;
input logic i_pipeline__i_gprs__rd_wen;
input logic i_pipeline__i_gprs__rd_wide;
input logic [4:0] i_pipeline__i_gprs__rd_addr;
input logic [31:0] i_pipeline__i_gprs__rd_wdata;
input logic [31:0] i_pipeline__i_gprs__rd_wdata_hi;
input logic [31:0] i_pipeline__i_gprs__rs3_data_t0;
input logic [4:0] i_pipeline__i_gprs__rs3_addr_t0;
input logic [31:0] i_pipeline__i_gprs__rs2_data_t0;
input logic [4:0] i_pipeline__i_gprs__rs2_addr_t0;
input logic [31:0] i_pipeline__i_gprs__rs1_data_t0;
input logic [4:0] i_pipeline__i_gprs__rs1_addr_t0;
input logic i_pipeline__i_gprs__rd_wide_t0;
input logic i_pipeline__i_gprs__rd_wen_t0;
input logic [31:0] i_pipeline__i_gprs__rd_wdata_hi_t0;
input logic [31:0] i_pipeline__i_gprs__rd_wdata_t0;
input logic [4:0] i_pipeline__i_gprs__rd_addr_t0;
input logic [31:0] i_pipeline__i_gprs__gprs_10__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_10_;
input logic [31:0] i_pipeline__i_gprs__gprs_11__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_11_;
input logic [31:0] i_pipeline__i_gprs__gprs_12__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_12_;
input logic [31:0] i_pipeline__i_gprs__gprs_13__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_13_;
input logic [31:0] i_pipeline__i_gprs__gprs_14__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_14_;
input logic [31:0] i_pipeline__i_gprs__gprs_15__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_15_;
input logic [31:0] i_pipeline__i_gprs__gprs_16__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_16_;
input logic [31:0] i_pipeline__i_gprs__gprs_17__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_17_;
input logic [31:0] i_pipeline__i_gprs__gprs_18__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_18_;
input logic [31:0] i_pipeline__i_gprs__gprs_19__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_19_;
input logic [31:0] i_pipeline__i_gprs__gprs_1__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_1_;
input logic [31:0] i_pipeline__i_gprs__gprs_20__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_20_;
input logic [31:0] i_pipeline__i_gprs__gprs_21__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_21_;
input logic [31:0] i_pipeline__i_gprs__gprs_22__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_22_;
input logic [31:0] i_pipeline__i_gprs__gprs_23__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_23_;
input logic [31:0] i_pipeline__i_gprs__gprs_24__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_24_;
input logic [31:0] i_pipeline__i_gprs__gprs_25__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_25_;
input logic [31:0] i_pipeline__i_gprs__gprs_26__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_26_;
input logic [31:0] i_pipeline__i_gprs__gprs_27__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_27_;
input logic [31:0] i_pipeline__i_gprs__gprs_28__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_28_;
input logic [31:0] i_pipeline__i_gprs__gprs_29__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_29_;
input logic [31:0] i_pipeline__i_gprs__gprs_2__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_2_;
input logic [31:0] i_pipeline__i_gprs__gprs_30__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_30_;
input logic [31:0] i_pipeline__i_gprs__gprs_31__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_31_;
input logic [31:0] i_pipeline__i_gprs__gprs_3__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_3_;
input logic [31:0] i_pipeline__i_gprs__gprs_4__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_4_;
input logic [31:0] i_pipeline__i_gprs__gprs_5__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_5_;
input logic [31:0] i_pipeline__i_gprs__gprs_6__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_6_;
input logic [31:0] i_pipeline__i_gprs__gprs_7__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_7_;
input logic [31:0] i_pipeline__i_gprs__gprs_8__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_8_;
input logic [31:0] i_pipeline__i_gprs__gprs_9__t0;
input logic [31:0] i_pipeline__i_gprs__gprs_9_;
input logic [31:0] i_pipeline__i_gprs__rd_wdata_odd_t0;
input logic [31:0] i_pipeline__i_gprs__rd_wdata_odd;
input logic i_pipeline__i_gprs__rd_wen_even_t0;
input logic i_pipeline__i_gprs__rd_wen_even;
input logic i_pipeline__i_gprs__rd_wen_odd_t0;
input logic i_pipeline__i_gprs__rd_wen_odd;
input logic i_pipeline__i_pipeline_s0_fetch__g_clk;
input logic i_pipeline__i_pipeline_s0_fetch__g_resetn;
input logic i_pipeline__i_pipeline_s0_fetch__cf_req;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__cf_target;
input logic i_pipeline__i_pipeline_s0_fetch__cf_ack;
input logic i_pipeline__i_pipeline_s0_fetch__imem_req;
input logic i_pipeline__i_pipeline_s0_fetch__imem_wen;
input logic [3:0] i_pipeline__i_pipeline_s0_fetch__imem_strb;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__imem_wdata;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__imem_addr;
input logic i_pipeline__i_pipeline_s0_fetch__imem_gnt;
input logic i_pipeline__i_pipeline_s0_fetch__imem_ack;
input logic i_pipeline__i_pipeline_s0_fetch__imem_recv;
input logic i_pipeline__i_pipeline_s0_fetch__imem_error;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__imem_rdata;
input logic i_pipeline__i_pipeline_s0_fetch__s0_flush;
input logic i_pipeline__i_pipeline_s0_fetch__s1_busy;
input logic i_pipeline__i_pipeline_s0_fetch__s1_valid;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__s1_data;
input logic i_pipeline__i_pipeline_s0_fetch__s1_error;
input logic i_pipeline__i_pipeline_s0_fetch__s1_valid_t0;
input logic i_pipeline__i_pipeline_s0_fetch__s1_error_t0;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__s1_data_t0;
input logic i_pipeline__i_pipeline_s0_fetch__s1_busy_t0;
input logic i_pipeline__i_pipeline_s0_fetch__s0_flush_t0;
input logic i_pipeline__i_pipeline_s0_fetch__imem_wen_t0;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__imem_wdata_t0;
input logic [3:0] i_pipeline__i_pipeline_s0_fetch__imem_strb_t0;
input logic i_pipeline__i_pipeline_s0_fetch__imem_req_t0;
input logic i_pipeline__i_pipeline_s0_fetch__imem_recv_t0;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__imem_rdata_t0;
input logic i_pipeline__i_pipeline_s0_fetch__imem_gnt_t0;
input logic i_pipeline__i_pipeline_s0_fetch__imem_error_t0;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__imem_addr_t0;
input logic i_pipeline__i_pipeline_s0_fetch__imem_ack_t0;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__cf_target_t0;
input logic i_pipeline__i_pipeline_s0_fetch__cf_req_t0;
input logic i_pipeline__i_pipeline_s0_fetch__cf_ack_t0;
input logic i_pipeline__i_pipeline_s0_fetch__allow_new_mem_req_t0;
input logic i_pipeline__i_pipeline_s0_fetch__allow_new_mem_req;
input logic i_pipeline__i_pipeline_s0_fetch__buf_16_t0;
input logic i_pipeline__i_pipeline_s0_fetch__buf_16;
input logic i_pipeline__i_pipeline_s0_fetch__buf_32_t0;
input logic i_pipeline__i_pipeline_s0_fetch__buf_32;
input logic [2:0] i_pipeline__i_pipeline_s0_fetch__buf_depth_t0;
input logic [2:0] i_pipeline__i_pipeline_s0_fetch__buf_depth;
input logic i_pipeline__i_pipeline_s0_fetch__buf_out_2_t0;
input logic i_pipeline__i_pipeline_s0_fetch__buf_out_2;
input logic i_pipeline__i_pipeline_s0_fetch__buf_out_4_t0;
input logic i_pipeline__i_pipeline_s0_fetch__buf_out_4;
input logic i_pipeline__i_pipeline_s0_fetch__buf_ready_t0;
input logic i_pipeline__i_pipeline_s0_fetch__buf_ready;
input logic i_pipeline__i_pipeline_s0_fetch__cf_change_t0;
input logic i_pipeline__i_pipeline_s0_fetch__cf_change;
input logic i_pipeline__i_pipeline_s0_fetch__drop_response_t0;
input logic i_pipeline__i_pipeline_s0_fetch__drop_response;
input logic i_pipeline__i_pipeline_s0_fetch__f_2byte_t0;
input logic i_pipeline__i_pipeline_s0_fetch__f_2byte;
input logic i_pipeline__i_pipeline_s0_fetch__f_4byte_t0;
input logic i_pipeline__i_pipeline_s0_fetch__f_4byte;
input logic i_pipeline__i_pipeline_s0_fetch__fetch_misaligned_t0;
input logic i_pipeline__i_pipeline_s0_fetch__fetch_misaligned;
input logic [2:0] i_pipeline__i_pipeline_s0_fetch__ignore_rsps_t0;
input logic [2:0] i_pipeline__i_pipeline_s0_fetch__ignore_rsps;
input logic i_pipeline__i_pipeline_s0_fetch__incomplete_instr_t0;
input logic i_pipeline__i_pipeline_s0_fetch__incomplete_instr;
input logic i_pipeline__i_pipeline_s0_fetch__n_fetch_misaligned_t0;
input logic i_pipeline__i_pipeline_s0_fetch__n_fetch_misaligned;
input logic [2:0] i_pipeline__i_pipeline_s0_fetch__n_ignore_rsps_t0;
input logic [2:0] i_pipeline__i_pipeline_s0_fetch__n_ignore_rsps;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__n_imem_addr_t0;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__n_imem_addr;
input logic i_pipeline__i_pipeline_s0_fetch__n_imem_req_t0;
input logic i_pipeline__i_pipeline_s0_fetch__n_imem_req;
input logic [2:0] i_pipeline__i_pipeline_s0_fetch__n_reqs_outstanding_t0;
input logic [2:0] i_pipeline__i_pipeline_s0_fetch__n_reqs_outstanding;
input logic i_pipeline__i_pipeline_s0_fetch__new_mem_req_t0;
input logic i_pipeline__i_pipeline_s0_fetch__new_mem_req;
input logic i_pipeline__i_pipeline_s0_fetch__progress_imem_addr_t0;
input logic i_pipeline__i_pipeline_s0_fetch__progress_imem_addr;
input logic [2:0] i_pipeline__i_pipeline_s0_fetch__reqs_outstanding_t0;
input logic [2:0] i_pipeline__i_pipeline_s0_fetch__reqs_outstanding;
input logic i_pipeline__i_pipeline_s0_fetch__rsp_recv_t0;
input logic i_pipeline__i_pipeline_s0_fetch__rsp_recv;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__g_clk;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__g_resetn;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__flush;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_4byte;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_2byte;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_err;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_in;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_ready;
input logic [2:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_depth;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_16;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_32;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out_2;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out_4;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_err;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_valid;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_ready;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_16_t0;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_32_t0;
input logic [2:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_depth_t0;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_err_t0;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out_t0;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out_2_t0;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_out_4_t0;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_ready_t0;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buf_valid_t0;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_2byte_t0;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_4byte_t0;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_err_t0;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_in_t0;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__f_ready_t0;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__flush_t0;
input logic [3:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buffer_err_t0;
input logic [3:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buffer_err;
input logic [63:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buffer_t0;
input logic [63:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__buffer;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__eat_2_t0;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__eat_2;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__eat_4_t0;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__eat_4;
input logic [2:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__insert_at_t0;
input logic [2:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__insert_at;
input logic [2:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_bdepth_t0;
input logic [2:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_bdepth;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_d_t0;
input logic [31:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_d;
input logic [3:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_err_t0;
input logic [3:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_err;
input logic [63:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_or_in_t0;
input logic [63:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_or_in;
input logic [63:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_shf_out_t0;
input logic [63:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_shf_out;
input logic [63:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer_t0;
input logic [63:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_buffer;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_err_in_t0;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_err_in;
input logic [3:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_err_or_in_t0;
input logic [3:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_err_or_in;
input logic [3:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_err_shf_out_t0;
input logic [3:0] i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__n_err_shf_out;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__update_buffer_t0;
input logic i_pipeline__i_pipeline_s0_fetch__i_core_fetch_buffer__update_buffer;
input logic i_pipeline__i_pipeline_s1_decode__g_clk;
input logic i_pipeline__i_pipeline_s1_decode__g_resetn;
input logic i_pipeline__i_pipeline_s1_decode__s1_valid;
input logic i_pipeline__i_pipeline_s1_decode__s1_busy;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s1_data;
input logic i_pipeline__i_pipeline_s1_decode__s1_error;
input logic i_pipeline__i_pipeline_s1_decode__s1_flush;
input logic i_pipeline__i_pipeline_s1_decode__s1_bubble;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__s1_rs1_addr;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__s1_rs2_addr;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__s1_rs3_addr;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s1_rs1_rdata;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s1_rs2_rdata;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s1_rs3_rdata;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__leak_prng;
input logic [12:0] i_pipeline__i_pipeline_s1_decode__leak_lkgcfg;
input logic i_pipeline__i_pipeline_s1_decode__s1_leak_fence;
input logic i_pipeline__i_pipeline_s1_decode__cf_req;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__cf_target;
input logic i_pipeline__i_pipeline_s1_decode__cf_ack;
input logic i_pipeline__i_pipeline_s1_decode__s2_valid;
input logic i_pipeline__i_pipeline_s1_decode__s2_busy;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__s2_rd;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s2_opr_a;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s2_opr_b;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s2_opr_c;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__s2_uop;
input logic [7:0] i_pipeline__i_pipeline_s1_decode__s2_fu;
input logic [2:0] i_pipeline__i_pipeline_s1_decode__s2_pw;
input logic i_pipeline__i_pipeline_s1_decode__s2_trap;
input logic [1:0] i_pipeline__i_pipeline_s1_decode__s2_size;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s2_instr;
input logic i_pipeline__i_pipeline_s1_decode__s2_valid_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__s2_uop_t0;
input logic i_pipeline__i_pipeline_s1_decode__s2_trap_t0;
input logic [1:0] i_pipeline__i_pipeline_s1_decode__s2_size_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__s2_rd_t0;
input logic [2:0] i_pipeline__i_pipeline_s1_decode__s2_pw_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s2_opr_c_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s2_opr_b_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s2_opr_a_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s2_instr_t0;
input logic [7:0] i_pipeline__i_pipeline_s1_decode__s2_fu_t0;
input logic i_pipeline__i_pipeline_s1_decode__s2_busy_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s1_rs3_rdata_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__s1_rs3_addr_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s1_rs2_rdata_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__s1_rs2_addr_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s1_rs1_rdata_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__s1_rs1_addr_t0;
input logic i_pipeline__i_pipeline_s1_decode__s1_leak_fence_t0;
input logic i_pipeline__i_pipeline_s1_decode__s1_flush_t0;
input logic i_pipeline__i_pipeline_s1_decode__s1_bubble_t0;
input logic [12:0] i_pipeline__i_pipeline_s1_decode__leak_lkgcfg_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__leak_prng_t0;
input logic i_pipeline__i_pipeline_s1_decode__s1_valid_t0;
input logic i_pipeline__i_pipeline_s1_decode__s1_error_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s1_data_t0;
input logic i_pipeline__i_pipeline_s1_decode__s1_busy_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__cf_target_t0;
input logic i_pipeline__i_pipeline_s1_decode__cf_req_t0;
input logic i_pipeline__i_pipeline_s1_decode__cf_ack_t0;
input logic i_pipeline__i_pipeline_s1_decode__cfu_no_rd_t0;
input logic i_pipeline__i_pipeline_s1_decode__cfu_no_rd;
input logic i_pipeline__i_pipeline_s1_decode__clr_rd_lsb_t0;
input logic i_pipeline__i_pipeline_s1_decode__clr_rd_lsb;
input logic i_pipeline__i_pipeline_s1_decode__csr_no_read_t0;
input logic i_pipeline__i_pipeline_s1_decode__csr_no_read;
input logic i_pipeline__i_pipeline_s1_decode__csr_no_write_t0;
input logic i_pipeline__i_pipeline_s1_decode__csr_no_write;
input logic i_pipeline__i_pipeline_s1_decode__csr_op_t0;
input logic i_pipeline__i_pipeline_s1_decode__csr_op;
input logic i_pipeline__i_pipeline_s1_decode__dec_add_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_add;
input logic i_pipeline__i_pipeline_s1_decode__dec_addi_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_addi;
input logic i_pipeline__i_pipeline_s1_decode__dec_and_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_and;
input logic i_pipeline__i_pipeline_s1_decode__dec_andi_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_andi;
input logic i_pipeline__i_pipeline_s1_decode__dec_auipc_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_auipc;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_bdep_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_bdep;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_bext_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_bext;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_clmul_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_clmul;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_clmulh_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_clmulh;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_clmulr_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_clmulr;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_cmov_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_cmov;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_fsl_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_fsl;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_fsr_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_fsr;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_fsri_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_fsri;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_grev_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_grev;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_grevi_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_grevi;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_ror_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_ror;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_rori_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_b_rori;
input logic i_pipeline__i_pipeline_s1_decode__dec_beq_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_beq;
input logic i_pipeline__i_pipeline_s1_decode__dec_bge_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_bge;
input logic i_pipeline__i_pipeline_s1_decode__dec_bgeu_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_bgeu;
input logic i_pipeline__i_pipeline_s1_decode__dec_blt_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_blt;
input logic i_pipeline__i_pipeline_s1_decode__dec_bltu_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_bltu;
input logic i_pipeline__i_pipeline_s1_decode__dec_bne_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_bne;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_add_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_add;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_addi16sp_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_addi16sp;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_addi4spn_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_addi4spn;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_addi_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_addi;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_and_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_and;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_andi_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_andi;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_beqz_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_beqz;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_bnez_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_bnez;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_ebreak_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_ebreak;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_j_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_j;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_jal_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_jal;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_jalr_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_jalr;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_jr_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_jr;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_li_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_li;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_lui_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_lui;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_lw_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_lw;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_lwsp_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_lwsp;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_mv_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_mv;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_nop_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_nop;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_or_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_or;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_slli_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_slli;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_srai_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_srai;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_srli_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_srli;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_sub_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_sub;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_sw_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_sw;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_swsp_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_swsp;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_xor_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_c_xor;
input logic i_pipeline__i_pipeline_s1_decode__dec_csrrc_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_csrrc;
input logic i_pipeline__i_pipeline_s1_decode__dec_csrrci_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_csrrci;
input logic i_pipeline__i_pipeline_s1_decode__dec_csrrs_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_csrrs;
input logic i_pipeline__i_pipeline_s1_decode__dec_csrrsi_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_csrrsi;
input logic i_pipeline__i_pipeline_s1_decode__dec_csrrw_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_csrrw;
input logic i_pipeline__i_pipeline_s1_decode__dec_csrrwi_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_csrrwi;
input logic i_pipeline__i_pipeline_s1_decode__dec_div_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_div;
input logic i_pipeline__i_pipeline_s1_decode__dec_divu_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_divu;
input logic i_pipeline__i_pipeline_s1_decode__dec_ebreak_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_ebreak;
input logic i_pipeline__i_pipeline_s1_decode__dec_ecall_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_ecall;
input logic i_pipeline__i_pipeline_s1_decode__dec_fence_i_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_fence_i;
input logic i_pipeline__i_pipeline_s1_decode__dec_fence_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_fence;
input logic i_pipeline__i_pipeline_s1_decode__dec_jal_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_jal;
input logic i_pipeline__i_pipeline_s1_decode__dec_jalr_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_jalr;
input logic i_pipeline__i_pipeline_s1_decode__dec_lb_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_lb;
input logic i_pipeline__i_pipeline_s1_decode__dec_lbu_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_lbu;
input logic i_pipeline__i_pipeline_s1_decode__dec_lh_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_lh;
input logic i_pipeline__i_pipeline_s1_decode__dec_lhu_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_lhu;
input logic i_pipeline__i_pipeline_s1_decode__dec_lui_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_lui;
input logic i_pipeline__i_pipeline_s1_decode__dec_lw_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_lw;
input logic i_pipeline__i_pipeline_s1_decode__dec_mret_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_mret;
input logic i_pipeline__i_pipeline_s1_decode__dec_mul_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_mul;
input logic i_pipeline__i_pipeline_s1_decode__dec_mulh_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_mulh;
input logic i_pipeline__i_pipeline_s1_decode__dec_mulhsu_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_mulhsu;
input logic i_pipeline__i_pipeline_s1_decode__dec_mulhu_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_mulhu;
input logic i_pipeline__i_pipeline_s1_decode__dec_or_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_or;
input logic i_pipeline__i_pipeline_s1_decode__dec_ori_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_ori;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__dec_rd_16_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__dec_rd_16;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__dec_rd_32_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__dec_rd_32;
input logic i_pipeline__i_pipeline_s1_decode__dec_rem_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_rem;
input logic i_pipeline__i_pipeline_s1_decode__dec_remu_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_remu;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__dec_rs1_16_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__dec_rs1_16;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__dec_rs2_16_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__dec_rs2_16;
input logic i_pipeline__i_pipeline_s1_decode__dec_sb_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_sb;
input logic i_pipeline__i_pipeline_s1_decode__dec_sh_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_sh;
input logic i_pipeline__i_pipeline_s1_decode__dec_sll_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_sll;
input logic i_pipeline__i_pipeline_s1_decode__dec_slli_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_slli;
input logic i_pipeline__i_pipeline_s1_decode__dec_slt_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_slt;
input logic i_pipeline__i_pipeline_s1_decode__dec_slti_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_slti;
input logic i_pipeline__i_pipeline_s1_decode__dec_sltiu_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_sltiu;
input logic i_pipeline__i_pipeline_s1_decode__dec_sltu_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_sltu;
input logic i_pipeline__i_pipeline_s1_decode__dec_sra_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_sra;
input logic i_pipeline__i_pipeline_s1_decode__dec_srai_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_srai;
input logic i_pipeline__i_pipeline_s1_decode__dec_srl_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_srl;
input logic i_pipeline__i_pipeline_s1_decode__dec_srli_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_srli;
input logic i_pipeline__i_pipeline_s1_decode__dec_sub_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_sub;
input logic i_pipeline__i_pipeline_s1_decode__dec_sw_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_sw;
input logic i_pipeline__i_pipeline_s1_decode__dec_wfi_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_wfi;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_aesmix_dec_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_aesmix_dec;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_aesmix_enc_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_aesmix_enc;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_dec_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_dec;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_decrot_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_decrot;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_enc_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_enc;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_encrot_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_aessub_encrot;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_bop_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_bop;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_b_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_b;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_bu_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_bu;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_h_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_h;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_hu_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_hu;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_w_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_ldr_w;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_lkgfence_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_lkgfence;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_lut_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_lut;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_macc_1_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_macc_1;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_madd_3_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_madd_3;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_mmul_3_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_mmul_3;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_mror_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_mror;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_msub_3_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_msub_3;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_padd_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_padd;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_pclmul_h_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_pclmul_h;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_pclmul_l_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_pclmul_l;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_pmul_h_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_pmul_h;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_pmul_l_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_pmul_l;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_pror_i_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_pror_i;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_pror_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_pror;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_psll_i_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_psll_i;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_psll_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_psll;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_psrl_i_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_psrl_i;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_psrl_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_psrl;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_psub_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_psub;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_rngsamp_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_rngsamp;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_rngseed_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_rngseed;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_rngtest_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_rngtest;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s0_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s1_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s1;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s2_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s2;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s3_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha256_s3;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_x1_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_x1;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_x2_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_x2;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_x4_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_x4;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_xy_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_xy;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_yx_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_sha3_yx;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_str_b_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_str_b;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_str_h_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_str_h;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_str_w_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xc_str_w;
input logic i_pipeline__i_pipeline_s1_decode__dec_xor_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xor;
input logic i_pipeline__i_pipeline_s1_decode__dec_xori_t0;
input logic i_pipeline__i_pipeline_s1_decode__dec_xori;
input logic i_pipeline__i_pipeline_s1_decode__instr_16bit_t0;
input logic i_pipeline__i_pipeline_s1_decode__instr_16bit;
input logic i_pipeline__i_pipeline_s1_decode__invalid_instr_t0;
input logic i_pipeline__i_pipeline_s1_decode__invalid_instr;
input logic i_pipeline__i_pipeline_s1_decode__leak_stall_t0;
input logic i_pipeline__i_pipeline_s1_decode__leak_stall;
input logic i_pipeline__i_pipeline_s1_decode__lf_count_ld_t0;
input logic i_pipeline__i_pipeline_s1_decode__lf_count_ld;
input logic [1:0] i_pipeline__i_pipeline_s1_decode__lf_count_t0;
input logic [1:0] i_pipeline__i_pipeline_s1_decode__lf_count;
input logic i_pipeline__i_pipeline_s1_decode__lsu_no_rd_t0;
input logic i_pipeline__i_pipeline_s1_decode__lsu_no_rd;
input logic [1:0] i_pipeline__i_pipeline_s1_decode__lsu_width_t0;
input logic [1:0] i_pipeline__i_pipeline_s1_decode__lsu_width;
input logic [1:0] i_pipeline__i_pipeline_s1_decode__n_lf_count_t0;
input logic [1:0] i_pipeline__i_pipeline_s1_decode__n_lf_count;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__n_program_counter_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__n_program_counter;
input logic [7:0] i_pipeline__i_pipeline_s1_decode__n_s2_fu_t0;
input logic [7:0] i_pipeline__i_pipeline_s1_decode__n_s2_fu;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__n_s2_imm_pc_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__n_s2_imm_pc;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__n_s2_imm_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__n_s2_imm;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__n_s2_instr_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__n_s2_instr;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__n_s2_opr_a_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__n_s2_opr_a;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__n_s2_opr_b_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__n_s2_opr_b;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__n_s2_opr_c_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__n_s2_opr_c;
input logic [2:0] i_pipeline__i_pipeline_s1_decode__n_s2_pw_t0;
input logic [2:0] i_pipeline__i_pipeline_s1_decode__n_s2_pw;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__n_s2_rd_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__n_s2_rd;
input logic i_pipeline__i_pipeline_s1_decode__n_s2_trap_t0;
input logic i_pipeline__i_pipeline_s1_decode__n_s2_trap;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__n_s2_uop_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__n_s2_uop;
input logic i_pipeline__i_pipeline_s1_decode__n_s2_valid_t0;
input logic i_pipeline__i_pipeline_s1_decode__n_s2_valid;
input logic i_pipeline__i_pipeline_s1_decode__opra_flush_t0;
input logic i_pipeline__i_pipeline_s1_decode__opra_flush;
input logic i_pipeline__i_pipeline_s1_decode__opra_ld_en_t0;
input logic i_pipeline__i_pipeline_s1_decode__opra_ld_en;
input logic i_pipeline__i_pipeline_s1_decode__opra_src_csri_t0;
input logic i_pipeline__i_pipeline_s1_decode__opra_src_csri;
input logic i_pipeline__i_pipeline_s1_decode__opra_src_rs1_t0;
input logic i_pipeline__i_pipeline_s1_decode__opra_src_rs1;
input logic i_pipeline__i_pipeline_s1_decode__opra_src_zero_t0;
input logic i_pipeline__i_pipeline_s1_decode__opra_src_zero;
input logic i_pipeline__i_pipeline_s1_decode__oprb_flush_t0;
input logic i_pipeline__i_pipeline_s1_decode__oprb_flush;
input logic i_pipeline__i_pipeline_s1_decode__oprb_ld_en_t0;
input logic i_pipeline__i_pipeline_s1_decode__oprb_ld_en;
input logic i_pipeline__i_pipeline_s1_decode__oprb_rs2_shf_1_t0;
input logic i_pipeline__i_pipeline_s1_decode__oprb_rs2_shf_1;
input logic i_pipeline__i_pipeline_s1_decode__oprb_rs2_shf_2_t0;
input logic i_pipeline__i_pipeline_s1_decode__oprb_rs2_shf_2;
input logic i_pipeline__i_pipeline_s1_decode__oprb_src_imm_t0;
input logic i_pipeline__i_pipeline_s1_decode__oprb_src_imm;
input logic i_pipeline__i_pipeline_s1_decode__oprb_src_rs2_t0;
input logic i_pipeline__i_pipeline_s1_decode__oprb_src_rs2;
input logic i_pipeline__i_pipeline_s1_decode__oprb_src_zero_t0;
input logic i_pipeline__i_pipeline_s1_decode__oprb_src_zero;
input logic i_pipeline__i_pipeline_s1_decode__oprc_flush_t0;
input logic i_pipeline__i_pipeline_s1_decode__oprc_flush;
input logic i_pipeline__i_pipeline_s1_decode__oprc_ld_en_t0;
input logic i_pipeline__i_pipeline_s1_decode__oprc_ld_en;
input logic i_pipeline__i_pipeline_s1_decode__oprc_src_pcim_t0;
input logic i_pipeline__i_pipeline_s1_decode__oprc_src_pcim;
input logic i_pipeline__i_pipeline_s1_decode__oprc_src_rs2_t0;
input logic i_pipeline__i_pipeline_s1_decode__oprc_src_rs2;
input logic i_pipeline__i_pipeline_s1_decode__oprc_src_rs3_t0;
input logic i_pipeline__i_pipeline_s1_decode__oprc_src_rs3;
input logic [55:0] i_pipeline__i_pipeline_s1_decode__p_in_t0;
input logic [55:0] i_pipeline__i_pipeline_s1_decode__p_in;
input logic [55:0] i_pipeline__i_pipeline_s1_decode__p_mr_t0;
input logic [55:0] i_pipeline__i_pipeline_s1_decode__p_mr;
input logic [55:0] i_pipeline__i_pipeline_s1_decode__p_out_t0;
input logic [55:0] i_pipeline__i_pipeline_s1_decode__p_out;
input logic i_pipeline__i_pipeline_s1_decode__p_s2_busy_t0;
input logic i_pipeline__i_pipeline_s1_decode__p_s2_busy;
input logic i_pipeline__i_pipeline_s1_decode__packed_instruction_t0;
input logic i_pipeline__i_pipeline_s1_decode__packed_instruction;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__pc_plus_imm_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__pc_plus_imm;
input logic i_pipeline__i_pipeline_s1_decode__pipe_progress_t0;
input logic i_pipeline__i_pipeline_s1_decode__pipe_progress;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__program_counter_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__program_counter;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s1_rs2_shf_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__s1_rs2_shf;
input logic [5:0] i_pipeline__i_pipeline_s1_decode__trap_cause_t0;
input logic [5:0] i_pipeline__i_pipeline_s1_decode__trap_cause;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__uop_alu_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__uop_alu;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__uop_asi_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__uop_asi;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__uop_bit_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__uop_bit;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__uop_cfu_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__uop_cfu;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__uop_csr_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__uop_csr;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__uop_lsu_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__uop_lsu;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__uop_mul_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__uop_mul;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__uop_rng_t0;
input logic [4:0] i_pipeline__i_pipeline_s1_decode__uop_rng;
input logic i_pipeline__i_pipeline_s1_decode__use_imm32_b_t0;
input logic i_pipeline__i_pipeline_s1_decode__use_imm32_b;
input logic i_pipeline__i_pipeline_s1_decode__use_imm32_i_t0;
input logic i_pipeline__i_pipeline_s1_decode__use_imm32_i;
input logic i_pipeline__i_pipeline_s1_decode__use_imm32_s_t0;
input logic i_pipeline__i_pipeline_s1_decode__use_imm32_s;
input logic i_pipeline__i_pipeline_s1_decode__use_imm32_u_t0;
input logic i_pipeline__i_pipeline_s1_decode__use_imm32_u;
input logic i_pipeline__i_pipeline_s1_decode__use_imm_csr_t0;
input logic i_pipeline__i_pipeline_s1_decode__use_imm_csr;
input logic i_pipeline__i_pipeline_s1_decode__use_imm_sha3_t0;
input logic i_pipeline__i_pipeline_s1_decode__use_imm_sha3;
input logic i_pipeline__i_pipeline_s1_decode__use_imm_shfi_t0;
input logic i_pipeline__i_pipeline_s1_decode__use_imm_shfi;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__g_clk;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__g_resetn;
input logic [55:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_data;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_valid;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_busy;
input logic [55:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__mr_data;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__flush;
input logic [55:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__flush_dat;
input logic [55:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_data;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_valid;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_busy;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__flush_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_valid_t0;
input logic [55:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_data_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__o_busy_t0;
input logic [55:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__mr_data_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_valid_t0;
input logic [55:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_data_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__i_busy_t0;
input logic [55:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__flush_dat_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__genblk1__progress_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg__genblk1__progress;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__g_clk;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__g_resetn;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_data;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_valid;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_busy;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__mr_data;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__flush;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__flush_dat;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_data;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_valid;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_busy;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__flush_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_data_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__o_busy_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__mr_data_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_data_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__i_busy_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__flush_dat_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__genblk1__progress_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_a__genblk1__progress;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__g_clk;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__g_resetn;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_data;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_valid;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_busy;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__mr_data;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__flush;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__flush_dat;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_data;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_valid;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_busy;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__flush_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_data_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__o_busy_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__mr_data_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_data_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__i_busy_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__flush_dat_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__genblk1__progress_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_b__genblk1__progress;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__g_clk;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__g_resetn;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_data;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_valid;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_busy;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__mr_data;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__flush;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__flush_dat;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_data;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_valid;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_busy;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__flush_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_data_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__o_busy_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__mr_data_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_data_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__i_busy_t0;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__flush_dat_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__genblk1__progress_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_decode_pipereg_opr_c__genblk1__progress;
input logic i_pipeline__i_pipeline_s1_decode__i_frv_leak__g_clk;
input logic i_pipeline__i_pipeline_s1_decode__i_frv_leak__g_resetn;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_frv_leak__leak_prng;
input logic i_pipeline__i_pipeline_s1_decode__i_frv_leak__leak_fence;
input logic [31:0] i_pipeline__i_pipeline_s1_decode__i_frv_leak__leak_prng_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_frv_leak__leak_fence_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_frv_leak__genblk1__genblk1__n_prng_lsb_t0;
input logic i_pipeline__i_pipeline_s1_decode__i_frv_leak__genblk1__genblk1__n_prng_lsb;
input logic i_pipeline__i_pipeline_s2_execute__g_clk;
input logic i_pipeline__i_pipeline_s2_execute__g_resetn;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__s2_rd;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__s2_opr_a;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__s2_opr_b;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__s2_opr_c;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__s2_uop;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__s2_fu;
input logic [2:0] i_pipeline__i_pipeline_s2_execute__s2_pw;
input logic i_pipeline__i_pipeline_s2_execute__s2_trap;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__s2_size;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__s2_instr;
input logic i_pipeline__i_pipeline_s2_execute__s2_busy;
input logic i_pipeline__i_pipeline_s2_execute__s2_valid;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__leak_prng;
input logic [12:0] i_pipeline__i_pipeline_s2_execute__leak_lkgcfg;
input logic i_pipeline__i_pipeline_s2_execute__rng_req_valid;
input logic [2:0] i_pipeline__i_pipeline_s2_execute__rng_req_op;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__rng_req_data;
input logic i_pipeline__i_pipeline_s2_execute__rng_req_ready;
input logic i_pipeline__i_pipeline_s2_execute__rng_rsp_valid;
input logic [2:0] i_pipeline__i_pipeline_s2_execute__rng_rsp_status;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__rng_rsp_data;
input logic i_pipeline__i_pipeline_s2_execute__rng_rsp_ready;
input logic i_pipeline__i_pipeline_s2_execute__uxcrypto_ct;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__uxcrypto_b0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__uxcrypto_b1;
input logic i_pipeline__i_pipeline_s2_execute__flush;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__fwd_s2_rd;
input logic i_pipeline__i_pipeline_s2_execute__fwd_s2_wide;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__fwd_s2_wdata;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__fwd_s2_wdata_hi;
input logic i_pipeline__i_pipeline_s2_execute__fwd_s2_load;
input logic i_pipeline__i_pipeline_s2_execute__fwd_s2_csr;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__s3_rd;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__s3_opr_a;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__s3_opr_b;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__s3_uop;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__s3_fu;
input logic i_pipeline__i_pipeline_s2_execute__s3_trap;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__s3_size;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__s3_instr;
input logic i_pipeline__i_pipeline_s2_execute__s3_busy;
input logic i_pipeline__i_pipeline_s2_execute__s3_valid;
input logic i_pipeline__i_pipeline_s2_execute__flush_t0;
input logic i_pipeline__i_pipeline_s2_execute__s2_valid_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__s2_uop_t0;
input logic i_pipeline__i_pipeline_s2_execute__s2_trap_t0;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__s2_size_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__s2_rd_t0;
input logic [2:0] i_pipeline__i_pipeline_s2_execute__s2_pw_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__s2_opr_c_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__s2_opr_b_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__s2_opr_a_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__s2_instr_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__s2_fu_t0;
input logic i_pipeline__i_pipeline_s2_execute__s2_busy_t0;
input logic [12:0] i_pipeline__i_pipeline_s2_execute__leak_lkgcfg_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__leak_prng_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__rng_req_data_t0;
input logic [2:0] i_pipeline__i_pipeline_s2_execute__rng_req_op_t0;
input logic i_pipeline__i_pipeline_s2_execute__rng_req_ready_t0;
input logic i_pipeline__i_pipeline_s2_execute__rng_req_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__rng_rsp_data_t0;
input logic i_pipeline__i_pipeline_s2_execute__rng_rsp_ready_t0;
input logic [2:0] i_pipeline__i_pipeline_s2_execute__rng_rsp_status_t0;
input logic i_pipeline__i_pipeline_s2_execute__rng_rsp_valid_t0;
input logic i_pipeline__i_pipeline_s2_execute__fwd_s2_csr_t0;
input logic i_pipeline__i_pipeline_s2_execute__fwd_s2_load_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__fwd_s2_rd_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__fwd_s2_wdata_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__fwd_s2_wdata_hi_t0;
input logic i_pipeline__i_pipeline_s2_execute__fwd_s2_wide_t0;
input logic i_pipeline__i_pipeline_s2_execute__s3_busy_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__s3_fu_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__s3_instr_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__s3_opr_a_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__s3_opr_b_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__s3_rd_t0;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__s3_size_t0;
input logic i_pipeline__i_pipeline_s2_execute__s3_trap_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__s3_uop_t0;
input logic i_pipeline__i_pipeline_s2_execute__s3_valid_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__uxcrypto_b0_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__uxcrypto_b1_t0;
input logic i_pipeline__i_pipeline_s2_execute__uxcrypto_ct_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__alu_add_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__alu_add_result;
input logic i_pipeline__i_pipeline_s2_execute__alu_eq_t0;
input logic i_pipeline__i_pipeline_s2_execute__alu_eq;
input logic i_pipeline__i_pipeline_s2_execute__alu_lt_t0;
input logic i_pipeline__i_pipeline_s2_execute__alu_lt;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_add_t0;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_add;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_and_t0;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_and;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_cmp_t0;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_cmp;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_or_t0;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_or;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_rot_t0;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_rot;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_shf_arith_t0;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_shf_arith;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_shf_left_t0;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_shf_left;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_shf_t0;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_shf;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_sub_t0;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_sub;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_unsigned_t0;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_unsigned;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_xor_t0;
input logic i_pipeline__i_pipeline_s2_execute__alu_op_xor;
input logic i_pipeline__i_pipeline_s2_execute__alu_ready_t0;
input logic i_pipeline__i_pipeline_s2_execute__alu_ready;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__alu_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__alu_result;
input logic i_pipeline__i_pipeline_s2_execute__asi_done_t0;
input logic i_pipeline__i_pipeline_s2_execute__asi_done;
input logic i_pipeline__i_pipeline_s2_execute__asi_finished_t0;
input logic i_pipeline__i_pipeline_s2_execute__asi_finished;
input logic i_pipeline__i_pipeline_s2_execute__asi_flush_aesmix_t0;
input logic i_pipeline__i_pipeline_s2_execute__asi_flush_aesmix;
input logic i_pipeline__i_pipeline_s2_execute__asi_flush_aessub_t0;
input logic i_pipeline__i_pipeline_s2_execute__asi_flush_aessub;
input logic i_pipeline__i_pipeline_s2_execute__asi_ready_t0;
input logic i_pipeline__i_pipeline_s2_execute__asi_ready;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__asi_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__asi_result;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__bitw_bop_lut_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__bitw_bop_lut;
input logic i_pipeline__i_pipeline_s2_execute__bitw_bop_t0;
input logic i_pipeline__i_pipeline_s2_execute__bitw_bop;
input logic i_pipeline__i_pipeline_s2_execute__bitw_cmov_t0;
input logic i_pipeline__i_pipeline_s2_execute__bitw_cmov;
input logic i_pipeline__i_pipeline_s2_execute__bitw_flush_t0;
input logic i_pipeline__i_pipeline_s2_execute__bitw_flush;
input logic i_pipeline__i_pipeline_s2_execute__bitw_fsl_t0;
input logic i_pipeline__i_pipeline_s2_execute__bitw_fsl;
input logic i_pipeline__i_pipeline_s2_execute__bitw_fsr_t0;
input logic i_pipeline__i_pipeline_s2_execute__bitw_fsr;
input logic i_pipeline__i_pipeline_s2_execute__bitw_gpr_wide_t0;
input logic i_pipeline__i_pipeline_s2_execute__bitw_gpr_wide;
input logic i_pipeline__i_pipeline_s2_execute__bitw_lut_t0;
input logic i_pipeline__i_pipeline_s2_execute__bitw_lut;
input logic i_pipeline__i_pipeline_s2_execute__bitw_ready_t0;
input logic i_pipeline__i_pipeline_s2_execute__bitw_ready;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__bitw_result_wide_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__bitw_result_wide;
input logic i_pipeline__i_pipeline_s2_execute__cfu_cond_t0;
input logic i_pipeline__i_pipeline_s2_execute__cfu_cond;
input logic i_pipeline__i_pipeline_s2_execute__cfu_cond_taken_t0;
input logic i_pipeline__i_pipeline_s2_execute__cfu_cond_taken;
input logic i_pipeline__i_pipeline_s2_execute__cfu_jalr_t0;
input logic i_pipeline__i_pipeline_s2_execute__cfu_jalr;
input logic i_pipeline__i_pipeline_s2_execute__cond_beq_t0;
input logic i_pipeline__i_pipeline_s2_execute__cond_beq;
input logic i_pipeline__i_pipeline_s2_execute__cond_bge_t0;
input logic i_pipeline__i_pipeline_s2_execute__cond_bge;
input logic i_pipeline__i_pipeline_s2_execute__cond_bgeu_t0;
input logic i_pipeline__i_pipeline_s2_execute__cond_bgeu;
input logic i_pipeline__i_pipeline_s2_execute__cond_blt_t0;
input logic i_pipeline__i_pipeline_s2_execute__cond_blt;
input logic i_pipeline__i_pipeline_s2_execute__cond_bltu_t0;
input logic i_pipeline__i_pipeline_s2_execute__cond_bltu;
input logic i_pipeline__i_pipeline_s2_execute__cond_bne_t0;
input logic i_pipeline__i_pipeline_s2_execute__cond_bne;
input logic i_pipeline__i_pipeline_s2_execute__imul_clmul_r_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_clmul_r;
input logic i_pipeline__i_pipeline_s2_execute__imul_clmul_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_clmul;
input logic i_pipeline__i_pipeline_s2_execute__imul_div_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_div;
input logic i_pipeline__i_pipeline_s2_execute__imul_divu_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_divu;
input logic i_pipeline__i_pipeline_s2_execute__imul_flush_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_flush;
input logic i_pipeline__i_pipeline_s2_execute__imul_gpr_wide_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_gpr_wide;
input logic i_pipeline__i_pipeline_s2_execute__imul_macc_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_macc;
input logic i_pipeline__i_pipeline_s2_execute__imul_madd_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_madd;
input logic i_pipeline__i_pipeline_s2_execute__imul_mmul_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_mmul;
input logic i_pipeline__i_pipeline_s2_execute__imul_msub_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_msub;
input logic i_pipeline__i_pipeline_s2_execute__imul_mul_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_mul;
input logic i_pipeline__i_pipeline_s2_execute__imul_mulhsu_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_mulhsu;
input logic i_pipeline__i_pipeline_s2_execute__imul_mulhu_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_mulhu;
input logic i_pipeline__i_pipeline_s2_execute__imul_pclmul_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_pclmul;
input logic i_pipeline__i_pipeline_s2_execute__imul_pmul_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_pmul;
input logic i_pipeline__i_pipeline_s2_execute__imul_pw_16_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_pw_16;
input logic i_pipeline__i_pipeline_s2_execute__imul_pw_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_pw_2;
input logic i_pipeline__i_pipeline_s2_execute__imul_pw_32_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_pw_32;
input logic i_pipeline__i_pipeline_s2_execute__imul_pw_4_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_pw_4;
input logic i_pipeline__i_pipeline_s2_execute__imul_pw_8_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_pw_8;
input logic i_pipeline__i_pipeline_s2_execute__imul_ready_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_ready;
input logic i_pipeline__i_pipeline_s2_execute__imul_rem_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_rem;
input logic i_pipeline__i_pipeline_s2_execute__imul_remu_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_remu;
input logic i_pipeline__i_pipeline_s2_execute__imul_result_hi_t0;
input logic i_pipeline__i_pipeline_s2_execute__imul_result_hi;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__imul_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__imul_result;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__imul_result_wide_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__imul_result_wide;
input logic i_pipeline__i_pipeline_s2_execute__leak_fence_t0;
input logic i_pipeline__i_pipeline_s2_execute__leak_fence;
input logic i_pipeline__i_pipeline_s2_execute__lsu_load_t0;
input logic i_pipeline__i_pipeline_s2_execute__lsu_load;
input logic i_pipeline__i_pipeline_s2_execute__lsu_store_t0;
input logic i_pipeline__i_pipeline_s2_execute__lsu_store;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_cfu_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_cfu;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_mul_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_mul;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_rng_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__n_s3_opr_a_rng;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__n_s3_opr_b_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__n_s3_opr_b;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__n_s3_uop_cfu_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__n_s3_uop_cfu;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__n_s3_uop_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__n_s3_uop;
input logic i_pipeline__i_pipeline_s2_execute__opra_flush_t0;
input logic i_pipeline__i_pipeline_s2_execute__opra_flush;
input logic i_pipeline__i_pipeline_s2_execute__opra_ld_en_t0;
input logic i_pipeline__i_pipeline_s2_execute__opra_ld_en;
input logic i_pipeline__i_pipeline_s2_execute__oprb_flush_t0;
input logic i_pipeline__i_pipeline_s2_execute__oprb_flush;
input logic i_pipeline__i_pipeline_s2_execute__oprb_ld_en_t0;
input logic i_pipeline__i_pipeline_s2_execute__oprb_ld_en;
input logic i_pipeline__i_pipeline_s2_execute__p_busy_t0;
input logic i_pipeline__i_pipeline_s2_execute__p_busy;
input logic i_pipeline__i_pipeline_s2_execute__p_valid_t0;
input logic i_pipeline__i_pipeline_s2_execute__p_valid;
input logic [52:0] i_pipeline__i_pipeline_s2_execute__pipe_reg_out_t0;
input logic [52:0] i_pipeline__i_pipeline_s2_execute__pipe_reg_out;
input logic i_pipeline__i_pipeline_s2_execute__rng_if_ready_t0;
input logic i_pipeline__i_pipeline_s2_execute__rng_if_ready;
input logic i_pipeline__i_pipeline_s2_execute__rng_ready_t0;
input logic i_pipeline__i_pipeline_s2_execute__rng_ready;
input logic i_pipeline__i_pipeline_s2_execute__rng_uop_samp_t0;
input logic i_pipeline__i_pipeline_s2_execute__rng_uop_samp;
input logic i_pipeline__i_pipeline_s2_execute__rng_uop_seed_t0;
input logic i_pipeline__i_pipeline_s2_execute__rng_uop_seed;
input logic i_pipeline__i_pipeline_s2_execute__rng_uop_test_t0;
input logic i_pipeline__i_pipeline_s2_execute__rng_uop_test;
input logic i_pipeline__i_pipeline_s2_execute__rng_valid_t0;
input logic i_pipeline__i_pipeline_s2_execute__rng_valid;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__g_clk;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__g_resetn;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_valid;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_flush;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_ready;
input logic [2:0] i_pipeline__i_pipeline_s2_execute__i_alu__alu_pw;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_add;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_sub;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_xor;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_or;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_and;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_rot;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf_left;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf_arith;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_cmp;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_unsigned;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_lt;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_eq;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__alu_add_result;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__alu_lhs;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__alu_rhs;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__alu_result;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__alu_add_result_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_eq_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_flush_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__alu_lhs_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_lt_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_add_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_and_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_cmp_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_or_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_rot_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf_arith_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_shf_left_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_sub_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_unsigned_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_op_xor_t0;
input logic [2:0] i_pipeline__i_pipeline_s2_execute__i_alu__alu_pw_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_ready_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__alu_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__alu_rhs_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_valid_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_lt_signed_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_lt_signed;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_lt_unsigned_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__alu_lt_unsigned;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__bw_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__bw_result;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__out_adder_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__out_adder;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__out_bw_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__out_bw;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__out_shift_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__out_shift;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_alu__pw_d_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_alu__pw_d;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__shift_arith_mask_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__shift_arith_mask;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__shift_arith_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__shift_arith;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__shift_out_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__shift_out;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__shift_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__shift_result;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__lhs;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__rhs;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__pw;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__cin;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__sub;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__c_en;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__c_out;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__result;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__c_en_t0;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__c_out_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__cin_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__lhs_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__pw_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__rhs_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__sub_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__carry_mask_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__carry_mask;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_0___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_0___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_0___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_0___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_10___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_10___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_10___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_10___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_11___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_11___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_11___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_11___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_11___force_carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_11___force_carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_12___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_12___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_12___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_12___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_13___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_13___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_13___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_13___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_13___force_carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_13___force_carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_14___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_14___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_14___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_14___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_15___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_15___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_15___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_15___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_15___force_carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_15___force_carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_16___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_16___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_16___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_16___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_17___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_17___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_17___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_17___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_18___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_18___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_18___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_18___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_19___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_19___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_19___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_19___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_1___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_1___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_1___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_1___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_20___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_20___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_20___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_20___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_21___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_21___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_21___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_21___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_22___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_22___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_22___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_22___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_23___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_23___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_23___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_23___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_23___force_carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_23___force_carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_24___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_24___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_24___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_24___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_25___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_25___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_25___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_25___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_26___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_26___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_26___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_26___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_27___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_27___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_27___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_27___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_28___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_28___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_28___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_28___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_29___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_29___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_29___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_29___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_2___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_2___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_2___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_2___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_30___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_30___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_30___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_30___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_31___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_31___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_31___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_31___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_3___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_3___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_3___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_3___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_4___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_4___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_4___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_4___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_5___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_5___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_5___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_5___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_6___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_6___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_6___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_6___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_7___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_7___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_7___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_7___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_8___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_8___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_8___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_8___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_9___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_9___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_9___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__genblk1_9___carry;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__rhs_m_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_addsub__rhs_m;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__crs1;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__shamt;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__pw;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__shift;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__rotate;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__left;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__right;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__result;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__pw_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__crs1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__left_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__right_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__rotate_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__shamt_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__shift_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_16_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_16;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_32_left_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_32_left;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_32_right_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l16_32_right;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_16_left_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_16_left;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_16_right_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_16_right;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_2_left_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_2_left;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_2_right_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_2_right;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_16_left_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_16_left;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_16_right_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_16_right;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_2_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_2;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_4_left_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_4_left;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_4_right_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_4_right;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l2;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_16_left_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_16_left;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_16_right_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_16_right;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_2_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_2;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_8_left_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_8_left;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_8_right_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_8_right;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l4;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_16_left_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_16_left;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_16_right_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_16_right;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_2_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_2;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__l8;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_16;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_2;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_32_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_32;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_4;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_l_8;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_16;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_2;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_32_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_32;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_4;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l16_r_8;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_16;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_2;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_32_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_32;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_4;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_l_8;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_16;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_2;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_32_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_32;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_4;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l1_r_8;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_2;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_16;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_32_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_32;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_4;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_l_8;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_16;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_32_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_32;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_4;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l2_r_8;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_16;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_2;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_32_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_32;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_4;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_l_8;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_16;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_2;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_32_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_32;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_4;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l4_r_8;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_16;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_2;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_32_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_32;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_4;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_l_8;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_16;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_2;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_32_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_32;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_4;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_alu__i_p_shfrot__ld_l8_r_8;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__g_clk;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__g_resetn;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__asi_valid;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__asi_ready;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_aessub;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_aesmix;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_data;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_asi__asi_uop;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__asi_rs1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__asi_rs2;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__i_asi__asi_shamt;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__asi_result;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_aesmix_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_aessub_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__asi_flush_data_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__asi_ready_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__asi_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__asi_rs1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__asi_rs2_t0;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__i_asi__asi_shamt_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_asi__asi_uop_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__asi_valid_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_ready_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_ready;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_rs1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_rs1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_rs2_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__aes_mix_rs2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_ready_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_ready;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_rs1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_rs1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_rs2_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__aes_sub_rs2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_aes_mix_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_aes_mix;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_aes_sub_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_aes_sub;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_aes_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_aes;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_x1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_x1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_x2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_x2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_x4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_x4;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_xy_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_xy;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_yx_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__insn_sha3_yx;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__result_aesmix_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__result_aesmix;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__result_aessub_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__result_aessub;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__result_sha2_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__result_sha2;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__result_sha3_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__result_sha3;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__sha2_rs1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__sha2_rs1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__clock;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__reset;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__flush;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__flush_data;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__valid;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__rs1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__rs2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__enc;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__ready;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__result;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__flush_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__result_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__ready_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__rs1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__rs2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__flush_data_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__enc_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d0_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d1_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d1;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d2_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d2;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d3_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__d3;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e0_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e1_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e1;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e2_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e2;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e3_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__e3;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__b_0_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__b_0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__b_1_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__b_1;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__b_2_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__b_2;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__b_3_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__b_3;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_0_lhs_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_0_lhs;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_0_out_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_0_out;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_1_lhs_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_1_lhs;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_1_out_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_1_out;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_2_lhs_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_2_lhs;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_2_out_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_2_out;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_3_lhs_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_3_lhs;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_3_out_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_3_out;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_byte_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__dec_byte;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_byte_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_byte;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x0_in_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x0_in;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x1_in_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x1_in;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x2_in_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x2_in;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x2_out_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x2_out;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x3_in_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x3_in;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x3_out_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__enc_x3_out;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__fsm_0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__fsm_0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__fsm_1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__fsm_1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__fsm_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__fsm_2;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__fsm_t0;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__fsm;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__n_fsm_t0;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aesmix__genblk1__n_fsm;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__clock;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__reset;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__flush;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__flush_data;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__valid;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rs1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rs2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__enc;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rot;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__ready;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__result;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__flush_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__result_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__ready_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rs1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rs2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__flush_data_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__enc_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__rot_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__b_0_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__b_0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__b_1_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__b_1;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__b_2_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__b_2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__fsm_0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__fsm_0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__fsm_1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__fsm_1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__fsm_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__fsm_2;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__fsm_t0;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__fsm;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__n_fsm_t0;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__n_fsm;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_in_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_in;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_out_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_out;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__in;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__inv;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__in_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__inv_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out_fwd_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out_fwd;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out_inv_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__out_inv;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__in;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__out;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__in_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__out_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s4;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s5_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s5;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s6_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s6;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s7_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__s7;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t10_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t10;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t11_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t11;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t12_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t12;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t13_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t13;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t14_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t14;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t15_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t15;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t16;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t17_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t17;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t18_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t18;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t19_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t19;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t20_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t20;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t21_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t21;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t22_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t22;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t23_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t23;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t24_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t24;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t25_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t25;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t26_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t26;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t27_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t27;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t28_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t28;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t29_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t29;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t30_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t30;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t31_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t31;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t32_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t32;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t33_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t33;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t34_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t34;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t35_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t35;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t36_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t36;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t37_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t37;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t38_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t38;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t39_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t39;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t40_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t40;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t41_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t41;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t42_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t42;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t43_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t43;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t44_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t44;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t45_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t45;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t4;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t5_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t5;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t6_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t6;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t7_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t7;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t8;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t9_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__t9;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc10_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc10;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc11_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc11;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc12_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc12;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc13_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc13;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc14_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc14;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc16;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc17_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc17;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc18_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc18;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc20_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc20;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc21_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc21;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc26_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc26;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc4;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc5_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc5;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc6_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc6;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc7_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc7;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc8;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc9_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__tc9;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y10_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y10;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y11_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y11;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y12_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y12;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y13_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y13;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y14_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y14;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y15_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y15;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y16;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y17_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y17;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y18_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y18;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y19_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y19;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y20_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y20;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y21_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y21;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y4;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y5_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y5;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y6_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y6;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y7_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y7;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y8;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y9_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__y9;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z10_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z10;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z11_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z11;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z12_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z12;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z13_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z13;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z14_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z14;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z15_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z15;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z16;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z17_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z17;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z4;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z5_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z5;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z6_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z6;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z7_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z7;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z8;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z9_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_fwd__z9;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__in;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__out;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__in_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__out_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__aa_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__aa;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab20_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab20;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab21_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab21;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab22_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab22;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab23_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab23;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ab3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd4;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd5_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd5;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd6_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__abcd6;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ah_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ah;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__al_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__al;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__bb_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__bb;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__bh_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__bh;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__bl_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__bl;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__cp4;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__d3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__dd_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__dd;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__dh_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__dh;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__dl_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__dl;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p4;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p6_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p6;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p7_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__p7;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph01_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph01;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph02_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph02;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph03_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph03;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph11_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph11;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph12_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph12;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph13_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__ph13;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl01_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl01;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl02_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl02;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl03_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl03;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl11_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl11;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl12_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl12;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl13_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pl13;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pr1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pr1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pr2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pr2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pr3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__pr3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__qr1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__qr1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__qr2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__qr2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__qr3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__qr3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r10_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r10;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r11_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r11;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r4;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r5_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r5;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r6_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r6;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r7_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r7;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r8;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r9_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__r9;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rr1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rr1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rr2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rr2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rtl0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rtl0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rtl1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rtl1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rtl2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__rtl2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s4;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s5_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s5;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s6_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s6;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s7_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__s7;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sa0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sa0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sa1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sa1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sb0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sb0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sb1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sb1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sd0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sd0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sd1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__sd1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__t01_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__t01;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__t02_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__t02;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv10_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv10;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv11_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv11;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv12_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv12;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv13_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv13;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv4;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv5_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv5;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv6_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv6;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv7_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv7;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv8;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv9_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__tinv9;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__vr1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__vr1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__vr2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__vr2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__vr3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__vr3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__wr1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__wr1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__wr2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__wr2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__wr3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__wr3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x11_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x11;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x13_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x13;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x14_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x14;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x16;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x18_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x18;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x19_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__x19;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y3;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y4;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y5_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y5;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y6_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y6;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y7_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_aessub__genblk1__sbox_0__i_sbox_inv__y7;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__rs1;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__ss;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__result;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__rs1_t0;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__ss_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s0_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s0_result;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s1_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s1_result;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s2_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s2_result;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s2;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s3_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s3_result;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha256__s3;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__rs1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__rs2;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shamt;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_xy;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x1;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x2;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x4;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_yx;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__result;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__result_t0;
input logic [1:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shamt_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__rs1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__rs2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_x4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_xy_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__f_yx_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__in_x_plus_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__in_x_plus;
input logic [6:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__in_y_plus_t0;
input logic [6:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__in_y_plus;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_in_lhs_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_in_lhs;
input logic [6:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_in_rhs_t0;
input logic [6:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_in_rhs;
input logic [2:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_out_lhs_t0;
input logic [2:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_out_lhs;
input logic [2:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_out_rhs_t0;
input logic [2:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__lut_out_rhs;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__result_sum_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__result_sum;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shf_1_t0;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shf_1;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shf_2_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__shf_2;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__sum_rhs_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_asi__i_xc_sha3__sum_rhs;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__g_clk;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__g_resetn;
input logic [52:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_data;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_valid;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_busy;
input logic [52:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__mr_data;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__flush;
input logic [52:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__flush_dat;
input logic [52:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_data;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_valid;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_busy;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__flush_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_valid_t0;
input logic [52:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_data_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__o_busy_t0;
input logic [52:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__mr_data_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_valid_t0;
input logic [52:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_data_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__i_busy_t0;
input logic [52:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__flush_dat_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__genblk1__progress_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg__genblk1__progress;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__g_clk;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__g_resetn;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_data;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_valid;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_busy;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__mr_data;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__flush;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__flush_dat;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_data;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_valid;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_busy;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__flush_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_data_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__o_busy_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__mr_data_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_data_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__i_busy_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__flush_dat_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__genblk1__progress_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_a__genblk1__progress;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__g_clk;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__g_resetn;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_data;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_valid;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_busy;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__mr_data;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__flush;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__flush_dat;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_data;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_valid;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_busy;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__flush_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_data_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__o_busy_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__mr_data_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_data_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__i_busy_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__flush_dat_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__genblk1__progress_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_execute_pipe_reg_opr_b__genblk1__progress;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs2;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs3;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__bop_lut;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__flush;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__valid;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_fsl;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_fsr;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_mror;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_cmov;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_lut;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_bop;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__ready;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__flush_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__ready_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rs3_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__bop_lut_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_bop_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_cmov_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_fsl_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_fsr_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_lut_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__uop_mror_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__r_in_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__r_in;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__r_out_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__r_out;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__ramt_t0;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__ramt;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_bop_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_bop;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_cmov_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_cmov;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_fsl_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_fsl;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_lut_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__result_lut;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_0_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_1_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_1;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_2_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_2;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_3_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_3;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_4_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_4;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_5_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rt_5;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rword_l_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__rword_l;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs2;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs3;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__result;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs2_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk2__i_b_lut__crs3_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rd;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rs1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rs2;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__lut;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__result;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rs1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rs2_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__lut_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_bitwise__genblk3__i_b_bop__rd_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__g_clk;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__g_resetn;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__flush;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__pipeline_progress;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__valid;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rs1;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_valid;
input logic [2:0] i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_op;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_data;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_ready;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_valid;
input logic [2:0] i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_status;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_data;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_ready;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_test;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_seed;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_samp;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_rngif__result;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__ready;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__flush_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_rngif__result_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__ready_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rs1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__valid_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__pipeline_progress_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_data_t0;
input logic [2:0] i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_op_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_ready_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_req_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_data_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_ready_t0;
input logic [2:0] i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_status_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__rng_rsp_valid_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_samp_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_seed_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__uop_test_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__n_req_done_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__n_req_done;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__req_done_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__req_done;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__status_healthy_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_frv_rngif__status_healthy;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__clock;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__resetn;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs2;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs3;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__flush;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__flush_data;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__valid;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_div;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_divu;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_rem;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_remu;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mul;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mulu;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mulsu;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_clmul;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_pmul;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_pclmul;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_madd;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_msub;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_macc;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mmul;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_32;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_16;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_8;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_4;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_2;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__result;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__ready;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__flush_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mul_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__result_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_32_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__pw_8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__ready_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__rs3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_macc_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_madd_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mmul_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_msub_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__flush_data_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_clmul_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_div_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_divu_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mulsu_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_mulu_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_pclmul_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_pmul_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_rem_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__uop_remu_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__acc_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__acc;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__arg_0_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__arg_0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__arg_1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__arg_1;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__count_en_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__count_en;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__count_t0;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__count;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__do_mulu_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__do_mulu;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__fsm_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__fsm;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__insn_divrem_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__insn_divrem;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__insn_long_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__insn_long;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__insn_mdr_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__insn_mdr;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__ld_long_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__ld_long;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__ld_mdr_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__ld_mdr;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__ld_on_init_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__ld_on_init;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_n_acc_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_n_acc;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_n_carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_n_carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_cin_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_cin;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_lhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_lhs;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_rhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_rhs;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_sub_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_padd_sub;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_ready_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_ready;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_result_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__long_result;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_acc_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_acc;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_arg_0_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_arg_0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_arg_1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_n_arg_1;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_cen_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_cen;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_cin_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_cin;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_lhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_lhs;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_rhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_rhs;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_sub_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_padd_sub;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_ready_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_ready;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_result_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__mdr_result;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_acc_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_acc;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_arg_0_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_arg_0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_carry;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_count_t0;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_count;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_fsm_t0;
input logic [7:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__n_fsm;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_cen_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_cen;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_cin_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_cin;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_cout_t0;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_cout;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_lhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_lhs;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_result;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_rhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_rhs;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_sub_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__padd_sub;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__reg_ld_en_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__reg_ld_en;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__clock;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__resetn;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs2;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs3;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__flush;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__valid;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_div;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_divu;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_rem;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_remu;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mul;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mulu;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mulsu;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_clmul;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_pmul;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_pclmul;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_32;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_16;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_8;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_4;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_2;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__count;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__acc;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_1;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_acc;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_arg_0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_arg_1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_lhs;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_rhs;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_sub;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cin;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cen;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cout;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_result;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__result;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__ready;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__flush_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__result_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__acc_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_0_t0;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__count_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_acc_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_arg_0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cen_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cin_t0;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_cout_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_lhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_rhs_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__padd_sub_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_32_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pw_8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__ready_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs2_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__n_arg_1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__valid_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_clmul_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_div_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_divu_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mul_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mulsu_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_mulu_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_pclmul_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_pmul_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_rem_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__do_remu_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rs3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_sel_neg_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_sel_neg;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_sel_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__arg_sel;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_n_acc_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_n_acc;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_n_arg_0_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_n_arg_0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_outsign_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_outsign;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_ready_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_ready;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_signed_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__div_signed;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__divrem_result_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__divrem_result;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_carryless_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_carryless;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_lhs_sign_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_lhs_sign;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_n_acc_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_n_acc;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_n_arg_0_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_n_arg_0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_cen_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_cen;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_cin_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_cin;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_lhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_lhs;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_rhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_rhs;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_sub_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_padd_sub;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_ready_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__mul_ready;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_n_acc_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_n_acc;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_n_arg_0_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_n_arg_0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_cen_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_cen;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_lhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_lhs;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_rhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_rhs;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_sub_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_padd_sub;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_ready_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_ready;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_result_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__pmul_result;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rem_outsign_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__rem_outsign;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__result_div_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__result_div;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__result_rem_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__result_rem;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__route_div_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__route_div;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__route_mul_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__route_mul;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__route_pmul_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__route_pmul;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__rs1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__rs2;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__count;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__acc;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__arg_0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__carryless;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_16;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_8;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_4;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_2;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_lhs;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_rhs;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_sub;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_cen;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_cout;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_result;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__n_acc;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__n_arg_0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__result;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__ready;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__result_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__acc_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__arg_0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__carryless_t0;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__count_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__n_acc_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__n_arg_0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_cen_t0;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_cout_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_lhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_rhs_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_sub_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pw_8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__ready_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__rs1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__rs2_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_mask_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__padd_mask;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pmul_result_0_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_malu_pmul__pmul_result_0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__clock;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__resetn;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__rs1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__rs2;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__valid;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__op_signed;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__flush;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__count;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__acc;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__arg_0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__arg_1;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_acc;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_arg_0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_arg_1;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__ready;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__flush_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__acc_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__arg_0_t0;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__count_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_acc_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_arg_0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__ready_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__rs1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__rs2_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__arg_1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__n_arg_1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__op_signed_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__valid_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__div_less_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__div_less;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__div_run_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__div_run;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__div_start_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__div_start;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__divisor_start_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__divisor_start;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__qmask_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__qmask;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__signed_lhs_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__signed_lhs;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__signed_rhs_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__signed_rhs;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__sub_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_divrem__sub_result;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rs1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rs2;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__count;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__acc;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__arg_0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__carryless;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_32;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_16;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_8;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_4;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_2;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__lhs_sign;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rhs_sign;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_lhs;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_rhs;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_sub;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cin;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cen;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cout;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_result;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__n_acc;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__n_arg_0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__ready;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__acc_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__arg_0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__carryless_t0;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__count_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__lhs_sign_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__n_acc_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__n_arg_0_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cen_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cin_t0;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_cout_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_lhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_rhs_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__padd_sub_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_16_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_32_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_4_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__pw_8_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__ready_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rhs_sign_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rs1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__rs2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_32_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_32;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_lhs_t0;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_lhs;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_rhs_t0;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_malu_muldivrem__i_xc_malu_mul__add_rhs;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__lhs;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__rhs;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__pw;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__cin;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__sub;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__c_en;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__c_out;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__result;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__c_en_t0;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__c_out_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__cin_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__lhs_t0;
input logic [4:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__pw_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__rhs_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__sub_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__carry_mask_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__carry_mask;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_0___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_0___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_0___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_0___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_10___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_10___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_10___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_10___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_11___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_11___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_11___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_11___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_11___force_carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_11___force_carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_12___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_12___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_12___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_12___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_13___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_13___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_13___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_13___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_13___force_carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_13___force_carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_14___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_14___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_14___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_14___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_15___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_15___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_15___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_15___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_15___force_carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_15___force_carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_16___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_16___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_16___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_16___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_17___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_17___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_17___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_17___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_18___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_18___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_18___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_18___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_19___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_19___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_19___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_19___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_1___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_1___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_1___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_1___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_20___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_20___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_20___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_20___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_21___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_21___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_21___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_21___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_22___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_22___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_22___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_22___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_23___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_23___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_23___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_23___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_23___force_carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_23___force_carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_24___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_24___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_24___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_24___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_25___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_25___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_25___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_25___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_26___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_26___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_26___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_26___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_27___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_27___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_27___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_27___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_28___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_28___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_28___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_28___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_29___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_29___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_29___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_29___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_2___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_2___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_2___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_2___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_30___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_30___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_30___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_30___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_31___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_31___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_31___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_31___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_3___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_3___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_3___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_3___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_4___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_4___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_4___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_4___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_5___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_5___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_5___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_5___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_6___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_6___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_6___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_6___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_7___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_7___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_7___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_7___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_8___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_8___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_8___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_8___carry;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_9___c_in_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_9___c_in;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_9___carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__genblk1_9___carry;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__rhs_m_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_p_addsub__rhs_m;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs1;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs2;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs3;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_init;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mdr;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_msub_1;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_macc_1;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mmul_1;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mmul_2;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_done;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__acc;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__carry;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__count;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_lhs;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_rhs;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_cin;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_sub;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_cout;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_result;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_madd;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_msub;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_macc;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_mmul;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__n_carry;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__n_acc;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__result;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__ready;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__result_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__acc_t0;
input logic [5:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__count_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__n_acc_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_cin_t0;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_cout_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_lhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_result_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_rhs_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__padd_sub_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__ready_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs1_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs2_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__rs3_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_done_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_init_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_macc_1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mdr_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mmul_1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_mmul_2_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__fsm_msub_1_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__n_carry_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_macc_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_madd_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_mmul_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__uop_msub_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_lhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_lhs;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_n_acc_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_n_acc;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_rhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__macc_rhs;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_lhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_lhs;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_n_acc_t0;
input logic [63:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_n_acc;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_rhs_t0;
input logic [31:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__mmul_rhs;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__msub_lhs_t0;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__msub_lhs;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__msub_rhs_t0;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__msub_rhs;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__result_acc_t0;
input logic i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__result_acc;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__sub_result_t0;
input logic [32:0] i_pipeline__i_pipeline_s2_execute__i_xc_malu__i_xc_malu_long__sub_result;
input logic i_pipeline__i_pipeline_s3_memory__g_clk;
input logic i_pipeline__i_pipeline_s3_memory__g_resetn;
input logic i_pipeline__i_pipeline_s3_memory__flush;
input logic [4:0] i_pipeline__i_pipeline_s3_memory__s3_rd;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__s3_opr_a;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__s3_opr_b;
input logic [4:0] i_pipeline__i_pipeline_s3_memory__s3_uop;
input logic [7:0] i_pipeline__i_pipeline_s3_memory__s3_fu;
input logic i_pipeline__i_pipeline_s3_memory__s3_trap;
input logic [1:0] i_pipeline__i_pipeline_s3_memory__s3_size;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__s3_instr;
input logic i_pipeline__i_pipeline_s3_memory__s3_busy;
input logic i_pipeline__i_pipeline_s3_memory__s3_valid;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__leak_prng;
input logic [12:0] i_pipeline__i_pipeline_s3_memory__leak_lkgcfg;
input logic i_pipeline__i_pipeline_s3_memory__leak_fence_unc0;
input logic i_pipeline__i_pipeline_s3_memory__leak_fence_unc1;
input logic i_pipeline__i_pipeline_s3_memory__leak_fence_unc2;
input logic [4:0] i_pipeline__i_pipeline_s3_memory__fwd_s3_rd;
input logic i_pipeline__i_pipeline_s3_memory__fwd_s3_wide;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__fwd_s3_wdata;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__fwd_s3_wdata_hi;
input logic i_pipeline__i_pipeline_s3_memory__fwd_s3_load;
input logic i_pipeline__i_pipeline_s3_memory__fwd_s3_csr;
input logic i_pipeline__i_pipeline_s3_memory__hold_lsu_req;
input logic i_pipeline__i_pipeline_s3_memory__mmio_en;
input logic i_pipeline__i_pipeline_s3_memory__mmio_wen;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__mmio_addr;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__mmio_wdata;
input logic i_pipeline__i_pipeline_s3_memory__dmem_req;
input logic i_pipeline__i_pipeline_s3_memory__dmem_wen;
input logic [3:0] i_pipeline__i_pipeline_s3_memory__dmem_strb;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__dmem_wdata;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__dmem_addr;
input logic i_pipeline__i_pipeline_s3_memory__dmem_gnt;
input logic [4:0] i_pipeline__i_pipeline_s3_memory__s4_rd;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__s4_opr_a;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__s4_opr_b;
input logic [4:0] i_pipeline__i_pipeline_s3_memory__s4_uop;
input logic [7:0] i_pipeline__i_pipeline_s3_memory__s4_fu;
input logic i_pipeline__i_pipeline_s3_memory__s4_trap;
input logic [1:0] i_pipeline__i_pipeline_s3_memory__s4_size;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__s4_instr;
input logic i_pipeline__i_pipeline_s3_memory__s4_busy;
input logic i_pipeline__i_pipeline_s3_memory__s4_valid;
input logic i_pipeline__i_pipeline_s3_memory__flush_t0;
input logic [12:0] i_pipeline__i_pipeline_s3_memory__leak_lkgcfg_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__leak_prng_t0;
input logic i_pipeline__i_pipeline_s3_memory__mmio_wen_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__mmio_wdata_t0;
input logic i_pipeline__i_pipeline_s3_memory__mmio_en_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__mmio_addr_t0;
input logic i_pipeline__i_pipeline_s3_memory__s3_busy_t0;
input logic [7:0] i_pipeline__i_pipeline_s3_memory__s3_fu_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__s3_instr_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__s3_opr_a_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__s3_opr_b_t0;
input logic [4:0] i_pipeline__i_pipeline_s3_memory__s3_rd_t0;
input logic [1:0] i_pipeline__i_pipeline_s3_memory__s3_size_t0;
input logic i_pipeline__i_pipeline_s3_memory__s3_trap_t0;
input logic [4:0] i_pipeline__i_pipeline_s3_memory__s3_uop_t0;
input logic i_pipeline__i_pipeline_s3_memory__s3_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__dmem_addr_t0;
input logic i_pipeline__i_pipeline_s3_memory__dmem_gnt_t0;
input logic i_pipeline__i_pipeline_s3_memory__dmem_req_t0;
input logic [3:0] i_pipeline__i_pipeline_s3_memory__dmem_strb_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__dmem_wdata_t0;
input logic i_pipeline__i_pipeline_s3_memory__dmem_wen_t0;
input logic i_pipeline__i_pipeline_s3_memory__hold_lsu_req_t0;
input logic i_pipeline__i_pipeline_s3_memory__fwd_s3_csr_t0;
input logic i_pipeline__i_pipeline_s3_memory__fwd_s3_load_t0;
input logic [4:0] i_pipeline__i_pipeline_s3_memory__fwd_s3_rd_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__fwd_s3_wdata_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__fwd_s3_wdata_hi_t0;
input logic i_pipeline__i_pipeline_s3_memory__fwd_s3_wide_t0;
input logic i_pipeline__i_pipeline_s3_memory__leak_fence_unc0_t0;
input logic i_pipeline__i_pipeline_s3_memory__leak_fence_unc1_t0;
input logic i_pipeline__i_pipeline_s3_memory__leak_fence_unc2_t0;
input logic i_pipeline__i_pipeline_s3_memory__s4_busy_t0;
input logic [7:0] i_pipeline__i_pipeline_s3_memory__s4_fu_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__s4_instr_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__s4_opr_a_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__s4_opr_b_t0;
input logic [4:0] i_pipeline__i_pipeline_s3_memory__s4_rd_t0;
input logic [1:0] i_pipeline__i_pipeline_s3_memory__s4_size_t0;
input logic i_pipeline__i_pipeline_s3_memory__s4_trap_t0;
input logic [4:0] i_pipeline__i_pipeline_s3_memory__s4_uop_t0;
input logic i_pipeline__i_pipeline_s3_memory__s4_valid_t0;
input logic i_pipeline__i_pipeline_s3_memory__bitw_gpr_wide_t0;
input logic i_pipeline__i_pipeline_s3_memory__bitw_gpr_wide;
input logic i_pipeline__i_pipeline_s3_memory__imul_gpr_wide_t0;
input logic i_pipeline__i_pipeline_s3_memory__imul_gpr_wide;
input logic i_pipeline__i_pipeline_s3_memory__leak_fence_t0;
input logic i_pipeline__i_pipeline_s3_memory__leak_fence;
input logic i_pipeline__i_pipeline_s3_memory__lsu_a_error_t0;
input logic i_pipeline__i_pipeline_s3_memory__lsu_a_error;
input logic i_pipeline__i_pipeline_s3_memory__lsu_byte_t0;
input logic i_pipeline__i_pipeline_s3_memory__lsu_byte;
input logic [5:0] i_pipeline__i_pipeline_s3_memory__lsu_cause_t0;
input logic [5:0] i_pipeline__i_pipeline_s3_memory__lsu_cause;
input logic i_pipeline__i_pipeline_s3_memory__lsu_half_t0;
input logic i_pipeline__i_pipeline_s3_memory__lsu_half;
input logic i_pipeline__i_pipeline_s3_memory__lsu_mmio_t0;
input logic i_pipeline__i_pipeline_s3_memory__lsu_mmio;
input logic i_pipeline__i_pipeline_s3_memory__lsu_ready_t0;
input logic i_pipeline__i_pipeline_s3_memory__lsu_ready;
input logic i_pipeline__i_pipeline_s3_memory__lsu_word_t0;
input logic i_pipeline__i_pipeline_s3_memory__lsu_word;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__n_s4_opr_a_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__n_s4_opr_a;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__n_s4_opr_b_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__n_s4_opr_b;
input logic [4:0] i_pipeline__i_pipeline_s3_memory__n_s4_rd_t0;
input logic [4:0] i_pipeline__i_pipeline_s3_memory__n_s4_rd;
input logic i_pipeline__i_pipeline_s3_memory__n_s4_trap_t0;
input logic i_pipeline__i_pipeline_s3_memory__n_s4_trap;
input logic i_pipeline__i_pipeline_s3_memory__opra_flush_t0;
input logic i_pipeline__i_pipeline_s3_memory__opra_flush;
input logic i_pipeline__i_pipeline_s3_memory__opra_ld_en_t0;
input logic i_pipeline__i_pipeline_s3_memory__opra_ld_en;
input logic i_pipeline__i_pipeline_s3_memory__oprb_flush_t0;
input logic i_pipeline__i_pipeline_s3_memory__oprb_flush;
input logic i_pipeline__i_pipeline_s3_memory__oprb_ld_en_t0;
input logic i_pipeline__i_pipeline_s3_memory__oprb_ld_en;
input logic i_pipeline__i_pipeline_s3_memory__p_busy_t0;
input logic i_pipeline__i_pipeline_s3_memory__p_busy;
input logic i_pipeline__i_pipeline_s3_memory__p_valid_t0;
input logic i_pipeline__i_pipeline_s3_memory__p_valid;
input logic [52:0] i_pipeline__i_pipeline_s3_memory__pipe_reg_out_t0;
input logic [52:0] i_pipeline__i_pipeline_s3_memory__pipe_reg_out;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__g_clk;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__g_resetn;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_valid;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_a_error;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_ready;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_mmio;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__pipe_prog;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_addr;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_wdata;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_load;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_store;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_byte;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_half;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_word;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_signed;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__hold_lsu_req;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_en;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_wen;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_addr;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_wdata;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_req;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_wen;
input logic [3:0] i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_strb;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_wdata;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_addr;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_gnt;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_wen_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_wdata_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_en_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_addr_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_load_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_store_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_addr_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_gnt_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_req_t0;
input logic [3:0] i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_strb_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_wdata_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_wen_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__hold_lsu_req_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_a_error_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_addr_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_byte_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_half_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_mmio_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_ready_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_signed_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_wdata_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_word_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__pipe_prog_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_txn_done_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__dmem_txn_done;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_finished_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__lsu_finished;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_done_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__mmio_done;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__n_lsu_finished_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__n_lsu_finished;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__n_mmio_done_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_lsu__n_mmio_done;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__g_clk;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__g_resetn;
input logic [52:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_data;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_valid;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_busy;
input logic [52:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__mr_data;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__flush;
input logic [52:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__flush_dat;
input logic [52:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_data;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_valid;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_busy;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__flush_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_valid_t0;
input logic [52:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_data_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__o_busy_t0;
input logic [52:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__mr_data_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_valid_t0;
input logic [52:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_data_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__i_busy_t0;
input logic [52:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__flush_dat_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__genblk1__progress_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg__genblk1__progress;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__g_clk;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__g_resetn;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_data;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_valid;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_busy;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__mr_data;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__flush;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__flush_dat;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_data;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_valid;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_busy;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__flush_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_data_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__o_busy_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__mr_data_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_data_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__i_busy_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__flush_dat_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__genblk1__progress_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_a__genblk1__progress;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__g_clk;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__g_resetn;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_data;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_valid;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_busy;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__mr_data;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__flush;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__flush_dat;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_data;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_valid;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_busy;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__flush_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_data_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__o_busy_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__mr_data_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_valid_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_data_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__i_busy_t0;
input logic [31:0] i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__flush_dat_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__genblk1__progress_t0;
input logic i_pipeline__i_pipeline_s3_memory__i_mem_pipereg_opr_b__genblk1__progress;
input logic i_pipeline__i_pipeline_s4_writeback__g_clk;
input logic i_pipeline__i_pipeline_s4_writeback__g_resetn;
input logic [4:0] i_pipeline__i_pipeline_s4_writeback__s4_rd;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__s4_opr_a;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__s4_opr_b;
input logic [4:0] i_pipeline__i_pipeline_s4_writeback__s4_uop;
input logic [7:0] i_pipeline__i_pipeline_s4_writeback__s4_fu;
input logic i_pipeline__i_pipeline_s4_writeback__s4_trap;
input logic [1:0] i_pipeline__i_pipeline_s4_writeback__s4_size;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__s4_instr;
input logic i_pipeline__i_pipeline_s4_writeback__s4_busy;
input logic i_pipeline__i_pipeline_s4_writeback__s4_valid;
input logic [4:0] i_pipeline__i_pipeline_s4_writeback__fwd_s4_rd;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__fwd_s4_wdata;
input logic i_pipeline__i_pipeline_s4_writeback__fwd_s4_load;
input logic i_pipeline__i_pipeline_s4_writeback__fwd_s4_csr;
input logic i_pipeline__i_pipeline_s4_writeback__gpr_wen;
input logic i_pipeline__i_pipeline_s4_writeback__gpr_wide;
input logic [4:0] i_pipeline__i_pipeline_s4_writeback__gpr_rd;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__gpr_wdata;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__gpr_wdata_hi;
input logic i_pipeline__i_pipeline_s4_writeback__int_trap_req;
input logic [5:0] i_pipeline__i_pipeline_s4_writeback__int_trap_cause;
input logic i_pipeline__i_pipeline_s4_writeback__int_trap_ack;
input logic i_pipeline__i_pipeline_s4_writeback__trap_cpu;
input logic i_pipeline__i_pipeline_s4_writeback__trap_int;
input logic [5:0] i_pipeline__i_pipeline_s4_writeback__trap_cause;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__trap_mtval;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__trap_pc;
input logic i_pipeline__i_pipeline_s4_writeback__exec_mret;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__csr_mepc;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__csr_mtvec;
input logic i_pipeline__i_pipeline_s4_writeback__vector_intrs;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__trs_pc;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__trs_instr;
input logic i_pipeline__i_pipeline_s4_writeback__trs_valid;
input logic i_pipeline__i_pipeline_s4_writeback__csr_en;
input logic i_pipeline__i_pipeline_s4_writeback__csr_wr;
input logic i_pipeline__i_pipeline_s4_writeback__csr_wr_set;
input logic i_pipeline__i_pipeline_s4_writeback__csr_wr_clr;
input logic [11:0] i_pipeline__i_pipeline_s4_writeback__csr_addr;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__csr_wdata;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__csr_rdata;
input logic i_pipeline__i_pipeline_s4_writeback__csr_error;
input logic i_pipeline__i_pipeline_s4_writeback__cf_req;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__cf_target;
input logic i_pipeline__i_pipeline_s4_writeback__cf_ack;
input logic i_pipeline__i_pipeline_s4_writeback__hold_lsu_req;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__mmio_rdata;
input logic i_pipeline__i_pipeline_s4_writeback__mmio_error;
input logic i_pipeline__i_pipeline_s4_writeback__dmem_recv;
input logic i_pipeline__i_pipeline_s4_writeback__dmem_ack;
input logic i_pipeline__i_pipeline_s4_writeback__dmem_error;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__dmem_rdata;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__cf_target_t0;
input logic i_pipeline__i_pipeline_s4_writeback__cf_req_t0;
input logic i_pipeline__i_pipeline_s4_writeback__cf_ack_t0;
input logic i_pipeline__i_pipeline_s4_writeback__int_trap_req_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__mmio_rdata_t0;
input logic i_pipeline__i_pipeline_s4_writeback__mmio_error_t0;
input logic [5:0] i_pipeline__i_pipeline_s4_writeback__int_trap_cause_t0;
input logic i_pipeline__i_pipeline_s4_writeback__int_trap_ack_t0;
input logic [5:0] i_pipeline__i_pipeline_s4_writeback__trap_cause_t0;
input logic i_pipeline__i_pipeline_s4_writeback__hold_lsu_req_t0;
input logic i_pipeline__i_pipeline_s4_writeback__s4_busy_t0;
input logic [7:0] i_pipeline__i_pipeline_s4_writeback__s4_fu_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__s4_instr_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__s4_opr_a_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__s4_opr_b_t0;
input logic [4:0] i_pipeline__i_pipeline_s4_writeback__s4_rd_t0;
input logic [1:0] i_pipeline__i_pipeline_s4_writeback__s4_size_t0;
input logic i_pipeline__i_pipeline_s4_writeback__s4_trap_t0;
input logic [4:0] i_pipeline__i_pipeline_s4_writeback__s4_uop_t0;
input logic i_pipeline__i_pipeline_s4_writeback__s4_valid_t0;
input logic [11:0] i_pipeline__i_pipeline_s4_writeback__csr_addr_t0;
input logic i_pipeline__i_pipeline_s4_writeback__csr_en_t0;
input logic i_pipeline__i_pipeline_s4_writeback__csr_error_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__csr_mepc_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__csr_mtvec_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__csr_rdata_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__csr_wdata_t0;
input logic i_pipeline__i_pipeline_s4_writeback__csr_wr_t0;
input logic i_pipeline__i_pipeline_s4_writeback__csr_wr_clr_t0;
input logic i_pipeline__i_pipeline_s4_writeback__csr_wr_set_t0;
input logic i_pipeline__i_pipeline_s4_writeback__dmem_ack_t0;
input logic i_pipeline__i_pipeline_s4_writeback__dmem_error_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__dmem_rdata_t0;
input logic i_pipeline__i_pipeline_s4_writeback__dmem_recv_t0;
input logic i_pipeline__i_pipeline_s4_writeback__exec_mret_t0;
input logic i_pipeline__i_pipeline_s4_writeback__fwd_s4_csr_t0;
input logic i_pipeline__i_pipeline_s4_writeback__fwd_s4_load_t0;
input logic [4:0] i_pipeline__i_pipeline_s4_writeback__fwd_s4_rd_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__fwd_s4_wdata_t0;
input logic [4:0] i_pipeline__i_pipeline_s4_writeback__gpr_rd_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__gpr_wdata_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__gpr_wdata_hi_t0;
input logic i_pipeline__i_pipeline_s4_writeback__gpr_wen_t0;
input logic i_pipeline__i_pipeline_s4_writeback__gpr_wide_t0;
input logic i_pipeline__i_pipeline_s4_writeback__trap_cpu_t0;
input logic i_pipeline__i_pipeline_s4_writeback__trap_int_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__trap_mtval_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__trap_pc_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__trs_instr_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__trs_pc_t0;
input logic i_pipeline__i_pipeline_s4_writeback__trs_valid_t0;
input logic i_pipeline__i_pipeline_s4_writeback__vector_intrs_t0;
input logic i_pipeline__i_pipeline_s4_writeback__cf_req_noint_t0;
input logic i_pipeline__i_pipeline_s4_writeback__cf_req_noint;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__cf_target_noint_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__cf_target_noint;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_busy_t0;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_busy;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_cf_taken_t0;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_cf_taken;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_done_t0;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_done;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_ebreak_t0;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_ebreak;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_ecall_t0;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_ecall;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_finish_now_t0;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_finish_now;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__cfu_gpr_wdata_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__cfu_gpr_wdata;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_gpr_wen_t0;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_gpr_wen;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_mret_t0;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_mret;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_tgt_trap_t0;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_tgt_trap;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_trap_t0;
input logic i_pipeline__i_pipeline_s4_writeback__cfu_trap;
input logic i_pipeline__i_pipeline_s4_writeback__csr_done_t0;
input logic i_pipeline__i_pipeline_s4_writeback__csr_done;
input logic i_pipeline__i_pipeline_s4_writeback__csr_gpr_wen_t0;
input logic i_pipeline__i_pipeline_s4_writeback__csr_gpr_wen;
input logic i_pipeline__i_pipeline_s4_writeback__csr_read_t0;
input logic i_pipeline__i_pipeline_s4_writeback__csr_read;
input logic i_pipeline__i_pipeline_s4_writeback__dmem_error_seen_t0;
input logic i_pipeline__i_pipeline_s4_writeback__dmem_error_seen;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_b_error_t0;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_b_error;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_busy_t0;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_busy;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_byte_t0;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_byte;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_gpr_wen_t0;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_gpr_wen;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_half_t0;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_half;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_load_t0;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_load;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_mmio_t0;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_mmio;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_rsp_seen_t0;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_rsp_seen;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_store_t0;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_store;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_txn_recv_t0;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_txn_recv;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_word_t0;
input logic i_pipeline__i_pipeline_s4_writeback__lsu_word;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__mem_rdata_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__mem_rdata;
input logic i_pipeline__i_pipeline_s4_writeback__n_cfu_done_t0;
input logic i_pipeline__i_pipeline_s4_writeback__n_cfu_done;
input logic i_pipeline__i_pipeline_s4_writeback__n_csr_done_t0;
input logic i_pipeline__i_pipeline_s4_writeback__n_csr_done;
input logic i_pipeline__i_pipeline_s4_writeback__n_dmem_error_seen_t0;
input logic i_pipeline__i_pipeline_s4_writeback__n_dmem_error_seen;
input logic i_pipeline__i_pipeline_s4_writeback__n_lsu_rsp_seen_t0;
input logic i_pipeline__i_pipeline_s4_writeback__n_lsu_rsp_seen;
input logic i_pipeline__i_pipeline_s4_writeback__pipe_progress_t0;
input logic i_pipeline__i_pipeline_s4_writeback__pipe_progress;
input logic [7:0] i_pipeline__i_pipeline_s4_writeback__rdata_b0_t0;
input logic [7:0] i_pipeline__i_pipeline_s4_writeback__rdata_b0;
input logic [7:0] i_pipeline__i_pipeline_s4_writeback__rdata_b1_t0;
input logic [7:0] i_pipeline__i_pipeline_s4_writeback__rdata_b1;
input logic [15:0] i_pipeline__i_pipeline_s4_writeback__rdata_h1_t0;
input logic [15:0] i_pipeline__i_pipeline_s4_writeback__rdata_h1;
input logic i_pipeline__i_pipeline_s4_writeback__rng_gpr_wen_t0;
input logic i_pipeline__i_pipeline_s4_writeback__rng_gpr_wen;
input logic i_pipeline__i_pipeline_s4_writeback__trap_int_pending_t0;
input logic i_pipeline__i_pipeline_s4_writeback__trap_int_pending;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__trap_target_addr_t0;
input logic [31:0] i_pipeline__i_pipeline_s4_writeback__trap_target_addr;
input logic [7:0] i_pipeline__i_pipeline_s4_writeback__trap_vector_offset_t0;
input logic [7:0] i_pipeline__i_pipeline_s4_writeback__trap_vector_offset;


`include `PROPERTIES_FILE

endmodule
