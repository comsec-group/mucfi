bind picorv32 picorv32_fpv picorv32_fpv_bind (
.clk(
  clk),
.resetn(
  resetn),
.trap(
  trap),
.mem_valid(
  mem_valid),
.mem_instr(
  mem_instr),
.mem_ready(
  mem_ready),
.mem_addr(
  mem_addr),
.mem_wdata(
  mem_wdata),
.mem_wstrb(
  mem_wstrb),
.mem_rdata(
  mem_rdata),
.mem_la_read(
  mem_la_read),
.mem_la_write(
  mem_la_write),
.mem_la_addr(
  mem_la_addr),
.mem_la_wdata(
  mem_la_wdata),
.mem_la_wstrb(
  mem_la_wstrb),
.pcpi_valid(
  pcpi_valid),
.pcpi_insn(
  pcpi_insn),
.pcpi_rs1(
  pcpi_rs1),
.pcpi_rs2(
  pcpi_rs2),
.pcpi_wr(
  pcpi_wr),
.pcpi_rd(
  pcpi_rd),
.pcpi_wait(
  pcpi_wait),
.pcpi_ready(
  pcpi_ready),
.irq(
  irq),
.eoi(
  eoi),
.rvfi_valid(
  rvfi_valid),
.rvfi_order(
  rvfi_order),
.rvfi_insn(
  rvfi_insn),
.rvfi_trap(
  rvfi_trap),
.rvfi_halt(
  rvfi_halt),
.rvfi_intr(
  rvfi_intr),
.rvfi_mode(
  rvfi_mode),
.rvfi_ixl(
  rvfi_ixl),
.rvfi_rs1_addr(
  rvfi_rs1_addr),
.rvfi_rs2_addr(
  rvfi_rs2_addr),
.rvfi_rs1_rdata(
  rvfi_rs1_rdata),
.rvfi_rs2_rdata(
  rvfi_rs2_rdata),
.rvfi_rd_addr(
  rvfi_rd_addr),
.rvfi_rd_wdata(
  rvfi_rd_wdata),
.rvfi_pc_rdata(
  rvfi_pc_rdata),
.rvfi_pc_wdata(
  rvfi_pc_wdata),
.rvfi_mem_addr(
  rvfi_mem_addr),
.rvfi_mem_rmask(
  rvfi_mem_rmask),
.rvfi_mem_wmask(
  rvfi_mem_wmask),
.rvfi_mem_rdata(
  rvfi_mem_rdata),
.rvfi_mem_wdata(
  rvfi_mem_wdata),
.rvfi_csr_mcycle_rmask(
  rvfi_csr_mcycle_rmask),
.rvfi_csr_mcycle_wmask(
  rvfi_csr_mcycle_wmask),
.rvfi_csr_mcycle_rdata(
  rvfi_csr_mcycle_rdata),
.rvfi_csr_mcycle_wdata(
  rvfi_csr_mcycle_wdata),
.rvfi_csr_minstret_rmask(
  rvfi_csr_minstret_rmask),
.rvfi_csr_minstret_wmask(
  rvfi_csr_minstret_wmask),
.rvfi_csr_minstret_rdata(
  rvfi_csr_minstret_rdata),
.rvfi_csr_minstret_wdata(
  rvfi_csr_minstret_wdata),
.trace_valid(
  trace_valid),
.trace_data(
  trace_data),
.trap_t0(
  trap_t0),
.trace_valid_t0(
  trace_valid_t0),
.trace_data_t0(
  trace_data_t0),
.rvfi_valid_t0(
  rvfi_valid_t0),
.rvfi_trap_t0(
  rvfi_trap_t0),
.rvfi_rs2_rdata_t0(
  rvfi_rs2_rdata_t0),
.rvfi_rs2_addr_t0(
  rvfi_rs2_addr_t0),
.rvfi_rs1_rdata_t0(
  rvfi_rs1_rdata_t0),
.rvfi_rs1_addr_t0(
  rvfi_rs1_addr_t0),
.rvfi_rd_wdata_t0(
  rvfi_rd_wdata_t0),
.rvfi_rd_addr_t0(
  rvfi_rd_addr_t0),
.rvfi_pc_wdata_t0(
  rvfi_pc_wdata_t0),
.rvfi_pc_rdata_t0(
  rvfi_pc_rdata_t0),
.rvfi_order_t0(
  rvfi_order_t0),
.rvfi_mode_t0(
  rvfi_mode_t0),
.rvfi_mem_wmask_t0(
  rvfi_mem_wmask_t0),
.rvfi_mem_wdata_t0(
  rvfi_mem_wdata_t0),
.rvfi_mem_rmask_t0(
  rvfi_mem_rmask_t0),
.rvfi_mem_rdata_t0(
  rvfi_mem_rdata_t0),
.rvfi_mem_addr_t0(
  rvfi_mem_addr_t0),
.rvfi_ixl_t0(
  rvfi_ixl_t0),
.rvfi_intr_t0(
  rvfi_intr_t0),
.rvfi_insn_t0(
  rvfi_insn_t0),
.rvfi_halt_t0(
  rvfi_halt_t0),
.rvfi_csr_minstret_wmask_t0(
  rvfi_csr_minstret_wmask_t0),
.rvfi_csr_minstret_wdata_t0(
  rvfi_csr_minstret_wdata_t0),
.rvfi_csr_minstret_rmask_t0(
  rvfi_csr_minstret_rmask_t0),
.rvfi_csr_minstret_rdata_t0(
  rvfi_csr_minstret_rdata_t0),
.rvfi_csr_mcycle_wmask_t0(
  rvfi_csr_mcycle_wmask_t0),
.rvfi_csr_mcycle_wdata_t0(
  rvfi_csr_mcycle_wdata_t0),
.rvfi_csr_mcycle_rmask_t0(
  rvfi_csr_mcycle_rmask_t0),
.rvfi_csr_mcycle_rdata_t0(
  rvfi_csr_mcycle_rdata_t0),
.mem_wstrb_t0(
  mem_wstrb_t0),
.mem_wdata_t0(
  mem_wdata_t0),
.mem_valid_t0(
  mem_valid_t0),
.mem_ready_t0(
  mem_ready_t0),
.mem_rdata_t0(
  mem_rdata_t0),
.mem_la_wstrb_t0(
  mem_la_wstrb_t0),
.mem_la_write_t0(
  mem_la_write_t0),
.mem_la_wdata_t0(
  mem_la_wdata_t0),
.mem_la_read_t0(
  mem_la_read_t0),
.mem_la_addr_t0(
  mem_la_addr_t0),
.mem_instr_t0(
  mem_instr_t0),
.mem_addr_t0(
  mem_addr_t0),
.irq_t0(
  irq_t0),
.eoi_t0(
  eoi_t0),
.pcpi_insn_t0(
  pcpi_insn_t0),
.pcpi_rd_t0(
  pcpi_rd_t0),
.pcpi_ready_t0(
  pcpi_ready_t0),
.pcpi_rs1_t0(
  pcpi_rs1_t0),
.pcpi_rs2_t0(
  pcpi_rs2_t0),
.pcpi_valid_t0(
  pcpi_valid_t0),
.pcpi_wait_t0(
  pcpi_wait_t0),
.pcpi_wr_t0(
  pcpi_wr_t0),
.alu_add_sub(
  alu_add_sub),
.alu_add_sub_t0(
  alu_add_sub_t0),
.alu_eq(
  alu_eq),
.alu_lts(
  alu_lts),
.alu_ltu(
  alu_ltu),
.alu_out(
  alu_out),
.alu_out_0(
  alu_out_0),
.alu_out_q(
  alu_out_q),
.alu_out_q_t0(
  alu_out_q_t0),
.alu_out_t0(
  alu_out_t0),
.cached_insn_opcode(
  cached_insn_opcode),
.cached_insn_opcode_t0(
  cached_insn_opcode_t0),
.cached_insn_rs1(
  cached_insn_rs1),
.cached_insn_rs1_t0(
  cached_insn_rs1_t0),
.cached_insn_rs2(
  cached_insn_rs2),
.cached_insn_rs2_t0(
  cached_insn_rs2_t0),
.count_cycle(
  count_cycle),
.count_cycle_t0(
  count_cycle_t0),
.count_instr(
  count_instr),
.count_instr_t0(
  count_instr_t0),
.cpu_state(
  cpu_state),
.cpuregs_0_(
  \cpuregs[0] ),
.cpuregs_0__t0(
  \cpuregs[0]_t0 ),
.cpuregs_10_(
  \cpuregs[10] ),
.cpuregs_10__t0(
  \cpuregs[10]_t0 ),
.cpuregs_11_(
  \cpuregs[11] ),
.cpuregs_11__t0(
  \cpuregs[11]_t0 ),
.cpuregs_12_(
  \cpuregs[12] ),
.cpuregs_12__t0(
  \cpuregs[12]_t0 ),
.cpuregs_13_(
  \cpuregs[13] ),
.cpuregs_13__t0(
  \cpuregs[13]_t0 ),
.cpuregs_14_(
  \cpuregs[14] ),
.cpuregs_14__t0(
  \cpuregs[14]_t0 ),
.cpuregs_15_(
  \cpuregs[15] ),
.cpuregs_15__t0(
  \cpuregs[15]_t0 ),
.cpuregs_16_(
  \cpuregs[16] ),
.cpuregs_16__t0(
  \cpuregs[16]_t0 ),
.cpuregs_17_(
  \cpuregs[17] ),
.cpuregs_17__t0(
  \cpuregs[17]_t0 ),
.cpuregs_18_(
  \cpuregs[18] ),
.cpuregs_18__t0(
  \cpuregs[18]_t0 ),
.cpuregs_19_(
  \cpuregs[19] ),
.cpuregs_19__t0(
  \cpuregs[19]_t0 ),
.cpuregs_1_(
  \cpuregs[1] ),
.cpuregs_1__t0(
  \cpuregs[1]_t0 ),
.cpuregs_20_(
  \cpuregs[20] ),
.cpuregs_20__t0(
  \cpuregs[20]_t0 ),
.cpuregs_21_(
  \cpuregs[21] ),
.cpuregs_21__t0(
  \cpuregs[21]_t0 ),
.cpuregs_22_(
  \cpuregs[22] ),
.cpuregs_22__t0(
  \cpuregs[22]_t0 ),
.cpuregs_23_(
  \cpuregs[23] ),
.cpuregs_23__t0(
  \cpuregs[23]_t0 ),
.cpuregs_24_(
  \cpuregs[24] ),
.cpuregs_24__t0(
  \cpuregs[24]_t0 ),
.cpuregs_25_(
  \cpuregs[25] ),
.cpuregs_25__t0(
  \cpuregs[25]_t0 ),
.cpuregs_26_(
  \cpuregs[26] ),
.cpuregs_26__t0(
  \cpuregs[26]_t0 ),
.cpuregs_27_(
  \cpuregs[27] ),
.cpuregs_27__t0(
  \cpuregs[27]_t0 ),
.cpuregs_28_(
  \cpuregs[28] ),
.cpuregs_28__t0(
  \cpuregs[28]_t0 ),
.cpuregs_29_(
  \cpuregs[29] ),
.cpuregs_29__t0(
  \cpuregs[29]_t0 ),
.cpuregs_2_(
  \cpuregs[2] ),
.cpuregs_2__t0(
  \cpuregs[2]_t0 ),
.cpuregs_30_(
  \cpuregs[30] ),
.cpuregs_30__t0(
  \cpuregs[30]_t0 ),
.cpuregs_31_(
  \cpuregs[31] ),
.cpuregs_31__t0(
  \cpuregs[31]_t0 ),
.cpuregs_3_(
  \cpuregs[3] ),
.cpuregs_3__t0(
  \cpuregs[3]_t0 ),
.cpuregs_4_(
  \cpuregs[4] ),
.cpuregs_4__t0(
  \cpuregs[4]_t0 ),
.cpuregs_5_(
  \cpuregs[5] ),
.cpuregs_5__t0(
  \cpuregs[5]_t0 ),
.cpuregs_6_(
  \cpuregs[6] ),
.cpuregs_6__t0(
  \cpuregs[6]_t0 ),
.cpuregs_7_(
  \cpuregs[7] ),
.cpuregs_7__t0(
  \cpuregs[7]_t0 ),
.cpuregs_8_(
  \cpuregs[8] ),
.cpuregs_8__t0(
  \cpuregs[8]_t0 ),
.cpuregs_9_(
  \cpuregs[9] ),
.cpuregs_9__t0(
  \cpuregs[9]_t0 ),
.cpuregs_rs1(
  cpuregs_rs1),
.cpuregs_rs1_t0(
  cpuregs_rs1_t0),
.cpuregs_rs2(
  cpuregs_rs2),
.cpuregs_rs2_t0(
  cpuregs_rs2_t0),
.cpuregs_wrdata(
  cpuregs_wrdata),
.cpuregs_wrdata_t0(
  cpuregs_wrdata_t0),
.cpuregs_write(
  cpuregs_write),
.dbg_insn_opcode(
  dbg_insn_opcode),
.dbg_insn_opcode_t0(
  dbg_insn_opcode_t0),
.dbg_insn_rs1(
  dbg_insn_rs1),
.dbg_insn_rs1_t0(
  dbg_insn_rs1_t0),
.dbg_insn_rs2(
  dbg_insn_rs2),
.dbg_insn_rs2_t0(
  dbg_insn_rs2_t0),
.dbg_next(
  dbg_next),
.dbg_rs1val(
  dbg_rs1val),
.dbg_rs1val_t0(
  dbg_rs1val_t0),
.dbg_rs1val_valid(
  dbg_rs1val_valid),
.dbg_rs2val(
  dbg_rs2val),
.dbg_rs2val_t0(
  dbg_rs2val_t0),
.dbg_rs2val_valid(
  dbg_rs2val_valid),
.dbg_valid_insn(
  dbg_valid_insn),
.decoded_imm(
  decoded_imm),
.decoded_imm_j(
  decoded_imm_j),
.decoded_imm_j_reg_10_(
  \decoded_imm_j_reg[10] ),
.decoded_imm_j_reg_11_(
  \decoded_imm_j_reg[11] ),
.decoded_imm_j_reg_4_(
  \decoded_imm_j_reg[4] ),
.decoded_imm_j_reg_5_(
  \decoded_imm_j_reg[5] ),
.decoded_imm_j_reg_6_(
  \decoded_imm_j_reg[6] ),
.decoded_imm_j_reg_7_(
  \decoded_imm_j_reg[7] ),
.decoded_imm_j_t0(
  decoded_imm_j_t0),
.decoded_imm_j_t0_reg_10_(
  \decoded_imm_j_t0_reg[10] ),
.decoded_imm_j_t0_reg_11_(
  \decoded_imm_j_t0_reg[11] ),
.decoded_imm_j_t0_reg_4_(
  \decoded_imm_j_t0_reg[4] ),
.decoded_imm_j_t0_reg_5_(
  \decoded_imm_j_t0_reg[5] ),
.decoded_imm_j_t0_reg_6_(
  \decoded_imm_j_t0_reg[6] ),
.decoded_imm_j_t0_reg_7_(
  \decoded_imm_j_t0_reg[7] ),
.decoded_imm_t0(
  decoded_imm_t0),
.decoded_rd(
  decoded_rd),
.decoded_rd_t0(
  decoded_rd_t0),
.decoded_rs1(
  decoded_rs1),
.decoded_rs1_t0(
  decoded_rs1_t0),
.decoded_rs2(
  decoded_rs2),
.decoded_rs2_t0(
  decoded_rs2_t0),
.decoder_pseudo_trigger(
  decoder_pseudo_trigger),
.decoder_pseudo_trigger_q(
  decoder_pseudo_trigger_q),
.decoder_trigger(
  decoder_trigger),
.decoder_trigger_q(
  decoder_trigger_q),
.instr_add(
  instr_add),
.instr_addi(
  instr_addi),
.instr_and(
  instr_and),
.instr_andi(
  instr_andi),
.instr_auipc(
  instr_auipc),
.instr_beq(
  instr_beq),
.instr_bge(
  instr_bge),
.instr_bgeu(
  instr_bgeu),
.instr_blt(
  instr_blt),
.instr_bltu(
  instr_bltu),
.instr_bne(
  instr_bne),
.instr_ecall_ebreak(
  instr_ecall_ebreak),
.instr_fence(
  instr_fence),
.instr_jal(
  instr_jal),
.instr_jalr(
  instr_jalr),
.instr_lb(
  instr_lb),
.instr_lbu(
  instr_lbu),
.instr_lh(
  instr_lh),
.instr_lhu(
  instr_lhu),
.instr_lui(
  instr_lui),
.instr_lw(
  instr_lw),
.instr_or(
  instr_or),
.instr_ori(
  instr_ori),
.instr_rdcycle(
  instr_rdcycle),
.instr_rdcycleh(
  instr_rdcycleh),
.instr_rdinstr(
  instr_rdinstr),
.instr_rdinstrh(
  instr_rdinstrh),
.instr_sb(
  instr_sb),
.instr_sh(
  instr_sh),
.instr_sll(
  instr_sll),
.instr_slli(
  instr_slli),
.instr_slt(
  instr_slt),
.instr_slti(
  instr_slti),
.instr_sltiu(
  instr_sltiu),
.instr_sltu(
  instr_sltu),
.instr_sra(
  instr_sra),
.instr_srai(
  instr_srai),
.instr_srl(
  instr_srl),
.instr_srli(
  instr_srli),
.instr_sub(
  instr_sub),
.instr_sw(
  instr_sw),
.instr_trap(
  instr_trap),
.instr_xor(
  instr_xor),
.instr_xori(
  instr_xori),
.is_alu_reg_imm(
  is_alu_reg_imm),
.is_alu_reg_reg(
  is_alu_reg_reg),
.is_beq_bne_blt_bge_bltu_bgeu(
  is_beq_bne_blt_bge_bltu_bgeu),
.is_compare(
  is_compare),
.is_jalr_addi_slti_sltiu_xori_ori_andi(
  is_jalr_addi_slti_sltiu_xori_ori_andi),
.is_lb_lh_lw_lbu_lhu(
  is_lb_lh_lw_lbu_lhu),
.is_lui_auipc_jal(
  is_lui_auipc_jal),
.is_rdcycle_rdcycleh_rdinstr_rdinstrh(
  is_rdcycle_rdcycleh_rdinstr_rdinstrh),
.is_sb_sh_sw(
  is_sb_sh_sw),
.is_sll_srl_sra(
  is_sll_srl_sra),
.is_slli_srli_srai(
  is_slli_srli_srai),
.is_slti_blt_slt(
  is_slti_blt_slt),
.is_sltiu_bltu_sltu(
  is_sltiu_bltu_sltu),
.latched_branch(
  latched_branch),
.latched_is_lb(
  latched_is_lb),
.latched_is_lh(
  latched_is_lh),
.latched_rd(
  latched_rd),
.latched_rd_t0(
  latched_rd_t0),
.latched_stalu(
  latched_stalu),
.latched_store(
  latched_store),
.launch_next_insn(
  launch_next_insn),
.mem_do_prefetch(
  mem_do_prefetch),
.mem_do_rdata(
  mem_do_rdata),
.mem_do_rinst(
  mem_do_rinst),
.mem_do_wdata(
  mem_do_wdata),
.mem_done(
  mem_done),
.mem_rdata_latched(
  mem_rdata_latched),
.mem_rdata_latched_t0(
  mem_rdata_latched_t0),
.mem_rdata_q(
  mem_rdata_q),
.mem_rdata_q_t0(
  mem_rdata_q_t0),
.mem_rdata_word(
  mem_rdata_word),
.mem_rdata_word_t0(
  mem_rdata_word_t0),
.mem_state(
  mem_state),
.mem_wordsize(
  mem_wordsize),
.mem_xfer(
  mem_xfer),
.next_insn_opcode(
  next_insn_opcode),
.next_insn_opcode_t0(
  next_insn_opcode_t0),
.next_pc(
  next_pc),
.next_pc_t0(
  next_pc_t0),
.pcpi_div_rd(
  pcpi_div_rd),
.pcpi_div_rd_t0(
  pcpi_div_rd_t0),
.pcpi_div_ready(
  pcpi_div_ready),
.pcpi_div_ready_t0(
  pcpi_div_ready_t0),
.pcpi_div_wait(
  pcpi_div_wait),
.pcpi_div_wait_t0(
  pcpi_div_wait_t0),
.pcpi_div_wr(
  pcpi_div_wr),
.pcpi_div_wr_t0(
  pcpi_div_wr_t0),
.pcpi_int_rd(
  pcpi_int_rd),
.pcpi_int_rd_t0(
  pcpi_int_rd_t0),
.pcpi_int_ready(
  pcpi_int_ready),
.pcpi_int_wait(
  pcpi_int_wait),
.pcpi_int_wr(
  pcpi_int_wr),
.pcpi_mul_rd(
  pcpi_mul_rd),
.pcpi_mul_rd_t0(
  pcpi_mul_rd_t0),
.pcpi_mul_ready(
  pcpi_mul_ready),
.pcpi_mul_ready_t0(
  pcpi_mul_ready_t0),
.pcpi_mul_wait(
  pcpi_mul_wait),
.pcpi_mul_wait_t0(
  pcpi_mul_wait_t0),
.pcpi_mul_wr(
  pcpi_mul_wr),
.pcpi_mul_wr_t0(
  pcpi_mul_wr_t0),
.pcpi_timeout(
  pcpi_timeout),
.pcpi_timeout_counter(
  pcpi_timeout_counter),
.q_insn_rs1(
  q_insn_rs1),
.q_insn_rs1_t0(
  q_insn_rs1_t0),
.q_insn_rs2(
  q_insn_rs2),
.q_insn_rs2_t0(
  q_insn_rs2_t0),
.reg_next_pc(
  reg_next_pc),
.reg_next_pc_t0(
  reg_next_pc_t0),
.reg_out(
  reg_out),
.reg_out_t0(
  reg_out_t0),
.reg_pc(
  reg_pc),
.reg_pc_t0(
  reg_pc_t0),
.reg_sh(
  reg_sh),
.genblk1__genblk1__pcpi_mul__clk(
  \genblk1.genblk1.pcpi_mul .clk),
.genblk1__genblk1__pcpi_mul__resetn(
  \genblk1.genblk1.pcpi_mul .resetn),
.genblk1__genblk1__pcpi_mul__pcpi_valid(
  \genblk1.genblk1.pcpi_mul .pcpi_valid),
.genblk1__genblk1__pcpi_mul__pcpi_insn(
  \genblk1.genblk1.pcpi_mul .pcpi_insn),
.genblk1__genblk1__pcpi_mul__pcpi_rs1(
  \genblk1.genblk1.pcpi_mul .pcpi_rs1),
.genblk1__genblk1__pcpi_mul__pcpi_rs2(
  \genblk1.genblk1.pcpi_mul .pcpi_rs2),
.genblk1__genblk1__pcpi_mul__pcpi_wr(
  \genblk1.genblk1.pcpi_mul .pcpi_wr),
.genblk1__genblk1__pcpi_mul__pcpi_rd(
  \genblk1.genblk1.pcpi_mul .pcpi_rd),
.genblk1__genblk1__pcpi_mul__pcpi_wait(
  \genblk1.genblk1.pcpi_mul .pcpi_wait),
.genblk1__genblk1__pcpi_mul__pcpi_ready(
  \genblk1.genblk1.pcpi_mul .pcpi_ready),
.genblk1__genblk1__pcpi_mul__pcpi_insn_t0(
  \genblk1.genblk1.pcpi_mul .pcpi_insn_t0),
.genblk1__genblk1__pcpi_mul__pcpi_rd_t0(
  \genblk1.genblk1.pcpi_mul .pcpi_rd_t0),
.genblk1__genblk1__pcpi_mul__pcpi_ready_t0(
  \genblk1.genblk1.pcpi_mul .pcpi_ready_t0),
.genblk1__genblk1__pcpi_mul__pcpi_rs1_t0(
  \genblk1.genblk1.pcpi_mul .pcpi_rs1_t0),
.genblk1__genblk1__pcpi_mul__pcpi_rs2_t0(
  \genblk1.genblk1.pcpi_mul .pcpi_rs2_t0),
.genblk1__genblk1__pcpi_mul__pcpi_valid_t0(
  \genblk1.genblk1.pcpi_mul .pcpi_valid_t0),
.genblk1__genblk1__pcpi_mul__pcpi_wait_t0(
  \genblk1.genblk1.pcpi_mul .pcpi_wait_t0),
.genblk1__genblk1__pcpi_mul__pcpi_wr_t0(
  \genblk1.genblk1.pcpi_mul .pcpi_wr_t0),
.genblk1__genblk1__pcpi_mul__instr_any_mul(
  \genblk1.genblk1.pcpi_mul .instr_any_mul),
.genblk1__genblk1__pcpi_mul__instr_any_mulh(
  \genblk1.genblk1.pcpi_mul .instr_any_mulh),
.genblk1__genblk1__pcpi_mul__instr_mul(
  \genblk1.genblk1.pcpi_mul .instr_mul),
.genblk1__genblk1__pcpi_mul__instr_mulh(
  \genblk1.genblk1.pcpi_mul .instr_mulh),
.genblk1__genblk1__pcpi_mul__instr_mulhsu(
  \genblk1.genblk1.pcpi_mul .instr_mulhsu),
.genblk1__genblk1__pcpi_mul__instr_mulhu(
  \genblk1.genblk1.pcpi_mul .instr_mulhu),
.genblk1__genblk1__pcpi_mul__instr_rs1_signed(
  \genblk1.genblk1.pcpi_mul .instr_rs1_signed),
.genblk1__genblk1__pcpi_mul__mul_counter(
  \genblk1.genblk1.pcpi_mul .mul_counter),
.genblk1__genblk1__pcpi_mul__mul_finish(
  \genblk1.genblk1.pcpi_mul .mul_finish),
.genblk1__genblk1__pcpi_mul__mul_start(
  \genblk1.genblk1.pcpi_mul .mul_start),
.genblk1__genblk1__pcpi_mul__mul_waiting(
  \genblk1.genblk1.pcpi_mul .mul_waiting),
.genblk1__genblk1__pcpi_mul__next_rd(
  \genblk1.genblk1.pcpi_mul .next_rd),
.genblk1__genblk1__pcpi_mul__next_rd_t0(
  \genblk1.genblk1.pcpi_mul .next_rd_t0),
.genblk1__genblk1__pcpi_mul__next_rdt(
  \genblk1.genblk1.pcpi_mul .next_rdt),
.genblk1__genblk1__pcpi_mul__next_rdt_t0(
  \genblk1.genblk1.pcpi_mul .next_rdt_t0),
.genblk1__genblk1__pcpi_mul__pcpi_wait_q(
  \genblk1.genblk1.pcpi_mul .pcpi_wait_q),
.genblk1__genblk1__pcpi_mul__rd(
  \genblk1.genblk1.pcpi_mul .rd),
.genblk1__genblk1__pcpi_mul__rd_t0(
  \genblk1.genblk1.pcpi_mul .rd_t0),
.genblk1__genblk1__pcpi_mul__rdx(
  \genblk1.genblk1.pcpi_mul .rdx),
.genblk1__genblk1__pcpi_mul__rdx_t0(
  \genblk1.genblk1.pcpi_mul .rdx_t0),
.genblk1__genblk1__pcpi_mul__rs1(
  \genblk1.genblk1.pcpi_mul .rs1),
.genblk1__genblk1__pcpi_mul__rs2(
  \genblk1.genblk1.pcpi_mul .rs2),
.genblk1__genblk1__pcpi_mul__rs2_t0(
  \genblk1.genblk1.pcpi_mul .rs2_t0),
.genblk1__genblk1__pcpi_mul__this_rs2(
  \genblk1.genblk1.pcpi_mul .this_rs2),
.genblk1__genblk1__pcpi_mul__this_rs2_t0(
  \genblk1.genblk1.pcpi_mul .this_rs2_t0),
.genblk2__pcpi_div__clk(
  \genblk2.pcpi_div .clk),
.genblk2__pcpi_div__resetn(
  \genblk2.pcpi_div .resetn),
.genblk2__pcpi_div__pcpi_valid(
  \genblk2.pcpi_div .pcpi_valid),
.genblk2__pcpi_div__pcpi_insn(
  \genblk2.pcpi_div .pcpi_insn),
.genblk2__pcpi_div__pcpi_rs1(
  \genblk2.pcpi_div .pcpi_rs1),
.genblk2__pcpi_div__pcpi_rs2(
  \genblk2.pcpi_div .pcpi_rs2),
.genblk2__pcpi_div__pcpi_wr(
  \genblk2.pcpi_div .pcpi_wr),
.genblk2__pcpi_div__pcpi_rd(
  \genblk2.pcpi_div .pcpi_rd),
.genblk2__pcpi_div__pcpi_wait(
  \genblk2.pcpi_div .pcpi_wait),
.genblk2__pcpi_div__pcpi_ready(
  \genblk2.pcpi_div .pcpi_ready),
.genblk2__pcpi_div__pcpi_insn_t0(
  \genblk2.pcpi_div .pcpi_insn_t0),
.genblk2__pcpi_div__pcpi_rd_t0(
  \genblk2.pcpi_div .pcpi_rd_t0),
.genblk2__pcpi_div__pcpi_ready_t0(
  \genblk2.pcpi_div .pcpi_ready_t0),
.genblk2__pcpi_div__pcpi_rs1_t0(
  \genblk2.pcpi_div .pcpi_rs1_t0),
.genblk2__pcpi_div__pcpi_rs2_t0(
  \genblk2.pcpi_div .pcpi_rs2_t0),
.genblk2__pcpi_div__pcpi_valid_t0(
  \genblk2.pcpi_div .pcpi_valid_t0),
.genblk2__pcpi_div__pcpi_wait_t0(
  \genblk2.pcpi_div .pcpi_wait_t0),
.genblk2__pcpi_div__pcpi_wr_t0(
  \genblk2.pcpi_div .pcpi_wr_t0),
.genblk2__pcpi_div__dividend(
  \genblk2.pcpi_div .dividend),
.genblk2__pcpi_div__dividend_t0(
  \genblk2.pcpi_div .dividend_t0),
.genblk2__pcpi_div__divisor(
  \genblk2.pcpi_div .divisor),
.genblk2__pcpi_div__divisor_t0(
  \genblk2.pcpi_div .divisor_t0),
.genblk2__pcpi_div__instr_any_div_rem(
  \genblk2.pcpi_div .instr_any_div_rem),
.genblk2__pcpi_div__instr_div(
  \genblk2.pcpi_div .instr_div),
.genblk2__pcpi_div__instr_divu(
  \genblk2.pcpi_div .instr_divu),
.genblk2__pcpi_div__instr_rem(
  \genblk2.pcpi_div .instr_rem),
.genblk2__pcpi_div__instr_remu(
  \genblk2.pcpi_div .instr_remu),
.genblk2__pcpi_div__outsign(
  \genblk2.pcpi_div .outsign),
.genblk2__pcpi_div__pcpi_wait_q(
  \genblk2.pcpi_div .pcpi_wait_q),
.genblk2__pcpi_div__quotient(
  \genblk2.pcpi_div .quotient),
.genblk2__pcpi_div__quotient_msk(
  \genblk2.pcpi_div .quotient_msk),
.genblk2__pcpi_div__quotient_msk_t0(
  \genblk2.pcpi_div .quotient_msk_t0),
.genblk2__pcpi_div__quotient_t0(
  \genblk2.pcpi_div .quotient_t0),
.genblk2__pcpi_div__running(
  \genblk2.pcpi_div .running),
.genblk2__pcpi_div__start(
  \genblk2.pcpi_div .start),
._1626_(
  _1626_),
._1868_(
  _1868_),
._1870_(
  _1870_),
._1871_(
  _1871_),
._1874_(
  _1874_),
._1886_(
  _1886_),
.genblk1__genblk1__pcpi_mul___820_(
  \genblk1.genblk1.pcpi_mul ._820_)
);
