`include "formal/assumptions/kronos_core_di_asm.sv"
`include "formal/assumptions/kronos_core_ti_asm.sv"
