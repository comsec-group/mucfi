`include "formal/assumptions/picorv32_di_asm.sv"
`include "formal/assumptions/picorv32_ti_asm.sv"
