    asm_no_taint_top_data_ack_t0: assume property(data_ack_t0 == 0);
    asm_no_taint_top_data_rd_data_t0: assume property(data_rd_data_t0 == 0);
    asm_no_taint_top_external_interrupt_t0: assume property(external_interrupt_t0 == 0);
    asm_no_taint_top_instr_ack_t0: assume property(instr_ack_t0 == 0);
    asm_no_taint_top_instr_data_t0: assume property(instr_data_t0 == 0);
    asm_no_taint_top_software_interrupt_t0: assume property(software_interrupt_t0 == 0);
    asm_no_taint_top_timer_interrupt_t0: assume property(timer_interrupt_t0 == 0);