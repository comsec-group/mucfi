module \$paramod$34601000fe8707ce2501f5ed778e152043201712\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _00_;
wire [6:0] _01_;
wire [6:0] _02_;
wire [6:0] _03_;
wire [6:0] _04_;
wire [6:0] _05_;
wire [6:0] _06_;
wire [6:0] _07_;
wire [6:0] _08_;
/* src = "generated/sv2v_out.v:14871.13-14871.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14875.28-14875.37" */
output [6:0] rd_data_o;
reg [6:0] rd_data_o;
/* cellift = 32'd1 */
output [6:0] rd_data_o_t0;
reg [6:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14876.14-14876.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14872.13-14872.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14873.27-14873.36" */
input [6:0] wr_data_i;
wire [6:0] wr_data_i;
/* cellift = 32'd1 */
input [6:0] wr_data_i_t0;
wire [6:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14874.13-14874.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _00_ = ~ wr_en_i;
assign _08_ = wr_data_i ^ rd_data_o;
assign _04_ = wr_data_i_t0 | rd_data_o_t0;
assign _05_ = _08_ | _04_;
assign _01_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _02_ = { _00_, _00_, _00_, _00_, _00_, _00_, _00_ } & rd_data_o_t0;
assign _03_ = _05_ & { wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0 };
assign _06_ = _01_ | _02_;
assign _07_ = _06_ | _03_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$34601000fe8707ce2501f5ed778e152043201712\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 7'h00;
else rd_data_o_t0 <= _07_;
/* src = "generated/sv2v_out.v:14878.2-14882.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$34601000fe8707ce2501f5ed778e152043201712\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 7'h00;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$410b37fbfbfa994790f1902c150d2be939cadb3b\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _00_;
wire [2:0] _01_;
wire [2:0] _02_;
wire [2:0] _03_;
wire [2:0] _04_;
wire [2:0] _05_;
wire [2:0] _06_;
wire [2:0] _07_;
wire [2:0] _08_;
/* src = "generated/sv2v_out.v:14871.13-14871.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14875.28-14875.37" */
output [2:0] rd_data_o;
reg [2:0] rd_data_o;
/* cellift = 32'd1 */
output [2:0] rd_data_o_t0;
reg [2:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14876.14-14876.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14872.13-14872.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14873.27-14873.36" */
input [2:0] wr_data_i;
wire [2:0] wr_data_i;
/* cellift = 32'd1 */
input [2:0] wr_data_i_t0;
wire [2:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14874.13-14874.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _00_ = ~ wr_en_i;
assign _08_ = wr_data_i ^ rd_data_o;
assign _04_ = wr_data_i_t0 | rd_data_o_t0;
assign _05_ = _08_ | _04_;
assign _01_ = { wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _02_ = { _00_, _00_, _00_ } & rd_data_o_t0;
assign _03_ = _05_ & { wr_en_i_t0, wr_en_i_t0, wr_en_i_t0 };
assign _06_ = _01_ | _02_;
assign _07_ = _06_ | _03_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$410b37fbfbfa994790f1902c150d2be939cadb3b\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 3'h0;
else rd_data_o_t0 <= _07_;
/* src = "generated/sv2v_out.v:14878.2-14882.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$410b37fbfbfa994790f1902c150d2be939cadb3b\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 3'h4;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_flop (clk_i, rst_ni, d_i, q_o, d_i_t0, q_o_t0);
/* src = "generated/sv2v_out.v:24647.8-24647.13" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:24649.22-24649.25" */
input [3:0] d_i;
wire [3:0] d_i;
/* cellift = 32'd1 */
input [3:0] d_i_t0;
wire [3:0] d_i_t0;
/* src = "generated/sv2v_out.v:24650.28-24650.31" */
output [3:0] q_o;
wire [3:0] q_o;
/* cellift = 32'd1 */
output [3:0] q_o_t0;
wire [3:0] q_o_t0;
/* src = "generated/sv2v_out.v:24648.8-24648.14" */
input rst_ni;
wire rst_ni;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:24668.6-24673.5" */
\$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_generic_flop  \gen_generic.u_impl_generic  (
.clk_i(clk_i),
.d_i(d_i),
.d_i_t0(d_i_t0),
.q_o(q_o),
.q_o_t0(q_o_t0),
.rst_ni(rst_ni)
);
endmodule

module \$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_generic_flop (clk_i, rst_ni, d_i, q_o, d_i_t0, q_o_t0);
/* src = "generated/sv2v_out.v:24907.8-24907.13" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:24909.22-24909.25" */
input [3:0] d_i;
wire [3:0] d_i;
/* cellift = 32'd1 */
input [3:0] d_i_t0;
wire [3:0] d_i_t0;
/* src = "generated/sv2v_out.v:24910.27-24910.30" */
output [3:0] q_o;
reg [3:0] q_o;
/* cellift = 32'd1 */
output [3:0] q_o_t0;
reg [3:0] q_o_t0;
/* src = "generated/sv2v_out.v:24908.8-24908.14" */
input rst_ni;
wire rst_ni;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_generic_flop  */
/* PC_TAINT_INFO STATE_NAME q_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) q_o_t0 <= 4'h0;
else q_o_t0 <= d_i_t0;
/* src = "generated/sv2v_out.v:24911.2-24915.15" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_generic_flop  */
/* PC_TAINT_INFO STATE_NAME q_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) q_o <= 4'ha;
else q_o <= d_i;
endmodule

module \$paramod$4f46e25470a27719ee9ca03cee1a0827eff766f7\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _00_;
wire [31:0] _01_;
wire [31:0] _02_;
wire [31:0] _03_;
wire [31:0] _04_;
wire [31:0] _05_;
wire [31:0] _06_;
wire [31:0] _07_;
wire [31:0] _08_;
/* src = "generated/sv2v_out.v:14871.13-14871.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14875.28-14875.37" */
output [31:0] rd_data_o;
reg [31:0] rd_data_o;
/* cellift = 32'd1 */
output [31:0] rd_data_o_t0;
reg [31:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14876.14-14876.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14872.13-14872.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14873.27-14873.36" */
input [31:0] wr_data_i;
wire [31:0] wr_data_i;
/* cellift = 32'd1 */
input [31:0] wr_data_i_t0;
wire [31:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14874.13-14874.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _00_ = ~ wr_en_i;
assign _08_ = wr_data_i ^ rd_data_o;
assign _04_ = wr_data_i_t0 | rd_data_o_t0;
assign _05_ = _08_ | _04_;
assign _01_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _02_ = { _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_ } & rd_data_o_t0;
assign _03_ = _05_ & { wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0 };
assign _06_ = _01_ | _02_;
assign _07_ = _06_ | _03_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$4f46e25470a27719ee9ca03cee1a0827eff766f7\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 32'd0;
else rd_data_o_t0 <= _07_;
/* src = "generated/sv2v_out.v:14878.2-14882.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$4f46e25470a27719ee9ca03cee1a0827eff766f7\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 32'd1;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$501c60d7519704ee720c78ef16ad88cf05835059\ibex_dummy_instr (clk_i, rst_ni, dummy_instr_en_i, dummy_instr_mask_i, dummy_instr_seed_en_i, dummy_instr_seed_i, fetch_valid_i, id_in_ready_i, insert_dummy_instr_o, dummy_instr_data_o, insert_dummy_instr_o_t0, id_in_ready_i_t0, fetch_valid_i_t0, dummy_instr_seed_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_mask_i_t0, dummy_instr_en_i_t0, dummy_instr_data_o_t0);
/* src = "generated/sv2v_out.v:15851.25-15851.57" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15851.25-15851.57" */
wire _001_;
wire [4:0] _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire [4:0] _007_;
wire [1:0] _008_;
wire _009_;
wire [1:0] _010_;
wire _011_;
wire _012_;
wire [2:0] _013_;
wire [4:0] _014_;
wire [2:0] _015_;
wire _016_;
wire _017_;
wire _018_;
wire [4:0] _019_;
wire _020_;
wire _021_;
wire _022_;
wire [4:0] _023_;
wire [4:0] _024_;
wire [4:0] _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire [4:0] _035_;
wire [4:0] _036_;
wire [4:0] _037_;
wire [31:0] _038_;
wire [31:0] _039_;
wire [31:0] _040_;
wire [1:0] _041_;
wire [2:0] _042_;
wire [2:0] _043_;
wire [4:0] _044_;
wire [4:0] _045_;
wire _046_;
wire _047_;
wire _048_;
wire [1:0] _049_;
wire [4:0] _050_;
wire [4:0] _051_;
wire [4:0] _052_;
wire _053_;
wire [4:0] _054_;
wire _055_;
wire _056_;
wire _057_;
wire [4:0] _058_;
wire [4:0] _059_;
wire [4:0] _060_;
wire [4:0] _061_;
wire [31:0] _062_;
wire [31:0] _063_;
wire [31:0] _064_;
wire [31:0] _065_;
wire [2:0] _066_;
wire [4:0] _067_;
wire _068_;
wire [4:0] _069_;
wire [4:0] _070_;
wire [4:0] _071_;
wire [31:0] _072_;
wire _073_;
wire _074_;
wire _075_;
wire [4:0] _076_;
wire [4:0] _077_;
wire [2:0] _078_;
/* cellift = 32'd1 */
wire [2:0] _079_;
/* src = "generated/sv2v_out.v:15857.50-15857.84" */
wire _080_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15857.50-15857.84" */
wire _081_;
/* src = "generated/sv2v_out.v:15851.62-15851.96" */
wire _082_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15851.62-15851.96" */
wire _083_;
wire _084_;
/* cellift = 32'd1 */
wire _085_;
wire _086_;
wire _087_;
/* cellift = 32'd1 */
wire _088_;
/* src = "generated/sv2v_out.v:15794.13-15794.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:15810.13-15810.24" */
wire [4:0] dummy_cnt_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15810.13-15810.24" */
wire [4:0] dummy_cnt_d_t0;
/* src = "generated/sv2v_out.v:15812.7-15812.19" */
wire dummy_cnt_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15812.7-15812.19" */
wire dummy_cnt_en_t0;
/* src = "generated/sv2v_out.v:15808.13-15808.27" */
wire [4:0] dummy_cnt_incr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15808.13-15808.27" */
wire [4:0] dummy_cnt_incr_t0;
/* src = "generated/sv2v_out.v:15811.12-15811.23" */
reg [4:0] dummy_cnt_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15811.12-15811.23" */
reg [4:0] dummy_cnt_q_t0;
/* src = "generated/sv2v_out.v:15809.13-15809.32" */
wire [4:0] dummy_cnt_threshold;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15809.13-15809.32" */
wire [4:0] dummy_cnt_threshold_t0;
/* src = "generated/sv2v_out.v:15803.21-15803.39" */
output [31:0] dummy_instr_data_o;
wire [31:0] dummy_instr_data_o;
/* cellift = 32'd1 */
output [31:0] dummy_instr_data_o_t0;
wire [31:0] dummy_instr_data_o_t0;
/* src = "generated/sv2v_out.v:15796.13-15796.29" */
input dummy_instr_en_i;
wire dummy_instr_en_i;
/* cellift = 32'd1 */
input dummy_instr_en_i_t0;
wire dummy_instr_en_i_t0;
/* src = "generated/sv2v_out.v:15797.19-15797.37" */
input [2:0] dummy_instr_mask_i;
wire [2:0] dummy_instr_mask_i;
/* cellift = 32'd1 */
input [2:0] dummy_instr_mask_i_t0;
wire [2:0] dummy_instr_mask_i_t0;
/* src = "generated/sv2v_out.v:15820.14-15820.32" */
wire [31:0] dummy_instr_seed_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15820.14-15820.32" */
wire [31:0] dummy_instr_seed_d_t0;
/* src = "generated/sv2v_out.v:15798.13-15798.34" */
input dummy_instr_seed_en_i;
wire dummy_instr_seed_en_i;
/* cellift = 32'd1 */
input dummy_instr_seed_en_i_t0;
wire dummy_instr_seed_en_i_t0;
/* src = "generated/sv2v_out.v:15799.20-15799.38" */
input [31:0] dummy_instr_seed_i;
wire [31:0] dummy_instr_seed_i;
/* cellift = 32'd1 */
input [31:0] dummy_instr_seed_i_t0;
wire [31:0] dummy_instr_seed_i_t0;
/* src = "generated/sv2v_out.v:15819.13-15819.31" */
reg [31:0] dummy_instr_seed_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15819.13-15819.31" */
reg [31:0] dummy_instr_seed_q_t0;
/* src = "generated/sv2v_out.v:15817.12-15817.24" */
wire [2:0] dummy_opcode;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15817.12-15817.24" */
wire [2:0] dummy_opcode_t0;
/* src = "generated/sv2v_out.v:15816.12-15816.21" */
wire [6:0] dummy_set;
/* src = "generated/sv2v_out.v:15800.13-15800.26" */
input fetch_valid_i;
wire fetch_valid_i;
/* cellift = 32'd1 */
input fetch_valid_i_t0;
wire fetch_valid_i_t0;
/* src = "generated/sv2v_out.v:15801.13-15801.26" */
input id_in_ready_i;
wire id_in_ready_i;
/* cellift = 32'd1 */
input id_in_ready_i_t0;
wire id_in_ready_i_t0;
/* src = "generated/sv2v_out.v:15802.14-15802.34" */
output insert_dummy_instr_o;
wire insert_dummy_instr_o;
/* cellift = 32'd1 */
output insert_dummy_instr_o_t0;
wire insert_dummy_instr_o_t0;
/* src = "generated/sv2v_out.v:15807.14-15807.23" */
wire [16:0] lfsr_data;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15807.14-15807.23" */
wire [16:0] lfsr_data_t0;
/* src = "generated/sv2v_out.v:15813.7-15813.14" */
wire lfsr_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15813.7-15813.14" */
wire lfsr_en_t0;
/* src = "generated/sv2v_out.v:15795.13-15795.19" */
input rst_ni;
wire rst_ni;
assign dummy_cnt_incr = dummy_cnt_q + /* src = "generated/sv2v_out.v:15849.26-15849.58" */ 5'h01;
assign lfsr_en = insert_dummy_instr_o & /* src = "generated/sv2v_out.v:15821.19-15821.53" */ id_in_ready_i;
assign dummy_cnt_threshold = lfsr_data[4:0] & /* src = "generated/sv2v_out.v:15848.31-15848.93" */ { dummy_instr_mask_i, 2'h3 };
assign _000_ = dummy_instr_en_i & /* src = "generated/sv2v_out.v:15851.25-15851.57" */ id_in_ready_i;
assign dummy_cnt_en = _000_ & /* src = "generated/sv2v_out.v:15851.24-15851.97" */ _082_;
assign insert_dummy_instr_o = dummy_instr_en_i & /* src = "generated/sv2v_out.v:15857.30-15857.85" */ _080_;
assign _002_ = ~ dummy_cnt_q_t0;
assign _019_ = dummy_cnt_q & _002_;
assign _076_ = _019_ + 5'h01;
assign _052_ = dummy_cnt_q | dummy_cnt_q_t0;
assign _077_ = _052_ + 5'h01;
assign _070_ = _076_ ^ _077_;
assign dummy_cnt_incr_t0 = _070_ | dummy_cnt_q_t0;
assign _003_ = ~ dummy_cnt_en;
assign _004_ = ~ dummy_instr_seed_en_i;
assign _071_ = dummy_cnt_d ^ dummy_cnt_q;
assign _072_ = dummy_instr_seed_d ^ dummy_instr_seed_q;
assign _058_ = dummy_cnt_d_t0 | dummy_cnt_q_t0;
assign _062_ = dummy_instr_seed_d_t0 | dummy_instr_seed_q_t0;
assign _059_ = _071_ | _058_;
assign _063_ = _072_ | _062_;
assign _035_ = { dummy_cnt_en, dummy_cnt_en, dummy_cnt_en, dummy_cnt_en, dummy_cnt_en } & dummy_cnt_d_t0;
assign _038_ = { dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i, dummy_instr_seed_en_i } & dummy_instr_seed_d_t0;
assign _036_ = { _003_, _003_, _003_, _003_, _003_ } & dummy_cnt_q_t0;
assign _039_ = { _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_ } & dummy_instr_seed_q_t0;
assign _037_ = _059_ & { dummy_cnt_en_t0, dummy_cnt_en_t0, dummy_cnt_en_t0, dummy_cnt_en_t0, dummy_cnt_en_t0 };
assign _040_ = _063_ & { dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_seed_en_i_t0 };
assign _060_ = _035_ | _036_;
assign _064_ = _038_ | _039_;
assign _061_ = _060_ | _037_;
assign _065_ = _064_ | _040_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$501c60d7519704ee720c78ef16ad88cf05835059\ibex_dummy_instr  */
/* PC_TAINT_INFO STATE_NAME dummy_cnt_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_cnt_q_t0 <= 5'h00;
else dummy_cnt_q_t0 <= _061_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$501c60d7519704ee720c78ef16ad88cf05835059\ibex_dummy_instr  */
/* PC_TAINT_INFO STATE_NAME dummy_instr_seed_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_instr_seed_q_t0 <= 32'd0;
else dummy_instr_seed_q_t0 <= _065_;
assign _020_ = insert_dummy_instr_o_t0 & id_in_ready_i;
assign _023_ = lfsr_data_t0[4:0] & { dummy_instr_mask_i, 2'h3 };
assign _026_ = dummy_instr_en_i_t0 & id_in_ready_i;
assign _029_ = _001_ & _082_;
assign _032_ = dummy_instr_en_i_t0 & _080_;
assign _021_ = id_in_ready_i_t0 & insert_dummy_instr_o;
assign _024_ = { dummy_instr_mask_i_t0, 2'h0 } & lfsr_data[4:0];
assign _027_ = id_in_ready_i_t0 & dummy_instr_en_i;
assign _030_ = _083_ & _000_;
assign _033_ = _081_ & dummy_instr_en_i;
assign _022_ = insert_dummy_instr_o_t0 & id_in_ready_i_t0;
assign _025_ = lfsr_data_t0[4:0] & { dummy_instr_mask_i_t0, 2'h0 };
assign _028_ = dummy_instr_en_i_t0 & id_in_ready_i_t0;
assign _031_ = _001_ & _083_;
assign _034_ = dummy_instr_en_i_t0 & _081_;
assign _053_ = _020_ | _021_;
assign _054_ = _023_ | _024_;
assign _055_ = _026_ | _027_;
assign _056_ = _029_ | _030_;
assign _057_ = _032_ | _033_;
assign lfsr_en_t0 = _053_ | _022_;
assign dummy_cnt_threshold_t0 = _054_ | _025_;
assign _001_ = _055_ | _028_;
assign dummy_cnt_en_t0 = _056_ | _031_;
assign insert_dummy_instr_o_t0 = _057_ | _034_;
assign _005_ = | { dummy_cnt_q_t0, dummy_cnt_threshold_t0 };
assign _006_ = | lfsr_data_t0[16:15];
assign _067_ = dummy_cnt_q_t0 | dummy_cnt_threshold_t0;
assign _007_ = ~ _067_;
assign _008_ = ~ lfsr_data_t0[16:15];
assign _044_ = dummy_cnt_q & _007_;
assign _049_ = lfsr_data[16:15] & _008_;
assign _045_ = dummy_cnt_threshold & _007_;
assign _073_ = _044_ == _045_;
assign _074_ = _049_ == _008_;
assign _075_ = _049_ == { _008_[1], 1'h0 };
assign _081_ = _073_ & _005_;
assign _085_ = _074_ & _006_;
assign _079_[2] = _075_ & _006_;
/* src = "generated/sv2v_out.v:15852.2-15856.31" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$501c60d7519704ee720c78ef16ad88cf05835059\ibex_dummy_instr  */
/* PC_TAINT_INFO STATE_NAME dummy_cnt_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_cnt_q <= 5'h00;
else if (dummy_cnt_en) dummy_cnt_q <= dummy_cnt_d;
/* src = "generated/sv2v_out.v:15823.2-15827.45" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$501c60d7519704ee720c78ef16ad88cf05835059\ibex_dummy_instr  */
/* PC_TAINT_INFO STATE_NAME dummy_instr_seed_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_instr_seed_q <= 32'd0;
else if (dummy_instr_seed_en_i) dummy_instr_seed_q <= dummy_instr_seed_d;
assign _009_ = | { _085_, _088_ };
assign _010_ = ~ { _088_, _085_ };
assign _041_ = { _087_, _084_ } & _010_;
assign _011_ = ! _041_;
assign _012_ = ! _049_;
assign dummy_instr_data_o_t0[25] = _011_ & _009_;
assign _088_ = _012_ & _006_;
assign _013_ = ~ { _084_, _084_, _084_ };
assign _014_ = ~ { insert_dummy_instr_o, insert_dummy_instr_o, insert_dummy_instr_o, insert_dummy_instr_o, insert_dummy_instr_o };
assign _066_ = { _085_, _085_, _085_ } | _013_;
assign _069_ = { insert_dummy_instr_o_t0, insert_dummy_instr_o_t0, insert_dummy_instr_o_t0, insert_dummy_instr_o_t0, insert_dummy_instr_o_t0 } | _014_;
assign _042_ = { _079_[2], 2'h0 } & _066_;
assign _050_ = dummy_cnt_incr_t0 & _069_;
assign _043_ = { _085_, _085_, _085_ } & _015_;
assign _051_ = { insert_dummy_instr_o_t0, insert_dummy_instr_o_t0, insert_dummy_instr_o_t0, insert_dummy_instr_o_t0, insert_dummy_instr_o_t0 } & dummy_cnt_incr;
assign dummy_opcode_t0 = _043_ | _042_;
assign dummy_cnt_d_t0 = _051_ | _050_;
assign _015_ = ~ _078_;
assign _018_ = | { _087_, _084_ };
assign _016_ = ~ fetch_valid_i;
assign _017_ = ~ insert_dummy_instr_o;
assign _046_ = fetch_valid_i_t0 & _017_;
assign _047_ = insert_dummy_instr_o_t0 & _016_;
assign _048_ = fetch_valid_i_t0 & insert_dummy_instr_o_t0;
assign _068_ = _046_ | _047_;
assign _083_ = _068_ | _048_;
assign _078_ = _086_ ? 3'h4 : 3'h0;
assign dummy_opcode = _084_ ? 3'h7 : _078_;
assign dummy_set = _018_ ? 7'h00 : 7'h01;
assign dummy_instr_seed_d_t0 = dummy_instr_seed_q_t0 | dummy_instr_seed_i_t0;
assign _080_ = dummy_cnt_q == /* src = "generated/sv2v_out.v:15857.50-15857.84" */ dummy_cnt_threshold;
assign _082_ = fetch_valid_i | /* src = "generated/sv2v_out.v:15851.62-15851.96" */ insert_dummy_instr_o;
assign _084_ = lfsr_data[16:15] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15859.3-15880.10" */ 2'h3;
assign _086_ = lfsr_data[16:15] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15859.3-15880.10" */ 2'h2;
assign _087_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15859.3-15880.10" */ lfsr_data[16:15];
assign dummy_cnt_d = insert_dummy_instr_o ? /* src = "generated/sv2v_out.v:15850.24-15850.73" */ 5'h00 : dummy_cnt_incr;
assign dummy_instr_seed_d = dummy_instr_seed_q ^ /* src = "generated/sv2v_out.v:15822.30-15822.69" */ dummy_instr_seed_i;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:15834.4-15842.3" */
\$paramod$5fd3ce2f8a67228d339c5f62898ff83b3c2a14f0\prim_lfsr  lfsr_i (
.clk_i(clk_i),
.entropy_i(8'h00),
.entropy_i_t0(8'h00),
.lfsr_en_i(lfsr_en),
.lfsr_en_i_t0(lfsr_en_t0),
.rst_ni(rst_ni),
.seed_en_i(dummy_instr_seed_en_i),
.seed_en_i_t0(dummy_instr_seed_en_i_t0),
.seed_i(dummy_instr_seed_d),
.seed_i_t0(dummy_instr_seed_d_t0),
.state_o(lfsr_data),
.state_o_t0(lfsr_data_t0)
);
assign _079_[1:0] = 2'h0;
assign dummy_instr_data_o = { dummy_set, lfsr_data[14:5], dummy_opcode, 12'h033 };
assign { dummy_instr_data_o_t0[31:26], dummy_instr_data_o_t0[24:0] } = { 6'h00, lfsr_data_t0[14:5], dummy_opcode_t0, 12'h000 };
endmodule

module \$paramod$5714e31d82f2b8816750797f158ebea69a089104\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _00_;
wire [5:0] _01_;
wire [5:0] _02_;
wire [5:0] _03_;
wire [5:0] _04_;
wire [5:0] _05_;
wire [5:0] _06_;
wire [5:0] _07_;
wire [5:0] _08_;
/* src = "generated/sv2v_out.v:14871.13-14871.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14875.28-14875.37" */
output [5:0] rd_data_o;
reg [5:0] rd_data_o;
/* cellift = 32'd1 */
output [5:0] rd_data_o_t0;
reg [5:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14876.14-14876.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14872.13-14872.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14873.27-14873.36" */
input [5:0] wr_data_i;
wire [5:0] wr_data_i;
/* cellift = 32'd1 */
input [5:0] wr_data_i_t0;
wire [5:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14874.13-14874.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _00_ = ~ wr_en_i;
assign _08_ = wr_data_i ^ rd_data_o;
assign _04_ = wr_data_i_t0 | rd_data_o_t0;
assign _05_ = _08_ | _04_;
assign _01_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _02_ = { _00_, _00_, _00_, _00_, _00_, _00_ } & rd_data_o_t0;
assign _03_ = _05_ & { wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0 };
assign _06_ = _01_ | _02_;
assign _07_ = _06_ | _03_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$5714e31d82f2b8816750797f158ebea69a089104\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 6'h00;
else rd_data_o_t0 <= _07_;
/* src = "generated/sv2v_out.v:14878.2-14882.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$5714e31d82f2b8816750797f158ebea69a089104\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 6'h10;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$5c0dc9f9e0551018f7d8916b4fcabdef94a17390\ibex_core (clk_i, rst_ni, hart_id_i, boot_addr_i, instr_req_o, instr_gnt_i, instr_rvalid_i, instr_addr_o, instr_rdata_i, instr_err_i, data_req_o, data_gnt_i, data_rvalid_i, data_we_o, data_be_o, data_addr_o, data_wdata_o, data_rdata_i, data_err_i, dummy_instr_id_o, dummy_instr_wb_o
, rf_raddr_a_o, rf_raddr_b_o, rf_waddr_wb_o, rf_we_wb_o, rf_wdata_wb_ecc_o, rf_rdata_a_ecc_i, rf_rdata_b_ecc_i, ic_tag_req_o, ic_tag_write_o, ic_tag_addr_o, ic_tag_wdata_o, ic_tag_rdata_i, ic_data_req_o, ic_data_write_o, ic_data_addr_o, ic_data_wdata_o, ic_data_rdata_i, ic_scr_key_valid_i, ic_scr_key_req_o, irq_software_i, irq_timer_i
, irq_external_i, irq_fast_i, irq_nm_i, irq_pending_o, debug_req_i, crash_dump_o, double_fault_seen_o, fetch_enable_i, alert_minor_o, alert_major_internal_o, alert_major_bus_o, core_busy_o, rf_raddr_b_o_t0, rf_raddr_a_o_t0, data_we_o_t0, data_req_o_t0, debug_req_i_t0, ic_tag_write_o_t0, ic_tag_wdata_o_t0, ic_tag_req_o_t0, ic_tag_rdata_i_t0
, ic_tag_addr_o_t0, ic_scr_key_valid_i_t0, ic_scr_key_req_o_t0, ic_data_write_o_t0, ic_data_wdata_o_t0, ic_data_req_o_t0, ic_data_rdata_i_t0, ic_data_addr_o_t0, dummy_instr_id_o_t0, boot_addr_i_t0, instr_rvalid_i_t0, instr_req_o_t0, instr_rdata_i_t0, instr_gnt_i_t0, instr_err_i_t0, instr_addr_o_t0, irq_nm_i_t0, data_addr_o_t0, data_be_o_t0, data_gnt_i_t0, data_rdata_i_t0
, data_rvalid_i_t0, data_wdata_o_t0, dummy_instr_wb_o_t0, rf_waddr_wb_o_t0, rf_we_wb_o_t0, double_fault_seen_o_t0, hart_id_i_t0, irq_external_i_t0, irq_fast_i_t0, irq_pending_o_t0, irq_software_i_t0, irq_timer_i_t0, alert_major_bus_o_t0, alert_major_internal_o_t0, alert_minor_o_t0, core_busy_o_t0, crash_dump_o_t0, data_err_i_t0, fetch_enable_i_t0, rf_rdata_a_ecc_i_t0, rf_rdata_b_ecc_i_t0
, rf_wdata_wb_ecc_o_t0);
/* src = "generated/sv2v_out.v:13414.30-13414.54" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13414.30-13414.54" */
wire _001_;
/* src = "generated/sv2v_out.v:13415.30-13415.54" */
wire _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13415.30-13415.54" */
wire _003_;
wire _004_;
wire [3:0] _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire [2:0] _012_;
wire [2:0] _013_;
wire [2:0] _014_;
wire [2:0] _015_;
wire [1:0] _016_;
wire [1:0] _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire [3:0] _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire [2:0] _076_;
wire [2:0] _077_;
wire [2:0] _078_;
wire [2:0] _079_;
wire [1:0] _080_;
wire [1:0] _081_;
wire [11:0] _082_;
wire [11:0] _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire [11:0] _097_;
wire _098_;
/* src = "generated/sv2v_out.v:13141.41-13141.56" */
wire _099_;
/* src = "generated/sv2v_out.v:13414.58-13414.75" */
wire _100_;
/* src = "generated/sv2v_out.v:13415.58-13415.75" */
wire _101_;
/* src = "generated/sv2v_out.v:13416.47-13416.80" */
wire _102_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13416.47-13416.80" */
wire _103_;
/* src = "generated/sv2v_out.v:13440.35-13440.70" */
wire _104_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13440.35-13440.70" */
wire _105_;
/* src = "generated/sv2v_out.v:13441.30-13441.78" */
wire _106_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13441.30-13441.78" */
wire _107_;
/* src = "generated/sv2v_out.v:13053.30-13053.81" */
wire _108_;
/* src = "generated/sv2v_out.v:13053.30-13053.81" */
wire _109_;
/* src = "generated/sv2v_out.v:13414.30-13414.43" */
wire _110_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13414.30-13414.43" */
wire _111_;
/* src = "generated/sv2v_out.v:13415.30-13415.43" */
wire _112_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13415.30-13415.43" */
wire _113_;
/* src = "generated/sv2v_out.v:12874.14-12874.31" */
output alert_major_bus_o;
wire alert_major_bus_o;
/* cellift = 32'd1 */
output alert_major_bus_o_t0;
wire alert_major_bus_o_t0;
/* src = "generated/sv2v_out.v:12873.14-12873.36" */
output alert_major_internal_o;
wire alert_major_internal_o;
/* cellift = 32'd1 */
output alert_major_internal_o_t0;
wire alert_major_internal_o_t0;
/* src = "generated/sv2v_out.v:12872.14-12872.27" */
output alert_minor_o;
wire alert_minor_o;
/* cellift = 32'd1 */
output alert_minor_o_t0;
wire alert_minor_o_t0;
/* src = "generated/sv2v_out.v:12951.14-12951.33" */
wire [31:0] alu_adder_result_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12951.14-12951.33" */
wire [31:0] alu_adder_result_ex_t0;
/* src = "generated/sv2v_out.v:12947.14-12947.30" */
wire [31:0] alu_operand_a_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12947.14-12947.30" */
wire [31:0] alu_operand_a_ex_t0;
/* src = "generated/sv2v_out.v:12948.14-12948.30" */
wire [31:0] alu_operand_b_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12948.14-12948.30" */
wire [31:0] alu_operand_b_ex_t0;
/* src = "generated/sv2v_out.v:12946.13-12946.28" */
wire [6:0] alu_operator_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12946.13-12946.28" */
wire [6:0] alu_operator_ex_t0;
/* src = "generated/sv2v_out.v:12825.20-12825.31" */
input [31:0] boot_addr_i;
wire [31:0] boot_addr_i;
/* cellift = 32'd1 */
input [31:0] boot_addr_i_t0;
wire [31:0] boot_addr_i_t0;
/* src = "generated/sv2v_out.v:12924.7-12924.22" */
wire branch_decision;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12924.7-12924.22" */
wire branch_decision_t0;
/* src = "generated/sv2v_out.v:12923.14-12923.30" */
wire [31:0] branch_target_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12923.14-12923.30" */
wire [31:0] branch_target_ex_t0;
/* src = "generated/sv2v_out.v:12949.14-12949.26" */
wire [31:0] bt_a_operand;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12949.14-12949.26" */
wire [31:0] bt_a_operand_t0;
/* src = "generated/sv2v_out.v:12950.14-12950.26" */
wire [31:0] bt_b_operand;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12950.14-12950.26" */
wire [31:0] bt_b_operand_t0;
/* src = "generated/sv2v_out.v:12822.13-12822.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:12875.20-12875.31" */
output [3:0] core_busy_o;
wire [3:0] core_busy_o;
/* cellift = 32'd1 */
output [3:0] core_busy_o_t0;
wire [3:0] core_busy_o_t0;
/* src = "generated/sv2v_out.v:13433.14-13433.30" */
wire [31:0] crash_dump_mtval;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13433.14-13433.30" */
wire [31:0] crash_dump_mtval_t0;
/* src = "generated/sv2v_out.v:12869.22-12869.34" */
output [159:0] crash_dump_o;
wire [159:0] crash_dump_o;
/* cellift = 32'd1 */
output [159:0] crash_dump_o_t0;
wire [159:0] crash_dump_o_t0;
/* src = "generated/sv2v_out.v:12962.7-12962.17" */
wire csr_access;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12962.7-12962.17" */
wire csr_access_t0;
/* src = "generated/sv2v_out.v:12965.14-12965.22" */
wire [11:0] csr_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12965.14-12965.22" */
wire [11:0] csr_addr_t0;
/* src = "generated/sv2v_out.v:12993.14-12993.22" */
wire [31:0] csr_depc;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12993.14-12993.22" */
wire [31:0] csr_depc_t0;
/* src = "generated/sv2v_out.v:12992.14-12992.22" */
wire [31:0] csr_mepc;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12992.14-12992.22" */
wire [31:0] csr_mepc_t0;
/* src = "generated/sv2v_out.v:12991.7-12991.22" */
wire csr_mstatus_mie;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12991.7-12991.22" */
wire csr_mstatus_mie_t0;
/* src = "generated/sv2v_out.v:13008.7-13008.21" */
wire csr_mstatus_tw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13008.7-13008.21" */
wire csr_mstatus_tw_t0;
/* src = "generated/sv2v_out.v:13007.14-13007.23" */
wire [31:0] csr_mtval;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13007.14-13007.23" */
wire [31:0] csr_mtval_t0;
/* src = "generated/sv2v_out.v:13006.14-13006.23" */
wire [31:0] csr_mtvec;
/* src = "generated/sv2v_out.v:13005.7-13005.21" */
wire csr_mtvec_init;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13005.7-13005.21" */
wire csr_mtvec_init_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13006.14-13006.23" */
wire [31:0] csr_mtvec_t0;
/* src = "generated/sv2v_out.v:12963.13-12963.19" */
wire [1:0] csr_op;
/* src = "generated/sv2v_out.v:12964.7-12964.16" */
wire csr_op_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12964.7-12964.16" */
wire csr_op_en_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12963.13-12963.19" */
wire [1:0] csr_op_t0;
/* src = "generated/sv2v_out.v:12994.36-12994.48" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135" */
wire [135:0] csr_pmp_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12994.36-12994.48" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135" */
wire [135:0] csr_pmp_addr_t0;
/* src = "generated/sv2v_out.v:12995.35-12995.46" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23" */
wire [23:0] csr_pmp_cfg;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12995.35-12995.46" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23" */
wire [23:0] csr_pmp_cfg_t0;
/* src = "generated/sv2v_out.v:12996.13-12996.28" */
/* unused_bits = "0 1 2" */
wire [2:0] csr_pmp_mseccfg;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12996.13-12996.28" */
/* unused_bits = "0 1 2" */
wire [2:0] csr_pmp_mseccfg_t0;
/* src = "generated/sv2v_out.v:12966.14-12966.23" */
wire [31:0] csr_rdata;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12966.14-12966.23" */
wire [31:0] csr_rdata_t0;
/* src = "generated/sv2v_out.v:13003.7-13003.26" */
wire csr_restore_dret_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13003.7-13003.26" */
wire csr_restore_dret_id_t0;
/* src = "generated/sv2v_out.v:13002.7-13002.26" */
wire csr_restore_mret_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13002.7-13002.26" */
wire csr_restore_mret_id_t0;
/* src = "generated/sv2v_out.v:13004.7-13004.21" */
wire csr_save_cause;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13004.7-13004.21" */
wire csr_save_cause_t0;
/* src = "generated/sv2v_out.v:13000.7-13000.18" */
wire csr_save_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13000.7-13000.18" */
wire csr_save_id_t0;
/* src = "generated/sv2v_out.v:12999.7-12999.18" */
wire csr_save_if;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12999.7-12999.18" */
wire csr_save_if_t0;
/* src = "generated/sv2v_out.v:13001.7-13001.18" */
wire csr_save_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13001.7-13001.18" */
wire csr_save_wb_t0;
/* src = "generated/sv2v_out.v:12907.7-12907.21" */
wire csr_shadow_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12907.7-12907.21" */
wire csr_shadow_err_t0;
/* src = "generated/sv2v_out.v:12925.7-12925.16" */
wire ctrl_busy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12925.7-12925.16" */
wire ctrl_busy_t0;
/* src = "generated/sv2v_out.v:12837.21-12837.32" */
output [31:0] data_addr_o;
wire [31:0] data_addr_o;
/* cellift = 32'd1 */
output [31:0] data_addr_o_t0;
wire [31:0] data_addr_o_t0;
/* src = "generated/sv2v_out.v:12836.20-12836.29" */
output [3:0] data_be_o;
wire [3:0] data_be_o;
/* cellift = 32'd1 */
output [3:0] data_be_o_t0;
wire [3:0] data_be_o_t0;
/* src = "generated/sv2v_out.v:12840.13-12840.23" */
input data_err_i;
wire data_err_i;
/* cellift = 32'd1 */
input data_err_i_t0;
wire data_err_i_t0;
/* src = "generated/sv2v_out.v:12833.13-12833.23" */
input data_gnt_i;
wire data_gnt_i;
/* cellift = 32'd1 */
input data_gnt_i_t0;
wire data_gnt_i_t0;
/* src = "generated/sv2v_out.v:12898.7-12898.22" */
wire data_ind_timing;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12898.7-12898.22" */
wire data_ind_timing_t0;
/* src = "generated/sv2v_out.v:12839.34-12839.46" */
input [38:0] data_rdata_i;
wire [38:0] data_rdata_i;
/* cellift = 32'd1 */
input [38:0] data_rdata_i_t0;
wire [38:0] data_rdata_i_t0;
/* src = "generated/sv2v_out.v:12832.14-12832.24" */
output data_req_o;
wire data_req_o;
/* cellift = 32'd1 */
output data_req_o_t0;
wire data_req_o_t0;
/* src = "generated/sv2v_out.v:12834.13-12834.26" */
input data_rvalid_i;
wire data_rvalid_i;
/* cellift = 32'd1 */
input data_rvalid_i_t0;
wire data_rvalid_i_t0;
/* src = "generated/sv2v_out.v:12838.35-12838.47" */
output [38:0] data_wdata_o;
wire [38:0] data_wdata_o;
/* cellift = 32'd1 */
output [38:0] data_wdata_o_t0;
wire [38:0] data_wdata_o_t0;
/* src = "generated/sv2v_out.v:12835.14-12835.23" */
output data_we_o;
wire data_we_o;
/* cellift = 32'd1 */
output data_we_o_t0;
wire data_we_o_t0;
/* src = "generated/sv2v_out.v:13013.13-13013.24" */
wire [2:0] debug_cause;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13013.13-13013.24" */
wire [2:0] debug_cause_t0;
/* src = "generated/sv2v_out.v:13014.7-13014.21" */
wire debug_csr_save;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13014.7-13014.21" */
wire debug_csr_save_t0;
/* src = "generated/sv2v_out.v:13016.7-13016.20" */
wire debug_ebreakm;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13016.7-13016.20" */
wire debug_ebreakm_t0;
/* src = "generated/sv2v_out.v:13017.7-13017.20" */
wire debug_ebreaku;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13017.7-13017.20" */
wire debug_ebreaku_t0;
/* src = "generated/sv2v_out.v:13011.7-13011.17" */
wire debug_mode;
/* src = "generated/sv2v_out.v:13012.7-13012.26" */
wire debug_mode_entering;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13012.7-13012.26" */
wire debug_mode_entering_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13011.7-13011.17" */
wire debug_mode_t0;
/* src = "generated/sv2v_out.v:12868.13-12868.24" */
input debug_req_i;
wire debug_req_i;
/* cellift = 32'd1 */
input debug_req_i_t0;
wire debug_req_i_t0;
/* src = "generated/sv2v_out.v:13015.7-13015.24" */
wire debug_single_step;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13015.7-13015.24" */
wire debug_single_step_t0;
/* src = "generated/sv2v_out.v:12954.7-12954.16" */
wire div_en_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12954.7-12954.16" */
wire div_en_ex_t0;
/* src = "generated/sv2v_out.v:12956.7-12956.17" */
wire div_sel_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12956.7-12956.17" */
wire div_sel_ex_t0;
/* src = "generated/sv2v_out.v:12870.14-12870.33" */
output double_fault_seen_o;
wire double_fault_seen_o;
/* cellift = 32'd1 */
output double_fault_seen_o_t0;
wire double_fault_seen_o_t0;
/* src = "generated/sv2v_out.v:12899.7-12899.21" */
wire dummy_instr_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12899.7-12899.21" */
wire dummy_instr_en_t0;
/* src = "generated/sv2v_out.v:12841.14-12841.30" */
output dummy_instr_id_o;
wire dummy_instr_id_o;
/* cellift = 32'd1 */
output dummy_instr_id_o_t0;
wire dummy_instr_id_o_t0;
/* src = "generated/sv2v_out.v:12900.13-12900.29" */
wire [2:0] dummy_instr_mask;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12900.13-12900.29" */
wire [2:0] dummy_instr_mask_t0;
/* src = "generated/sv2v_out.v:12902.14-12902.30" */
wire [31:0] dummy_instr_seed;
/* src = "generated/sv2v_out.v:12901.7-12901.26" */
wire dummy_instr_seed_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12901.7-12901.26" */
wire dummy_instr_seed_en_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12902.14-12902.30" */
wire [31:0] dummy_instr_seed_t0;
/* src = "generated/sv2v_out.v:12842.14-12842.30" */
output dummy_instr_wb_o;
wire dummy_instr_wb_o;
/* cellift = 32'd1 */
output dummy_instr_wb_o_t0;
wire dummy_instr_wb_o_t0;
/* src = "generated/sv2v_out.v:12982.7-12982.12" */
wire en_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12982.7-12982.12" */
wire en_wb_t0;
/* src = "generated/sv2v_out.v:12976.7-12976.15" */
wire ex_valid;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12976.7-12976.15" */
wire ex_valid_t0;
/* src = "generated/sv2v_out.v:12915.13-12915.22" */
wire [6:0] exc_cause;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12915.13-12915.22" */
wire [6:0] exc_cause_t0;
/* src = "generated/sv2v_out.v:12914.13-12914.26" */
wire [1:0] exc_pc_mux_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12914.13-12914.26" */
wire [1:0] exc_pc_mux_id_t0;
/* src = "generated/sv2v_out.v:12871.19-12871.33" */
input [3:0] fetch_enable_i;
wire [3:0] fetch_enable_i;
/* cellift = 32'd1 */
input [3:0] fetch_enable_i_t0;
wire [3:0] fetch_enable_i_t0;
/* src = "generated/sv2v_out.v:13042.16-13042.29" */
wire [11:0] \g_core_busy_secure.busy_bits_buf ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13042.16-13042.29" */
wire [11:0] \g_core_busy_secure.busy_bits_buf_t0 ;
/* src = "generated/sv2v_out.v:13567.15-13567.33" */
/* unused_bits = "0 1" */
wire [1:0] \g_no_pmp.unused_priv_lvl_ls ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13567.15-13567.33" */
/* unused_bits = "0 1" */
wire [1:0] \g_no_pmp.unused_priv_lvl_ls_t0 ;
/* src = "generated/sv2v_out.v:13396.15-13396.27" */
wire [1:0] \gen_regfile_ecc.rf_ecc_err_a ;
/* src = "generated/sv2v_out.v:13398.9-13398.24" */
wire \gen_regfile_ecc.rf_ecc_err_a_id ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13398.9-13398.24" */
wire \gen_regfile_ecc.rf_ecc_err_a_id_t0 ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13396.15-13396.27" */
wire [1:0] \gen_regfile_ecc.rf_ecc_err_a_t0 ;
/* src = "generated/sv2v_out.v:13397.15-13397.27" */
wire [1:0] \gen_regfile_ecc.rf_ecc_err_b ;
/* src = "generated/sv2v_out.v:13399.9-13399.24" */
wire \gen_regfile_ecc.rf_ecc_err_b_id ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13399.9-13399.24" */
wire \gen_regfile_ecc.rf_ecc_err_b_id_t0 ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13397.15-13397.27" */
wire [1:0] \gen_regfile_ecc.rf_ecc_err_b_t0 ;
/* src = "generated/sv2v_out.v:12824.20-12824.29" */
input [31:0] hart_id_i;
wire [31:0] hart_id_i;
/* cellift = 32'd1 */
input [31:0] hart_id_i_t0;
wire [31:0] hart_id_i_t0;
/* src = "generated/sv2v_out.v:12857.42-12857.56" */
output [7:0] ic_data_addr_o;
wire [7:0] ic_data_addr_o;
/* cellift = 32'd1 */
output [7:0] ic_data_addr_o_t0;
wire [7:0] ic_data_addr_o_t0;
/* src = "generated/sv2v_out.v:12859.58-12859.73" */
input [127:0] ic_data_rdata_i;
wire [127:0] ic_data_rdata_i;
/* cellift = 32'd1 */
input [127:0] ic_data_rdata_i_t0;
wire [127:0] ic_data_rdata_i_t0;
/* src = "generated/sv2v_out.v:12855.20-12855.33" */
output [1:0] ic_data_req_o;
wire [1:0] ic_data_req_o;
/* cellift = 32'd1 */
output [1:0] ic_data_req_o_t0;
wire [1:0] ic_data_req_o_t0;
/* src = "generated/sv2v_out.v:12858.34-12858.49" */
output [63:0] ic_data_wdata_o;
wire [63:0] ic_data_wdata_o;
/* cellift = 32'd1 */
output [63:0] ic_data_wdata_o_t0;
wire [63:0] ic_data_wdata_o_t0;
/* src = "generated/sv2v_out.v:12856.14-12856.29" */
output ic_data_write_o;
wire ic_data_write_o;
/* cellift = 32'd1 */
output ic_data_write_o_t0;
wire ic_data_write_o_t0;
/* src = "generated/sv2v_out.v:12861.14-12861.30" */
output ic_scr_key_req_o;
wire ic_scr_key_req_o;
/* cellift = 32'd1 */
output ic_scr_key_req_o_t0;
wire ic_scr_key_req_o_t0;
/* src = "generated/sv2v_out.v:12860.13-12860.31" */
input ic_scr_key_valid_i;
wire ic_scr_key_valid_i;
/* cellift = 32'd1 */
input ic_scr_key_valid_i_t0;
wire ic_scr_key_valid_i_t0;
/* src = "generated/sv2v_out.v:12852.42-12852.55" */
output [7:0] ic_tag_addr_o;
wire [7:0] ic_tag_addr_o;
/* cellift = 32'd1 */
output [7:0] ic_tag_addr_o_t0;
wire [7:0] ic_tag_addr_o_t0;
/* src = "generated/sv2v_out.v:12854.57-12854.71" */
input [43:0] ic_tag_rdata_i;
wire [43:0] ic_tag_rdata_i;
/* cellift = 32'd1 */
input [43:0] ic_tag_rdata_i_t0;
wire [43:0] ic_tag_rdata_i_t0;
/* src = "generated/sv2v_out.v:12850.20-12850.32" */
output [1:0] ic_tag_req_o;
wire [1:0] ic_tag_req_o;
/* cellift = 32'd1 */
output [1:0] ic_tag_req_o_t0;
wire [1:0] ic_tag_req_o_t0;
/* src = "generated/sv2v_out.v:12853.33-12853.47" */
output [21:0] ic_tag_wdata_o;
wire [21:0] ic_tag_wdata_o;
/* cellift = 32'd1 */
output [21:0] ic_tag_wdata_o_t0;
wire [21:0] ic_tag_wdata_o_t0;
/* src = "generated/sv2v_out.v:12851.14-12851.28" */
output ic_tag_write_o;
wire ic_tag_write_o;
/* cellift = 32'd1 */
output ic_tag_write_o_t0;
wire ic_tag_write_o_t0;
/* src = "generated/sv2v_out.v:12903.7-12903.20" */
wire icache_enable;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12903.7-12903.20" */
wire icache_enable_t0;
/* src = "generated/sv2v_out.v:12904.7-12904.19" */
wire icache_inval;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12904.7-12904.19" */
wire icache_inval_t0;
/* src = "generated/sv2v_out.v:12975.7-12975.18" */
wire id_in_ready;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12975.7-12975.18" */
wire id_in_ready_t0;
/* src = "generated/sv2v_out.v:12926.7-12926.14" */
wire if_busy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12926.7-12926.14" */
wire if_busy_t0;
/* src = "generated/sv2v_out.v:12891.7-12891.24" */
wire illegal_c_insn_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12891.7-12891.24" */
wire illegal_c_insn_id_t0;
/* src = "generated/sv2v_out.v:12968.7-12968.26" */
wire illegal_csr_insn_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12968.7-12968.26" */
wire illegal_csr_insn_id_t0;
/* src = "generated/sv2v_out.v:13034.7-13034.22" */
/* unused_bits = "0" */
wire illegal_insn_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13034.7-13034.22" */
/* unused_bits = "0" */
wire illegal_insn_id_t0;
/* src = "generated/sv2v_out.v:12895.14-12895.26" */
wire [67:0] imd_val_d_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12895.14-12895.26" */
wire [67:0] imd_val_d_ex_t0;
/* src = "generated/sv2v_out.v:12896.14-12896.26" */
wire [67:0] imd_val_q_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12896.14-12896.26" */
wire [67:0] imd_val_q_ex_t0;
/* src = "generated/sv2v_out.v:12897.13-12897.26" */
wire [1:0] imd_val_we_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12897.13-12897.26" */
wire [1:0] imd_val_we_ex_t0;
/* src = "generated/sv2v_out.v:12829.21-12829.33" */
output [31:0] instr_addr_o;
wire [31:0] instr_addr_o;
/* cellift = 32'd1 */
output [31:0] instr_addr_o_t0;
wire [31:0] instr_addr_o_t0;
/* src = "generated/sv2v_out.v:12888.7-12888.24" */
wire instr_bp_taken_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12888.7-12888.24" */
wire instr_bp_taken_id_t0;
/* src = "generated/sv2v_out.v:13020.7-13020.20" */
/* unused_bits = "0" */
wire instr_done_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13020.7-13020.20" */
/* unused_bits = "0" */
wire instr_done_wb_t0;
/* src = "generated/sv2v_out.v:12831.13-12831.24" */
input instr_err_i;
wire instr_err_i;
/* cellift = 32'd1 */
input instr_err_i_t0;
wire instr_err_i_t0;
/* src = "generated/sv2v_out.v:12981.7-12981.17" */
wire instr_exec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12981.7-12981.17" */
wire instr_exec_t0;
/* src = "generated/sv2v_out.v:12889.7-12889.22" */
wire instr_fetch_err;
/* src = "generated/sv2v_out.v:12890.7-12890.28" */
wire instr_fetch_err_plus2;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12890.7-12890.28" */
wire instr_fetch_err_plus2_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12889.7-12889.22" */
wire instr_fetch_err_t0;
/* src = "generated/sv2v_out.v:12908.7-12908.27" */
wire instr_first_cycle_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12908.7-12908.27" */
wire instr_first_cycle_id_t0;
/* src = "generated/sv2v_out.v:12827.13-12827.24" */
input instr_gnt_i;
wire instr_gnt_i;
/* cellift = 32'd1 */
input instr_gnt_i_t0;
wire instr_gnt_i_t0;
/* src = "generated/sv2v_out.v:13019.7-13019.20" */
/* unused_bits = "0" */
wire instr_id_done;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13019.7-13019.20" */
/* unused_bits = "0" */
wire instr_id_done_t0;
/* src = "generated/sv2v_out.v:12916.7-12916.21" */
wire instr_intg_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12916.7-12916.21" */
wire instr_intg_err_t0;
/* src = "generated/sv2v_out.v:12886.7-12886.29" */
wire instr_is_compressed_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12886.7-12886.29" */
wire instr_is_compressed_id_t0;
/* src = "generated/sv2v_out.v:12882.7-12882.19" */
/* unused_bits = "0" */
wire instr_new_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12882.7-12882.19" */
/* unused_bits = "0" */
wire instr_new_id_t0;
/* src = "generated/sv2v_out.v:12887.7-12887.26" */
wire instr_perf_count_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12887.7-12887.26" */
wire instr_perf_count_id_t0;
/* src = "generated/sv2v_out.v:12884.14-12884.32" */
wire [31:0] instr_rdata_alu_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12884.14-12884.32" */
wire [31:0] instr_rdata_alu_id_t0;
/* src = "generated/sv2v_out.v:12885.14-12885.30" */
wire [15:0] instr_rdata_c_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12885.14-12885.30" */
wire [15:0] instr_rdata_c_id_t0;
/* src = "generated/sv2v_out.v:12830.34-12830.47" */
input [38:0] instr_rdata_i;
wire [38:0] instr_rdata_i;
/* cellift = 32'd1 */
input [38:0] instr_rdata_i_t0;
wire [38:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:12883.14-12883.28" */
wire [31:0] instr_rdata_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12883.14-12883.28" */
wire [31:0] instr_rdata_id_t0;
/* src = "generated/sv2v_out.v:12980.7-12980.22" */
wire instr_req_gated;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12980.7-12980.22" */
wire instr_req_gated_t0;
/* src = "generated/sv2v_out.v:12979.7-12979.20" */
wire instr_req_int;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12979.7-12979.20" */
wire instr_req_int_t0;
/* src = "generated/sv2v_out.v:12826.14-12826.25" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:12828.13-12828.27" */
input instr_rvalid_i;
wire instr_rvalid_i;
/* cellift = 32'd1 */
input instr_rvalid_i_t0;
wire instr_rvalid_i_t0;
/* src = "generated/sv2v_out.v:12983.13-12983.26" */
wire [1:0] instr_type_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12983.13-12983.26" */
wire [1:0] instr_type_wb_t0;
/* src = "generated/sv2v_out.v:12909.7-12909.24" */
wire instr_valid_clear;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12909.7-12909.24" */
wire instr_valid_clear_t0;
/* src = "generated/sv2v_out.v:12881.7-12881.21" */
wire instr_valid_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12881.7-12881.21" */
wire instr_valid_id_t0;
/* src = "generated/sv2v_out.v:12864.13-12864.27" */
input irq_external_i;
wire irq_external_i;
/* cellift = 32'd1 */
input irq_external_i_t0;
wire irq_external_i_t0;
/* src = "generated/sv2v_out.v:12865.20-12865.30" */
input [14:0] irq_fast_i;
wire [14:0] irq_fast_i;
/* cellift = 32'd1 */
input [14:0] irq_fast_i_t0;
wire [14:0] irq_fast_i_t0;
/* src = "generated/sv2v_out.v:12866.13-12866.21" */
input irq_nm_i;
wire irq_nm_i;
/* cellift = 32'd1 */
input irq_nm_i_t0;
wire irq_nm_i_t0;
/* src = "generated/sv2v_out.v:12867.14-12867.27" */
output irq_pending_o;
wire irq_pending_o;
/* cellift = 32'd1 */
output irq_pending_o_t0;
wire irq_pending_o_t0;
/* src = "generated/sv2v_out.v:12862.13-12862.27" */
input irq_software_i;
wire irq_software_i;
/* cellift = 32'd1 */
input irq_software_i_t0;
wire irq_software_i_t0;
/* src = "generated/sv2v_out.v:12863.13-12863.24" */
input irq_timer_i;
wire irq_timer_i;
/* cellift = 32'd1 */
input irq_timer_i_t0;
wire irq_timer_i_t0;
/* src = "generated/sv2v_out.v:12990.14-12990.18" */
wire [17:0] irqs;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12990.14-12990.18" */
wire [17:0] irqs_t0;
/* src = "generated/sv2v_out.v:12921.7-12921.24" */
wire lsu_addr_incr_req;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12921.7-12921.24" */
wire lsu_addr_incr_req_t0;
/* src = "generated/sv2v_out.v:12922.14-12922.27" */
wire [31:0] lsu_addr_last;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12922.14-12922.27" */
wire [31:0] lsu_addr_last_t0;
/* src = "generated/sv2v_out.v:12927.7-12927.15" */
wire lsu_busy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12927.7-12927.15" */
wire lsu_busy_t0;
/* src = "generated/sv2v_out.v:12917.7-12917.19" */
wire lsu_load_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12917.7-12917.19" */
wire lsu_load_err_t0;
/* src = "generated/sv2v_out.v:12919.7-12919.29" */
wire lsu_load_resp_intg_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12919.7-12919.29" */
wire lsu_load_resp_intg_err_t0;
/* src = "generated/sv2v_out.v:12972.7-12972.14" */
wire lsu_req;
/* src = "generated/sv2v_out.v:12974.7-12974.19" */
wire lsu_req_done;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12974.7-12974.19" */
wire lsu_req_done_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12972.7-12972.14" */
wire lsu_req_t0;
/* src = "generated/sv2v_out.v:12978.7-12978.19" */
wire lsu_resp_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12978.7-12978.19" */
wire lsu_resp_err_t0;
/* src = "generated/sv2v_out.v:12977.7-12977.21" */
wire lsu_resp_valid;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12977.7-12977.21" */
wire lsu_resp_valid_t0;
/* src = "generated/sv2v_out.v:12971.7-12971.19" */
wire lsu_sign_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12971.7-12971.19" */
wire lsu_sign_ext_t0;
/* src = "generated/sv2v_out.v:12918.7-12918.20" */
wire lsu_store_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12918.7-12918.20" */
wire lsu_store_err_t0;
/* src = "generated/sv2v_out.v:12920.7-12920.30" */
wire lsu_store_resp_intg_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12920.7-12920.30" */
wire lsu_store_resp_intg_err_t0;
/* src = "generated/sv2v_out.v:12970.13-12970.21" */
wire [1:0] lsu_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12970.13-12970.21" */
wire [1:0] lsu_type_t0;
/* src = "generated/sv2v_out.v:12973.14-12973.23" */
wire [31:0] lsu_wdata;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12973.14-12973.23" */
wire [31:0] lsu_wdata_t0;
/* src = "generated/sv2v_out.v:12969.7-12969.13" */
wire lsu_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12969.7-12969.13" */
wire lsu_we_t0;
/* src = "generated/sv2v_out.v:12953.7-12953.17" */
wire mult_en_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12953.7-12953.17" */
wire mult_en_ex_t0;
/* src = "generated/sv2v_out.v:12955.7-12955.18" */
wire mult_sel_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12955.7-12955.18" */
wire mult_sel_ex_t0;
/* src = "generated/sv2v_out.v:12959.14-12959.34" */
wire [31:0] multdiv_operand_a_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12959.14-12959.34" */
wire [31:0] multdiv_operand_a_ex_t0;
/* src = "generated/sv2v_out.v:12960.14-12960.34" */
wire [31:0] multdiv_operand_b_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12960.14-12960.34" */
wire [31:0] multdiv_operand_b_ex_t0;
/* src = "generated/sv2v_out.v:12957.13-12957.32" */
wire [1:0] multdiv_operator_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12957.13-12957.32" */
wire [1:0] multdiv_operator_ex_t0;
/* src = "generated/sv2v_out.v:12961.7-12961.23" */
wire multdiv_ready_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12961.7-12961.23" */
wire multdiv_ready_id_t0;
/* src = "generated/sv2v_out.v:12958.13-12958.35" */
wire [1:0] multdiv_signed_mode_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12958.13-12958.35" */
wire [1:0] multdiv_signed_mode_ex_t0;
/* src = "generated/sv2v_out.v:12989.7-12989.15" */
wire nmi_mode;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12989.7-12989.15" */
wire nmi_mode_t0;
/* src = "generated/sv2v_out.v:12912.14-12912.28" */
wire [31:0] nt_branch_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12912.14-12912.28" */
wire [31:0] nt_branch_addr_t0;
/* src = "generated/sv2v_out.v:12911.7-12911.27" */
wire nt_branch_mispredict;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12911.7-12911.27" */
wire nt_branch_mispredict_t0;
/* src = "generated/sv2v_out.v:12986.7-12986.26" */
wire outstanding_load_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12986.7-12986.26" */
wire outstanding_load_wb_t0;
/* src = "generated/sv2v_out.v:12987.7-12987.27" */
wire outstanding_store_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12987.7-12987.27" */
wire outstanding_store_wb_t0;
/* src = "generated/sv2v_out.v:12893.14-12893.19" */
wire [31:0] pc_id /* verilator public */;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12893.14-12893.19" */
wire [31:0] pc_id_t0 /* verilator public */;
/* src = "generated/sv2v_out.v:12892.14-12892.19" */
wire [31:0] pc_if;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12892.14-12892.19" */
wire [31:0] pc_if_t0;
/* src = "generated/sv2v_out.v:12906.7-12906.24" */
wire pc_mismatch_alert;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12906.7-12906.24" */
wire pc_mismatch_alert_t0;
/* src = "generated/sv2v_out.v:12913.13-12913.22" */
wire [2:0] pc_mux_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12913.13-12913.22" */
wire [2:0] pc_mux_id_t0;
/* src = "generated/sv2v_out.v:12910.7-12910.13" */
wire pc_set;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12910.7-12910.13" */
wire pc_set_t0;
/* src = "generated/sv2v_out.v:12894.14-12894.19" */
wire [31:0] pc_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12894.14-12894.19" */
wire [31:0] pc_wb_t0;
/* src = "generated/sv2v_out.v:13030.7-13030.18" */
wire perf_branch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13030.7-13030.18" */
wire perf_branch_t0;
/* src = "generated/sv2v_out.v:13028.7-13028.20" */
wire perf_div_wait;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13028.7-13028.20" */
wire perf_div_wait_t0;
/* src = "generated/sv2v_out.v:13026.7-13026.22" */
wire perf_dside_wait;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13026.7-13026.22" */
wire perf_dside_wait_t0;
/* src = "generated/sv2v_out.v:13022.7-13022.35" */
wire perf_instr_ret_compressed_wb;
/* src = "generated/sv2v_out.v:13024.7-13024.40" */
wire perf_instr_ret_compressed_wb_spec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13024.7-13024.40" */
wire perf_instr_ret_compressed_wb_spec_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13022.7-13022.35" */
wire perf_instr_ret_compressed_wb_t0;
/* src = "generated/sv2v_out.v:13021.7-13021.24" */
wire perf_instr_ret_wb;
/* src = "generated/sv2v_out.v:13023.7-13023.29" */
wire perf_instr_ret_wb_spec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13023.7-13023.29" */
wire perf_instr_ret_wb_spec_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13021.7-13021.24" */
wire perf_instr_ret_wb_t0;
/* src = "generated/sv2v_out.v:13025.7-13025.22" */
wire perf_iside_wait;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13025.7-13025.22" */
wire perf_iside_wait_t0;
/* src = "generated/sv2v_out.v:13029.7-13029.16" */
wire perf_jump;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13029.7-13029.16" */
wire perf_jump_t0;
/* src = "generated/sv2v_out.v:13032.7-13032.16" */
wire perf_load;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13032.7-13032.16" */
wire perf_load_t0;
/* src = "generated/sv2v_out.v:13027.7-13027.20" */
wire perf_mul_wait;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13027.7-13027.20" */
wire perf_mul_wait_t0;
/* src = "generated/sv2v_out.v:13033.7-13033.17" */
wire perf_store;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13033.7-13033.17" */
wire perf_store_t0;
/* src = "generated/sv2v_out.v:13031.7-13031.19" */
wire perf_tbranch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13031.7-13031.19" */
wire perf_tbranch_t0;
/* src = "generated/sv2v_out.v:13009.13-13009.25" */
wire [1:0] priv_mode_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13009.13-13009.25" */
wire [1:0] priv_mode_id_t0;
/* src = "generated/sv2v_out.v:12984.7-12984.15" */
wire ready_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12984.7-12984.15" */
wire ready_wb_t0;
/* src = "generated/sv2v_out.v:12952.14-12952.23" */
wire [31:0] result_ex;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12952.14-12952.23" */
wire [31:0] result_ex_t0;
/* src = "generated/sv2v_out.v:12940.7-12940.22" */
wire rf_ecc_err_comb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12940.7-12940.22" */
wire rf_ecc_err_comb_t0;
/* src = "generated/sv2v_out.v:12843.20-12843.32" */
output [4:0] rf_raddr_a_o;
wire [4:0] rf_raddr_a_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_a_o_t0;
wire [4:0] rf_raddr_a_o_t0;
/* src = "generated/sv2v_out.v:12844.20-12844.32" */
output [4:0] rf_raddr_b_o;
wire [4:0] rf_raddr_b_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_b_o_t0;
wire [4:0] rf_raddr_b_o_t0;
/* src = "generated/sv2v_out.v:12944.7-12944.23" */
wire rf_rd_a_wb_match;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12944.7-12944.23" */
wire rf_rd_a_wb_match_t0;
/* src = "generated/sv2v_out.v:12945.7-12945.23" */
wire rf_rd_b_wb_match;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12945.7-12945.23" */
wire rf_rd_b_wb_match_t0;
/* src = "generated/sv2v_out.v:12848.38-12848.54" */
input [38:0] rf_rdata_a_ecc_i;
wire [38:0] rf_rdata_a_ecc_i;
/* cellift = 32'd1 */
input [38:0] rf_rdata_a_ecc_i_t0;
wire [38:0] rf_rdata_a_ecc_i_t0;
/* src = "generated/sv2v_out.v:12849.38-12849.54" */
input [38:0] rf_rdata_b_ecc_i;
wire [38:0] rf_rdata_b_ecc_i;
/* cellift = 32'd1 */
input [38:0] rf_rdata_b_ecc_i_t0;
wire [38:0] rf_rdata_b_ecc_i_t0;
/* src = "generated/sv2v_out.v:12932.7-12932.15" */
wire rf_ren_a;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12932.7-12932.15" */
wire rf_ren_a_t0;
/* src = "generated/sv2v_out.v:12933.7-12933.15" */
wire rf_ren_b;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12933.7-12933.15" */
wire rf_ren_b_t0;
/* src = "generated/sv2v_out.v:12941.13-12941.24" */
wire [4:0] rf_waddr_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12941.13-12941.24" */
wire [4:0] rf_waddr_id_t0;
/* src = "generated/sv2v_out.v:12845.20-12845.33" */
output [4:0] rf_waddr_wb_o;
wire [4:0] rf_waddr_wb_o;
/* cellift = 32'd1 */
output [4:0] rf_waddr_wb_o_t0;
wire [4:0] rf_waddr_wb_o_t0;
/* src = "generated/sv2v_out.v:12936.14-12936.29" */
wire [31:0] rf_wdata_fwd_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12936.14-12936.29" */
wire [31:0] rf_wdata_fwd_wb_t0;
/* src = "generated/sv2v_out.v:12942.14-12942.25" */
wire [31:0] rf_wdata_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12942.14-12942.25" */
wire [31:0] rf_wdata_id_t0;
/* src = "generated/sv2v_out.v:12937.14-12937.26" */
wire [31:0] rf_wdata_lsu;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12937.14-12937.26" */
wire [31:0] rf_wdata_lsu_t0;
/* src = "generated/sv2v_out.v:12935.14-12935.25" */
wire [31:0] rf_wdata_wb;
/* src = "generated/sv2v_out.v:12847.39-12847.56" */
output [38:0] rf_wdata_wb_ecc_o;
wire [38:0] rf_wdata_wb_ecc_o;
/* cellift = 32'd1 */
output [38:0] rf_wdata_wb_ecc_o_t0;
wire [38:0] rf_wdata_wb_ecc_o_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12935.14-12935.25" */
wire [31:0] rf_wdata_wb_t0;
/* src = "generated/sv2v_out.v:12943.7-12943.15" */
wire rf_we_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12943.7-12943.15" */
wire rf_we_id_t0;
/* src = "generated/sv2v_out.v:12939.7-12939.16" */
wire rf_we_lsu;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12939.7-12939.16" */
wire rf_we_lsu_t0;
/* src = "generated/sv2v_out.v:12846.14-12846.24" */
output rf_we_wb_o;
wire rf_we_wb_o;
/* cellift = 32'd1 */
output rf_we_wb_o_t0;
wire rf_we_wb_o_t0;
/* src = "generated/sv2v_out.v:12985.7-12985.18" */
wire rf_write_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12985.7-12985.18" */
wire rf_write_wb_t0;
/* src = "generated/sv2v_out.v:12823.13-12823.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:13018.7-13018.20" */
wire trigger_match;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13018.7-13018.20" */
wire trigger_match_t0;
assign perf_iside_wait = id_in_ready & /* src = "generated/sv2v_out.v:13141.27-13141.56" */ _099_;
assign instr_req_gated = instr_req_int & /* src = "generated/sv2v_out.v:13144.29-13144.84" */ instr_exec;
assign _000_ = _110_ & /* src = "generated/sv2v_out.v:13414.30-13414.54" */ rf_ren_a;
assign \gen_regfile_ecc.rf_ecc_err_a_id  = _000_ & /* src = "generated/sv2v_out.v:13414.29-13414.75" */ _100_;
assign _002_ = _112_ & /* src = "generated/sv2v_out.v:13415.30-13415.54" */ rf_ren_b;
assign \gen_regfile_ecc.rf_ecc_err_b_id  = _002_ & /* src = "generated/sv2v_out.v:13415.29-13415.75" */ _101_;
assign rf_ecc_err_comb = instr_valid_id & /* src = "generated/sv2v_out.v:13416.29-13416.81" */ _102_;
assign _036_ = id_in_ready_t0 & _099_;
assign _039_ = instr_req_int_t0 & instr_exec;
assign _042_ = _111_ & rf_ren_a;
assign _045_ = _001_ & _100_;
assign _048_ = _113_ & rf_ren_b;
assign _051_ = _003_ & _101_;
assign _054_ = instr_valid_id_t0 & _102_;
assign _037_ = instr_valid_id_t0 & id_in_ready;
assign _040_ = instr_exec_t0 & instr_req_int;
assign _043_ = rf_ren_a_t0 & _110_;
assign _046_ = rf_rd_a_wb_match_t0 & _000_;
assign _049_ = rf_ren_b_t0 & _112_;
assign _052_ = rf_rd_b_wb_match_t0 & _002_;
assign _055_ = _103_ & instr_valid_id;
assign _038_ = id_in_ready_t0 & instr_valid_id_t0;
assign _041_ = instr_req_int_t0 & instr_exec_t0;
assign _044_ = _111_ & rf_ren_a_t0;
assign _047_ = _001_ & rf_rd_a_wb_match_t0;
assign _050_ = _113_ & rf_ren_b_t0;
assign _053_ = _003_ & rf_rd_b_wb_match_t0;
assign _056_ = instr_valid_id_t0 & _103_;
assign _084_ = _036_ | _037_;
assign _085_ = _039_ | _040_;
assign _086_ = _042_ | _043_;
assign _087_ = _045_ | _046_;
assign _088_ = _048_ | _049_;
assign _089_ = _051_ | _052_;
assign _090_ = _054_ | _055_;
assign perf_iside_wait_t0 = _084_ | _038_;
assign instr_req_gated_t0 = _085_ | _041_;
assign _001_ = _086_ | _044_;
assign \gen_regfile_ecc.rf_ecc_err_a_id_t0  = _087_ | _047_;
assign _003_ = _088_ | _050_;
assign \gen_regfile_ecc.rf_ecc_err_b_id_t0  = _089_ | _053_;
assign rf_ecc_err_comb_t0 = _090_ | _056_;
assign _004_ = | fetch_enable_i_t0;
assign _005_ = ~ fetch_enable_i_t0;
assign _057_ = fetch_enable_i & _005_;
assign _098_ = _057_ == { 1'h0, _005_[2], 1'h0, _005_[0] };
assign instr_exec_t0 = _098_ & _004_;
assign _006_ = | \g_core_busy_secure.busy_bits_buf_t0 [2:0];
assign _007_ = | \g_core_busy_secure.busy_bits_buf_t0 [8:6];
assign _008_ = | \g_core_busy_secure.busy_bits_buf_t0 [5:3];
assign _009_ = | \g_core_busy_secure.busy_bits_buf_t0 [11:9];
assign _010_ = | \gen_regfile_ecc.rf_ecc_err_a_t0 ;
assign _011_ = | \gen_regfile_ecc.rf_ecc_err_b_t0 ;
assign _012_ = ~ \g_core_busy_secure.busy_bits_buf_t0 [2:0];
assign _013_ = ~ \g_core_busy_secure.busy_bits_buf_t0 [8:6];
assign _014_ = ~ \g_core_busy_secure.busy_bits_buf_t0 [5:3];
assign _015_ = ~ \g_core_busy_secure.busy_bits_buf_t0 [11:9];
assign _016_ = ~ \gen_regfile_ecc.rf_ecc_err_a_t0 ;
assign _017_ = ~ \gen_regfile_ecc.rf_ecc_err_b_t0 ;
assign _076_ = \g_core_busy_secure.busy_bits_buf [2:0] & _012_;
assign _077_ = \g_core_busy_secure.busy_bits_buf [8:6] & _013_;
assign _078_ = \g_core_busy_secure.busy_bits_buf [5:3] & _014_;
assign _079_ = \g_core_busy_secure.busy_bits_buf [11:9] & _015_;
assign _080_ = \gen_regfile_ecc.rf_ecc_err_a  & _016_;
assign _081_ = \gen_regfile_ecc.rf_ecc_err_b  & _017_;
assign _018_ = ! _076_;
assign _019_ = ! _077_;
assign _020_ = ! _078_;
assign _021_ = ! _079_;
assign _022_ = ! _080_;
assign _023_ = ! _081_;
assign core_busy_o_t0[0] = _018_ & _006_;
assign core_busy_o_t0[2] = _019_ & _007_;
assign core_busy_o_t0[1] = _020_ & _008_;
assign core_busy_o_t0[3] = _021_ & _009_;
assign _111_ = _022_ & _010_;
assign _113_ = _023_ & _011_;
assign _097_ = { csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0 } | { csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access, csr_access };
assign _082_ = alu_operand_b_ex_t0[11:0] & _097_;
assign _083_ = { csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0, csr_access_t0 } & alu_operand_b_ex[11:0];
assign csr_addr_t0 = _083_ | _082_;
assign _024_ = ~ lsu_load_err;
assign _025_ = ~ \gen_regfile_ecc.rf_ecc_err_a_id ;
assign _026_ = ~ rf_ecc_err_comb;
assign _027_ = ~ _104_;
assign _028_ = ~ lsu_load_resp_intg_err;
assign _029_ = ~ _106_;
assign _030_ = ~ lsu_store_err;
assign _031_ = ~ \gen_regfile_ecc.rf_ecc_err_b_id ;
assign _032_ = ~ pc_mismatch_alert;
assign _033_ = ~ csr_shadow_err;
assign _034_ = ~ lsu_store_resp_intg_err;
assign _035_ = ~ instr_intg_err;
assign _058_ = lsu_load_err_t0 & _030_;
assign _061_ = \gen_regfile_ecc.rf_ecc_err_a_id_t0  & _031_;
assign _064_ = rf_ecc_err_comb_t0 & _032_;
assign _067_ = _105_ & _033_;
assign _070_ = lsu_load_resp_intg_err_t0 & _034_;
assign _073_ = _107_ & _035_;
assign _059_ = lsu_store_err_t0 & _024_;
assign _062_ = \gen_regfile_ecc.rf_ecc_err_b_id_t0  & _025_;
assign _065_ = pc_mismatch_alert_t0 & _026_;
assign _068_ = csr_shadow_err_t0 & _027_;
assign _071_ = lsu_store_resp_intg_err_t0 & _028_;
assign _074_ = instr_intg_err_t0 & _029_;
assign _060_ = lsu_load_err_t0 & lsu_store_err_t0;
assign _063_ = \gen_regfile_ecc.rf_ecc_err_a_id_t0  & \gen_regfile_ecc.rf_ecc_err_b_id_t0 ;
assign _066_ = rf_ecc_err_comb_t0 & pc_mismatch_alert_t0;
assign _069_ = _105_ & csr_shadow_err_t0;
assign _072_ = lsu_load_resp_intg_err_t0 & lsu_store_resp_intg_err_t0;
assign _075_ = _107_ & instr_intg_err_t0;
assign _091_ = _058_ | _059_;
assign _092_ = _061_ | _062_;
assign _093_ = _064_ | _065_;
assign _094_ = _067_ | _068_;
assign _095_ = _070_ | _071_;
assign _096_ = _073_ | _074_;
assign lsu_resp_err_t0 = _091_ | _060_;
assign _103_ = _092_ | _063_;
assign _105_ = _093_ | _066_;
assign alert_major_internal_o_t0 = _094_ | _069_;
assign _107_ = _095_ | _072_;
assign alert_major_bus_o_t0 = _096_ | _075_;
assign instr_exec = fetch_enable_i == /* src = "generated/sv2v_out.v:13145.24-13145.61" */ 4'h5;
assign core_busy_o[1] = ! /* src = "generated/sv2v_out.v:13053.30-13053.81" */ _108_;
assign core_busy_o[3] = ! /* src = "generated/sv2v_out.v:13053.30-13053.81" */ _109_;
assign _099_ = ~ /* src = "generated/sv2v_out.v:13141.41-13141.56" */ instr_valid_id;
assign _100_ = ~ /* src = "generated/sv2v_out.v:13414.58-13414.75" */ rf_rd_a_wb_match;
assign _101_ = ~ /* src = "generated/sv2v_out.v:13415.58-13415.75" */ rf_rd_b_wb_match;
assign lsu_resp_err = lsu_load_err | /* src = "generated/sv2v_out.v:13315.24-13315.52" */ lsu_store_err;
assign _102_ = \gen_regfile_ecc.rf_ecc_err_a_id  | /* src = "generated/sv2v_out.v:13416.47-13416.80" */ \gen_regfile_ecc.rf_ecc_err_b_id ;
assign _104_ = rf_ecc_err_comb | /* src = "generated/sv2v_out.v:13440.35-13440.70" */ pc_mismatch_alert;
assign alert_major_internal_o = _104_ | /* src = "generated/sv2v_out.v:13440.34-13440.88" */ csr_shadow_err;
assign _106_ = lsu_load_resp_intg_err | /* src = "generated/sv2v_out.v:13441.30-13441.78" */ lsu_store_resp_intg_err;
assign alert_major_bus_o = _106_ | /* src = "generated/sv2v_out.v:13441.29-13441.96" */ instr_intg_err;
assign core_busy_o[0] = | /* src = "generated/sv2v_out.v:13050.30-13050.80" */ \g_core_busy_secure.busy_bits_buf [2:0];
assign core_busy_o[2] = | /* src = "generated/sv2v_out.v:13050.30-13050.80" */ \g_core_busy_secure.busy_bits_buf [8:6];
assign _108_ = | /* src = "generated/sv2v_out.v:13053.30-13053.81" */ \g_core_busy_secure.busy_bits_buf [5:3];
assign _109_ = | /* src = "generated/sv2v_out.v:13053.30-13053.81" */ \g_core_busy_secure.busy_bits_buf [11:9];
assign _110_ = | /* src = "generated/sv2v_out.v:13414.30-13414.43" */ \gen_regfile_ecc.rf_ecc_err_a ;
assign _112_ = | /* src = "generated/sv2v_out.v:13415.30-13415.43" */ \gen_regfile_ecc.rf_ecc_err_b ;
assign csr_addr = csr_access ? /* src = "generated/sv2v_out.v:13447.34-13447.88" */ alu_operand_b_ex[11:0] : 12'h000;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13463.4-13535.3" */
\$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers  cs_registers_i (
.boot_addr_i(boot_addr_i),
.boot_addr_i_t0(boot_addr_i_t0),
.branch_i(perf_branch),
.branch_i_t0(perf_branch_t0),
.branch_taken_i(perf_tbranch),
.branch_taken_i_t0(perf_tbranch_t0),
.clk_i(clk_i),
.csr_access_i(csr_access),
.csr_access_i_t0(csr_access_t0),
.csr_addr_i(csr_addr),
.csr_addr_i_t0(csr_addr_t0),
.csr_depc_o(csr_depc),
.csr_depc_o_t0(csr_depc_t0),
.csr_mcause_i(exc_cause),
.csr_mcause_i_t0(exc_cause_t0),
.csr_mepc_o(csr_mepc),
.csr_mepc_o_t0(csr_mepc_t0),
.csr_mstatus_mie_o(csr_mstatus_mie),
.csr_mstatus_mie_o_t0(csr_mstatus_mie_t0),
.csr_mstatus_tw_o(csr_mstatus_tw),
.csr_mstatus_tw_o_t0(csr_mstatus_tw_t0),
.csr_mtval_i(csr_mtval),
.csr_mtval_i_t0(csr_mtval_t0),
.csr_mtval_o(crash_dump_mtval),
.csr_mtval_o_t0(crash_dump_mtval_t0),
.csr_mtvec_init_i(csr_mtvec_init),
.csr_mtvec_init_i_t0(csr_mtvec_init_t0),
.csr_mtvec_o(csr_mtvec),
.csr_mtvec_o_t0(csr_mtvec_t0),
.csr_op_en_i(csr_op_en),
.csr_op_en_i_t0(csr_op_en_t0),
.csr_op_i(csr_op),
.csr_op_i_t0(csr_op_t0),
.csr_pmp_addr_o(csr_pmp_addr),
.csr_pmp_addr_o_t0(csr_pmp_addr_t0),
.csr_pmp_cfg_o(csr_pmp_cfg),
.csr_pmp_cfg_o_t0(csr_pmp_cfg_t0),
.csr_pmp_mseccfg_o(csr_pmp_mseccfg),
.csr_pmp_mseccfg_o_t0(csr_pmp_mseccfg_t0),
.csr_rdata_o(csr_rdata),
.csr_rdata_o_t0(csr_rdata_t0),
.csr_restore_dret_i(csr_restore_dret_id),
.csr_restore_dret_i_t0(csr_restore_dret_id_t0),
.csr_restore_mret_i(csr_restore_mret_id),
.csr_restore_mret_i_t0(csr_restore_mret_id_t0),
.csr_save_cause_i(csr_save_cause),
.csr_save_cause_i_t0(csr_save_cause_t0),
.csr_save_id_i(csr_save_id),
.csr_save_id_i_t0(csr_save_id_t0),
.csr_save_if_i(csr_save_if),
.csr_save_if_i_t0(csr_save_if_t0),
.csr_save_wb_i(csr_save_wb),
.csr_save_wb_i_t0(csr_save_wb_t0),
.csr_shadow_err_o(csr_shadow_err),
.csr_shadow_err_o_t0(csr_shadow_err_t0),
.csr_wdata_i(alu_operand_a_ex),
.csr_wdata_i_t0(alu_operand_a_ex_t0),
.data_ind_timing_o(data_ind_timing),
.data_ind_timing_o_t0(data_ind_timing_t0),
.debug_cause_i(debug_cause),
.debug_cause_i_t0(debug_cause_t0),
.debug_csr_save_i(debug_csr_save),
.debug_csr_save_i_t0(debug_csr_save_t0),
.debug_ebreakm_o(debug_ebreakm),
.debug_ebreakm_o_t0(debug_ebreakm_t0),
.debug_ebreaku_o(debug_ebreaku),
.debug_ebreaku_o_t0(debug_ebreaku_t0),
.debug_mode_entering_i(debug_mode_entering),
.debug_mode_entering_i_t0(debug_mode_entering_t0),
.debug_mode_i(debug_mode),
.debug_mode_i_t0(debug_mode_t0),
.debug_single_step_o(debug_single_step),
.debug_single_step_o_t0(debug_single_step_t0),
.div_wait_i(perf_div_wait),
.div_wait_i_t0(perf_div_wait_t0),
.double_fault_seen_o(double_fault_seen_o),
.double_fault_seen_o_t0(double_fault_seen_o_t0),
.dside_wait_i(perf_dside_wait),
.dside_wait_i_t0(perf_dside_wait_t0),
.dummy_instr_en_o(dummy_instr_en),
.dummy_instr_en_o_t0(dummy_instr_en_t0),
.dummy_instr_mask_o(dummy_instr_mask),
.dummy_instr_mask_o_t0(dummy_instr_mask_t0),
.dummy_instr_seed_en_o(dummy_instr_seed_en),
.dummy_instr_seed_en_o_t0(dummy_instr_seed_en_t0),
.dummy_instr_seed_o(dummy_instr_seed),
.dummy_instr_seed_o_t0(dummy_instr_seed_t0),
.hart_id_i(hart_id_i),
.hart_id_i_t0(hart_id_i_t0),
.ic_scr_key_valid_i(ic_scr_key_valid_i),
.ic_scr_key_valid_i_t0(ic_scr_key_valid_i_t0),
.icache_enable_o(icache_enable),
.icache_enable_o_t0(icache_enable_t0),
.illegal_csr_insn_o(illegal_csr_insn_id),
.illegal_csr_insn_o_t0(illegal_csr_insn_id_t0),
.instr_ret_compressed_i(perf_instr_ret_compressed_wb),
.instr_ret_compressed_i_t0(perf_instr_ret_compressed_wb_t0),
.instr_ret_compressed_spec_i(perf_instr_ret_compressed_wb_spec),
.instr_ret_compressed_spec_i_t0(perf_instr_ret_compressed_wb_spec_t0),
.instr_ret_i(perf_instr_ret_wb),
.instr_ret_i_t0(perf_instr_ret_wb_t0),
.instr_ret_spec_i(perf_instr_ret_wb_spec),
.instr_ret_spec_i_t0(perf_instr_ret_wb_spec_t0),
.irq_external_i(irq_external_i),
.irq_external_i_t0(irq_external_i_t0),
.irq_fast_i(irq_fast_i),
.irq_fast_i_t0(irq_fast_i_t0),
.irq_pending_o(irq_pending_o),
.irq_pending_o_t0(irq_pending_o_t0),
.irq_software_i(irq_software_i),
.irq_software_i_t0(irq_software_i_t0),
.irq_timer_i(irq_timer_i),
.irq_timer_i_t0(irq_timer_i_t0),
.irqs_o(irqs),
.irqs_o_t0(irqs_t0),
.iside_wait_i(perf_iside_wait),
.iside_wait_i_t0(perf_iside_wait_t0),
.jump_i(perf_jump),
.jump_i_t0(perf_jump_t0),
.mem_load_i(perf_load),
.mem_load_i_t0(perf_load_t0),
.mem_store_i(perf_store),
.mem_store_i_t0(perf_store_t0),
.mul_wait_i(perf_mul_wait),
.mul_wait_i_t0(perf_mul_wait_t0),
.nmi_mode_i(nmi_mode),
.nmi_mode_i_t0(nmi_mode_t0),
.pc_id_i(pc_id),
.pc_id_i_t0(pc_id_t0),
.pc_if_i(pc_if),
.pc_if_i_t0(pc_if_t0),
.pc_wb_i(pc_wb),
.pc_wb_i_t0(pc_wb_t0),
.priv_mode_id_o(priv_mode_id),
.priv_mode_id_o_t0(priv_mode_id_t0),
.priv_mode_lsu_o(\g_no_pmp.unused_priv_lvl_ls ),
.priv_mode_lsu_o_t0(\g_no_pmp.unused_priv_lvl_ls_t0 ),
.rst_ni(rst_ni),
.trigger_match_o(trigger_match),
.trigger_match_o_t0(trigger_match_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13285.4-13312.3" */
\$paramod$a308247794889ee6093207090edbf289adef8be1\ibex_ex_block  ex_block_i (
.alu_adder_result_ex_o(alu_adder_result_ex),
.alu_adder_result_ex_o_t0(alu_adder_result_ex_t0),
.alu_instr_first_cycle_i(instr_first_cycle_id),
.alu_instr_first_cycle_i_t0(instr_first_cycle_id_t0),
.alu_operand_a_i(alu_operand_a_ex),
.alu_operand_a_i_t0(alu_operand_a_ex_t0),
.alu_operand_b_i(alu_operand_b_ex),
.alu_operand_b_i_t0(alu_operand_b_ex_t0),
.alu_operator_i(alu_operator_ex),
.alu_operator_i_t0(alu_operator_ex_t0),
.branch_decision_o(branch_decision),
.branch_decision_o_t0(branch_decision_t0),
.branch_target_o(branch_target_ex),
.branch_target_o_t0(branch_target_ex_t0),
.bt_a_operand_i(bt_a_operand),
.bt_a_operand_i_t0(bt_a_operand_t0),
.bt_b_operand_i(bt_b_operand),
.bt_b_operand_i_t0(bt_b_operand_t0),
.clk_i(clk_i),
.data_ind_timing_i(data_ind_timing),
.data_ind_timing_i_t0(data_ind_timing_t0),
.div_en_i(div_en_ex),
.div_en_i_t0(div_en_ex_t0),
.div_sel_i(div_sel_ex),
.div_sel_i_t0(div_sel_ex_t0),
.ex_valid_o(ex_valid),
.ex_valid_o_t0(ex_valid_t0),
.imd_val_d_o(imd_val_d_ex),
.imd_val_d_o_t0(imd_val_d_ex_t0),
.imd_val_q_i(imd_val_q_ex),
.imd_val_q_i_t0(imd_val_q_ex_t0),
.imd_val_we_o(imd_val_we_ex),
.imd_val_we_o_t0(imd_val_we_ex_t0),
.mult_en_i(mult_en_ex),
.mult_en_i_t0(mult_en_ex_t0),
.mult_sel_i(mult_sel_ex),
.mult_sel_i_t0(mult_sel_ex_t0),
.multdiv_operand_a_i(multdiv_operand_a_ex),
.multdiv_operand_a_i_t0(multdiv_operand_a_ex_t0),
.multdiv_operand_b_i(multdiv_operand_b_ex),
.multdiv_operand_b_i_t0(multdiv_operand_b_ex_t0),
.multdiv_operator_i(multdiv_operator_ex),
.multdiv_operator_i_t0(multdiv_operator_ex_t0),
.multdiv_ready_id_i(multdiv_ready_id),
.multdiv_ready_id_i_t0(multdiv_ready_id_t0),
.multdiv_signed_mode_i(multdiv_signed_mode_ex),
.multdiv_signed_mode_i_t0(multdiv_signed_mode_ex_t0),
.result_ex_o(result_ex),
.result_ex_o_t0(result_ex_t0),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13043.36-13046.5" */
\$paramod\prim_buf\Width=32'00000000000000000000000000001100  \g_core_busy_secure.u_fetch_enable_buf  (
.in_i({ ctrl_busy, if_busy, lsu_busy, ctrl_busy, if_busy, lsu_busy, ctrl_busy, if_busy, lsu_busy, ctrl_busy, if_busy, lsu_busy }),
.in_i_t0({ ctrl_busy_t0, if_busy_t0, lsu_busy_t0, ctrl_busy_t0, if_busy_t0, lsu_busy_t0, ctrl_busy_t0, if_busy_t0, lsu_busy_t0, ctrl_busy_t0, if_busy_t0, lsu_busy_t0 }),
.out_o(\g_core_busy_secure.busy_bits_buf ),
.out_o_t0(\g_core_busy_secure.busy_bits_buf_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13404.30-13407.5" */
prim_secded_inv_39_32_dec \gen_regfile_ecc.regfile_ecc_dec_a  (
.data_i(rf_rdata_a_ecc_i),
.data_i_t0(rf_rdata_a_ecc_i_t0),
.err_o(\gen_regfile_ecc.rf_ecc_err_a ),
.err_o_t0(\gen_regfile_ecc.rf_ecc_err_a_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13408.30-13411.5" */
prim_secded_inv_39_32_dec \gen_regfile_ecc.regfile_ecc_dec_b  (
.data_i(rf_rdata_b_ecc_i),
.data_i_t0(rf_rdata_b_ecc_i_t0),
.err_o(\gen_regfile_ecc.rf_ecc_err_b ),
.err_o_t0(\gen_regfile_ecc.rf_ecc_err_b_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13400.30-13403.5" */
prim_secded_inv_39_32_enc \gen_regfile_ecc.regfile_ecc_enc  (
.data_i(rf_wdata_wb),
.data_i_t0(rf_wdata_wb_t0),
.data_o(rf_wdata_wb_ecc_o),
.data_o_t0(rf_wdata_wb_ecc_o_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13163.4-13279.3" */
\$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  id_stage_i (
.alu_operand_a_ex_o(alu_operand_a_ex),
.alu_operand_a_ex_o_t0(alu_operand_a_ex_t0),
.alu_operand_b_ex_o(alu_operand_b_ex),
.alu_operand_b_ex_o_t0(alu_operand_b_ex_t0),
.alu_operator_ex_o(alu_operator_ex),
.alu_operator_ex_o_t0(alu_operator_ex_t0),
.branch_decision_i(branch_decision),
.branch_decision_i_t0(branch_decision_t0),
.bt_a_operand_o(bt_a_operand),
.bt_a_operand_o_t0(bt_a_operand_t0),
.bt_b_operand_o(bt_b_operand),
.bt_b_operand_o_t0(bt_b_operand_t0),
.clk_i(clk_i),
.csr_access_o(csr_access),
.csr_access_o_t0(csr_access_t0),
.csr_mstatus_mie_i(csr_mstatus_mie),
.csr_mstatus_mie_i_t0(csr_mstatus_mie_t0),
.csr_mstatus_tw_i(csr_mstatus_tw),
.csr_mstatus_tw_i_t0(csr_mstatus_tw_t0),
.csr_mtval_o(csr_mtval),
.csr_mtval_o_t0(csr_mtval_t0),
.csr_op_en_o(csr_op_en),
.csr_op_en_o_t0(csr_op_en_t0),
.csr_op_o(csr_op),
.csr_op_o_t0(csr_op_t0),
.csr_rdata_i(csr_rdata),
.csr_rdata_i_t0(csr_rdata_t0),
.csr_restore_dret_id_o(csr_restore_dret_id),
.csr_restore_dret_id_o_t0(csr_restore_dret_id_t0),
.csr_restore_mret_id_o(csr_restore_mret_id),
.csr_restore_mret_id_o_t0(csr_restore_mret_id_t0),
.csr_save_cause_o(csr_save_cause),
.csr_save_cause_o_t0(csr_save_cause_t0),
.csr_save_id_o(csr_save_id),
.csr_save_id_o_t0(csr_save_id_t0),
.csr_save_if_o(csr_save_if),
.csr_save_if_o_t0(csr_save_if_t0),
.csr_save_wb_o(csr_save_wb),
.csr_save_wb_o_t0(csr_save_wb_t0),
.ctrl_busy_o(ctrl_busy),
.ctrl_busy_o_t0(ctrl_busy_t0),
.data_ind_timing_i(data_ind_timing),
.data_ind_timing_i_t0(data_ind_timing_t0),
.debug_cause_o(debug_cause),
.debug_cause_o_t0(debug_cause_t0),
.debug_csr_save_o(debug_csr_save),
.debug_csr_save_o_t0(debug_csr_save_t0),
.debug_ebreakm_i(debug_ebreakm),
.debug_ebreakm_i_t0(debug_ebreakm_t0),
.debug_ebreaku_i(debug_ebreaku),
.debug_ebreaku_i_t0(debug_ebreaku_t0),
.debug_mode_entering_o(debug_mode_entering),
.debug_mode_entering_o_t0(debug_mode_entering_t0),
.debug_mode_o(debug_mode),
.debug_mode_o_t0(debug_mode_t0),
.debug_req_i(debug_req_i),
.debug_req_i_t0(debug_req_i_t0),
.debug_single_step_i(debug_single_step),
.debug_single_step_i_t0(debug_single_step_t0),
.div_en_ex_o(div_en_ex),
.div_en_ex_o_t0(div_en_ex_t0),
.div_sel_ex_o(div_sel_ex),
.div_sel_ex_o_t0(div_sel_ex_t0),
.en_wb_o(en_wb),
.en_wb_o_t0(en_wb_t0),
.ex_valid_i(ex_valid),
.ex_valid_i_t0(ex_valid_t0),
.exc_cause_o(exc_cause),
.exc_cause_o_t0(exc_cause_t0),
.exc_pc_mux_o(exc_pc_mux_id),
.exc_pc_mux_o_t0(exc_pc_mux_id_t0),
.icache_inval_o(icache_inval),
.icache_inval_o_t0(icache_inval_t0),
.id_in_ready_o(id_in_ready),
.id_in_ready_o_t0(id_in_ready_t0),
.illegal_c_insn_i(illegal_c_insn_id),
.illegal_c_insn_i_t0(illegal_c_insn_id_t0),
.illegal_csr_insn_i(illegal_csr_insn_id),
.illegal_csr_insn_i_t0(illegal_csr_insn_id_t0),
.illegal_insn_o(illegal_insn_id),
.illegal_insn_o_t0(illegal_insn_id_t0),
.imd_val_d_ex_i(imd_val_d_ex),
.imd_val_d_ex_i_t0(imd_val_d_ex_t0),
.imd_val_q_ex_o(imd_val_q_ex),
.imd_val_q_ex_o_t0(imd_val_q_ex_t0),
.imd_val_we_ex_i(imd_val_we_ex),
.imd_val_we_ex_i_t0(imd_val_we_ex_t0),
.instr_bp_taken_i(instr_bp_taken_id),
.instr_bp_taken_i_t0(instr_bp_taken_id_t0),
.instr_exec_i(instr_exec),
.instr_exec_i_t0(instr_exec_t0),
.instr_fetch_err_i(instr_fetch_err),
.instr_fetch_err_i_t0(instr_fetch_err_t0),
.instr_fetch_err_plus2_i(instr_fetch_err_plus2),
.instr_fetch_err_plus2_i_t0(instr_fetch_err_plus2_t0),
.instr_first_cycle_id_o(instr_first_cycle_id),
.instr_first_cycle_id_o_t0(instr_first_cycle_id_t0),
.instr_id_done_o(instr_id_done),
.instr_id_done_o_t0(instr_id_done_t0),
.instr_is_compressed_i(instr_is_compressed_id),
.instr_is_compressed_i_t0(instr_is_compressed_id_t0),
.instr_perf_count_id_o(instr_perf_count_id),
.instr_perf_count_id_o_t0(instr_perf_count_id_t0),
.instr_rdata_alu_i(instr_rdata_alu_id),
.instr_rdata_alu_i_t0(instr_rdata_alu_id_t0),
.instr_rdata_c_i(instr_rdata_c_id),
.instr_rdata_c_i_t0(instr_rdata_c_id_t0),
.instr_rdata_i(instr_rdata_id),
.instr_rdata_i_t0(instr_rdata_id_t0),
.instr_req_o(instr_req_int),
.instr_req_o_t0(instr_req_int_t0),
.instr_type_wb_o(instr_type_wb),
.instr_type_wb_o_t0(instr_type_wb_t0),
.instr_valid_clear_o(instr_valid_clear),
.instr_valid_clear_o_t0(instr_valid_clear_t0),
.instr_valid_i(instr_valid_id),
.instr_valid_i_t0(instr_valid_id_t0),
.irq_nm_i(irq_nm_i),
.irq_nm_i_t0(irq_nm_i_t0),
.irq_pending_i(irq_pending_o),
.irq_pending_i_t0(irq_pending_o_t0),
.irqs_i(irqs),
.irqs_i_t0(irqs_t0),
.lsu_addr_incr_req_i(lsu_addr_incr_req),
.lsu_addr_incr_req_i_t0(lsu_addr_incr_req_t0),
.lsu_addr_last_i(lsu_addr_last),
.lsu_addr_last_i_t0(lsu_addr_last_t0),
.lsu_load_err_i(lsu_load_err),
.lsu_load_err_i_t0(lsu_load_err_t0),
.lsu_load_resp_intg_err_i(lsu_load_resp_intg_err),
.lsu_load_resp_intg_err_i_t0(lsu_load_resp_intg_err_t0),
.lsu_req_done_i(lsu_req_done),
.lsu_req_done_i_t0(lsu_req_done_t0),
.lsu_req_o(lsu_req),
.lsu_req_o_t0(lsu_req_t0),
.lsu_resp_valid_i(lsu_resp_valid),
.lsu_resp_valid_i_t0(lsu_resp_valid_t0),
.lsu_sign_ext_o(lsu_sign_ext),
.lsu_sign_ext_o_t0(lsu_sign_ext_t0),
.lsu_store_err_i(lsu_store_err),
.lsu_store_err_i_t0(lsu_store_err_t0),
.lsu_store_resp_intg_err_i(lsu_store_resp_intg_err),
.lsu_store_resp_intg_err_i_t0(lsu_store_resp_intg_err_t0),
.lsu_type_o(lsu_type),
.lsu_type_o_t0(lsu_type_t0),
.lsu_wdata_o(lsu_wdata),
.lsu_wdata_o_t0(lsu_wdata_t0),
.lsu_we_o(lsu_we),
.lsu_we_o_t0(lsu_we_t0),
.mult_en_ex_o(mult_en_ex),
.mult_en_ex_o_t0(mult_en_ex_t0),
.mult_sel_ex_o(mult_sel_ex),
.mult_sel_ex_o_t0(mult_sel_ex_t0),
.multdiv_operand_a_ex_o(multdiv_operand_a_ex),
.multdiv_operand_a_ex_o_t0(multdiv_operand_a_ex_t0),
.multdiv_operand_b_ex_o(multdiv_operand_b_ex),
.multdiv_operand_b_ex_o_t0(multdiv_operand_b_ex_t0),
.multdiv_operator_ex_o(multdiv_operator_ex),
.multdiv_operator_ex_o_t0(multdiv_operator_ex_t0),
.multdiv_ready_id_o(multdiv_ready_id),
.multdiv_ready_id_o_t0(multdiv_ready_id_t0),
.multdiv_signed_mode_ex_o(multdiv_signed_mode_ex),
.multdiv_signed_mode_ex_o_t0(multdiv_signed_mode_ex_t0),
.nmi_mode_o(nmi_mode),
.nmi_mode_o_t0(nmi_mode_t0),
.nt_branch_addr_o(nt_branch_addr),
.nt_branch_addr_o_t0(nt_branch_addr_t0),
.nt_branch_mispredict_o(nt_branch_mispredict),
.nt_branch_mispredict_o_t0(nt_branch_mispredict_t0),
.outstanding_load_wb_i(outstanding_load_wb),
.outstanding_load_wb_i_t0(outstanding_load_wb_t0),
.outstanding_store_wb_i(outstanding_store_wb),
.outstanding_store_wb_i_t0(outstanding_store_wb_t0),
.pc_id_i(pc_id),
.pc_id_i_t0(pc_id_t0),
.pc_mux_o(pc_mux_id),
.pc_mux_o_t0(pc_mux_id_t0),
.pc_set_o(pc_set),
.pc_set_o_t0(pc_set_t0),
.perf_branch_o(perf_branch),
.perf_branch_o_t0(perf_branch_t0),
.perf_div_wait_o(perf_div_wait),
.perf_div_wait_o_t0(perf_div_wait_t0),
.perf_dside_wait_o(perf_dside_wait),
.perf_dside_wait_o_t0(perf_dside_wait_t0),
.perf_jump_o(perf_jump),
.perf_jump_o_t0(perf_jump_t0),
.perf_mul_wait_o(perf_mul_wait),
.perf_mul_wait_o_t0(perf_mul_wait_t0),
.perf_tbranch_o(perf_tbranch),
.perf_tbranch_o_t0(perf_tbranch_t0),
.priv_mode_i(priv_mode_id),
.priv_mode_i_t0(priv_mode_id_t0),
.ready_wb_i(ready_wb),
.ready_wb_i_t0(ready_wb_t0),
.result_ex_i(result_ex),
.result_ex_i_t0(result_ex_t0),
.rf_raddr_a_o(rf_raddr_a_o),
.rf_raddr_a_o_t0(rf_raddr_a_o_t0),
.rf_raddr_b_o(rf_raddr_b_o),
.rf_raddr_b_o_t0(rf_raddr_b_o_t0),
.rf_rd_a_wb_match_o(rf_rd_a_wb_match),
.rf_rd_a_wb_match_o_t0(rf_rd_a_wb_match_t0),
.rf_rd_b_wb_match_o(rf_rd_b_wb_match),
.rf_rd_b_wb_match_o_t0(rf_rd_b_wb_match_t0),
.rf_rdata_a_i(rf_rdata_a_ecc_i[31:0]),
.rf_rdata_a_i_t0(rf_rdata_a_ecc_i_t0[31:0]),
.rf_rdata_b_i(rf_rdata_b_ecc_i[31:0]),
.rf_rdata_b_i_t0(rf_rdata_b_ecc_i_t0[31:0]),
.rf_ren_a_o(rf_ren_a),
.rf_ren_a_o_t0(rf_ren_a_t0),
.rf_ren_b_o(rf_ren_b),
.rf_ren_b_o_t0(rf_ren_b_t0),
.rf_waddr_id_o(rf_waddr_id),
.rf_waddr_id_o_t0(rf_waddr_id_t0),
.rf_waddr_wb_i(rf_waddr_wb_o),
.rf_waddr_wb_i_t0(rf_waddr_wb_o_t0),
.rf_wdata_fwd_wb_i(rf_wdata_fwd_wb),
.rf_wdata_fwd_wb_i_t0(rf_wdata_fwd_wb_t0),
.rf_wdata_id_o(rf_wdata_id),
.rf_wdata_id_o_t0(rf_wdata_id_t0),
.rf_we_id_o(rf_we_id),
.rf_we_id_o_t0(rf_we_id_t0),
.rf_write_wb_i(rf_write_wb),
.rf_write_wb_i_t0(rf_write_wb_t0),
.rst_ni(rst_ni),
.trigger_match_i(trigger_match),
.trigger_match_i_t0(trigger_match_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13079.4-13140.3" */
\$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  if_stage_i (
.boot_addr_i(boot_addr_i),
.boot_addr_i_t0(boot_addr_i_t0),
.branch_target_ex_i(branch_target_ex),
.branch_target_ex_i_t0(branch_target_ex_t0),
.clk_i(clk_i),
.csr_depc_i(csr_depc),
.csr_depc_i_t0(csr_depc_t0),
.csr_mepc_i(csr_mepc),
.csr_mepc_i_t0(csr_mepc_t0),
.csr_mtvec_i(csr_mtvec),
.csr_mtvec_i_t0(csr_mtvec_t0),
.csr_mtvec_init_o(csr_mtvec_init),
.csr_mtvec_init_o_t0(csr_mtvec_init_t0),
.dummy_instr_en_i(dummy_instr_en),
.dummy_instr_en_i_t0(dummy_instr_en_t0),
.dummy_instr_id_o(dummy_instr_id_o),
.dummy_instr_id_o_t0(dummy_instr_id_o_t0),
.dummy_instr_mask_i(dummy_instr_mask),
.dummy_instr_mask_i_t0(dummy_instr_mask_t0),
.dummy_instr_seed_en_i(dummy_instr_seed_en),
.dummy_instr_seed_en_i_t0(dummy_instr_seed_en_t0),
.dummy_instr_seed_i(dummy_instr_seed),
.dummy_instr_seed_i_t0(dummy_instr_seed_t0),
.exc_cause(exc_cause),
.exc_cause_t0(exc_cause_t0),
.exc_pc_mux_i(exc_pc_mux_id),
.exc_pc_mux_i_t0(exc_pc_mux_id_t0),
.ic_data_addr_o(ic_data_addr_o),
.ic_data_addr_o_t0(ic_data_addr_o_t0),
.ic_data_rdata_i(ic_data_rdata_i),
.ic_data_rdata_i_t0(ic_data_rdata_i_t0),
.ic_data_req_o(ic_data_req_o),
.ic_data_req_o_t0(ic_data_req_o_t0),
.ic_data_wdata_o(ic_data_wdata_o),
.ic_data_wdata_o_t0(ic_data_wdata_o_t0),
.ic_data_write_o(ic_data_write_o),
.ic_data_write_o_t0(ic_data_write_o_t0),
.ic_scr_key_req_o(ic_scr_key_req_o),
.ic_scr_key_req_o_t0(ic_scr_key_req_o_t0),
.ic_scr_key_valid_i(ic_scr_key_valid_i),
.ic_scr_key_valid_i_t0(ic_scr_key_valid_i_t0),
.ic_tag_addr_o(ic_tag_addr_o),
.ic_tag_addr_o_t0(ic_tag_addr_o_t0),
.ic_tag_rdata_i(ic_tag_rdata_i),
.ic_tag_rdata_i_t0(ic_tag_rdata_i_t0),
.ic_tag_req_o(ic_tag_req_o),
.ic_tag_req_o_t0(ic_tag_req_o_t0),
.ic_tag_wdata_o(ic_tag_wdata_o),
.ic_tag_wdata_o_t0(ic_tag_wdata_o_t0),
.ic_tag_write_o(ic_tag_write_o),
.ic_tag_write_o_t0(ic_tag_write_o_t0),
.icache_ecc_error_o(alert_minor_o),
.icache_ecc_error_o_t0(alert_minor_o_t0),
.icache_enable_i(icache_enable),
.icache_enable_i_t0(icache_enable_t0),
.icache_inval_i(icache_inval),
.icache_inval_i_t0(icache_inval_t0),
.id_in_ready_i(id_in_ready),
.id_in_ready_i_t0(id_in_ready_t0),
.if_busy_o(if_busy),
.if_busy_o_t0(if_busy_t0),
.illegal_c_insn_id_o(illegal_c_insn_id),
.illegal_c_insn_id_o_t0(illegal_c_insn_id_t0),
.instr_addr_o(instr_addr_o),
.instr_addr_o_t0(instr_addr_o_t0),
.instr_bp_taken_o(instr_bp_taken_id),
.instr_bp_taken_o_t0(instr_bp_taken_id_t0),
.instr_bus_err_i(instr_err_i),
.instr_bus_err_i_t0(instr_err_i_t0),
.instr_fetch_err_o(instr_fetch_err),
.instr_fetch_err_o_t0(instr_fetch_err_t0),
.instr_fetch_err_plus2_o(instr_fetch_err_plus2),
.instr_fetch_err_plus2_o_t0(instr_fetch_err_plus2_t0),
.instr_gnt_i(instr_gnt_i),
.instr_gnt_i_t0(instr_gnt_i_t0),
.instr_intg_err_o(instr_intg_err),
.instr_intg_err_o_t0(instr_intg_err_t0),
.instr_is_compressed_id_o(instr_is_compressed_id),
.instr_is_compressed_id_o_t0(instr_is_compressed_id_t0),
.instr_new_id_o(instr_new_id),
.instr_new_id_o_t0(instr_new_id_t0),
.instr_rdata_alu_id_o(instr_rdata_alu_id),
.instr_rdata_alu_id_o_t0(instr_rdata_alu_id_t0),
.instr_rdata_c_id_o(instr_rdata_c_id),
.instr_rdata_c_id_o_t0(instr_rdata_c_id_t0),
.instr_rdata_i(instr_rdata_i),
.instr_rdata_i_t0(instr_rdata_i_t0),
.instr_rdata_id_o(instr_rdata_id),
.instr_rdata_id_o_t0(instr_rdata_id_t0),
.instr_req_o(instr_req_o),
.instr_req_o_t0(instr_req_o_t0),
.instr_rvalid_i(instr_rvalid_i),
.instr_rvalid_i_t0(instr_rvalid_i_t0),
.instr_valid_clear_i(instr_valid_clear),
.instr_valid_clear_i_t0(instr_valid_clear_t0),
.instr_valid_id_o(instr_valid_id),
.instr_valid_id_o_t0(instr_valid_id_t0),
.nt_branch_addr_i(nt_branch_addr),
.nt_branch_addr_i_t0(nt_branch_addr_t0),
.nt_branch_mispredict_i(nt_branch_mispredict),
.nt_branch_mispredict_i_t0(nt_branch_mispredict_t0),
.pc_id_o(pc_id),
.pc_id_o_t0(pc_id_t0),
.pc_if_o(pc_if),
.pc_if_o_t0(pc_if_t0),
.pc_mismatch_alert_o(pc_mismatch_alert),
.pc_mismatch_alert_o_t0(pc_mismatch_alert_t0),
.pc_mux_i(pc_mux_id),
.pc_mux_i_t0(pc_mux_id_t0),
.pc_set_i(pc_set),
.pc_set_i_t0(pc_set_t0),
.pmp_err_if_i(1'h0),
.pmp_err_if_i_t0(1'h0),
.pmp_err_if_plus2_i(1'h0),
.pmp_err_if_plus2_i_t0(1'h0),
.req_i(instr_req_gated),
.req_i_t0(instr_req_gated_t0),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13319.4-13351.3" */
\$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  load_store_unit_i (
.adder_result_ex_i(alu_adder_result_ex),
.adder_result_ex_i_t0(alu_adder_result_ex_t0),
.addr_incr_req_o(lsu_addr_incr_req),
.addr_incr_req_o_t0(lsu_addr_incr_req_t0),
.addr_last_o(lsu_addr_last),
.addr_last_o_t0(lsu_addr_last_t0),
.busy_o(lsu_busy),
.busy_o_t0(lsu_busy_t0),
.clk_i(clk_i),
.data_addr_o(data_addr_o),
.data_addr_o_t0(data_addr_o_t0),
.data_be_o(data_be_o),
.data_be_o_t0(data_be_o_t0),
.data_bus_err_i(data_err_i),
.data_bus_err_i_t0(data_err_i_t0),
.data_gnt_i(data_gnt_i),
.data_gnt_i_t0(data_gnt_i_t0),
.data_pmp_err_i(1'h0),
.data_pmp_err_i_t0(1'h0),
.data_rdata_i(data_rdata_i),
.data_rdata_i_t0(data_rdata_i_t0),
.data_req_o(data_req_o),
.data_req_o_t0(data_req_o_t0),
.data_rvalid_i(data_rvalid_i),
.data_rvalid_i_t0(data_rvalid_i_t0),
.data_wdata_o(data_wdata_o),
.data_wdata_o_t0(data_wdata_o_t0),
.data_we_o(data_we_o),
.data_we_o_t0(data_we_o_t0),
.load_err_o(lsu_load_err),
.load_err_o_t0(lsu_load_err_t0),
.load_resp_intg_err_o(lsu_load_resp_intg_err),
.load_resp_intg_err_o_t0(lsu_load_resp_intg_err_t0),
.lsu_rdata_o(rf_wdata_lsu),
.lsu_rdata_o_t0(rf_wdata_lsu_t0),
.lsu_rdata_valid_o(rf_we_lsu),
.lsu_rdata_valid_o_t0(rf_we_lsu_t0),
.lsu_req_done_o(lsu_req_done),
.lsu_req_done_o_t0(lsu_req_done_t0),
.lsu_req_i(lsu_req),
.lsu_req_i_t0(lsu_req_t0),
.lsu_resp_valid_o(lsu_resp_valid),
.lsu_resp_valid_o_t0(lsu_resp_valid_t0),
.lsu_sign_ext_i(lsu_sign_ext),
.lsu_sign_ext_i_t0(lsu_sign_ext_t0),
.lsu_type_i(lsu_type),
.lsu_type_i_t0(lsu_type_t0),
.lsu_wdata_i(lsu_wdata),
.lsu_wdata_i_t0(lsu_wdata_t0),
.lsu_we_i(lsu_we),
.lsu_we_i_t0(lsu_we_t0),
.perf_load_o(perf_load),
.perf_load_o_t0(perf_load_t0),
.perf_store_o(perf_store),
.perf_store_o_t0(perf_store_t0),
.rst_ni(rst_ni),
.store_err_o(lsu_store_err),
.store_err_o_t0(lsu_store_err_t0),
.store_resp_intg_err_o(lsu_store_resp_intg_err),
.store_resp_intg_err_o_t0(lsu_store_resp_intg_err_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:13356.4-13387.3" */
\$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'0\DummyInstructions=1'1  wb_stage_i (
.clk_i(clk_i),
.dummy_instr_id_i(dummy_instr_id_o),
.dummy_instr_id_i_t0(dummy_instr_id_o_t0),
.dummy_instr_wb_o(dummy_instr_wb_o),
.dummy_instr_wb_o_t0(dummy_instr_wb_o_t0),
.en_wb_i(en_wb),
.en_wb_i_t0(en_wb_t0),
.instr_done_wb_o(instr_done_wb),
.instr_done_wb_o_t0(instr_done_wb_t0),
.instr_is_compressed_id_i(instr_is_compressed_id),
.instr_is_compressed_id_i_t0(instr_is_compressed_id_t0),
.instr_perf_count_id_i(instr_perf_count_id),
.instr_perf_count_id_i_t0(instr_perf_count_id_t0),
.instr_type_wb_i(instr_type_wb),
.instr_type_wb_i_t0(instr_type_wb_t0),
.lsu_resp_err_i(lsu_resp_err),
.lsu_resp_err_i_t0(lsu_resp_err_t0),
.lsu_resp_valid_i(lsu_resp_valid),
.lsu_resp_valid_i_t0(lsu_resp_valid_t0),
.outstanding_load_wb_o(outstanding_load_wb),
.outstanding_load_wb_o_t0(outstanding_load_wb_t0),
.outstanding_store_wb_o(outstanding_store_wb),
.outstanding_store_wb_o_t0(outstanding_store_wb_t0),
.pc_id_i(pc_id),
.pc_id_i_t0(pc_id_t0),
.pc_wb_o(pc_wb),
.pc_wb_o_t0(pc_wb_t0),
.perf_instr_ret_compressed_wb_o(perf_instr_ret_compressed_wb),
.perf_instr_ret_compressed_wb_o_t0(perf_instr_ret_compressed_wb_t0),
.perf_instr_ret_compressed_wb_spec_o(perf_instr_ret_compressed_wb_spec),
.perf_instr_ret_compressed_wb_spec_o_t0(perf_instr_ret_compressed_wb_spec_t0),
.perf_instr_ret_wb_o(perf_instr_ret_wb),
.perf_instr_ret_wb_o_t0(perf_instr_ret_wb_t0),
.perf_instr_ret_wb_spec_o(perf_instr_ret_wb_spec),
.perf_instr_ret_wb_spec_o_t0(perf_instr_ret_wb_spec_t0),
.ready_wb_o(ready_wb),
.ready_wb_o_t0(ready_wb_t0),
.rf_waddr_id_i(rf_waddr_id),
.rf_waddr_id_i_t0(rf_waddr_id_t0),
.rf_waddr_wb_o(rf_waddr_wb_o),
.rf_waddr_wb_o_t0(rf_waddr_wb_o_t0),
.rf_wdata_fwd_wb_o(rf_wdata_fwd_wb),
.rf_wdata_fwd_wb_o_t0(rf_wdata_fwd_wb_t0),
.rf_wdata_id_i(rf_wdata_id),
.rf_wdata_id_i_t0(rf_wdata_id_t0),
.rf_wdata_lsu_i(rf_wdata_lsu),
.rf_wdata_lsu_i_t0(rf_wdata_lsu_t0),
.rf_wdata_wb_o(rf_wdata_wb),
.rf_wdata_wb_o_t0(rf_wdata_wb_t0),
.rf_we_id_i(rf_we_id),
.rf_we_id_i_t0(rf_we_id_t0),
.rf_we_lsu_i(rf_we_lsu),
.rf_we_lsu_i_t0(rf_we_lsu_t0),
.rf_we_wb_o(rf_we_wb_o),
.rf_we_wb_o_t0(rf_we_wb_o_t0),
.rf_write_wb_o(rf_write_wb),
.rf_write_wb_o_t0(rf_write_wb_t0),
.rst_ni(rst_ni)
);
assign crash_dump_o = { pc_id, pc_if, lsu_addr_last, csr_mepc, crash_dump_mtval };
assign crash_dump_o_t0 = { pc_id_t0, pc_if_t0, lsu_addr_last_t0, csr_mepc_t0, crash_dump_mtval_t0 };
endmodule

module \$paramod$5fd3ce2f8a67228d339c5f62898ff83b3c2a14f0\prim_lfsr (clk_i, rst_ni, seed_en_i, seed_i, lfsr_en_i, entropy_i, state_o, state_o_t0, seed_i_t0, seed_en_i_t0, lfsr_en_i_t0, entropy_i_t0);
wire _000_;
wire _001_;
wire _002_;
wire [2:0] _003_;
wire [31:0] _004_;
wire _005_;
wire _006_;
wire [31:0] _007_;
wire [31:0] _008_;
wire [17:0] _009_;
wire _010_;
/* cellift = 32'd1 */
wire _011_;
wire [31:0] _012_;
wire [31:0] _013_;
wire [31:0] _014_;
wire [2:0] _015_;
wire _016_;
wire _017_;
wire _018_;
wire [31:0] _019_;
wire [31:0] _020_;
wire [31:0] _021_;
wire [31:0] _022_;
wire [31:0] _023_;
wire [31:0] _024_;
wire [31:0] _025_;
wire [31:0] _026_;
wire [31:0] _027_;
wire [31:0] _028_;
wire _029_;
wire [31:0] _030_;
wire [31:0] _031_;
wire [31:0] _032_;
wire [31:0] _033_;
wire [31:0] _034_;
wire [31:0] _035_;
wire [31:0] _036_;
wire [31:0] _037_;
/* src = "generated/sv2v_out.v:25475.41-25475.60" */
wire _038_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25475.41-25475.60" */
wire _039_;
/* src = "generated/sv2v_out.v:25457.22-25457.29" */
wire _040_;
/* src = "generated/sv2v_out.v:25475.83-25475.119" */
wire [31:0] _041_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25475.83-25475.119" */
wire [31:0] _042_;
/* src = "generated/sv2v_out.v:25475.41-25475.120" */
wire [31:0] _043_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25475.41-25475.120" */
wire [31:0] _044_;
/* src = "generated/sv2v_out.v:25456.30-25456.90" */
wire [31:0] _045_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25456.30-25456.90" */
wire [31:0] _046_;
/* src = "generated/sv2v_out.v:25423.8-25423.13" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:25428.26-25428.35" */
input [7:0] entropy_i;
wire [7:0] entropy_i;
/* cellift = 32'd1 */
input [7:0] entropy_i_t0;
wire [7:0] entropy_i_t0;
/* src = "generated/sv2v_out.v:25435.22-25435.28" */
wire [31:0] lfsr_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25435.22-25435.28" */
wire [31:0] lfsr_d_t0;
/* src = "generated/sv2v_out.v:25427.8-25427.17" */
input lfsr_en_i;
wire lfsr_en_i;
/* cellift = 32'd1 */
input lfsr_en_i_t0;
wire lfsr_en_i_t0;
/* src = "generated/sv2v_out.v:25436.21-25436.27" */
reg [31:0] lfsr_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25436.21-25436.27" */
reg [31:0] lfsr_q_t0;
/* src = "generated/sv2v_out.v:25434.7-25434.13" */
wire lockup;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25434.7-25434.13" */
wire lockup_t0;
/* src = "generated/sv2v_out.v:25437.22-25437.37" */
wire [31:0] next_lfsr_state;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:25437.22-25437.37" */
wire [31:0] next_lfsr_state_t0;
/* src = "generated/sv2v_out.v:25424.8-25424.14" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:25425.8-25425.17" */
input seed_en_i;
wire seed_en_i;
/* cellift = 32'd1 */
input seed_en_i_t0;
wire seed_en_i_t0;
/* src = "generated/sv2v_out.v:25426.23-25426.29" */
input [31:0] seed_i;
wire [31:0] seed_i;
/* cellift = 32'd1 */
input [31:0] seed_i_t0;
wire [31:0] seed_i_t0;
/* src = "generated/sv2v_out.v:25429.33-25429.40" */
output [16:0] state_o;
wire [16:0] state_o;
/* cellift = 32'd1 */
output [16:0] state_o_t0;
wire [16:0] state_o_t0;
assign _000_ = ~ _010_;
assign _035_ = lfsr_d ^ lfsr_q;
assign _025_ = lfsr_d_t0 | lfsr_q_t0;
assign _026_ = _035_ | _025_;
assign _012_ = { _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_, _010_ } & lfsr_d_t0;
assign _013_ = { _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_, _000_ } & lfsr_q_t0;
assign _014_ = _026_ & { _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_, _011_ };
assign _027_ = _012_ | _013_;
assign _028_ = _027_ | _014_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$5fd3ce2f8a67228d339c5f62898ff83b3c2a14f0\prim_lfsr  */
/* PC_TAINT_INFO STATE_NAME lfsr_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) lfsr_q_t0 <= 32'd0;
else lfsr_q_t0 <= _028_;
/* src = "generated/sv2v_out.v:25554.2-25559.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$5fd3ce2f8a67228d339c5f62898ff83b3c2a14f0\prim_lfsr  */
/* PC_TAINT_INFO STATE_NAME lfsr_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) lfsr_q <= 32'd2891135988;
else if (_010_) lfsr_q <= lfsr_d;
assign _016_ = lfsr_en_i_t0 & lockup;
assign _017_ = lockup_t0 & lfsr_en_i;
assign _018_ = lfsr_en_i_t0 & lockup_t0;
assign _029_ = _016_ | _017_;
assign _039_ = _029_ | _018_;
assign _001_ = | { lfsr_en_i_t0, seed_en_i_t0, _039_ };
assign _002_ = | lfsr_q_t0;
assign _003_ = ~ { lfsr_en_i_t0, seed_en_i_t0, _039_ };
assign _004_ = ~ lfsr_q_t0;
assign _015_ = { lfsr_en_i, seed_en_i, _038_ } & _003_;
assign _019_ = lfsr_q & _004_;
assign _005_ = ! _015_;
assign _006_ = ! _019_;
assign _011_ = _005_ & _001_;
assign lockup_t0 = _006_ & _002_;
assign _007_ = ~ { _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_, _038_ };
assign _008_ = ~ { seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i };
assign _031_ = { _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_ } | _007_;
assign _032_ = { seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0 } | _008_;
assign _030_ = { lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0, lfsr_en_i_t0 } | { lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i, lfsr_en_i };
assign _033_ = { seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0 } | { seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i, seed_en_i };
assign _020_ = _042_ & _031_;
assign _022_ = _044_ & _032_;
assign _042_ = next_lfsr_state_t0 & _030_;
assign _023_ = seed_i_t0 & _033_;
assign _034_ = _022_ | _023_;
assign _037_ = _043_ ^ seed_i;
assign _021_ = { _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_, _039_ } & { _009_[17], _036_[30], _009_[16], _036_[28], _009_[15:14], _036_[25:23], _009_[13], _036_[21], _009_[12], _036_[19:18], _009_[11:10], _036_[15:14], _009_[9:7], _036_[10], _009_[6:1], _036_[3], _009_[0], _036_[1:0] };
assign _024_ = { seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0, seed_en_i_t0 } & _037_;
assign _044_ = _021_ | _020_;
assign lfsr_d_t0 = _024_ | _034_;
assign _010_ = | { lfsr_en_i, seed_en_i, _038_ };
assign _009_ = ~ { _041_[31], _041_[29], _041_[27:26], _041_[22], _041_[20], _041_[17:16], _041_[13:11], _041_[9:4], _041_[2] };
assign _046_ = { 24'h000000, entropy_i_t0 } | { lfsr_q_t0[0], 24'h000000, lfsr_q_t0[0], 1'h0, lfsr_q_t0[0], 1'h0, lfsr_q_t0[0], lfsr_q_t0[0], lfsr_q_t0[0] };
assign next_lfsr_state_t0 = _046_ | { 1'h0, lfsr_q_t0[31:1] };
assign _038_ = lfsr_en_i && /* src = "generated/sv2v_out.v:25475.41-25475.60" */ lockup;
assign lockup = ~ /* src = "generated/sv2v_out.v:25457.20-25457.30" */ _040_;
assign _040_ = | /* src = "generated/sv2v_out.v:25457.22-25457.29" */ lfsr_q;
assign { _041_[31], _036_[30], _041_[29], _036_[28], _041_[27:26], _036_[25:23], _041_[22], _036_[21], _041_[20], _036_[19:18], _041_[17:16], _036_[15:14], _041_[13:11], _036_[10], _041_[9:4], _036_[3], _041_[2], _036_[1:0] } = lfsr_en_i ? /* src = "generated/sv2v_out.v:25475.83-25475.119" */ next_lfsr_state : 32'hxxxxxxxx;
assign _043_ = _038_ ? /* src = "generated/sv2v_out.v:25475.41-25475.120" */ 32'd2891135988 : { _041_[31], _036_[30], _041_[29], _036_[28], _041_[27:26], _036_[25:23], _041_[22], _036_[21], _041_[20], _036_[19:18], _041_[17:16], _036_[15:14], _041_[13:11], _036_[10], _041_[9:4], _036_[3], _041_[2], _036_[1:0] };
assign lfsr_d = seed_en_i ? /* src = "generated/sv2v_out.v:25475.19-25475.121" */ seed_i : _043_;
assign _045_ = { 24'h000000, entropy_i } ^ /* src = "generated/sv2v_out.v:25456.30-25456.90" */ { lfsr_q[0], 24'h000000, lfsr_q[0], 1'h0, lfsr_q[0], 1'h0, lfsr_q[0], lfsr_q[0], lfsr_q[0] };
assign next_lfsr_state = _045_ ^ /* src = "generated/sv2v_out.v:25456.29-25456.107" */ { 1'h0, lfsr_q[31:1] };
assign { _036_[31], _036_[29], _036_[27:26], _036_[22], _036_[20], _036_[17:16], _036_[13:11], _036_[9:4], _036_[2] } = _009_;
assign { _041_[30], _041_[28], _041_[25:23], _041_[21], _041_[19:18], _041_[15:14], _041_[10], _041_[3], _041_[1:0] } = { _036_[30], _036_[28], _036_[25:23], _036_[21], _036_[19:18], _036_[15:14], _036_[10], _036_[3], _036_[1:0] };
assign state_o = { lfsr_q[21], lfsr_q[16], lfsr_q[5], lfsr_q[9], lfsr_q[12], lfsr_q[0], lfsr_q[19], lfsr_q[29], lfsr_q[4], lfsr_q[7], lfsr_q[1], lfsr_q[28], lfsr_q[10], lfsr_q[17], lfsr_q[22], lfsr_q[23], lfsr_q[13] };
assign state_o_t0 = { lfsr_q_t0[21], lfsr_q_t0[16], lfsr_q_t0[5], lfsr_q_t0[9], lfsr_q_t0[12], lfsr_q_t0[0], lfsr_q_t0[19], lfsr_q_t0[29], lfsr_q_t0[4], lfsr_q_t0[7], lfsr_q_t0[1], lfsr_q_t0[28], lfsr_q_t0[10], lfsr_q_t0[17], lfsr_q_t0[22], lfsr_q_t0[23], lfsr_q_t0[13] };
endmodule

module \$paramod$5ffe4cc9ba21eb548f33468a0c4a93d38de3dae5\ibex_decoder (clk_i, rst_ni, illegal_insn_o, ebrk_insn_o, mret_insn_o, dret_insn_o, ecall_insn_o, wfi_insn_o, jump_set_o, branch_taken_i, icache_inval_o, instr_first_cycle_i, instr_rdata_i, instr_rdata_alu_i, illegal_c_insn_i, imm_a_mux_sel_o, imm_b_mux_sel_o, bt_a_mux_sel_o, bt_b_mux_sel_o, imm_i_type_o, imm_s_type_o
, imm_b_type_o, imm_u_type_o, imm_j_type_o, zimm_rs1_type_o, rf_wdata_sel_o, rf_we_o, rf_raddr_a_o, rf_raddr_b_o, rf_waddr_o, rf_ren_a_o, rf_ren_b_o, alu_operator_o, alu_op_a_mux_sel_o, alu_op_b_mux_sel_o, alu_multicycle_o, mult_en_o, div_en_o, mult_sel_o, div_sel_o, multdiv_operator_o, multdiv_signed_mode_o
, csr_access_o, csr_op_o, data_req_o, data_we_o, data_type_o, data_sign_extension_o, jump_in_dec_o, branch_in_dec_o, zimm_rs1_type_o_t0, wfi_insn_o_t0, rf_we_o_t0, rf_wdata_sel_o_t0, rf_waddr_o_t0, rf_ren_b_o_t0, rf_raddr_b_o_t0, rf_ren_a_o_t0, multdiv_signed_mode_o_t0, rf_raddr_a_o_t0, multdiv_operator_o_t0, mult_sel_o_t0, mult_en_o_t0
, mret_insn_o_t0, div_sel_o_t0, div_en_o_t0, data_we_o_t0, data_type_o_t0, data_sign_extension_o_t0, data_req_o_t0, csr_op_o_t0, csr_access_o_t0, bt_b_mux_sel_o_t0, bt_a_mux_sel_o_t0, branch_taken_i_t0, branch_in_dec_o_t0, alu_operator_o_t0, alu_op_b_mux_sel_o_t0, alu_op_a_mux_sel_o_t0, alu_multicycle_o_t0, jump_set_o_t0, jump_in_dec_o_t0, instr_rdata_alu_i_t0, instr_first_cycle_i_t0
, imm_u_type_o_t0, imm_s_type_o_t0, imm_j_type_o_t0, imm_i_type_o_t0, imm_b_type_o_t0, imm_b_mux_sel_o_t0, imm_a_mux_sel_o_t0, illegal_insn_o_t0, illegal_c_insn_i_t0, icache_inval_o_t0, ecall_insn_o_t0, ebrk_insn_o_t0, dret_insn_o_t0, instr_rdata_i_t0);
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [6:0] _0000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [6:0] _0001_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [6:0] _0002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [6:0] _0003_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [6:0] _0004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [6:0] _0005_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0007_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [6:0] _0008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [6:0] _0009_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0011_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [6:0] _0012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [6:0] _0013_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0015_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0016_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0017_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0018_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0019_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0021_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0022_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0023_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0024_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0025_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0026_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0027_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0028_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0029_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0030_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0031_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0032_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0033_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0034_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0035_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0036_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0037_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0038_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0039_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0040_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0041_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire [1:0] _0042_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire [1:0] _0043_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire [1:0] _0044_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire [1:0] _0045_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire _0046_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire _0047_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0048_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0049_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0050_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0051_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0052_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0053_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0054_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0055_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0056_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire _0057_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire _0058_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [2:0] _0059_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0060_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0061_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0062_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0063_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0064_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire _0065_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire _0066_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire [1:0] _0067_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire [1:0] _0068_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire [1:0] _0069_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire [1:0] _0070_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0071_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0072_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0073_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0074_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0075_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [1:0] _0076_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0077_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0078_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire [1:0] _0079_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire [1:0] _0080_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire _0081_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire _0082_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0083_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0084_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0085_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0086_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0087_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0088_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0089_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0090_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [2:0] _0091_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0092_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0093_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire _0094_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire _0095_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire [1:0] _0096_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire [1:0] _0097_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire [1:0] _0098_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire [1:0] _0099_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0100_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0101_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0102_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [6:0] _0103_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [6:0] _0104_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0105_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [2:0] _0106_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [2:0] _0107_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [6:0] _0108_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [6:0] _0109_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0110_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0111_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [2:0] _0112_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [1:0] _0113_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [1:0] _0114_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire _0115_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0116_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0117_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [2:0] _0118_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [6:0] _0119_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [6:0] _0120_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [2:0] _0121_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [2:0] _0122_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [1:0] _0123_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [1:0] _0124_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0125_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0126_;
/* src = "generated/sv2v_out.v:15319.2-15770.5" */
wire [1:0] _0127_;
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0128_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15067.2-15318.5" */
wire _0129_;
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire _0139_;
wire _0140_;
wire _0141_;
wire [1:0] _0142_;
wire [2:0] _0143_;
wire [4:0] _0144_;
wire [9:0] _0145_;
wire [2:0] _0146_;
wire [6:0] _0147_;
wire [1:0] _0148_;
wire [11:0] _0149_;
wire [9:0] _0150_;
wire [4:0] _0151_;
wire [2:0] _0152_;
wire [6:0] _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire _0186_;
wire _0187_;
wire _0188_;
wire [1:0] _0189_;
wire [1:0] _0190_;
wire [2:0] _0191_;
wire [4:0] _0192_;
wire [3:0] _0193_;
wire [5:0] _0194_;
wire [3:0] _0195_;
wire [3:0] _0196_;
wire [1:0] _0197_;
wire [1:0] _0198_;
wire [2:0] _0199_;
wire [8:0] _0200_;
wire [2:0] _0201_;
wire [1:0] _0202_;
wire [5:0] _0203_;
wire [17:0] _0204_;
wire [1:0] _0205_;
wire [1:0] _0206_;
wire [1:0] _0207_;
wire [1:0] _0208_;
wire [2:0] _0209_;
wire [1:0] _0210_;
wire [2:0] _0211_;
wire [3:0] _0212_;
wire [2:0] _0213_;
wire [2:0] _0214_;
wire [5:0] _0215_;
wire [2:0] _0216_;
wire [3:0] _0217_;
wire [5:0] _0218_;
wire [4:0] _0219_;
wire [4:0] _0220_;
wire [1:0] _0221_;
wire [1:0] _0222_;
wire [5:0] _0223_;
wire _0224_;
wire _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire _0241_;
wire _0242_;
wire _0243_;
wire _0244_;
wire _0245_;
wire _0246_;
wire _0247_;
wire _0248_;
wire _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire [1:0] _0271_;
wire [1:0] _0272_;
wire [6:0] _0273_;
wire [6:0] _0274_;
wire [6:0] _0275_;
wire [6:0] _0276_;
wire [6:0] _0277_;
wire [6:0] _0278_;
wire [6:0] _0279_;
wire [6:0] _0280_;
wire [6:0] _0281_;
wire [6:0] _0282_;
wire [6:0] _0283_;
wire _0284_;
wire _0285_;
wire _0286_;
wire [1:0] _0287_;
wire [1:0] _0288_;
wire [1:0] _0289_;
wire [6:0] _0290_;
wire [6:0] _0291_;
wire [6:0] _0292_;
wire [6:0] _0293_;
wire [2:0] _0294_;
wire [2:0] _0295_;
wire [2:0] _0296_;
wire [2:0] _0297_;
wire [2:0] _0298_;
wire [1:0] _0299_;
wire [1:0] _0300_;
wire [1:0] _0301_;
wire [1:0] _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire [6:0] _0315_;
wire [6:0] _0316_;
wire [2:0] _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire [1:0] _0323_;
wire _0324_;
wire [1:0] _0325_;
wire _0326_;
wire _0327_;
wire [1:0] _0328_;
wire _0329_;
wire _0330_;
wire _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire _0335_;
wire _0336_;
wire _0337_;
wire [1:0] _0338_;
wire [1:0] _0339_;
wire [1:0] _0340_;
wire [3:0] _0341_;
wire _0342_;
wire [1:0] _0343_;
wire _0344_;
wire [2:0] _0345_;
wire [2:0] _0346_;
wire [1:0] _0347_;
wire [2:0] _0348_;
wire _0349_;
wire [1:0] _0350_;
wire _0351_;
wire _0352_;
wire _0353_;
wire _0354_;
wire _0355_;
wire _0356_;
wire _0357_;
wire _0358_;
wire _0359_;
wire _0360_;
wire _0361_;
wire _0362_;
wire _0363_;
wire _0364_;
wire _0365_;
wire _0366_;
wire _0367_;
/* cellift = 32'd1 */
wire _0368_;
wire _0369_;
/* cellift = 32'd1 */
wire _0370_;
wire _0371_;
/* cellift = 32'd1 */
wire _0372_;
wire _0373_;
/* cellift = 32'd1 */
wire _0374_;
wire _0375_;
/* cellift = 32'd1 */
wire _0376_;
wire _0377_;
/* cellift = 32'd1 */
wire _0378_;
wire _0379_;
/* cellift = 32'd1 */
wire _0380_;
wire _0381_;
/* cellift = 32'd1 */
wire _0382_;
wire _0383_;
/* cellift = 32'd1 */
wire _0384_;
wire _0385_;
wire _0386_;
/* cellift = 32'd1 */
wire _0387_;
wire _0388_;
wire _0389_;
/* cellift = 32'd1 */
wire _0390_;
wire _0391_;
/* cellift = 32'd1 */
wire _0392_;
wire _0393_;
/* cellift = 32'd1 */
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
/* cellift = 32'd1 */
wire _0398_;
wire _0399_;
/* cellift = 32'd1 */
wire _0400_;
wire _0401_;
/* cellift = 32'd1 */
wire _0402_;
wire _0403_;
/* cellift = 32'd1 */
wire _0404_;
wire _0405_;
/* cellift = 32'd1 */
wire _0406_;
wire _0407_;
/* cellift = 32'd1 */
wire _0408_;
wire _0409_;
/* cellift = 32'd1 */
wire _0410_;
wire _0411_;
wire _0412_;
/* cellift = 32'd1 */
wire _0413_;
wire [1:0] _0414_;
wire [1:0] _0415_;
wire [2:0] _0416_;
wire [4:0] _0417_;
wire [3:0] _0418_;
wire [5:0] _0419_;
wire [3:0] _0420_;
wire [3:0] _0421_;
wire [1:0] _0422_;
wire [1:0] _0423_;
wire [2:0] _0424_;
wire [8:0] _0425_;
wire [2:0] _0426_;
wire [1:0] _0427_;
wire [5:0] _0428_;
wire [17:0] _0429_;
wire [1:0] _0430_;
wire [1:0] _0431_;
wire [1:0] _0432_;
wire [1:0] _0433_;
wire [2:0] _0434_;
wire [1:0] _0435_;
wire [2:0] _0436_;
wire _0437_;
wire _0438_;
wire _0439_;
wire _0440_;
wire _0441_;
wire _0442_;
wire _0443_;
wire _0444_;
wire _0445_;
wire _0446_;
wire _0447_;
wire _0448_;
wire _0449_;
wire _0450_;
wire _0451_;
wire _0452_;
wire _0453_;
wire _0454_;
wire _0455_;
wire _0456_;
wire _0457_;
wire _0458_;
wire _0459_;
wire _0460_;
wire _0461_;
wire _0462_;
wire _0463_;
wire _0464_;
wire _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire _0469_;
wire _0470_;
wire _0471_;
wire _0472_;
wire [3:0] _0473_;
wire [2:0] _0474_;
wire [2:0] _0475_;
wire [5:0] _0476_;
wire [2:0] _0477_;
wire [3:0] _0478_;
wire [5:0] _0479_;
wire [1:0] _0480_;
wire [1:0] _0481_;
wire [6:0] _0482_;
wire [6:0] _0483_;
wire [6:0] _0484_;
wire [6:0] _0485_;
wire [6:0] _0486_;
wire [6:0] _0487_;
wire [6:0] _0488_;
wire [6:0] _0489_;
wire [6:0] _0490_;
wire [6:0] _0491_;
wire [6:0] _0492_;
wire [6:0] _0493_;
wire [6:0] _0494_;
wire [6:0] _0495_;
wire [6:0] _0496_;
wire [6:0] _0497_;
wire [6:0] _0498_;
wire [6:0] _0499_;
wire [6:0] _0500_;
wire [6:0] _0501_;
wire [6:0] _0502_;
wire [6:0] _0503_;
wire [6:0] _0504_;
wire [6:0] _0505_;
wire [6:0] _0506_;
wire [6:0] _0507_;
wire [6:0] _0508_;
wire [6:0] _0509_;
wire [6:0] _0510_;
wire [6:0] _0511_;
wire [6:0] _0512_;
wire [6:0] _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0517_;
wire _0518_;
wire _0519_;
wire _0520_;
wire [1:0] _0521_;
wire [1:0] _0522_;
wire [1:0] _0523_;
wire [1:0] _0524_;
wire [1:0] _0525_;
wire [1:0] _0526_;
wire [1:0] _0527_;
wire [1:0] _0528_;
wire [1:0] _0529_;
wire [1:0] _0530_;
wire [1:0] _0531_;
wire [1:0] _0532_;
wire [6:0] _0533_;
wire [6:0] _0534_;
wire [6:0] _0535_;
wire [6:0] _0536_;
wire [6:0] _0537_;
wire [6:0] _0538_;
wire [6:0] _0539_;
wire [6:0] _0540_;
wire [6:0] _0541_;
wire [6:0] _0542_;
wire [6:0] _0543_;
wire [6:0] _0544_;
wire [6:0] _0545_;
wire [2:0] _0546_;
wire [2:0] _0547_;
wire [2:0] _0548_;
wire [2:0] _0549_;
wire [2:0] _0550_;
wire [2:0] _0551_;
wire [2:0] _0552_;
wire [2:0] _0553_;
wire [2:0] _0554_;
wire [2:0] _0555_;
wire [2:0] _0556_;
wire [2:0] _0557_;
wire [2:0] _0558_;
wire [2:0] _0559_;
wire [2:0] _0560_;
wire [2:0] _0561_;
wire [1:0] _0562_;
wire [1:0] _0563_;
wire [1:0] _0564_;
wire [1:0] _0565_;
wire [1:0] _0566_;
wire [1:0] _0567_;
wire [1:0] _0568_;
wire [1:0] _0569_;
wire _0570_;
wire _0571_;
wire _0572_;
wire _0573_;
wire _0574_;
wire [1:0] _0575_;
wire [1:0] _0576_;
wire _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire _0596_;
wire _0597_;
wire _0598_;
wire _0599_;
wire _0600_;
wire _0601_;
wire _0602_;
wire _0603_;
wire _0604_;
wire _0605_;
wire _0606_;
wire _0607_;
wire _0608_;
wire _0609_;
wire _0610_;
wire _0611_;
wire _0612_;
wire _0613_;
wire _0614_;
wire _0615_;
wire _0616_;
wire _0617_;
wire _0618_;
wire _0619_;
wire _0620_;
wire _0621_;
wire [1:0] _0622_;
wire [4:0] _0623_;
wire [2:0] _0624_;
wire [4:0] _0625_;
wire _0626_;
wire _0627_;
wire _0628_;
wire _0629_;
wire _0630_;
wire _0631_;
wire _0632_;
wire _0633_;
wire _0634_;
wire [2:0] _0635_;
wire [4:0] _0636_;
wire [1:0] _0637_;
wire [1:0] _0638_;
wire [9:0] _0639_;
wire _0640_;
wire _0641_;
wire _0642_;
wire _0643_;
wire [6:0] _0644_;
wire [6:0] _0645_;
wire [6:0] _0646_;
wire [6:0] _0647_;
wire [2:0] _0648_;
wire [6:0] _0649_;
wire [6:0] _0650_;
wire [2:0] _0651_;
wire [2:0] _0652_;
wire [6:0] _0653_;
wire _0654_;
wire _0655_;
wire _0656_;
wire _0657_;
wire _0658_;
wire _0659_;
wire _0660_;
wire _0661_;
wire _0662_;
wire _0663_;
wire _0664_;
wire _0665_;
wire _0666_;
wire _0667_;
wire _0668_;
wire _0669_;
wire _0670_;
wire _0671_;
wire _0672_;
wire _0673_;
wire _0674_;
wire _0675_;
wire [1:0] _0676_;
wire _0677_;
wire _0678_;
wire [11:0] _0679_;
wire _0680_;
wire _0681_;
wire _0682_;
wire _0683_;
wire _0684_;
wire _0685_;
wire _0686_;
wire _0687_;
wire _0688_;
wire _0689_;
wire _0690_;
wire _0691_;
wire _0692_;
wire _0693_;
wire _0694_;
wire [1:0] _0695_;
wire [1:0] _0696_;
wire _0697_;
wire _0698_;
wire [9:0] _0699_;
wire _0700_;
wire _0701_;
wire [1:0] _0702_;
wire [1:0] _0703_;
wire [1:0] _0704_;
wire [1:0] _0705_;
wire _0706_;
wire _0707_;
wire [1:0] _0708_;
wire [4:0] _0709_;
wire _0710_;
wire _0711_;
wire [1:0] _0712_;
wire _0713_;
wire _0714_;
wire _0715_;
wire _0716_;
wire [5:0] _0717_;
wire [6:0] _0718_;
wire _0719_;
wire _0720_;
wire [1:0] _0721_;
wire [1:0] _0722_;
wire [1:0] _0723_;
wire [1:0] _0724_;
wire [1:0] _0725_;
wire [1:0] _0726_;
wire _0727_;
wire _0728_;
wire _0729_;
wire _0730_;
wire _0731_;
wire _0732_;
wire _0733_;
wire _0734_;
wire _0735_;
wire _0736_;
wire _0737_;
wire _0738_;
wire [1:0] _0739_;
wire [1:0] _0740_;
wire [1:0] _0741_;
wire [1:0] _0742_;
wire _0743_;
wire _0744_;
wire _0745_;
wire _0746_;
wire _0747_;
wire _0748_;
wire _0749_;
wire _0750_;
wire _0751_;
wire _0752_;
wire _0753_;
wire _0754_;
wire _0755_;
wire _0756_;
wire _0757_;
wire _0758_;
wire [1:0] _0759_;
wire [1:0] _0760_;
wire [6:0] _0761_;
wire [6:0] _0762_;
wire [6:0] _0763_;
wire [6:0] _0764_;
wire [6:0] _0765_;
wire [6:0] _0766_;
wire [6:0] _0767_;
wire [6:0] _0768_;
wire [6:0] _0769_;
wire [6:0] _0770_;
wire [6:0] _0771_;
wire [6:0] _0772_;
wire [6:0] _0773_;
wire [6:0] _0774_;
wire [6:0] _0775_;
wire [6:0] _0776_;
wire [6:0] _0777_;
wire [6:0] _0778_;
wire [6:0] _0779_;
wire [6:0] _0780_;
wire [6:0] _0781_;
wire [6:0] _0782_;
wire [6:0] _0783_;
wire [6:0] _0784_;
wire [6:0] _0785_;
wire [6:0] _0786_;
wire [6:0] _0787_;
wire [6:0] _0788_;
wire _0789_;
wire _0790_;
wire _0791_;
wire _0792_;
wire _0793_;
wire _0794_;
wire [1:0] _0795_;
wire [1:0] _0796_;
wire [1:0] _0797_;
wire [1:0] _0798_;
wire [1:0] _0799_;
wire [1:0] _0800_;
wire [1:0] _0801_;
wire [1:0] _0802_;
wire [1:0] _0803_;
wire [6:0] _0804_;
wire [6:0] _0805_;
wire [6:0] _0806_;
wire [6:0] _0807_;
wire [6:0] _0808_;
wire [6:0] _0809_;
wire [6:0] _0810_;
wire [6:0] _0811_;
wire [6:0] _0812_;
wire [6:0] _0813_;
wire [6:0] _0814_;
wire [2:0] _0815_;
wire [2:0] _0816_;
wire [2:0] _0817_;
wire [2:0] _0818_;
wire [2:0] _0819_;
wire [2:0] _0820_;
wire [2:0] _0821_;
wire [2:0] _0822_;
wire [2:0] _0823_;
wire [2:0] _0824_;
wire [2:0] _0825_;
wire [2:0] _0826_;
wire [2:0] _0827_;
wire [2:0] _0828_;
wire [1:0] _0829_;
wire [1:0] _0830_;
wire [1:0] _0831_;
wire [1:0] _0832_;
wire [1:0] _0833_;
wire [1:0] _0834_;
wire [1:0] _0835_;
wire [1:0] _0836_;
wire _0837_;
wire _0838_;
wire _0839_;
wire _0840_;
wire _0841_;
wire _0842_;
wire _0843_;
wire _0844_;
wire _0845_;
wire _0846_;
wire _0847_;
wire _0848_;
wire _0849_;
wire _0850_;
wire _0851_;
wire _0852_;
wire _0853_;
wire _0854_;
wire _0855_;
wire _0856_;
wire _0857_;
wire _0858_;
wire _0859_;
wire _0860_;
wire _0861_;
wire _0862_;
wire _0863_;
wire _0864_;
wire _0865_;
wire _0866_;
wire _0867_;
wire _0868_;
wire _0869_;
wire _0870_;
wire _0871_;
wire _0872_;
wire _0873_;
wire _0874_;
wire _0875_;
wire _0876_;
wire _0877_;
wire _0878_;
wire _0879_;
wire [6:0] _0880_;
wire [6:0] _0881_;
wire [6:0] _0882_;
wire [2:0] _0883_;
wire _0884_;
wire _0885_;
wire _0886_;
wire _0887_;
wire _0888_;
wire _0889_;
wire _0890_;
wire [1:0] _0891_;
wire _0892_;
wire [1:0] _0893_;
wire _0894_;
wire _0895_;
wire _0896_;
wire _0897_;
wire [1:0] _0898_;
wire [1:0] _0899_;
wire [1:0] _0900_;
wire [1:0] _0901_;
wire _0902_;
/* cellift = 32'd1 */
wire _0903_;
wire _0904_;
/* cellift = 32'd1 */
wire _0905_;
wire _0906_;
/* cellift = 32'd1 */
wire _0907_;
wire _0908_;
/* cellift = 32'd1 */
wire _0909_;
wire _0910_;
/* cellift = 32'd1 */
wire _0911_;
wire _0912_;
/* cellift = 32'd1 */
wire _0913_;
wire _0914_;
/* cellift = 32'd1 */
wire _0915_;
wire _0916_;
/* cellift = 32'd1 */
wire _0917_;
wire _0918_;
/* cellift = 32'd1 */
wire _0919_;
wire _0920_;
/* cellift = 32'd1 */
wire _0921_;
wire _0922_;
/* cellift = 32'd1 */
wire _0923_;
wire _0924_;
/* cellift = 32'd1 */
wire _0925_;
wire [1:0] _0926_;
wire [6:0] _0927_;
wire [6:0] _0928_;
wire [6:0] _0929_;
wire [6:0] _0930_;
wire [6:0] _0931_;
wire [6:0] _0932_;
wire [6:0] _0933_;
wire [6:0] _0934_;
wire [6:0] _0935_;
wire [6:0] _0936_;
wire [6:0] _0937_;
wire _0938_;
wire [1:0] _0939_;
wire [1:0] _0940_;
wire [1:0] _0941_;
wire [6:0] _0942_;
wire [6:0] _0943_;
wire [6:0] _0944_;
wire [6:0] _0945_;
wire [2:0] _0946_;
wire [2:0] _0947_;
wire [2:0] _0948_;
wire [2:0] _0949_;
wire [1:0] _0950_;
wire [1:0] _0951_;
wire _0952_;
wire [1:0] _0953_;
wire _0954_;
wire _0955_;
wire _0956_;
wire _0957_;
wire _0958_;
wire _0959_;
wire _0960_;
wire _0961_;
wire _0962_;
wire _0963_;
wire _0964_;
wire _0965_;
wire _0966_;
wire _0967_;
wire _0968_;
wire _0969_;
wire _0970_;
wire _0971_;
wire _0972_;
wire _0973_;
wire _0974_;
wire _0975_;
wire _0976_;
wire _0977_;
wire _0978_;
wire _0979_;
wire _0980_;
wire _0981_;
wire _0982_;
wire _0983_;
wire _0984_;
wire _0985_;
wire _0986_;
wire _0987_;
wire _0988_;
wire _0989_;
wire _0990_;
wire _0991_;
wire _0992_;
wire _0993_;
wire _0994_;
wire _0995_;
wire _0996_;
wire _0997_;
wire _0998_;
wire _0999_;
wire _1000_;
wire _1001_;
wire _1002_;
wire _1003_;
wire _1004_;
wire _1005_;
wire _1006_;
wire _1007_;
wire _1008_;
wire _1009_;
wire _1010_;
wire _1011_;
wire _1012_;
wire _1013_;
wire _1014_;
wire _1015_;
wire _1016_;
wire _1017_;
wire _1018_;
wire _1019_;
wire _1020_;
wire _1021_;
wire _1022_;
wire _1023_;
wire _1024_;
wire _1025_;
wire _1026_;
wire _1027_;
wire _1028_;
wire _1029_;
wire _1030_;
wire _1031_;
wire _1032_;
wire _1033_;
wire _1034_;
wire _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire [1:0] _1046_;
wire [6:0] _1047_;
wire [6:0] _1048_;
/* cellift = 32'd1 */
wire [6:0] _1049_;
wire [6:0] _1050_;
/* cellift = 32'd1 */
wire [6:0] _1051_;
wire [6:0] _1052_;
/* cellift = 32'd1 */
wire [6:0] _1053_;
wire [6:0] _1054_;
/* cellift = 32'd1 */
wire [6:0] _1055_;
wire [6:0] _1056_;
/* cellift = 32'd1 */
wire [6:0] _1057_;
wire [6:0] _1058_;
/* cellift = 32'd1 */
wire [6:0] _1059_;
wire [6:0] _1060_;
/* cellift = 32'd1 */
wire [6:0] _1061_;
wire [6:0] _1062_;
/* cellift = 32'd1 */
wire [6:0] _1063_;
wire [6:0] _1064_;
/* cellift = 32'd1 */
wire [6:0] _1065_;
wire [6:0] _1066_;
/* cellift = 32'd1 */
wire [6:0] _1067_;
wire [6:0] _1068_;
/* cellift = 32'd1 */
wire [6:0] _1069_;
wire [6:0] _1070_;
/* cellift = 32'd1 */
wire [6:0] _1071_;
wire [6:0] _1072_;
/* cellift = 32'd1 */
wire [6:0] _1073_;
wire [6:0] _1074_;
/* cellift = 32'd1 */
wire [6:0] _1075_;
wire [6:0] _1076_;
/* cellift = 32'd1 */
wire [6:0] _1077_;
wire [6:0] _1078_;
wire [6:0] _1079_;
wire [6:0] _1080_;
/* cellift = 32'd1 */
wire [6:0] _1081_;
wire _1082_;
/* cellift = 32'd1 */
wire _1083_;
wire _1084_;
/* cellift = 32'd1 */
wire _1085_;
wire [1:0] _1086_;
/* cellift = 32'd1 */
wire [1:0] _1087_;
wire [1:0] _1088_;
/* cellift = 32'd1 */
wire [1:0] _1089_;
wire [1:0] _1090_;
/* cellift = 32'd1 */
wire [1:0] _1091_;
wire [1:0] _1092_;
/* cellift = 32'd1 */
wire [1:0] _1093_;
wire [6:0] _1094_;
/* cellift = 32'd1 */
wire [6:0] _1095_;
wire [6:0] _1096_;
/* cellift = 32'd1 */
wire [6:0] _1097_;
/* cellift = 32'd1 */
wire [6:0] _1098_;
wire [6:0] _1099_;
/* cellift = 32'd1 */
wire [6:0] _1100_;
wire [2:0] _1101_;
/* cellift = 32'd1 */
wire [2:0] _1102_;
wire [2:0] _1103_;
/* cellift = 32'd1 */
wire [2:0] _1104_;
wire [2:0] _1105_;
/* cellift = 32'd1 */
wire [2:0] _1106_;
wire [2:0] _1107_;
/* cellift = 32'd1 */
wire [2:0] _1108_;
wire [2:0] _1109_;
/* cellift = 32'd1 */
wire [2:0] _1110_;
wire [1:0] _1111_;
/* cellift = 32'd1 */
wire [1:0] _1112_;
wire [1:0] _1113_;
/* cellift = 32'd1 */
wire [1:0] _1114_;
wire [1:0] _1115_;
/* cellift = 32'd1 */
wire [1:0] _1116_;
wire [1:0] _1117_;
wire [1:0] _1118_;
wire _1119_;
/* cellift = 32'd1 */
wire _1120_;
wire [1:0] _1121_;
/* cellift = 32'd1 */
wire [1:0] _1122_;
wire _1123_;
wire _1124_;
/* cellift = 32'd1 */
wire _1125_;
wire _1126_;
/* cellift = 32'd1 */
wire _1127_;
wire _1128_;
/* cellift = 32'd1 */
wire _1129_;
wire _1130_;
wire _1131_;
/* cellift = 32'd1 */
wire _1132_;
wire _1133_;
/* cellift = 32'd1 */
wire _1134_;
wire _1135_;
/* cellift = 32'd1 */
wire _1136_;
wire _1137_;
/* cellift = 32'd1 */
wire _1138_;
wire _1139_;
/* cellift = 32'd1 */
wire _1140_;
wire _1141_;
/* cellift = 32'd1 */
wire _1142_;
wire _1143_;
/* cellift = 32'd1 */
wire _1144_;
wire _1145_;
/* cellift = 32'd1 */
wire _1146_;
wire _1147_;
/* src = "generated/sv2v_out.v:15064.9-15064.23" */
wire _1148_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15064.9-15064.23" */
wire _1149_;
/* src = "generated/sv2v_out.v:15064.29-15064.43" */
wire _1150_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15064.29-15064.43" */
wire _1151_;
/* src = "generated/sv2v_out.v:15064.50-15064.74" */
wire _1152_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15064.50-15064.74" */
wire _1153_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15162.34-15162.55" */
wire _1154_;
/* src = "generated/sv2v_out.v:15214.9-15214.44" */
wire _1155_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15214.9-15214.44" */
wire _1156_;
/* src = "generated/sv2v_out.v:15524.16-15524.44" */
wire _1157_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15524.16-15524.44" */
wire _1158_;
/* src = "generated/sv2v_out.v:15526.16-15526.44" */
wire _1159_;
/* src = "generated/sv2v_out.v:15754.9-15754.35" */
wire _1160_;
/* src = "generated/sv2v_out.v:15064.7-15064.75" */
wire _1161_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15064.7-15064.75" */
wire _1162_;
/* src = "generated/sv2v_out.v:15064.8-15064.44" */
wire _1163_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15064.8-15064.44" */
wire _1164_;
/* src = "generated/sv2v_out.v:15288.10-15288.59" */
wire _1165_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15288.10-15288.59" */
wire _1166_;
/* src = "generated/sv2v_out.v:15110.9-15110.31" */
wire _1167_;
/* src = "generated/sv2v_out.v:15288.11-15288.32" */
wire _1168_;
/* src = "generated/sv2v_out.v:15288.38-15288.58" */
wire _1169_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15288.38-15288.58" */
wire _1170_;
wire _1171_;
/* cellift = 32'd1 */
wire _1172_;
wire _1173_;
wire _1174_;
/* cellift = 32'd1 */
wire _1175_;
wire _1176_;
/* cellift = 32'd1 */
wire _1177_;
wire _1178_;
/* cellift = 32'd1 */
wire _1179_;
wire _1180_;
/* cellift = 32'd1 */
wire _1181_;
wire _1182_;
/* cellift = 32'd1 */
wire _1183_;
wire _1184_;
/* cellift = 32'd1 */
wire _1185_;
wire _1186_;
/* cellift = 32'd1 */
wire _1187_;
wire _1188_;
/* cellift = 32'd1 */
wire _1189_;
wire _1190_;
/* cellift = 32'd1 */
wire _1191_;
wire _1192_;
/* cellift = 32'd1 */
wire _1193_;
wire _1194_;
/* cellift = 32'd1 */
wire _1195_;
wire _1196_;
wire _1197_;
/* cellift = 32'd1 */
wire _1198_;
wire _1199_;
wire _1200_;
/* cellift = 32'd1 */
wire _1201_;
wire _1202_;
/* cellift = 32'd1 */
wire _1203_;
wire _1204_;
wire _1205_;
/* cellift = 32'd1 */
wire _1206_;
wire _1207_;
/* cellift = 32'd1 */
wire _1208_;
wire _1209_;
/* cellift = 32'd1 */
wire _1210_;
wire _1211_;
/* cellift = 32'd1 */
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire _1216_;
/* cellift = 32'd1 */
wire _1217_;
wire _1218_;
wire _1219_;
/* cellift = 32'd1 */
wire _1220_;
wire _1221_;
/* cellift = 32'd1 */
wire _1222_;
wire _1223_;
/* cellift = 32'd1 */
wire _1224_;
wire _1225_;
/* cellift = 32'd1 */
wire _1226_;
wire _1227_;
/* cellift = 32'd1 */
wire _1228_;
wire _1229_;
/* cellift = 32'd1 */
wire _1230_;
wire _1231_;
/* cellift = 32'd1 */
wire _1232_;
wire _1233_;
wire _1234_;
/* cellift = 32'd1 */
wire _1235_;
wire _1236_;
wire _1237_;
/* cellift = 32'd1 */
wire _1238_;
wire _1239_;
wire _1240_;
wire _1241_;
wire _1242_;
wire _1243_;
wire _1244_;
wire _1245_;
/* cellift = 32'd1 */
wire _1246_;
wire _1247_;
/* cellift = 32'd1 */
wire _1248_;
wire _1249_;
/* cellift = 32'd1 */
wire _1250_;
wire _1251_;
/* cellift = 32'd1 */
wire _1252_;
wire _1253_;
/* cellift = 32'd1 */
wire _1254_;
wire _1255_;
/* cellift = 32'd1 */
wire _1256_;
wire _1257_;
wire _1258_;
/* cellift = 32'd1 */
wire _1259_;
wire _1260_;
/* cellift = 32'd1 */
wire _1261_;
wire [9:0] _1262_;
/* cellift = 32'd1 */
wire [9:0] _1263_;
wire _1264_;
/* cellift = 32'd1 */
wire _1265_;
wire _1266_;
/* cellift = 32'd1 */
wire _1267_;
wire _1268_;
/* cellift = 32'd1 */
wire _1269_;
wire [1:0] _1270_;
/* cellift = 32'd1 */
wire [1:0] _1271_;
wire _1272_;
/* cellift = 32'd1 */
wire _1273_;
/* unused_bits = "1 2" */
wire [5:0] _1274_;
/* cellift = 32'd1 */
/* unused_bits = "1 2" */
wire [5:0] _1275_;
wire _1276_;
/* cellift = 32'd1 */
wire _1277_;
wire _1278_;
wire _1279_;
wire _1280_;
wire _1281_;
wire _1282_;
/* cellift = 32'd1 */
wire _1283_;
wire _1284_;
/* cellift = 32'd1 */
wire _1285_;
wire _1286_;
/* cellift = 32'd1 */
wire _1287_;
wire _1288_;
/* cellift = 32'd1 */
wire _1289_;
/* src = "generated/sv2v_out.v:15162.34-15162.69" */
wire _1290_;
/* src = "generated/sv2v_out.v:14990.13-14990.29" */
output alu_multicycle_o;
wire alu_multicycle_o;
/* cellift = 32'd1 */
output alu_multicycle_o_t0;
wire alu_multicycle_o_t0;
/* src = "generated/sv2v_out.v:14988.19-14988.37" */
output [1:0] alu_op_a_mux_sel_o;
wire [1:0] alu_op_a_mux_sel_o;
/* cellift = 32'd1 */
output [1:0] alu_op_a_mux_sel_o_t0;
wire [1:0] alu_op_a_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:14989.13-14989.31" */
output alu_op_b_mux_sel_o;
wire alu_op_b_mux_sel_o;
/* cellift = 32'd1 */
output alu_op_b_mux_sel_o_t0;
wire alu_op_b_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:14987.19-14987.33" */
output [6:0] alu_operator_o;
wire [6:0] alu_operator_o;
/* cellift = 32'd1 */
output [6:0] alu_operator_o_t0;
wire [6:0] alu_operator_o_t0;
/* src = "generated/sv2v_out.v:15004.13-15004.28" */
output branch_in_dec_o;
wire branch_in_dec_o;
/* cellift = 32'd1 */
output branch_in_dec_o_t0;
wire branch_in_dec_o_t0;
/* src = "generated/sv2v_out.v:14964.13-14964.27" */
input branch_taken_i;
wire branch_taken_i;
/* cellift = 32'd1 */
input branch_taken_i_t0;
wire branch_taken_i_t0;
/* src = "generated/sv2v_out.v:14972.19-14972.33" */
output [1:0] bt_a_mux_sel_o;
wire [1:0] bt_a_mux_sel_o;
/* cellift = 32'd1 */
output [1:0] bt_a_mux_sel_o_t0;
wire [1:0] bt_a_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:14973.19-14973.33" */
output [2:0] bt_b_mux_sel_o;
wire [2:0] bt_b_mux_sel_o;
/* cellift = 32'd1 */
output [2:0] bt_b_mux_sel_o_t0;
wire [2:0] bt_b_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:14955.13-14955.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14997.13-14997.25" */
output csr_access_o;
wire csr_access_o;
/* cellift = 32'd1 */
output csr_access_o_t0;
wire csr_access_o_t0;
/* src = "generated/sv2v_out.v:15018.12-15018.18" */
wire [1:0] csr_op;
/* src = "generated/sv2v_out.v:14998.19-14998.27" */
output [1:0] csr_op_o;
wire [1:0] csr_op_o;
/* cellift = 32'd1 */
output [1:0] csr_op_o_t0;
wire [1:0] csr_op_o_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15018.12-15018.18" */
wire [1:0] csr_op_t0;
/* src = "generated/sv2v_out.v:14999.13-14999.23" */
output data_req_o;
wire data_req_o;
/* cellift = 32'd1 */
output data_req_o_t0;
wire data_req_o_t0;
/* src = "generated/sv2v_out.v:15002.13-15002.34" */
output data_sign_extension_o;
wire data_sign_extension_o;
/* cellift = 32'd1 */
output data_sign_extension_o_t0;
wire data_sign_extension_o_t0;
/* src = "generated/sv2v_out.v:15001.19-15001.30" */
output [1:0] data_type_o;
wire [1:0] data_type_o;
/* cellift = 32'd1 */
output [1:0] data_type_o_t0;
wire [1:0] data_type_o_t0;
/* src = "generated/sv2v_out.v:15000.13-15000.22" */
output data_we_o;
wire data_we_o;
/* cellift = 32'd1 */
output data_we_o_t0;
wire data_we_o_t0;
/* src = "generated/sv2v_out.v:14992.14-14992.22" */
output div_en_o;
wire div_en_o;
/* cellift = 32'd1 */
output div_en_o_t0;
wire div_en_o_t0;
/* src = "generated/sv2v_out.v:14994.13-14994.22" */
output div_sel_o;
wire div_sel_o;
/* cellift = 32'd1 */
output div_sel_o_t0;
wire div_sel_o_t0;
/* src = "generated/sv2v_out.v:14960.13-14960.24" */
output dret_insn_o;
wire dret_insn_o;
/* cellift = 32'd1 */
output dret_insn_o_t0;
wire dret_insn_o_t0;
/* src = "generated/sv2v_out.v:14958.13-14958.24" */
output ebrk_insn_o;
wire ebrk_insn_o;
/* cellift = 32'd1 */
output ebrk_insn_o_t0;
wire ebrk_insn_o_t0;
/* src = "generated/sv2v_out.v:14961.13-14961.25" */
output ecall_insn_o;
wire ecall_insn_o;
/* cellift = 32'd1 */
output ecall_insn_o_t0;
wire ecall_insn_o_t0;
/* src = "generated/sv2v_out.v:14965.13-14965.27" */
output icache_inval_o;
wire icache_inval_o;
/* cellift = 32'd1 */
output icache_inval_o_t0;
wire icache_inval_o_t0;
/* src = "generated/sv2v_out.v:14969.13-14969.29" */
input illegal_c_insn_i;
wire illegal_c_insn_i;
/* cellift = 32'd1 */
input illegal_c_insn_i_t0;
wire illegal_c_insn_i_t0;
/* src = "generated/sv2v_out.v:14957.14-14957.28" */
output illegal_insn_o;
wire illegal_insn_o;
/* cellift = 32'd1 */
output illegal_insn_o_t0;
wire illegal_insn_o_t0;
/* src = "generated/sv2v_out.v:14970.13-14970.28" */
output imm_a_mux_sel_o;
wire imm_a_mux_sel_o;
/* cellift = 32'd1 */
output imm_a_mux_sel_o_t0;
wire imm_a_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:14971.19-14971.34" */
output [2:0] imm_b_mux_sel_o;
wire [2:0] imm_b_mux_sel_o;
/* cellift = 32'd1 */
output [2:0] imm_b_mux_sel_o_t0;
wire [2:0] imm_b_mux_sel_o_t0;
/* src = "generated/sv2v_out.v:14976.21-14976.33" */
output [31:0] imm_b_type_o;
wire [31:0] imm_b_type_o;
/* cellift = 32'd1 */
output [31:0] imm_b_type_o_t0;
wire [31:0] imm_b_type_o_t0;
/* src = "generated/sv2v_out.v:14974.21-14974.33" */
output [31:0] imm_i_type_o;
wire [31:0] imm_i_type_o;
/* cellift = 32'd1 */
output [31:0] imm_i_type_o_t0;
wire [31:0] imm_i_type_o_t0;
/* src = "generated/sv2v_out.v:14978.21-14978.33" */
output [31:0] imm_j_type_o;
wire [31:0] imm_j_type_o;
/* cellift = 32'd1 */
output [31:0] imm_j_type_o_t0;
wire [31:0] imm_j_type_o_t0;
/* src = "generated/sv2v_out.v:14975.21-14975.33" */
output [31:0] imm_s_type_o;
wire [31:0] imm_s_type_o;
/* cellift = 32'd1 */
output [31:0] imm_s_type_o_t0;
wire [31:0] imm_s_type_o_t0;
/* src = "generated/sv2v_out.v:14977.21-14977.33" */
output [31:0] imm_u_type_o;
wire [31:0] imm_u_type_o;
/* cellift = 32'd1 */
output [31:0] imm_u_type_o_t0;
wire [31:0] imm_u_type_o_t0;
/* src = "generated/sv2v_out.v:14966.13-14966.32" */
input instr_first_cycle_i;
wire instr_first_cycle_i;
/* cellift = 32'd1 */
input instr_first_cycle_i_t0;
wire instr_first_cycle_i_t0;
/* src = "generated/sv2v_out.v:14968.20-14968.37" */
input [31:0] instr_rdata_alu_i;
wire [31:0] instr_rdata_alu_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_alu_i_t0;
wire [31:0] instr_rdata_alu_i_t0;
/* src = "generated/sv2v_out.v:14967.20-14967.33" */
input [31:0] instr_rdata_i;
wire [31:0] instr_rdata_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_i_t0;
wire [31:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:15003.13-15003.26" */
output jump_in_dec_o;
wire jump_in_dec_o;
/* cellift = 32'd1 */
output jump_in_dec_o_t0;
wire jump_in_dec_o_t0;
/* src = "generated/sv2v_out.v:14963.13-14963.23" */
output jump_set_o;
wire jump_set_o;
/* cellift = 32'd1 */
output jump_set_o_t0;
wire jump_set_o_t0;
/* src = "generated/sv2v_out.v:14959.13-14959.24" */
output mret_insn_o;
wire mret_insn_o;
/* cellift = 32'd1 */
output mret_insn_o_t0;
wire mret_insn_o_t0;
/* src = "generated/sv2v_out.v:14991.14-14991.23" */
output mult_en_o;
wire mult_en_o;
/* cellift = 32'd1 */
output mult_en_o_t0;
wire mult_en_o_t0;
/* src = "generated/sv2v_out.v:14993.13-14993.23" */
output mult_sel_o;
wire mult_sel_o;
/* cellift = 32'd1 */
output mult_sel_o_t0;
wire mult_sel_o_t0;
/* src = "generated/sv2v_out.v:14995.19-14995.37" */
output [1:0] multdiv_operator_o;
wire [1:0] multdiv_operator_o;
/* cellift = 32'd1 */
output [1:0] multdiv_operator_o_t0;
wire [1:0] multdiv_operator_o_t0;
/* src = "generated/sv2v_out.v:14996.19-14996.40" */
output [1:0] multdiv_signed_mode_o;
wire [1:0] multdiv_signed_mode_o;
/* cellift = 32'd1 */
output [1:0] multdiv_signed_mode_o_t0;
wire [1:0] multdiv_signed_mode_o_t0;
/* src = "generated/sv2v_out.v:14982.20-14982.32" */
output [4:0] rf_raddr_a_o;
wire [4:0] rf_raddr_a_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_a_o_t0;
wire [4:0] rf_raddr_a_o_t0;
/* src = "generated/sv2v_out.v:14983.20-14983.32" */
output [4:0] rf_raddr_b_o;
wire [4:0] rf_raddr_b_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_b_o_t0;
wire [4:0] rf_raddr_b_o_t0;
/* src = "generated/sv2v_out.v:14985.13-14985.23" */
output rf_ren_a_o;
wire rf_ren_a_o;
/* cellift = 32'd1 */
output rf_ren_a_o_t0;
wire rf_ren_a_o_t0;
/* src = "generated/sv2v_out.v:14986.13-14986.23" */
output rf_ren_b_o;
wire rf_ren_b_o;
/* cellift = 32'd1 */
output rf_ren_b_o_t0;
wire rf_ren_b_o_t0;
/* src = "generated/sv2v_out.v:14984.20-14984.30" */
output [4:0] rf_waddr_o;
wire [4:0] rf_waddr_o;
/* cellift = 32'd1 */
output [4:0] rf_waddr_o_t0;
wire [4:0] rf_waddr_o_t0;
/* src = "generated/sv2v_out.v:14980.13-14980.27" */
output rf_wdata_sel_o;
wire rf_wdata_sel_o;
/* cellift = 32'd1 */
output rf_wdata_sel_o_t0;
wire rf_wdata_sel_o_t0;
/* src = "generated/sv2v_out.v:14981.14-14981.21" */
output rf_we_o;
wire rf_we_o;
/* cellift = 32'd1 */
output rf_we_o_t0;
wire rf_we_o_t0;
/* src = "generated/sv2v_out.v:14956.13-14956.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14962.13-14962.23" */
output wfi_insn_o;
wire wfi_insn_o;
/* cellift = 32'd1 */
output wfi_insn_o_t0;
wire wfi_insn_o_t0;
/* src = "generated/sv2v_out.v:14979.21-14979.36" */
output [31:0] zimm_rs1_type_o;
wire [31:0] zimm_rs1_type_o;
/* cellift = 32'd1 */
output [31:0] zimm_rs1_type_o_t0;
wire [31:0] zimm_rs1_type_o_t0;
assign _0130_ = | csr_op_t0;
assign _0131_ = | { instr_rdata_i_t0[26], instr_rdata_i_t0[13:12] };
assign _0133_ = | { instr_rdata_alu_i_t0[31:25], instr_rdata_alu_i_t0[14:12] };
assign _0134_ = | instr_rdata_alu_i_t0[14:12];
assign _0135_ = | instr_rdata_alu_i_t0[6:0];
assign _0136_ = | instr_rdata_i_t0[13:12];
assign _0138_ = | { instr_rdata_i_t0[31:25], instr_rdata_i_t0[14:12] };
assign _0140_ = | instr_rdata_i_t0[14:12];
assign _0141_ = | instr_rdata_i_t0[6:0];
assign _0142_ = ~ csr_op_t0;
assign _0143_ = ~ { instr_rdata_i_t0[26], instr_rdata_i_t0[13:12] };
assign _0144_ = ~ instr_rdata_alu_i_t0[31:27];
assign _0145_ = ~ { instr_rdata_alu_i_t0[31:25], instr_rdata_alu_i_t0[14:12] };
assign _0146_ = ~ instr_rdata_alu_i_t0[14:12];
assign _0147_ = ~ instr_rdata_alu_i_t0[6:0];
assign _0148_ = ~ instr_rdata_i_t0[13:12];
assign _0150_ = ~ { instr_rdata_i_t0[31:25], instr_rdata_i_t0[14:12] };
assign _0151_ = ~ instr_rdata_i_t0[31:27];
assign _0153_ = ~ instr_rdata_i_t0[6:0];
assign _0622_ = csr_op & _0142_;
assign _0624_ = { instr_rdata_i[26], instr_rdata_i[13:12] } & _0143_;
assign _0625_ = instr_rdata_alu_i[31:27] & _0144_;
assign _0639_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } & _0145_;
assign _0648_ = instr_rdata_alu_i[14:12] & _0146_;
assign _0653_ = instr_rdata_alu_i[6:0] & _0147_;
assign _0699_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } & _0150_;
assign _0709_ = instr_rdata_i[31:27] & _0151_;
assign _0635_ = instr_rdata_i[14:12] & _0152_;
assign _0718_ = instr_rdata_i[6:0] & _0153_;
assign _0967_ = _0622_ == { _0142_[1], 1'h0 };
assign _0968_ = _0622_ == _0142_;
assign _0969_ = _0624_ == { _0143_[2], 1'h0, _0143_[0] };
assign _0970_ = _0625_ == { 1'h0, _0144_[3], 3'h0 };
assign _0971_ = _0639_ == { 1'h0, _0145_[8], 5'h00, _0145_[2], 1'h0, _0145_[0] };
assign _0972_ = _0639_ == { 7'h00, _0145_[2], 1'h0, _0145_[0] };
assign _0973_ = _0639_ == { 9'h000, _0145_[0] };
assign _0974_ = _0639_ == { 7'h00, _0145_[2:0] };
assign _0975_ = _0639_ == { 7'h00, _0145_[2:1], 1'h0 };
assign _0976_ = _0639_ == { 7'h00, _0145_[2], 2'h0 };
assign _0977_ = _0639_ == { 8'h00, _0145_[1], 1'h0 };
assign _0978_ = _0639_ == { 1'h0, _0145_[8], 8'h00 };
assign _0979_ = _0639_ == { 6'h00, _0145_[3:0] };
assign _0980_ = _0639_ == { 6'h00, _0145_[3:1], 1'h0 };
assign _0981_ = _0639_ == { 6'h00, _0145_[3:2], 1'h0, _0145_[0] };
assign _0982_ = _0639_ == { 6'h00, _0145_[3:2], 2'h0 };
assign _0983_ = _0639_ == { 6'h00, _0145_[3], 1'h0, _0145_[1:0] };
assign _0984_ = _0639_ == { 6'h00, _0145_[3], 1'h0, _0145_[1], 1'h0 };
assign _0985_ = _0639_ == { 6'h00, _0145_[3], 2'h0, _0145_[0] };
assign _0986_ = _0639_ == { 6'h00, _0145_[3], 3'h0 };
assign _0987_ = _0648_ == { 1'h0, _0146_[1:0] };
assign _0988_ = _0648_ == { 1'h0, _0146_[1], 1'h0 };
assign _0989_ = _0648_ == _0146_;
assign _0990_ = _0648_ == { _0146_[2:1], 1'h0 };
assign _0991_ = _0648_ == { _0146_[2], 1'h0, _0146_[0] };
assign _0992_ = _0648_ == { _0146_[2], 2'h0 };
assign _0993_ = _0648_ == { 2'h0, _0146_[0] };
assign _0994_ = _0653_ == { 2'h0, _0147_[4], 2'h0, _0147_[1:0] };
assign _0995_ = _0653_ == { 5'h00, _0147_[1:0] };
assign _0996_ = _0653_ == { 3'h0, _0147_[3:0] };
assign _0997_ = _0653_ == { 2'h0, _0147_[4], 1'h0, _0147_[2:0] };
assign _0998_ = _0653_ == { 1'h0, _0147_[5:4], 1'h0, _0147_[2:0] };
assign _0999_ = _0653_ == { 1'h0, _0147_[5], 3'h0, _0147_[1:0] };
assign _1000_ = _0653_ == { _0147_[6:5], 3'h0, _0147_[1:0] };
assign _1001_ = _0653_ == { _0147_[6:5], 2'h0, _0147_[2:0] };
assign _1002_ = _0653_ == { _0147_[6:5], 1'h0, _0147_[3:0] };
assign _1003_ = _0653_ == { 1'h0, _0147_[5:4], 2'h0, _0147_[1:0] };
assign _1004_ = _0653_ == { _0147_[6:4], 2'h0, _0147_[1:0] };
assign _1005_ = _0676_ == _0148_;
assign _1006_ = _0679_ == { 3'h0, _0149_[8], 5'h00, _0149_[2], 1'h0, _0149_[0] };
assign _1007_ = _0679_ == { 1'h0, _0149_[10:7], 1'h0, _0149_[5:4], 2'h0, _0149_[1], 1'h0 };
assign _1008_ = _0679_ == { 2'h0, _0149_[9:8], 6'h00, _0149_[1], 1'h0 };
assign _1009_ = _0679_ == { 11'h000, _0149_[0] };
assign _1010_ = _0699_ == { 6'h00, _0150_[3], 3'h0 };
assign _1011_ = _0699_ == { 1'h0, _0150_[8], 8'h00 };
assign _1012_ = _0699_ == { 8'h00, _0150_[1], 1'h0 };
assign _1013_ = _0699_ == { 8'h00, _0150_[1:0] };
assign _1014_ = _0699_ == { 7'h00, _0150_[2], 2'h0 };
assign _1015_ = _0699_ == { 7'h00, _0150_[2:1], 1'h0 };
assign _1016_ = _0699_ == { 7'h00, _0150_[2:0] };
assign _1017_ = _0699_ == { 9'h000, _0150_[0] };
assign _1018_ = _0699_ == { 7'h00, _0150_[2], 1'h0, _0150_[0] };
assign _1019_ = _0699_ == { 1'h0, _0150_[8], 5'h00, _0150_[2], 1'h0, _0150_[0] };
assign _1020_ = _0699_ == { 6'h00, _0150_[3:0] };
assign _1021_ = _0699_ == { 6'h00, _0150_[3:1], 1'h0 };
assign _1022_ = _0699_ == { 6'h00, _0150_[3:2], 1'h0, _0150_[0] };
assign _1023_ = _0699_ == { 6'h00, _0150_[3:2], 2'h0 };
assign _1024_ = _0699_ == { 6'h00, _0150_[3], 1'h0, _0150_[1:0] };
assign _1025_ = _0699_ == { 6'h00, _0150_[3], 1'h0, _0150_[1], 1'h0 };
assign _1026_ = _0699_ == { 6'h00, _0150_[3], 2'h0, _0150_[0] };
assign _1027_ = _0709_ == { 1'h0, _0151_[3], 3'h0 };
assign _1028_ = _0676_ == { _0148_[1], 1'h0 };
assign _1029_ = _0676_ == { 1'h0, _0148_[0] };
assign _1030_ = _0635_ == { 2'h0, _0152_[0] };
assign _1031_ = _0635_ == { _0152_[2], 2'h0 };
assign _1032_ = _0635_ == { _0152_[2], 1'h0, _0152_[0] };
assign _1033_ = _0635_ == { _0152_[2:1], 1'h0 };
assign _1034_ = _0635_ == _0152_;
assign _1035_ = _0718_ == { 2'h0, _0153_[4], 1'h0, _0153_[2:0] };
assign _1036_ = _0718_ == { 1'h0, _0153_[5:4], 1'h0, _0153_[2:0] };
assign _1037_ = _0718_ == { _0153_[6:5], 1'h0, _0153_[3:0] };
assign _1038_ = _0718_ == { 1'h0, _0153_[5:4], 2'h0, _0153_[1:0] };
assign _1039_ = _0718_ == { 2'h0, _0153_[4], 2'h0, _0153_[1:0] };
assign _1040_ = _0718_ == { 5'h00, _0153_[1:0] };
assign _1041_ = _0718_ == { 1'h0, _0153_[5], 3'h0, _0153_[1:0] };
assign _1042_ = _0718_ == { _0153_[6:5], 3'h0, _0153_[1:0] };
assign _1043_ = _0718_ == { _0153_[6:5], 2'h0, _0153_[2:0] };
assign _1044_ = _0718_ == { 3'h0, _0153_[3:0] };
assign _1045_ = _0718_ == { _0153_[6:4], 2'h0, _0153_[1:0] };
assign _1149_ = _0967_ & _0130_;
assign _1151_ = _0968_ & _0130_;
assign _1156_ = _0969_ & _0131_;
assign _0003_[5] = _0970_ & _0132_;
assign _1193_ = _0971_ & _0133_;
assign _1195_ = _0972_ & _0133_;
assign _1049_[3] = _0973_ & _0133_;
assign _1198_ = _0974_ & _0133_;
assign _1055_[0] = _0975_ & _0133_;
assign _1201_ = _0976_ & _0133_;
assign _1203_ = _0977_ & _0133_;
assign _1057_[5] = _0978_ & _0133_;
assign _1177_ = _0979_ & _0133_;
assign _1179_ = _0980_ & _0133_;
assign _1181_ = _0981_ & _0133_;
assign _1183_ = _0982_ & _0133_;
assign _1185_ = _0983_ & _0133_;
assign _1187_ = _0984_ & _0133_;
assign _1189_ = _0985_ & _0133_;
assign _1191_ = _0986_ & _0133_;
assign _1217_ = _0987_ & _0134_;
assign _1071_[5] = _0988_ & _0134_;
assign _1065_[2] = _0989_ & _0134_;
assign _1075_[0] = _0990_ & _0134_;
assign _1210_ = _0991_ & _0134_;
assign _1069_[5] = _0992_ & _0134_;
assign _0122_[2] = _0993_ & _0134_;
assign _1212_ = _0994_ & _0135_;
assign _1230_ = _0995_ & _0135_;
assign _1175_ = _0996_ & _0135_;
assign _1228_ = _0997_ & _0135_;
assign _1232_ = _0998_ & _0135_;
assign _1220_ = _0999_ & _0135_;
assign _1222_ = _1000_ & _0135_;
assign _1224_ = _1001_ & _0135_;
assign _1226_ = _1002_ & _0135_;
assign _1208_ = _1003_ & _0135_;
assign _1172_ = _1004_ & _0135_;
assign _1112_[0] = _1005_ & _0136_;
assign _0102_ = _1006_ & _0137_;
assign _0084_ = _1007_ & _0137_;
assign _0093_ = _1008_ & _0137_;
assign _0086_ = _1009_ & _0137_;
assign _1261_ = _1010_ & _0138_;
assign _1263_[1] = _1011_ & _0138_;
assign _1263_[2] = _1012_ & _0138_;
assign _1263_[3] = _1013_ & _0138_;
assign _1263_[4] = _1014_ & _0138_;
assign _1263_[5] = _1015_ & _0138_;
assign _1263_[6] = _1016_ & _0138_;
assign _1263_[7] = _1017_ & _0138_;
assign _1263_[8] = _1018_ & _0138_;
assign _1263_[9] = _1019_ & _0138_;
assign _1248_ = _1020_ & _0138_;
assign _1250_ = _1021_ & _0138_;
assign _1252_ = _1022_ & _0138_;
assign _1254_ = _1023_ & _0138_;
assign _1256_ = _1024_ & _0138_;
assign _1116_[0] = _1025_ & _0138_;
assign _1259_ = _1026_ & _0138_;
assign _1271_[1] = _1027_ & _0139_;
assign _1235_ = _1028_ & _0136_;
assign _1114_[0] = _1029_ & _0136_;
assign _0061_ = _1030_ & _0140_;
assign _1275_[3] = _1031_ & _0140_;
assign _1267_ = _1032_ & _0140_;
assign _1275_[4] = _1033_ & _0140_;
assign _1275_[5] = _1034_ & _0140_;
assign _1287_ = _1035_ & _0141_;
assign _1289_ = _1036_ & _0141_;
assign _1285_ = _1037_ & _0141_;
assign _1265_ = _1038_ & _0141_;
assign _1269_ = _1039_ & _0141_;
assign _1277_ = _1040_ & _0141_;
assign _0021_ = _1041_ & _0141_;
assign _0017_ = _1042_ & _0141_;
assign _1283_ = _1043_ & _0141_;
assign _1246_ = _1044_ & _0141_;
assign _1238_ = _1045_ & _0141_;
assign _0626_ = _1164_ & _1152_;
assign _0627_ = _1153_ & _1163_;
assign _0628_ = _1164_ & _1153_;
assign _0876_ = _0626_ | _0627_;
assign _1162_ = _0876_ | _0628_;
assign _0154_ = | { _0041_, _0061_ };
assign _0155_ = | { _1226_, _1228_ };
assign _0156_ = | { _0021_, _0017_, _1265_ };
assign _0157_ = | { _0086_, _0093_, _0084_, _0102_, _0088_ };
assign _0158_ = | { _1269_, _1287_, _1289_, _1265_ };
assign _0159_ = | { _0021_, _0017_, _1269_, _1277_, _1283_, _1265_ };
assign _0160_ = | { _1185_, _1187_, _1189_, _1191_ };
assign _0161_ = | { _1177_, _1179_, _1181_, _1183_ };
assign _0162_ = | { _1248_, _1250_ };
assign _0163_ = | { _1252_, _1254_ };
assign _0164_ = | { _1116_[0], _1256_, _1259_ };
assign _0165_ = | { _1185_, _1187_, _1189_, _1191_, _1177_, _1179_, _1181_, _1183_, _1206_ };
assign _0166_ = | { _1250_, _1254_, _1259_ };
assign _0167_ = | { _1232_, _1228_ };
assign _0168_ = | { _1232_, _1220_, _1224_, _1230_, _1226_, _1228_ };
assign _0169_ = | { _1116_[0], _1248_, _1250_, _1252_, _1254_, _1256_, _1259_, _1261_, _1263_ };
assign _0170_ = | { _1224_, _1222_ };
assign _0171_ = | { _1283_, _1285_ };
assign _0172_ = | { _0021_, _1277_ };
assign _0173_ = | { _0122_[2], _0058_ };
assign _0174_ = | { _1114_[0], _1112_[0], _1235_ };
assign _0175_ = | { _1114_[0], _1122_[1] };
assign _0176_ = | { _1114_[0], _1122_[1], _1235_ };
assign _0177_ = | { _0903_, _1195_, _1198_, _1049_[3] };
assign _0178_ = | { _0907_, _1065_[2], _1075_[0] };
assign _0179_ = | { _1210_, _1065_[2], _1075_[0] };
assign _0180_ = | { _1172_, _1212_, _1175_, _1208_, _1220_, _1230_ };
assign _0181_ = | { _1212_, _1175_, _1208_ };
assign _0182_ = | { _1175_, _1232_, _1220_, _1228_ };
assign _0183_ = | { _0923_, _1269_, _1287_, _1289_, _1285_, _1265_ };
assign _0184_ = | instr_rdata_i_t0[19:15];
assign _0132_ = | instr_rdata_alu_i_t0[31:27];
assign _0185_ = | instr_rdata_i_t0[11:7];
assign _0137_ = | instr_rdata_i_t0[31:20];
assign _0186_ = | _1271_;
assign _0187_ = | instr_rdata_i_t0[26:25];
assign _0139_ = | instr_rdata_i_t0[31:27];
assign _0188_ = | { _0041_, _1267_, _0061_, _1275_[5:3] };
assign _0189_ = ~ { _0061_, _0041_ };
assign _0190_ = ~ { _1228_, _1226_ };
assign _0191_ = ~ { _0017_, _0021_, _1265_ };
assign _0192_ = ~ { _0086_, _0093_, _0084_, _0102_, _0088_ };
assign _0193_ = ~ { _1289_, _1287_, _1269_, _1265_ };
assign _0194_ = ~ { _1283_, _0017_, _0021_, _1277_, _1269_, _1265_ };
assign _0195_ = ~ { _1191_, _1189_, _1187_, _1185_ };
assign _0196_ = ~ { _1183_, _1181_, _1179_, _1177_ };
assign _0197_ = ~ { _1250_, _1248_ };
assign _0198_ = ~ { _1254_, _1252_ };
assign _0199_ = ~ { _1259_, _1116_[0], _1256_ };
assign _0200_ = ~ { _1206_, _1191_, _1189_, _1187_, _1185_, _1183_, _1181_, _1179_, _1177_ };
assign _0201_ = ~ { _1259_, _1254_, _1250_ };
assign _0202_ = ~ { _1232_, _1228_ };
assign _0203_ = ~ { _1232_, _1230_, _1228_, _1226_, _1224_, _1220_ };
assign _0204_ = ~ { _1263_, _1261_, _1259_, _1116_[0], _1256_, _1254_, _1252_, _1250_, _1248_ };
assign _0205_ = ~ { _1224_, _1222_ };
assign _0206_ = ~ { _1285_, _1283_ };
assign _0207_ = ~ { _0021_, _1277_ };
assign _0208_ = ~ { _0122_[2], _0058_ };
assign _0209_ = ~ { _1114_[0], _1235_, _1112_[0] };
assign _0210_ = ~ { _1122_[1], _1114_[0] };
assign _0211_ = ~ { _1122_[1], _1114_[0], _1235_ };
assign _0212_ = ~ { _0903_, _1198_, _1049_[3], _1195_ };
assign _0213_ = ~ { _1075_[0], _1065_[2], _0907_ };
assign _0214_ = ~ { _1075_[0], _1065_[2], _1210_ };
assign _0215_ = ~ { _1230_, _1220_, _1212_, _1208_, _1175_, _1172_ };
assign _0216_ = ~ { _1212_, _1208_, _1175_ };
assign _0217_ = ~ { _1232_, _1228_, _1220_, _1175_ };
assign _0218_ = ~ { _0923_, _1289_, _1287_, _1285_, _1269_, _1265_ };
assign _0152_ = ~ instr_rdata_i_t0[14:12];
assign _0219_ = ~ instr_rdata_i_t0[19:15];
assign _0220_ = ~ instr_rdata_i_t0[11:7];
assign _0149_ = ~ instr_rdata_i_t0[31:20];
assign _0221_ = ~ _1271_;
assign _0222_ = ~ instr_rdata_i_t0[26:25];
assign _0223_ = ~ { _1275_[5:3], _1267_, _0061_, _0041_ };
assign _0414_ = { _1244_, _0336_ } & _0189_;
assign _0415_ = { _1227_, _1225_ } & _0190_;
assign _0416_ = { _1281_, _1279_, _1264_ } & _0191_;
assign _0417_ = { _1243_, _1242_, _1241_, _1240_, _1239_ } & _0192_;
assign _0418_ = { _1288_, _1286_, _1268_, _1264_ } & _0193_;
assign _0419_ = { _1282_, _1281_, _1279_, _1276_, _1268_, _1264_ } & _0194_;
assign _0420_ = { _1190_, _1188_, _1186_, _1184_ } & _0195_;
assign _0421_ = { _1182_, _1180_, _1178_, _1176_ } & _0196_;
assign _0422_ = { _1249_, _1247_ } & _0197_;
assign _0423_ = { _1253_, _1251_ } & _0198_;
assign _0424_ = { _1258_, _1257_, _1255_ } & _0199_;
assign _0425_ = { _1205_, _1190_, _1188_, _1186_, _1184_, _1182_, _1180_, _1178_, _1176_ } & _0200_;
assign _0426_ = { _1258_, _1253_, _1249_ } & _0201_;
assign _0427_ = { _1231_, _1227_ } & _0202_;
assign _0428_ = { _1231_, _1229_, _1227_, _1225_, _1223_, _1219_ } & _0203_;
assign _0429_ = { _1262_, _1260_, _1258_, _1257_, _1255_, _1253_, _1251_, _1249_, _1247_ } & _0204_;
assign _0430_ = { _1223_, _1221_ } & _0205_;
assign _0431_ = { _1284_, _1282_ } & _0206_;
assign _0432_ = { _1279_, _1276_ } & _0207_;
assign _0433_ = { _1173_, _1160_ } & _0208_;
assign _0434_ = { _1236_, _1234_, _1233_ } & _0209_;
assign _0435_ = { _1278_, _1236_ } & _0210_;
assign _0436_ = { _1278_, _1236_, _1234_ } & _0211_;
assign _0473_ = { _0902_, _1197_, _1196_, _1194_ } & _0212_;
assign _0474_ = { _1214_, _1213_, _0906_ } & _0213_;
assign _0475_ = { _1214_, _1213_, _1209_ } & _0214_;
assign _0476_ = { _1229_, _1219_, _1211_, _1207_, _1174_, _1171_ } & _0215_;
assign _0477_ = { _1211_, _1207_, _1174_ } & _0216_;
assign _0478_ = { _1231_, _1227_, _1219_, _1174_ } & _0217_;
assign _0479_ = { _0922_, _1288_, _1286_, _1284_, _1268_, _1264_ } & _0218_;
assign _0623_ = instr_rdata_i[19:15] & _0219_;
assign _0636_ = instr_rdata_i[11:7] & _0220_;
assign _0679_ = instr_rdata_i[31:20] & _0149_;
assign _0708_ = _1270_ & _0221_;
assign _0712_ = instr_rdata_i[26:25] & _0222_;
assign _0676_ = instr_rdata_i[13:12] & _0148_;
assign _0717_ = { _1274_[5:3], _1266_, _1244_, _0336_ } & _0223_;
assign _0224_ = ! _0414_;
assign _0225_ = ! _0415_;
assign _0226_ = ! _0416_;
assign _0227_ = ! _0417_;
assign _0228_ = ! _0418_;
assign _0229_ = ! _0419_;
assign _0230_ = ! _0420_;
assign _0231_ = ! _0421_;
assign _0232_ = ! _0422_;
assign _0233_ = ! _0423_;
assign _0234_ = ! _0424_;
assign _0235_ = ! _0425_;
assign _0236_ = ! _0426_;
assign _0237_ = ! _0427_;
assign _0238_ = ! _0428_;
assign _0239_ = ! _0429_;
assign _0240_ = ! _0430_;
assign _0241_ = ! _0431_;
assign _0242_ = ! _0432_;
assign _0243_ = ! _0433_;
assign _0244_ = ! _0434_;
assign _0245_ = ! _0435_;
assign _0246_ = ! _0436_;
assign _0247_ = ! _0473_;
assign _0248_ = ! _0474_;
assign _0249_ = ! _0475_;
assign _0250_ = ! _0476_;
assign _0251_ = ! _0477_;
assign _0252_ = ! _0478_;
assign _0253_ = ! _0479_;
assign _0254_ = ! _0623_;
assign _0255_ = ! _0625_;
assign _0256_ = ! _0635_;
assign _0257_ = ! _0636_;
assign _0258_ = ! _0639_;
assign _0259_ = ! _0648_;
assign _0260_ = ! _0679_;
assign _0261_ = ! _0699_;
assign _0262_ = ! _0708_;
assign _0263_ = ! _0712_;
assign _0264_ = ! _0709_;
assign _0265_ = ! _0676_;
assign _0266_ = ! _0717_;
assign _0033_ = _0224_ & _0154_;
assign _0387_ = _0225_ & _0155_;
assign rf_ren_b_o_t0 = _0226_ & _0156_;
assign _0037_ = _0227_ & _0157_;
assign _0390_ = _0228_ & _0158_;
assign _0394_ = _0229_ & _0159_;
assign _0095_ = _0230_ & _0160_;
assign _0082_ = _0231_ & _0161_;
assign _0398_ = _0232_ & _0162_;
assign _0400_ = _0233_ & _0163_;
assign _0402_ = _0234_ & _0164_;
assign _0404_ = _0235_ & _0165_;
assign _0406_ = _0236_ & _0166_;
assign _0408_ = _0237_ & _0167_;
assign _0410_ = _0238_ & _0168_;
assign _0031_ = _0239_ & _0169_;
assign _0413_ = _0240_ & _0170_;
assign _0392_ = _0241_ & _0171_;
assign _0019_ = _0242_ & _0172_;
assign _0013_[5] = _0243_ & _0173_;
assign _0078_ = _0244_ & _0174_;
assign _0368_ = _0245_ & _0175_;
assign _0370_ = _0246_ & _0176_;
assign _0372_ = _0247_ & _0177_;
assign _0374_ = _0248_ & _0178_;
assign _0376_ = _0249_ & _0179_;
assign _0378_ = _0250_ & _0180_;
assign _0380_ = _0251_ & _0181_;
assign _0382_ = _0252_ & _0182_;
assign _0384_ = _0253_ & _0183_;
assign _1153_ = _0254_ & _0184_;
assign _1158_ = _0255_ & _0132_;
assign _0041_ = _0256_ & _0140_;
assign _1170_ = _0257_ & _0185_;
assign _1206_ = _0258_ & _0133_;
assign _0058_ = _0259_ & _0134_;
assign _0088_ = _0260_ & _0137_;
assign _1263_[0] = _0261_ & _0138_;
assign _1273_ = _0262_ & _0186_;
assign _1154_ = _0263_ & _0187_;
assign _1271_[0] = _0264_ & _0139_;
assign _1122_[1] = _0265_ & _0136_;
assign _0090_ = _0266_ & _0188_;
assign _0267_ = ~ _1148_;
assign _0268_ = ~ _1168_;
assign _0269_ = ~ _1150_;
assign _0270_ = ~ _1169_;
assign _0629_ = _1149_ & _0269_;
assign _0632_ = _1153_ & _0270_;
assign _0630_ = _1151_ & _0267_;
assign _0633_ = _1170_ & _0268_;
assign _0631_ = _1149_ & _1151_;
assign _0634_ = _1153_ & _1170_;
assign _0877_ = _0629_ | _0630_;
assign _0878_ = _0632_ | _0633_;
assign _1164_ = _0877_ | _0631_;
assign _1166_ = _0878_ | _0634_;
assign _0271_ = ~ { _1160_, _1160_ };
assign _0272_ = ~ { _1173_, _1173_ };
assign _0273_ = ~ { _1194_, _1194_, _1194_, _1194_, _1194_, _1194_, _1194_ };
assign _0274_ = ~ { _0902_, _0902_, _0902_, _0902_, _0902_, _0902_, _0902_ };
assign _0275_ = ~ { _1202_, _1202_, _1202_, _1202_, _1202_, _1202_, _1202_ };
assign _0276_ = ~ { _0904_, _0904_, _0904_, _0904_, _0904_, _0904_, _0904_ };
assign _0277_ = ~ { _0371_, _0371_, _0371_, _0371_, _0371_, _0371_, _0371_ };
assign _0278_ = ~ { _1213_, _1213_, _1213_, _1213_, _1213_, _1213_, _1213_ };
assign _0279_ = ~ { _0906_, _0906_, _0906_, _0906_, _0906_, _0906_, _0906_ };
assign _0280_ = ~ { _0908_, _0908_, _0908_, _0908_, _0908_, _0908_, _0908_ };
assign _0281_ = ~ { _0373_, _0373_, _0373_, _0373_, _0373_, _0373_, _0373_ };
assign _0282_ = ~ { _0910_, _0910_, _0910_, _0910_, _0910_, _0910_, _0910_ };
assign _0283_ = ~ { _0375_, _0375_, _0375_, _0375_, _0375_, _0375_, _0375_ };
assign _0284_ = ~ _1207_;
assign _0285_ = ~ _1221_;
assign _0286_ = ~ _0912_;
assign _0287_ = ~ { _1171_, _1171_ };
assign _0288_ = ~ { _0386_, _0386_ };
assign _0289_ = ~ { _0377_, _0377_ };
assign _0290_ = ~ { _1207_, _1207_, _1207_, _1207_, _1207_, _1207_, _1207_ };
assign _0291_ = ~ { _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_ };
assign _0292_ = ~ { _0409_, _0409_, _0409_, _0409_, _0409_, _0409_, _0409_ };
assign _0293_ = ~ { _0379_, _0379_, _0379_, _0379_, _0379_, _0379_, _0379_ };
assign _0294_ = ~ { _0407_, _0407_, _0407_ };
assign _0295_ = ~ { _1174_, _1174_, _1174_ };
assign _0296_ = ~ { _1221_, _1221_, _1221_ };
assign _0297_ = ~ { _0914_, _0914_, _0914_ };
assign _0298_ = ~ { _0381_, _0381_, _0381_ };
assign _0299_ = ~ { _1236_, _1236_ };
assign _0300_ = ~ { _0916_, _0916_ };
assign _0301_ = ~ { _0405_, _0405_ };
assign _0302_ = ~ { _0918_, _0918_ };
assign _0303_ = ~ _1266_;
assign _0304_ = ~ _1234_;
assign _0305_ = ~ _1237_;
assign _0306_ = ~ _0920_;
assign _0307_ = ~ _1245_;
assign _0308_ = ~ _1264_;
assign _0309_ = ~ _0922_;
assign _0310_ = ~ _1276_;
assign _0311_ = ~ _1281_;
assign _0312_ = ~ _0924_;
assign _0313_ = ~ _0383_;
assign _0314_ = ~ instr_rdata_alu_i[26];
assign _0315_ = ~ { instr_rdata_alu_i[26], instr_rdata_alu_i[26], instr_rdata_alu_i[26], instr_rdata_alu_i[26], instr_rdata_alu_i[26], instr_rdata_alu_i[26], instr_rdata_alu_i[26] };
assign _0316_ = ~ { _1157_, _1157_, _1157_, _1157_, _1157_, _1157_, _1157_ };
assign _0317_ = ~ { instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i };
assign _0318_ = ~ illegal_insn_o;
assign _0319_ = ~ illegal_c_insn_i;
assign _0320_ = ~ instr_rdata_i[14];
assign _0321_ = ~ _1165_;
assign _0322_ = ~ _0336_;
assign _0323_ = ~ { _0336_, _0336_ };
assign _0324_ = ~ _1155_;
assign _0325_ = ~ { _1155_, _1155_ };
assign _0326_ = ~ instr_rdata_i[26];
assign _0327_ = ~ _1279_;
assign _0328_ = ~ { _1161_, _1161_ };
assign _0759_ = { _0058_, _0058_ } | _0271_;
assign _0760_ = { _0122_[2], _0122_[2] } | _0272_;
assign _0761_ = { _1195_, _1195_, _1195_, _1195_, _1195_, _1195_, _1195_ } | _0273_;
assign _0762_ = { _0903_, _0903_, _0903_, _0903_, _0903_, _0903_, _0903_ } | _0274_;
assign _0765_ = { _1203_, _1203_, _1203_, _1203_, _1203_, _1203_, _1203_ } | _0275_;
assign _0766_ = { _0905_, _0905_, _0905_, _0905_, _0905_, _0905_, _0905_ } | _0276_;
assign _0769_ = { _0372_, _0372_, _0372_, _0372_, _0372_, _0372_, _0372_ } | _0277_;
assign _0773_ = { _1065_[2], _1065_[2], _1065_[2], _1065_[2], _1065_[2], _1065_[2], _1065_[2] } | _0278_;
assign _0774_ = { _0907_, _0907_, _0907_, _0907_, _0907_, _0907_, _0907_ } | _0279_;
assign _0777_ = { _0909_, _0909_, _0909_, _0909_, _0909_, _0909_, _0909_ } | _0280_;
assign _0780_ = { _0374_, _0374_, _0374_, _0374_, _0374_, _0374_, _0374_ } | _0281_;
assign _0783_ = { _0911_, _0911_, _0911_, _0911_, _0911_, _0911_, _0911_ } | _0282_;
assign _0786_ = { _0376_, _0376_, _0376_, _0376_, _0376_, _0376_, _0376_ } | _0283_;
assign _0789_ = _1208_ | _0284_;
assign _0792_ = _0913_ | _0286_;
assign _0796_ = { _1172_, _1172_ } | _0287_;
assign _0800_ = { _0387_, _0387_ } | _0288_;
assign _0801_ = { _0378_, _0378_ } | _0289_;
assign _0804_ = { _1208_, _1208_, _1208_, _1208_, _1208_, _1208_, _1208_ } | _0290_;
assign _0807_ = { _1175_, _1175_, _1175_, _1175_, _1175_, _1175_, _1175_ } | _0291_;
assign _0811_ = { _0410_, _0410_, _0410_, _0410_, _0410_, _0410_, _0410_ } | _0292_;
assign _0812_ = { _0380_, _0380_, _0380_, _0380_, _0380_, _0380_, _0380_ } | _0293_;
assign _0815_ = { _0408_, _0408_, _0408_ } | _0294_;
assign _0816_ = { _1175_, _1175_, _1175_ } | _0295_;
assign _0819_ = { _1222_, _1222_, _1222_ } | _0296_;
assign _0823_ = { _0915_, _0915_, _0915_ } | _0297_;
assign _0826_ = { _0382_, _0382_, _0382_ } | _0298_;
assign _0829_ = { _1114_[0], _1114_[0] } | _0299_;
assign _0830_ = { _0917_, _0917_ } | _0300_;
assign _0833_ = { _0406_, _0406_ } | _0301_;
assign _0834_ = { _0919_, _0919_ } | _0302_;
assign _0838_ = _1267_ | _0303_;
assign _0841_ = _1235_ | _0304_;
assign _0844_ = _1238_ | _0305_;
assign _0847_ = _0921_ | _0306_;
assign _0850_ = _1246_ | _0307_;
assign _0856_ = _1265_ | _0308_;
assign _0859_ = _0923_ | _0309_;
assign _0862_ = _1277_ | _0310_;
assign _0866_ = _0017_ | _0311_;
assign _0869_ = _0925_ | _0312_;
assign _0872_ = _0384_ | _0313_;
assign _0879_ = instr_rdata_alu_i_t0[26] | _0314_;
assign _0880_ = { instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26] } | _0315_;
assign _0881_ = { _1158_, _1158_, _1158_, _1158_, _1158_, _1158_, _1158_ } | _0316_;
assign _0883_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0 } | _0317_;
assign _0885_ = illegal_insn_o_t0 | _0318_;
assign _0886_ = illegal_c_insn_i_t0 | _0319_;
assign _0887_ = _1166_ | _0321_;
assign _0888_ = _0041_ | _0322_;
assign _0891_ = { _0041_, _0041_ } | _0323_;
assign _0892_ = _1156_ | _0324_;
assign _0893_ = { _1156_, _1156_ } | _0325_;
assign _0895_ = instr_rdata_i_t0[26] | _0326_;
assign _0901_ = { _1162_, _1162_ } | _0328_;
assign _0763_ = { _0903_, _0903_, _0903_, _0903_, _0903_, _0903_, _0903_ } | { _0902_, _0902_, _0902_, _0902_, _0902_, _0902_, _0902_ };
assign _0767_ = { _0905_, _0905_, _0905_, _0905_, _0905_, _0905_, _0905_ } | { _0904_, _0904_, _0904_, _0904_, _0904_, _0904_, _0904_ };
assign _0770_ = { _0372_, _0372_, _0372_, _0372_, _0372_, _0372_, _0372_ } | { _0371_, _0371_, _0371_, _0371_, _0371_, _0371_, _0371_ };
assign _0772_ = { _1210_, _1210_, _1210_, _1210_, _1210_, _1210_, _1210_ } | { _1209_, _1209_, _1209_, _1209_, _1209_, _1209_, _1209_ };
assign _0775_ = { _0907_, _0907_, _0907_, _0907_, _0907_, _0907_, _0907_ } | { _0906_, _0906_, _0906_, _0906_, _0906_, _0906_, _0906_ };
assign _0778_ = { _0909_, _0909_, _0909_, _0909_, _0909_, _0909_, _0909_ } | { _0908_, _0908_, _0908_, _0908_, _0908_, _0908_, _0908_ };
assign _0781_ = { _0374_, _0374_, _0374_, _0374_, _0374_, _0374_, _0374_ } | { _0373_, _0373_, _0373_, _0373_, _0373_, _0373_, _0373_ };
assign _0784_ = { _0911_, _0911_, _0911_, _0911_, _0911_, _0911_, _0911_ } | { _0910_, _0910_, _0910_, _0910_, _0910_, _0910_, _0910_ };
assign _0787_ = { _0376_, _0376_, _0376_, _0376_, _0376_, _0376_, _0376_ } | { _0375_, _0375_, _0375_, _0375_, _0375_, _0375_, _0375_ };
assign _0790_ = _1208_ | _1207_;
assign _0791_ = _1222_ | _1221_;
assign _0793_ = _0913_ | _0912_;
assign _0795_ = { _1175_, _1175_ } | { _1174_, _1174_ };
assign _0797_ = { _1172_, _1172_ } | { _1171_, _1171_ };
assign _0799_ = { _0413_, _0413_ } | { _0412_, _0412_ };
assign _0802_ = { _0378_, _0378_ } | { _0377_, _0377_ };
assign _0805_ = { _1208_, _1208_, _1208_, _1208_, _1208_, _1208_, _1208_ } | { _1207_, _1207_, _1207_, _1207_, _1207_, _1207_, _1207_ };
assign _0808_ = { _1175_, _1175_, _1175_, _1175_, _1175_, _1175_, _1175_ } | { _1174_, _1174_, _1174_, _1174_, _1174_, _1174_, _1174_ };
assign _0810_ = { _1222_, _1222_, _1222_, _1222_, _1222_, _1222_, _1222_ } | { _1221_, _1221_, _1221_, _1221_, _1221_, _1221_, _1221_ };
assign _0813_ = { _0380_, _0380_, _0380_, _0380_, _0380_, _0380_, _0380_ } | { _0379_, _0379_, _0379_, _0379_, _0379_, _0379_, _0379_ };
assign _0817_ = { _1175_, _1175_, _1175_ } | { _1174_, _1174_, _1174_ };
assign _0820_ = { _1222_, _1222_, _1222_ } | { _1221_, _1221_, _1221_ };
assign _0822_ = { _1226_, _1226_, _1226_ } | { _1225_, _1225_, _1225_ };
assign _0824_ = { _0915_, _0915_, _0915_ } | { _0914_, _0914_, _0914_ };
assign _0827_ = { _0382_, _0382_, _0382_ } | { _0381_, _0381_, _0381_ };
assign _0831_ = { _0917_, _0917_ } | { _0916_, _0916_ };
assign _0835_ = { _0919_, _0919_ } | { _0918_, _0918_ };
assign _0837_ = _0061_ | _1244_;
assign _0839_ = _1267_ | _1266_;
assign _0842_ = _1235_ | _1234_;
assign _0845_ = _1238_ | _1237_;
assign _0846_ = _0392_ | _0391_;
assign _0848_ = _0921_ | _0920_;
assign _0851_ = _1246_ | _1245_;
assign _0855_ = _1269_ | _1268_;
assign _0857_ = _1265_ | _1264_;
assign _0860_ = _0923_ | _0922_;
assign _0863_ = _1277_ | _1276_;
assign _0865_ = _1283_ | _1282_;
assign _0867_ = _0017_ | _1281_;
assign _0870_ = _0925_ | _0924_;
assign _0873_ = _0384_ | _0383_;
assign _0882_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0 } | { instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i };
assign _0884_ = _1172_ | _1171_;
assign _0889_ = _0041_ | _0336_;
assign _0894_ = _1273_ | _1272_;
assign _0896_ = _1271_[0] | _1270_[0];
assign _0897_ = _0370_ | _0369_;
assign _0898_ = { _0019_, _0019_ } | { _0411_, _0411_ };
assign _0899_ = { _1265_, _1265_ } | { _1264_, _1264_ };
assign _0900_ = { _1238_, _1238_ } | { _1237_, _1237_ };
assign _0480_ = { _0058_, _0058_ } & _0760_;
assign _0482_ = { 3'h0, _1049_[3], _1049_[3], _1049_[3], 1'h0 } & _0761_;
assign _0484_ = _1051_ & _0762_;
assign _0487_ = { 1'h0, _1057_[5], 1'h0, _1057_[5], _1057_[5], 1'h0, _1057_[5] } & _0765_;
assign _0489_ = _1059_ & _0766_;
assign _0492_ = _1061_ & _0769_;
assign _0497_ = { 4'h0, _1065_[2], _1065_[2], _1065_[2] } & _0774_;
assign _0500_ = { 1'h0, _1071_[5], 1'h0, _1071_[5], 1'h0, _1071_[5], _1071_[5] } & _0777_;
assign _0503_ = _1073_ & _0780_;
assign _0506_ = { 6'h00, _1075_[0] } & _0773_;
assign _0508_ = { 1'h0, _0058_, _0058_, 3'h0, _0058_ } & _0783_;
assign _0511_ = _1081_ & _0786_;
assign _0514_ = instr_rdata_alu_i_t0[14] & _0789_;
assign _0518_ = _1085_ & _0792_;
assign _0523_ = _1087_ & _0796_;
assign _0528_ = _1091_ & _0800_;
assign _0530_ = _1093_ & _0801_;
assign _0533_ = _0120_ & _0804_;
assign _0536_ = _1095_ & _0807_;
assign _0541_ = _1098_ & _0811_;
assign _0543_ = _1100_ & _0812_;
assign _0546_ = { 2'h0, instr_rdata_alu_i_t0[14] } & _0815_;
assign _0548_ = _1102_ & _0816_;
assign _0551_ = { instr_first_cycle_i_t0, 1'h0, instr_first_cycle_i_t0 } & _0819_;
assign _0556_ = _1108_ & _0823_;
assign _0559_ = _1110_ & _0826_;
assign _0562_ = { 1'h0, _1114_[0] } & _0830_;
assign _0565_ = { 1'h0, _1116_[0] } & _0833_;
assign _0567_ = { 1'h0, _0402_ } & _0834_;
assign _0572_ = _1120_ & _0838_;
assign _0575_ = { _1122_[1], 1'h0 } & _0829_;
assign _0577_ = _0368_ & _0841_;
assign _0584_ = _1127_ & _0847_;
assign _0588_ = _1129_ & _0850_;
assign _0591_ = _0392_ & _0850_;
assign _0594_ = _0033_ & _0844_;
assign _0599_ = _1134_ & _0856_;
assign _0602_ = _1136_ & _0859_;
assign _0605_ = _0111_ & _0862_;
assign _0610_ = _1142_ & _0866_;
assign _0613_ = _1144_ & _0869_;
assign _0616_ = _1146_ & _0872_;
assign _0619_ = _0394_ & _0844_;
assign _0637_ = { instr_rdata_alu_i_t0[14], instr_rdata_alu_i_t0[14] } & _0759_;
assign _0640_ = _0082_ & _0879_;
assign _0642_ = _0095_ & _0879_;
assign _0644_ = _0009_ & _0880_;
assign _0646_ = { 1'h0, _0003_[5], 2'h0, _0003_[5], 2'h0 } & _0881_;
assign _0651_ = { branch_taken_i_t0, branch_taken_i_t0, branch_taken_i_t0 } & _0883_;
assign _0660_ = rf_wdata_sel_o_t0 & _0885_;
assign _0662_ = _0017_ & _0885_;
assign _0664_ = _0027_ & _0885_;
assign _0666_ = _0025_ & _0885_;
assign _0668_ = _0021_ & _0885_;
assign _0670_ = _0019_ & _0885_;
assign _0672_ = _0029_ & _0885_;
assign _0674_ = _0023_ & _0886_;
assign _0677_ = _0037_ & _0887_;
assign _0680_ = _0078_ & _0888_;
assign _0693_ = instr_rdata_i_t0[14] & _0888_;
assign _0695_ = _0080_ & _0891_;
assign _0700_ = _0031_ & _0892_;
assign _0702_ = _0099_ & _0893_;
assign _0704_ = _0097_ & _0893_;
assign _0710_ = _0011_ & _0895_;
assign _0741_ = csr_op_t0 & _0901_;
assign _0743_ = mult_sel_o_t0 & _0885_;
assign _0745_ = div_sel_o_t0 & _0885_;
assign _0485_ = { 3'h0, _0404_, 3'h0 } & _0763_;
assign _0490_ = { 6'h00, _1055_[0] } & _0767_;
assign _0493_ = _1053_ & _0770_;
assign _0495_ = _0001_ & _0772_;
assign _0498_ = _1063_ & _0775_;
assign _0501_ = { 1'h0, _1069_[5], 1'h0, _1069_[5], _1069_[5], _1069_[5], 1'h0 } & _0778_;
assign _0504_ = _1067_ & _0781_;
assign _0509_ = { 4'h0, _1069_[5], _1069_[5], _1069_[5] } & _0784_;
assign _0512_ = _1077_ & _0787_;
assign _0516_ = instr_first_cycle_i_t0 & _0791_;
assign _0519_ = _1083_ & _0793_;
assign _0521_ = _0114_ & _0795_;
assign _0524_ = _0124_ & _0797_;
assign _0526_ = { instr_first_cycle_i_t0, 1'h0 } & _0799_;
assign _0531_ = _1089_ & _0802_;
assign _0534_ = _0005_ & _0805_;
assign _0537_ = { 1'h0, _0013_[5], 1'h0, _0013_[5], _0013_[5], 2'h0 } & _0808_;
assign _0539_ = _0109_ & _0810_;
assign _0544_ = _1097_ & _0813_;
assign _0549_ = { _0122_[2], 1'h0, _0122_[2] } & _0817_;
assign _0552_ = _0107_ & _0820_;
assign _0554_ = { 2'h0, instr_first_cycle_i_t0 } & _0822_;
assign _0557_ = _1106_ & _0824_;
assign _0560_ = _1104_ & _0827_;
assign _0563_ = { 1'h0, _1112_[0] } & _0831_;
assign _0568_ = { 1'h0, _0398_ } & _0835_;
assign _0570_ = _0129_ & _0837_;
assign _0573_ = _0007_ & _0839_;
assign _0578_ = instr_rdata_i_t0[14] & _0842_;
assign _0580_ = _0041_ & _0845_;
assign _0582_ = instr_first_cycle_i_t0 & _0846_;
assign _0585_ = _1125_ & _0848_;
assign _0589_ = _0055_ & _0851_;
assign _0592_ = _0061_ & _0851_;
assign _0595_ = _0035_ & _0845_;
assign _0597_ = _0126_ & _0855_;
assign _0600_ = _0015_ & _0857_;
assign _0603_ = _1132_ & _0860_;
assign _0606_ = _0117_ & _0863_;
assign _0608_ = _0041_ & _0865_;
assign _0611_ = _0090_ & _0867_;
assign _0614_ = _1140_ & _0870_;
assign _0617_ = _1138_ & _0873_;
assign _0620_ = _0072_ & _0845_;
assign _0649_ = _0104_ & _0882_;
assign _0654_ = _0047_ & _0790_;
assign _0656_ = _0066_ & _0790_;
assign _0658_ = _0058_ & _0884_;
assign _0681_ = _0039_ & _0889_;
assign _0683_ = _0102_ & _0889_;
assign _0685_ = _0088_ & _0889_;
assign _0687_ = _0084_ & _0889_;
assign _0689_ = _0093_ & _0889_;
assign _0691_ = _0086_ & _0889_;
assign _0697_ = instr_first_cycle_i_t0 & _0837_;
assign _0706_ = _1154_ & _0894_;
assign _0713_ = _1154_ & _0896_;
assign _0715_ = instr_rdata_i_t0[14] & _0897_;
assign _0719_ = instr_rdata_i_t0[14] & _0863_;
assign _0721_ = _0045_ & _0898_;
assign _0723_ = _0070_ & _0899_;
assign _0725_ = _0068_ & _0899_;
assign _0728_ = _0075_ & _0845_;
assign _0730_ = _0053_ & _0845_;
assign _0732_ = _0049_ & _0845_;
assign _0734_ = _0064_ & _0845_;
assign _0736_ = _0051_ & _0845_;
assign _0739_ = _0043_ & _0900_;
assign _0764_ = _0484_ | _0485_;
assign _0768_ = _0489_ | _0490_;
assign _0771_ = _0492_ | _0493_;
assign _0776_ = _0497_ | _0498_;
assign _0779_ = _0500_ | _0501_;
assign _0782_ = _0503_ | _0504_;
assign _0785_ = _0508_ | _0509_;
assign _0788_ = _0511_ | _0512_;
assign _0794_ = _0518_ | _0519_;
assign _0798_ = _0523_ | _0524_;
assign _0803_ = _0530_ | _0531_;
assign _0806_ = _0533_ | _0534_;
assign _0809_ = _0536_ | _0537_;
assign _0814_ = _0543_ | _0544_;
assign _0818_ = _0548_ | _0549_;
assign _0821_ = _0551_ | _0552_;
assign _0825_ = _0556_ | _0557_;
assign _0828_ = _0559_ | _0560_;
assign _0832_ = _0562_ | _0563_;
assign _0836_ = _0567_ | _0568_;
assign _0840_ = _0572_ | _0573_;
assign _0843_ = _0577_ | _0578_;
assign _0849_ = _0584_ | _0585_;
assign _0852_ = _0588_ | _0589_;
assign _0853_ = _0591_ | _0592_;
assign _0854_ = _0594_ | _0595_;
assign _0858_ = _0599_ | _0600_;
assign _0861_ = _0602_ | _0603_;
assign _0864_ = _0605_ | _0606_;
assign _0868_ = _0610_ | _0611_;
assign _0871_ = _0613_ | _0614_;
assign _0874_ = _0616_ | _0617_;
assign _0875_ = _0619_ | _0620_;
assign _0890_ = _0680_ | _0681_;
assign _0928_ = _1050_ ^ _1047_;
assign _0930_ = _1058_ ^ _1054_;
assign _0931_ = _1060_ ^ _1052_;
assign _0932_ = _1064_ ^ _1062_;
assign _0933_ = _1070_ ^ _1068_;
assign _0934_ = _1072_ ^ _1066_;
assign _0936_ = _1079_ ^ _1078_;
assign _0937_ = _1080_ ^ _1076_;
assign _0938_ = _1084_ ^ _1082_;
assign _0939_ = _1086_ ^ _0123_;
assign _0941_ = _1092_ ^ _1088_;
assign _0942_ = _0119_ ^ _0004_;
assign _0943_ = _1094_ ^ _0012_;
assign _0945_ = _1099_ ^ _1096_;
assign _0946_ = _1101_ ^ _0121_;
assign _0947_ = _0091_ ^ _0106_;
assign _0948_ = _1107_ ^ _1105_;
assign _0949_ = _1109_ ^ _1103_;
assign _0950_ = _1113_ ^ _1111_;
assign _0951_ = _1118_ ^ _1117_;
assign _0952_ = _1119_ ^ _0006_;
assign _0954_ = _1123_ ^ _0105_;
assign _0955_ = _1126_ ^ _1124_;
assign _0956_ = _1128_ ^ _0054_;
assign _0957_ = _1130_ ^ _0060_;
assign _0958_ = _0032_ ^ _0034_;
assign _0959_ = _1133_ ^ _0014_;
assign _0960_ = _1135_ ^ _1131_;
assign _0961_ = _0110_ ^ _0116_;
assign _0962_ = _1141_ ^ _0089_;
assign _0963_ = _1143_ ^ _1139_;
assign _0964_ = _1145_ ^ _1137_;
assign _0965_ = _1147_ ^ _0071_;
assign _0966_ = _0077_ ^ _0038_;
assign _0481_ = { _0122_[2], _0122_[2] } & { _0342_, _0926_[0] };
assign _0483_ = { _1195_, _1195_, _1195_, _1195_, _1195_, _1195_, _1195_ } & { _0927_[6:4], _0347_[1], _0927_[2:1], _0347_[0] };
assign _0486_ = { _0903_, _0903_, _0903_, _0903_, _0903_, _0903_, _0903_ } & _0928_;
assign _0488_ = { _1203_, _1203_, _1203_, _1203_, _1203_, _1203_, _1203_ } & { _0929_[6], _0341_[3], _0929_[4], _0341_[2], _0929_[2], _0341_[1:0] };
assign _0491_ = { _0905_, _0905_, _0905_, _0905_, _0905_, _0905_, _0905_ } & _0930_;
assign _0494_ = { _0372_, _0372_, _0372_, _0372_, _0372_, _0372_, _0372_ } & _0931_;
assign _0496_ = { _1210_, _1210_, _1210_, _1210_, _1210_, _1210_, _1210_ } & { _0000_[6:4], _0339_[1], _0000_[2], _0339_[0], _0000_[0] };
assign _0499_ = { _0907_, _0907_, _0907_, _0907_, _0907_, _0907_, _0907_ } & _0932_;
assign _0502_ = { _0909_, _0909_, _0909_, _0909_, _0909_, _0909_, _0909_ } & _0933_;
assign _0505_ = { _0374_, _0374_, _0374_, _0374_, _0374_, _0374_, _0374_ } & _0934_;
assign _0507_ = { _1065_[2], _1065_[2], _1065_[2], _1065_[2], _1065_[2], _1065_[2], _1065_[2] } & { _0935_[6:5], _0345_, _0935_[1:0] };
assign _0510_ = { _0911_, _0911_, _0911_, _0911_, _0911_, _0911_, _0911_ } & _0936_;
assign _0513_ = { _0376_, _0376_, _0376_, _0376_, _0376_, _0376_, _0376_ } & _0937_;
assign _0515_ = _1208_ & _0115_;
assign _0517_ = _1222_ & instr_first_cycle_i;
assign _0520_ = _0913_ & _0938_;
assign _0522_ = { _1175_, _1175_ } & _0113_;
assign _0525_ = { _1172_, _1172_ } & _0939_;
assign _0527_ = { _0413_, _0413_ } & _0343_;
assign _0529_ = { _0387_, _0387_ } & { _0344_, _0940_[0] };
assign _0532_ = { _0378_, _0378_ } & _0941_;
assign _0535_ = { _1208_, _1208_, _1208_, _1208_, _1208_, _1208_, _1208_ } & _0942_;
assign _0538_ = { _1175_, _1175_, _1175_, _1175_, _1175_, _1175_, _1175_ } & _0943_;
assign _0540_ = { _1222_, _1222_, _1222_, _1222_, _1222_, _1222_, _1222_ } & { _0108_[6], _0346_[2], _0108_[4], _0346_[1:0], _0108_[1:0] };
assign _0542_ = { _0410_, _0410_, _0410_, _0410_, _0410_, _0410_, _0410_ } & _0944_;
assign _0545_ = { _0380_, _0380_, _0380_, _0380_, _0380_, _0380_, _0380_ } & _0945_;
assign _0547_ = { _0408_, _0408_, _0408_ } & { _0118_[2], _0350_ };
assign _0550_ = { _1175_, _1175_, _1175_ } & _0946_;
assign _0553_ = { _1222_, _1222_, _1222_ } & _0947_;
assign _0555_ = { _1226_, _1226_, _1226_ } & _0059_;
assign _0558_ = { _0915_, _0915_, _0915_ } & _0948_;
assign _0561_ = { _0382_, _0382_, _0382_ } & _0949_;
assign _0564_ = { _0917_, _0917_ } & _0950_;
assign _0566_ = { _0406_, _0406_ } & _0340_;
assign _0569_ = { _0919_, _0919_ } & _0951_;
assign _0571_ = _0061_ & _0128_;
assign _0574_ = _1267_ & _0952_;
assign _0576_ = { _1114_[0], _1114_[0] } & { _0953_[1], _0349_ };
assign _0579_ = _1235_ & _0954_;
assign _0581_ = _1238_ & _0336_;
assign _0583_ = _0392_ & _0073_;
assign _0586_ = _0921_ & _0955_;
assign _0587_ = _0392_ & _0062_;
assign _0590_ = _1246_ & _0956_;
assign _0593_ = _1246_ & _0957_;
assign _0596_ = _1238_ & _0958_;
assign _0598_ = _1269_ & _0125_;
assign _0601_ = _1265_ & _0959_;
assign _0604_ = _0923_ & _0960_;
assign _0607_ = _1277_ & _0961_;
assign _0609_ = _1283_ & _0333_;
assign _0612_ = _0017_ & _0962_;
assign _0615_ = _0925_ & _0963_;
assign _0618_ = _0384_ & _0964_;
assign _0621_ = _1238_ & _0965_;
assign _0638_ = { _0058_, _0058_ } & _0127_;
assign _0641_ = instr_rdata_alu_i_t0[26] & _0081_;
assign _0643_ = instr_rdata_alu_i_t0[26] & _0094_;
assign _0645_ = { instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26], instr_rdata_alu_i_t0[26] } & { _0008_[6], _0348_[2], _0008_[4], _0348_[1:0], _0008_[1:0] };
assign _0647_ = { _1158_, _1158_, _1158_, _1158_, _1158_, _1158_, _1158_ } & { _0002_[6:4], _0338_[1], _0002_[2:1], _0338_[0] };
assign _0650_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0 } & _0103_;
assign _0652_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0 } & _0112_;
assign _0655_ = _1208_ & _0046_;
assign _0657_ = _1208_ & _0065_;
assign _0659_ = _1172_ & _0337_;
assign _0661_ = illegal_insn_o_t0 & rf_wdata_sel_o;
assign _0663_ = illegal_insn_o_t0 & _0016_;
assign _0665_ = illegal_insn_o_t0 & _0026_;
assign _0667_ = illegal_insn_o_t0 & _0024_;
assign _0669_ = illegal_insn_o_t0 & _0020_;
assign _0671_ = illegal_insn_o_t0 & _0018_;
assign _0673_ = illegal_insn_o_t0 & _0028_;
assign _0675_ = illegal_c_insn_i_t0 & _0335_;
assign _0678_ = _1166_ & _0329_;
assign _0682_ = _0041_ & _0966_;
assign _0684_ = _0041_ & _0101_;
assign _0686_ = _0041_ & _0087_;
assign _0688_ = _0041_ & _0083_;
assign _0690_ = _0041_ & _0092_;
assign _0692_ = _0041_ & _0085_;
assign _0694_ = _0041_ & _0100_;
assign _0696_ = { _0041_, _0041_ } & _0079_;
assign _0698_ = _0061_ & _0062_;
assign _0701_ = _1156_ & _0332_;
assign _0703_ = { _1156_, _1156_ } & _0098_;
assign _0705_ = { _1156_, _1156_ } & _0096_;
assign _0707_ = _1273_ & _0330_;
assign _0711_ = instr_rdata_i_t0[26] & _0331_;
assign _0714_ = _1271_[0] & _0330_;
assign _0716_ = _0370_ & _0334_;
assign _0720_ = _1277_ & _0320_;
assign _0722_ = { _0019_, _0019_ } & _0044_;
assign _0724_ = { _1265_, _1265_ } & _0069_;
assign _0726_ = { _1265_, _1265_ } & _0067_;
assign _0727_ = _1238_ & _0040_;
assign _0729_ = _1238_ & _0074_;
assign _0731_ = _1238_ & _0052_;
assign _0733_ = _1238_ & _0048_;
assign _0735_ = _1238_ & _0063_;
assign _0737_ = _1238_ & _0050_;
assign _0738_ = _1246_ & _0054_;
assign _0740_ = { _1238_, _1238_ } & _0042_;
assign _0742_ = { _1162_, _1162_ } & csr_op;
assign _0744_ = illegal_insn_o_t0 & mult_sel_o;
assign _0746_ = illegal_insn_o_t0 & div_sel_o;
assign _0114_ = _0481_ | _0480_;
assign _1051_ = _0483_ | _0482_;
assign _1053_ = _0486_ | _0764_;
assign _1059_ = _0488_ | _0487_;
assign _1061_ = _0491_ | _0768_;
assign _0009_ = _0494_ | _0771_;
assign _1063_ = _0496_ | _0495_;
assign _1067_ = _0499_ | _0776_;
assign _1073_ = _0502_ | _0779_;
assign _0120_ = _0505_ | _0782_;
assign _1077_ = _0507_ | _0506_;
assign _1081_ = _0510_ | _0785_;
assign _0104_ = _0513_ | _0788_;
assign _1083_ = _0515_ | _0514_;
assign _1085_ = _0517_ | _0516_;
assign alu_op_b_mux_sel_o_t0 = _0520_ | _0794_;
assign _1087_ = _0522_ | _0521_;
assign _1089_ = _0525_ | _0798_;
assign _1091_ = _0527_ | _0526_;
assign _1093_ = _0529_ | _0528_;
assign alu_op_a_mux_sel_o_t0 = _0532_ | _0803_;
assign _1095_ = _0535_ | _0806_;
assign _1097_ = _0538_ | _0809_;
assign _1098_ = _0540_ | _0539_;
assign _1100_ = _0542_ | _0541_;
assign alu_operator_o_t0 = _0545_ | _0814_;
assign _1102_ = _0547_ | _0546_;
assign _1104_ = _0550_ | _0818_;
assign _1106_ = _0553_ | _0821_;
assign _1108_ = _0555_ | _0554_;
assign _1110_ = _0558_ | _0825_;
assign imm_b_mux_sel_o_t0 = _0561_ | _0828_;
assign _0080_ = _0564_ | _0832_;
assign _0099_ = _0566_ | _0565_;
assign _0097_ = _0569_ | _0836_;
assign _1120_ = _0571_ | _0570_;
assign _0126_ = _0574_ | _0840_;
assign _0045_ = _0576_ | _0575_;
assign _0117_ = _0579_ | _0843_;
assign _1125_ = _0581_ | _0580_;
assign _1127_ = _0583_ | _0582_;
assign _0029_ = _0586_ | _0849_;
assign _1129_ = _0587_ | _0582_;
assign _0027_ = _0590_ | _0852_;
assign _0025_ = _0593_ | _0853_;
assign _1132_ = _0596_ | _0854_;
assign _1134_ = _0598_ | _0597_;
assign _1136_ = _0601_ | _0858_;
assign _1138_ = _0604_ | _0861_;
assign _1140_ = _0607_ | _0864_;
assign _1142_ = _0609_ | _0608_;
assign _1144_ = _0612_ | _0868_;
assign _1146_ = _0615_ | _0871_;
assign _0023_ = _0618_ | _0874_;
assign rf_ren_a_o_t0 = _0621_ | _0875_;
assign _0124_ = _0638_ | _0637_;
assign _0047_ = _0641_ | _0640_;
assign _0066_ = _0643_ | _0642_;
assign _0005_ = _0645_ | _0644_;
assign _0001_ = _0647_ | _0646_;
assign _0109_ = _0650_ | _0649_;
assign _0107_ = _0652_ | _0651_;
assign div_sel_o_t0 = _0655_ | _0654_;
assign mult_sel_o_t0 = _0657_ | _0656_;
assign imm_a_mux_sel_o_t0 = _0659_ | _0658_;
assign csr_access_o_t0 = _0661_ | _0660_;
assign branch_in_dec_o_t0 = _0663_ | _0662_;
assign jump_set_o_t0 = _0665_ | _0664_;
assign jump_in_dec_o_t0 = _0667_ | _0666_;
assign data_we_o_t0 = _0669_ | _0668_;
assign data_req_o_t0 = _0671_ | _0670_;
assign rf_we_o_t0 = _0673_ | _0672_;
assign illegal_insn_o_t0 = _0675_ | _0674_;
assign _0039_ = _0678_ | _0677_;
assign _0035_ = _0682_ | _0890_;
assign _0075_ = _0684_ | _0683_;
assign _0053_ = _0686_ | _0685_;
assign _0049_ = _0688_ | _0687_;
assign _0064_ = _0690_ | _0689_;
assign _0051_ = _0692_ | _0691_;
assign _0072_ = _0694_ | _0693_;
assign _0043_ = _0696_ | _0695_;
assign _0055_ = _0698_ | _0697_;
assign _0015_ = _0701_ | _0700_;
assign _0070_ = _0703_ | _0702_;
assign _0068_ = _0705_ | _0704_;
assign _0011_ = _0707_ | _0706_;
assign _0007_ = _0711_ | _0710_;
assign _0129_ = _0714_ | _0713_;
assign _0111_ = _0716_ | _0715_;
assign data_sign_extension_o_t0 = _0720_ | _0719_;
assign data_type_o_t0 = _0722_ | _0721_;
assign multdiv_signed_mode_o_t0 = _0724_ | _0723_;
assign multdiv_operator_o_t0 = _0726_ | _0725_;
assign rf_wdata_sel_o_t0 = _0727_ | _0580_;
assign wfi_insn_o_t0 = _0729_ | _0728_;
assign ecall_insn_o_t0 = _0731_ | _0730_;
assign dret_insn_o_t0 = _0733_ | _0732_;
assign mret_insn_o_t0 = _0735_ | _0734_;
assign ebrk_insn_o_t0 = _0737_ | _0736_;
assign icache_inval_o_t0 = _0738_ | _0589_;
assign csr_op_t0 = _0740_ | _0739_;
assign csr_op_o_t0 = _0742_ | _0741_;
assign mult_en_o_t0 = _0744_ | _0743_;
assign div_en_o_t0 = _0746_ | _0745_;
assign _0331_ = ~ _0010_;
assign _0333_ = ~ _0056_;
assign _0334_ = ~ _0105_;
assign _0335_ = ~ _0022_;
assign _0337_ = ~ _0057_;
assign _0338_ = ~ { _0002_[3], _0002_[0] };
assign _0339_ = ~ { _0000_[3], _0000_[1] };
assign _0340_ = ~ _1115_;
assign _0341_ = ~ { _1056_[5], _1056_[3], _1056_[1:0] };
assign _0342_ = ~ _1046_[1];
assign _0343_ = ~ _0076_;
assign _0344_ = ~ _1090_[1];
assign _0345_ = ~ _1074_[4:2];
assign _0346_ = ~ { _0108_[5], _0108_[3:2] };
assign _0347_ = ~ { _1048_[3], _1048_[0] };
assign _0348_ = ~ { _0008_[5], _0008_[3:2] };
assign _0349_ = ~ _1121_[0];
assign _0350_ = ~ _0118_[1:0];
assign _0385_ = | { _0336_, _1244_ };
assign _0386_ = | { _1227_, _1225_ };
assign _0388_ = | { _1281_, _1279_, _1264_ };
assign _0329_ = | { _1243_, _1242_, _1241_, _1240_, _1239_ };
assign _0389_ = | { _1288_, _1286_, _1268_, _1264_ };
assign _0393_ = | { _1282_, _1281_, _1279_, _1276_, _1268_, _1264_ };
assign _0395_ = | { _1190_, _1188_, _1186_, _1184_ };
assign _0396_ = | { _1182_, _1180_, _1178_, _1176_ };
assign _0397_ = | { _1249_, _1247_ };
assign _0399_ = | { _1253_, _1251_ };
assign _0401_ = | { _1258_, _1257_, _1255_ };
assign _0403_ = | { _1205_, _1190_, _1188_, _1186_, _1184_, _1182_, _1180_, _1178_, _1176_ };
assign _0405_ = | { _1258_, _1253_, _1249_ };
assign _0407_ = | { _1231_, _1227_ };
assign _0409_ = | { _1231_, _1229_, _1227_, _1225_, _1223_, _1219_ };
assign _0332_ = | { _1262_, _1260_, _1258_, _1257_, _1255_, _1253_, _1251_, _1249_, _1247_ };
assign _0412_ = | { _1223_, _1221_ };
assign _0391_ = | { _1284_, _1282_ };
assign _0411_ = | { _1279_, _1276_ };
assign _0351_ = ~ _1192_;
assign _0352_ = ~ _1200_;
assign _0353_ = ~ _1173_;
assign _0354_ = ~ _1216_;
assign _0355_ = ~ _1219_;
assign _0356_ = ~ _1223_;
assign _0357_ = ~ _0399_;
assign _0358_ = ~ _0389_;
assign _0359_ = ~ _0403_;
assign _0360_ = ~ _1199_;
assign _0361_ = ~ _1209_;
assign _0362_ = ~ _1215_;
assign _0363_ = ~ _1233_;
assign _0364_ = ~ _0397_;
assign _0437_ = _1193_ & _0359_;
assign _0440_ = _1201_ & _0360_;
assign _0443_ = _0122_[2] & _0361_;
assign _0446_ = _1217_ & _0362_;
assign _0449_ = _0122_[2] & _0362_;
assign _0452_ = _1220_ & _0284_;
assign _0455_ = _1224_ & _0285_;
assign _0458_ = _1235_ & _0363_;
assign _0461_ = _0400_ & _0364_;
assign _0464_ = _0390_ & _0305_;
assign _0467_ = _1246_ & _0305_;
assign _0470_ = _0021_ & _0310_;
assign _0438_ = _0404_ & _0351_;
assign _0441_ = _1055_[0] & _0352_;
assign _0444_ = _1210_ & _0353_;
assign _0447_ = _1069_[5] & _0354_;
assign _0450_ = _1069_[5] & _0353_;
assign _0453_ = _1208_ & _0355_;
assign _0456_ = _1222_ & _0356_;
assign _0459_ = _1112_[0] & _0304_;
assign _0462_ = _0398_ & _0357_;
assign _0465_ = _1238_ & _0358_;
assign _0468_ = _1238_ & _0307_;
assign _0471_ = _1277_ & _0327_;
assign _0439_ = _1193_ & _0404_;
assign _0442_ = _1201_ & _1055_[0];
assign _0445_ = _0122_[2] & _1210_;
assign _0448_ = _1217_ & _1069_[5];
assign _0451_ = _0122_[2] & _1069_[5];
assign _0454_ = _1220_ & _1208_;
assign _0457_ = _1224_ & _1222_;
assign _0460_ = _1235_ & _1112_[0];
assign _0463_ = _0400_ & _0398_;
assign _0466_ = _0390_ & _1238_;
assign _0469_ = _1246_ & _1238_;
assign _0472_ = _0021_ & _1277_;
assign _0747_ = _0437_ | _0438_;
assign _0748_ = _0440_ | _0441_;
assign _0749_ = _0443_ | _0444_;
assign _0750_ = _0446_ | _0447_;
assign _0751_ = _0449_ | _0450_;
assign _0752_ = _0452_ | _0453_;
assign _0753_ = _0455_ | _0456_;
assign _0754_ = _0458_ | _0459_;
assign _0755_ = _0461_ | _0462_;
assign _0756_ = _0464_ | _0465_;
assign _0757_ = _0467_ | _0468_;
assign _0758_ = _0470_ | _0471_;
assign _0903_ = _0747_ | _0439_;
assign _0905_ = _0748_ | _0442_;
assign _0907_ = _0749_ | _0445_;
assign _0909_ = _0750_ | _0448_;
assign _0911_ = _0751_ | _0451_;
assign _0913_ = _0752_ | _0454_;
assign _0915_ = _0753_ | _0457_;
assign _0917_ = _0754_ | _0460_;
assign _0919_ = _0755_ | _0463_;
assign _0921_ = _0756_ | _0466_;
assign _0923_ = _0757_ | _0469_;
assign _0925_ = _0758_ | _0472_;
assign _0365_ = | { _1173_, _1160_ };
assign _0366_ = | { _1236_, _1234_, _1233_ };
assign _0367_ = | { _1278_, _1236_ };
assign _0369_ = | { _1278_, _1236_, _1234_ };
assign _0902_ = _1192_ | _0403_;
assign _0904_ = _1200_ | _1199_;
assign _0906_ = _1173_ | _1209_;
assign _0908_ = _1216_ | _1215_;
assign _0910_ = _1173_ | _1215_;
assign _0912_ = _1219_ | _1207_;
assign _0914_ = _1223_ | _1221_;
assign _0916_ = _1234_ | _1233_;
assign _0918_ = _0399_ | _0397_;
assign _0920_ = _0389_ | _1237_;
assign _0922_ = _1245_ | _1237_;
assign _0924_ = _1279_ | _1276_;
assign _0371_ = | { _0902_, _1197_, _1196_, _1194_ };
assign _0373_ = | { _1214_, _1213_, _0906_ };
assign _0375_ = | { _1214_, _1213_, _1209_ };
assign _0377_ = | { _1229_, _1219_, _1211_, _1207_, _1174_, _1171_ };
assign _0379_ = | { _1211_, _1207_, _1174_ };
assign _0381_ = | { _1231_, _1227_, _1219_, _1174_ };
assign _0383_ = | { _0922_, _1288_, _1286_, _1284_, _1268_, _1264_ };
assign { _1046_[1], _0926_[0] } = _1160_ ? 2'h0 : 2'h3;
assign _0113_ = _1173_ ? 2'h2 : { _1046_[1], _0926_[0] };
assign _1047_ = _0403_ ? 7'h00 : 7'h08;
assign { _0927_[6:4], _1048_[3], _0927_[2:1], _1048_[0] } = _1196_ ? 7'h0a : 7'h04;
assign _1050_ = _1194_ ? 7'h09 : { _0927_[6:4], _1048_[3], _0927_[2:1], _1048_[0] };
assign _1052_ = _0902_ ? _1047_ : _1050_;
assign _1054_ = _1199_ ? 7'h03 : 7'h02;
assign { _0929_[6], _1056_[5], _0929_[4], _1056_[3], _0929_[2], _1056_[1:0] } = _1204_ ? 7'h01 : 7'h2c;
assign _1058_ = _1202_ ? 7'h2b : { _0929_[6], _1056_[5], _0929_[4], _1056_[3], _0929_[2], _1056_[1:0] };
assign _1060_ = _0904_ ? _1054_ : _1058_;
assign _0008_ = _0371_ ? _1052_ : _1060_;
assign _1062_ = _1209_ ? _0000_ : 7'h0a;
assign _1064_ = _1213_ ? 7'h04 : 7'h03;
assign _1066_ = _0906_ ? _1062_ : _1064_;
assign _1068_ = _1215_ ? 7'h02 : 7'h2c;
assign _1070_ = _1218_ ? 7'h2b : 7'h00;
assign _1072_ = _0908_ ? _1068_ : _1070_;
assign _0119_ = _0373_ ? _1066_ : _1072_;
assign { _0935_[6:5], _1074_[4:2], _0935_[1:0] } = _1214_ ? 7'h1a : 7'h1b;
assign _1076_ = _1213_ ? 7'h1c : { _0935_[6:5], _1074_[4:2], _0935_[1:0] };
assign _1078_ = _1215_ ? 7'h19 : 7'h1e;
assign _1079_ = _1160_ ? 7'h1d : 7'h2c;
assign _1080_ = _0910_ ? _1078_ : _1079_;
assign _0103_ = _0375_ ? _1076_ : _1080_;
assign _1082_ = _1207_ ? 1'h0 : _0115_;
assign _1084_ = _1221_ ? _0073_ : 1'h1;
assign alu_op_b_mux_sel_o = _0912_ ? _1082_ : _1084_;
assign _1086_ = _1174_ ? _0113_ : 2'h0;
assign _1088_ = _1171_ ? _0123_ : _1086_;
assign { _1090_[1], _0940_[0] } = _0412_ ? _0076_ : 2'h3;
assign _1092_ = _0386_ ? 2'h2 : { _1090_[1], _0940_[0] };
assign alu_op_a_mux_sel_o = _0377_ ? _1088_ : _1092_;
assign _1094_ = _1207_ ? _0004_ : _0119_;
assign _1096_ = _1174_ ? _0012_ : _1094_;
assign _0944_ = _1221_ ? _0108_ : 7'h2c;
assign _1099_ = _0409_ ? 7'h00 : _0944_;
assign alu_operator_o = _0379_ ? _1096_ : _1099_;
assign _1101_ = _0407_ ? 3'h3 : _0118_;
assign _1103_ = _1174_ ? _0121_ : _1101_;
assign _1105_ = _1221_ ? _0106_ : _0091_;
assign _1107_ = _1225_ ? _0059_ : 3'h0;
assign _1109_ = _0914_ ? _1105_ : _1107_;
assign imm_b_mux_sel_o = _0381_ ? _1103_ : _1109_;
assign _1111_ = _1233_ ? 2'h3 : 2'h2;
assign _1113_ = _1236_ ? 2'h1 : 2'h0;
assign _0079_ = _0916_ ? _1111_ : _1113_;
assign _1115_ = _1257_ ? 2'h1 : 2'h0;
assign _0098_ = _0405_ ? 2'h3 : _1115_;
assign _1117_ = _0397_ ? 2'h3 : 2'h2;
assign _1118_ = _0401_ ? 2'h1 : 2'h0;
assign _0096_ = _0918_ ? _1117_ : _1118_;
assign _1119_ = _1244_ ? _0128_ : 1'h0;
assign _0125_ = _1266_ ? _0006_ : _1119_;
assign { _0953_[1], _1121_[0] } = _1278_ ? 2'h2 : 2'h0;
assign _0044_ = _1236_ ? 2'h1 : { _0953_[1], _1121_[0] };
assign _1123_ = _0367_ ? 1'h0 : 1'h1;
assign _0116_ = _1234_ ? _0105_ : _1123_;
assign _1124_ = _1237_ ? _0040_ : 1'h1;
assign _1126_ = _0391_ ? _0073_ : 1'h0;
assign _0028_ = _0920_ ? _1124_ : _1126_;
assign _1128_ = _0391_ ? _0062_ : 1'h0;
assign _0026_ = _1245_ ? _0054_ : _1128_;
assign _1130_ = _0391_ ? 1'h1 : 1'h0;
assign _0024_ = _1245_ ? _0060_ : _1130_;
assign _1131_ = _1237_ ? _0034_ : _0032_;
assign _1133_ = _1268_ ? _0125_ : 1'h0;
assign _1135_ = _1264_ ? _0014_ : _1133_;
assign _1137_ = _0922_ ? _1131_ : _1135_;
assign _1139_ = _1276_ ? _0116_ : _0110_;
assign _1141_ = _1282_ ? _0056_ : 1'h1;
assign _1143_ = _1281_ ? _0089_ : _1141_;
assign _1145_ = _0924_ ? _1139_ : _1143_;
assign _0022_ = _0383_ ? _1137_ : _1145_;
assign _1147_ = _0393_ ? 1'h1 : 1'h0;
assign rf_ren_a_o = _1237_ ? _0071_ : _1147_;
assign _1148_ = csr_op == /* src = "generated/sv2v_out.v:15064.9-15064.23" */ 2'h2;
assign _1150_ = csr_op == /* src = "generated/sv2v_out.v:15064.29-15064.43" */ 2'h3;
assign _1152_ = ! /* src = "generated/sv2v_out.v:15064.50-15064.74" */ instr_rdata_i[19:15];
assign _1155_ = { instr_rdata_i[26], instr_rdata_i[13:12] } == /* src = "generated/sv2v_out.v:15214.9-15214.44" */ 3'h5;
assign _1157_ = ! /* src = "generated/sv2v_out.v:15524.16-15524.44" */ instr_rdata_alu_i[31:27];
assign _1159_ = instr_rdata_alu_i[31:27] == /* src = "generated/sv2v_out.v:15526.16-15526.44" */ 5'h08;
assign _1161_ = _1163_ && /* src = "generated/sv2v_out.v:15064.7-15064.75" */ _1152_;
assign _1163_ = _1148_ || /* src = "generated/sv2v_out.v:15064.8-15064.44" */ _1150_;
assign _1165_ = _1168_ || /* src = "generated/sv2v_out.v:15288.10-15288.59" */ _1169_;
assign _1167_ = | /* src = "generated/sv2v_out.v:15110.9-15110.31" */ instr_rdata_i[14:12];
assign _1168_ = | /* src = "generated/sv2v_out.v:15288.11-15288.32" */ instr_rdata_i[19:15];
assign _1169_ = | /* src = "generated/sv2v_out.v:15288.38-15288.58" */ instr_rdata_i[11:7];
assign _0127_ = instr_rdata_alu_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15762.10-15762.23|generated/sv2v_out.v:15762.6-15765.33" */ 2'h3 : 2'h0;
assign _0123_ = _1160_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15754.9-15754.35|generated/sv2v_out.v:15754.5-15766.8" */ 2'h0 : _0127_;
assign _0057_ = _1160_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15754.9-15754.35|generated/sv2v_out.v:15754.5-15766.8" */ 1'h1 : 1'h0;
assign _0012_ = _0365_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15733.5-15752.12" */ 7'h00 : 7'h2c;
assign _0121_ = _1173_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15733.5-15752.12" */ 3'h5 : 3'h0;
assign _1192_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 10'h105;
assign _1194_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 10'h005;
assign _1196_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 10'h001;
assign _1197_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 10'h007;
assign _1199_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 10'h006;
assign _1200_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 10'h004;
assign _1202_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 10'h002;
assign _1204_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 10'h100;
assign _1205_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] };
assign _0081_ = _0396_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 1'h1 : 1'h0;
assign _1176_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 10'h00f;
assign _1178_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 10'h00e;
assign _1180_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 10'h00d;
assign _1182_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 10'h00c;
assign _0094_ = _0395_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 1'h1 : 1'h0;
assign _1184_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 10'h00b;
assign _1186_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 10'h00a;
assign _1188_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 10'h009;
assign _1190_ = { instr_rdata_alu_i[31:25], instr_rdata_alu_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15575.6-15730.13" */ 10'h008;
assign _0046_ = instr_rdata_alu_i[26] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15535.9-15535.22|generated/sv2v_out.v:15535.5-15730.13" */ 1'h0 : _0081_;
assign _0065_ = instr_rdata_alu_i[26] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15535.9-15535.22|generated/sv2v_out.v:15535.5-15730.13" */ 1'h0 : _0094_;
assign _0004_ = instr_rdata_alu_i[26] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15535.9-15535.22|generated/sv2v_out.v:15535.5-15730.13" */ 7'h2c : _0008_;
assign _0002_ = _1159_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15526.16-15526.44|generated/sv2v_out.v:15526.12-15527.30" */ 7'h08 : 7'h2c;
assign _0000_ = _1157_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15524.16-15524.44|generated/sv2v_out.v:15524.12-15527.30" */ 7'h09 : _0002_;
assign _1216_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15427.5-15530.12" */ 3'h3;
assign _1218_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15427.5-15530.12" */ 3'h2;
assign _0115_ = instr_rdata_alu_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15399.9-15399.23|generated/sv2v_out.v:15399.5-15402.8" */ 1'h0 : 1'h1;
assign _0118_ = instr_rdata_alu_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15399.9-15399.23|generated/sv2v_out.v:15399.5-15402.8" */ 3'h0 : 3'h1;
assign _0073_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15384.9-15384.28|generated/sv2v_out.v:15384.5-15393.8" */ 1'h0 : 1'h1;
assign _0108_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15384.9-15384.28|generated/sv2v_out.v:15384.5-15393.8" */ _0103_ : 7'h00;
assign _0106_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15384.9-15384.28|generated/sv2v_out.v:15384.5-15393.8" */ 3'h0 : _0112_;
assign _1213_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15370.5-15379.12" */ 3'h7;
assign _1214_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15370.5-15379.12" */ 3'h6;
assign _1209_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15370.5-15379.12" */ 3'h5;
assign _1215_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15370.5-15379.12" */ 3'h4;
assign _1173_ = instr_rdata_alu_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15370.5-15379.12" */ 3'h1;
assign _1160_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15370.5-15379.12" */ instr_rdata_alu_i[14:12];
assign _0091_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15356.9-15356.48|generated/sv2v_out.v:15356.5-15367.8" */ 3'h0 : 3'h5;
assign _0076_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15356.9-15356.48|generated/sv2v_out.v:15356.5-15367.8" */ 2'h0 : 2'h2;
assign _0059_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15338.9-15338.48|generated/sv2v_out.v:15338.5-15349.8" */ 3'h4 : 3'h5;
assign _1211_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15332.3-15769.10" */ 7'h13;
assign _1229_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15332.3-15769.10" */ 7'h03;
assign _1174_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15332.3-15769.10" */ 7'h0f;
assign _1227_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15332.3-15769.10" */ 7'h17;
assign _1231_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15332.3-15769.10" */ 7'h37;
assign _1219_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15332.3-15769.10" */ 7'h23;
assign _1221_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15332.3-15769.10" */ 7'h63;
assign _1223_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15332.3-15769.10" */ 7'h67;
assign _1225_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15332.3-15769.10" */ 7'h6f;
assign div_sel_o = _1207_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15332.3-15769.10" */ _0046_ : 1'h0;
assign mult_sel_o = _1207_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15332.3-15769.10" */ _0065_ : 1'h0;
assign _1207_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15332.3-15769.10" */ 7'h33;
assign imm_a_mux_sel_o = _1171_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15332.3-15769.10" */ _0057_ : 1'h1;
assign _1171_ = instr_rdata_alu_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15332.3-15769.10" */ 7'h73;
assign csr_access_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15309.7-15309.19|generated/sv2v_out.v:15309.3-15317.6" */ 1'h0 : rf_wdata_sel_o;
assign branch_in_dec_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15309.7-15309.19|generated/sv2v_out.v:15309.3-15317.6" */ 1'h0 : _0016_;
assign jump_set_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15309.7-15309.19|generated/sv2v_out.v:15309.3-15317.6" */ 1'h0 : _0026_;
assign jump_in_dec_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15309.7-15309.19|generated/sv2v_out.v:15309.3-15317.6" */ 1'h0 : _0024_;
assign data_we_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15309.7-15309.19|generated/sv2v_out.v:15309.3-15317.6" */ 1'h0 : _0020_;
assign data_req_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15309.7-15309.19|generated/sv2v_out.v:15309.3-15317.6" */ 1'h0 : _0018_;
assign rf_we_o = illegal_insn_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15309.7-15309.19|generated/sv2v_out.v:15309.3-15317.6" */ 1'h0 : _0028_;
assign illegal_insn_o = illegal_c_insn_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15307.7-15307.23|generated/sv2v_out.v:15307.3-15308.24" */ 1'h1 : _0022_;
assign _0077_ = _0366_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15297.6-15302.13" */ 1'h0 : 1'h1;
assign _1233_ = instr_rdata_i[13:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15297.6-15302.13" */ 2'h3;
assign _0100_ = instr_rdata_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15295.10-15295.20|generated/sv2v_out.v:15295.6-15296.25" */ 1'h0 : 1'h1;
assign _0038_ = _1165_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15288.10-15288.59|generated/sv2v_out.v:15288.6-15289.27" */ 1'h1 : _0036_;
assign _0087_ = _1239_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15280.6-15287.13" */ 1'h1 : 1'h0;
assign _0036_ = _0329_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15280.6-15287.13" */ 1'h0 : 1'h1;
assign _1239_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15280.6-15287.13" */ instr_rdata_i[31:20];
assign _0101_ = _1240_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15280.6-15287.13" */ 1'h1 : 1'h0;
assign _1240_ = instr_rdata_i[31:20] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15280.6-15287.13" */ 12'h105;
assign _0083_ = _1241_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15280.6-15287.13" */ 1'h1 : 1'h0;
assign _1241_ = instr_rdata_i[31:20] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15280.6-15287.13" */ 12'h7b2;
assign _0092_ = _1242_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15280.6-15287.13" */ 1'h1 : 1'h0;
assign _1242_ = instr_rdata_i[31:20] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15280.6-15287.13" */ 12'h302;
assign _0085_ = _1243_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15280.6-15287.13" */ 1'h1 : 1'h0;
assign _1243_ = instr_rdata_i[31:20] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15280.6-15287.13" */ 12'h001;
assign _0034_ = _0336_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15279.9-15279.31|generated/sv2v_out.v:15279.5-15304.8" */ _0038_ : _0077_;
assign _0074_ = _0336_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15279.9-15279.31|generated/sv2v_out.v:15279.5-15304.8" */ _0101_ : 1'h0;
assign _0052_ = _0336_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15279.9-15279.31|generated/sv2v_out.v:15279.5-15304.8" */ _0087_ : 1'h0;
assign _0048_ = _0336_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15279.9-15279.31|generated/sv2v_out.v:15279.5-15304.8" */ _0083_ : 1'h0;
assign _0063_ = _0336_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15279.9-15279.31|generated/sv2v_out.v:15279.5-15304.8" */ _0092_ : 1'h0;
assign _0050_ = _0336_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15279.9-15279.31|generated/sv2v_out.v:15279.5-15304.8" */ _0085_ : 1'h0;
assign _0071_ = _0336_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15279.9-15279.31|generated/sv2v_out.v:15279.5-15304.8" */ 1'h0 : _0100_;
assign _0040_ = _0336_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15279.9-15279.31|generated/sv2v_out.v:15279.5-15304.8" */ 1'h0 : 1'h1;
assign _0042_ = _0336_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15279.9-15279.31|generated/sv2v_out.v:15279.5-15304.8" */ 2'h0 : _0079_;
assign _0032_ = _0385_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15266.5-15277.12" */ 1'h0 : 1'h1;
assign _0060_ = _1244_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15266.5-15277.12" */ 1'h1 : 1'h0;
assign _0054_ = _1244_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15266.5-15277.12" */ _0062_ : 1'h0;
assign _0030_ = _0332_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 1'h0 : 1'h1;
assign _1260_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h008;
assign _1262_[0] = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ { instr_rdata_i[31:25], instr_rdata_i[14:12] };
assign _1262_[1] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h100;
assign _1262_[2] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h002;
assign _1262_[3] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h003;
assign _1262_[4] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h004;
assign _1262_[5] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h006;
assign _1262_[6] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h007;
assign _1262_[7] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h001;
assign _1262_[8] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h005;
assign _1262_[9] = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h105;
assign _1247_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h00f;
assign _1249_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h00e;
assign _1251_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h00d;
assign _1253_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h00c;
assign _1255_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h00b;
assign _1257_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h00a;
assign _1258_ = { instr_rdata_i[31:25], instr_rdata_i[14:12] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15217.6-15263.13" */ 10'h009;
assign _0014_ = _1155_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15214.9-15214.44|generated/sv2v_out.v:15214.5-15263.13" */ 1'h1 : _0030_;
assign _0069_ = _1155_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15214.9-15214.44|generated/sv2v_out.v:15214.5-15263.13" */ 2'h0 : _0098_;
assign _0067_ = _1155_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15214.9-15214.44|generated/sv2v_out.v:15214.5-15263.13" */ 2'h0 : _0096_;
assign _0010_ = _1272_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15182.8-15206.15" */ _1290_ : 1'h1;
assign _1272_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15182.8-15206.15" */ _1270_;
assign _1270_[1] = instr_rdata_i[31:27] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15182.8-15206.15" */ 5'h08;
assign _0006_ = instr_rdata_i[26] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15179.11-15179.20|generated/sv2v_out.v:15179.7-15206.15" */ 1'h1 : _0010_;
assign _0330_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15171.9-15175.16" */ instr_rdata_i[26:25];
assign _0128_ = _1270_[0] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15161.7-15177.14" */ _1290_ : 1'h1;
assign _1270_[0] = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15161.7-15177.14" */ instr_rdata_i[31:27];
assign _0105_ = instr_rdata_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15147.11-15147.20|generated/sv2v_out.v:15147.7-15148.28" */ 1'h1 : 1'h0;
assign _0110_ = _0369_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15130.5-15135.12" */ _0105_ : 1'h1;
assign _1234_ = instr_rdata_i[13:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15130.5-15135.12" */ 2'h2;
assign _1236_ = instr_rdata_i[13:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15130.5-15135.12" */ 2'h1;
assign _1278_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15130.5-15135.12" */ instr_rdata_i[13:12];
assign _0089_ = _1280_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15116.5-15119.12" */ 1'h0 : 1'h1;
assign _1280_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15116.5-15119.12" */ { _0336_, _1274_[5:3], _1266_, _1244_ };
assign _0336_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15116.5-15119.12" */ instr_rdata_i[14:12];
assign _1244_ = instr_rdata_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15116.5-15119.12" */ 3'h1;
assign _1274_[3] = instr_rdata_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15116.5-15119.12" */ 3'h4;
assign _1266_ = instr_rdata_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15116.5-15119.12" */ 3'h5;
assign _1274_[4] = instr_rdata_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15116.5-15119.12" */ 3'h6;
assign _1274_[5] = instr_rdata_i[14:12] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15116.5-15119.12" */ 3'h7;
assign _0056_ = _1167_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15110.9-15110.31|generated/sv2v_out.v:15110.5-15111.26" */ 1'h1 : 1'h0;
assign _0062_ = instr_first_cycle_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15104.9-15104.28|generated/sv2v_out.v:15104.5-15109.19" */ 1'h1 : 1'h0;
assign _1286_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ 7'h17;
assign _1288_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ 7'h37;
assign _1284_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ 7'h6f;
assign _0016_ = _1281_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ 1'h1 : 1'h0;
assign data_sign_extension_o = _1276_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ _0320_ : 1'h0;
assign data_type_o = _0411_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ _0044_ : 2'h0;
assign multdiv_signed_mode_o = _1264_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ _0069_ : 2'h0;
assign multdiv_operator_o = _1264_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ _0067_ : 2'h0;
assign rf_wdata_sel_o = _1237_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ _0040_ : 1'h0;
assign wfi_insn_o = _1237_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ _0074_ : 1'h0;
assign ecall_insn_o = _1237_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ _0052_ : 1'h0;
assign dret_insn_o = _1237_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ _0048_ : 1'h0;
assign mret_insn_o = _1237_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ _0063_ : 1'h0;
assign ebrk_insn_o = _1237_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ _0050_ : 1'h0;
assign rf_ren_b_o = _0388_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ 1'h1 : 1'h0;
assign _1264_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ 7'h33;
assign _1268_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ 7'h13;
assign _1276_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ 7'h03;
assign _1279_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ 7'h23;
assign _1281_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ 7'h63;
assign _1282_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ 7'h67;
assign icache_inval_o = _1245_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ _0054_ : 1'h0;
assign _1245_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ 7'h0f;
assign csr_op = _1237_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ _0042_ : 2'h0;
assign _1237_ = instr_rdata_i[6:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ 7'h73;
assign _0020_ = _1279_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ 1'h1 : 1'h0;
assign _0018_ = _0411_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:15092.3-15306.10" */ 1'h1 : 1'h0;
assign csr_op_o = _1161_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:15064.7-15064.75|generated/sv2v_out.v:15064.3-15065.20" */ 2'h0 : csr_op;
assign _1290_ = _0330_ ? /* src = "generated/sv2v_out.v:15183.45-15183.80" */ 1'h0 : 1'h1;
assign _0112_ = branch_taken_i ? /* src = "generated/sv2v_out.v:15391.25-15391.53" */ 3'h2 : 3'h5;
assign mult_en_o = illegal_insn_o ? /* src = "generated/sv2v_out.v:15771.22-15771.54" */ 1'h0 : mult_sel_o;
assign div_en_o = illegal_insn_o ? /* src = "generated/sv2v_out.v:15772.21-15772.52" */ 1'h0 : div_sel_o;
assign { _0003_[6], _0003_[4:0] } = { 3'h0, _0003_[5], 2'h0 };
assign { _0013_[6], _0013_[4:0] } = { 2'h0, _0013_[5], _0013_[5], 2'h0 };
assign _0122_[1:0] = { 1'h0, _0122_[2] };
assign _0926_[1] = _0342_;
assign { _0927_[3], _0927_[0] } = _0347_;
assign { _0929_[5], _0929_[3], _0929_[1:0] } = _0341_;
assign _0935_[4:2] = _0345_;
assign _0940_[1] = _0344_;
assign _0953_[0] = _0349_;
assign _1046_[0] = _0926_[0];
assign { _1048_[6:4], _1048_[2:1] } = { _0927_[6:4], _0927_[2:1] };
assign { _1049_[6:4], _1049_[2:0] } = { 3'h0, _1049_[3], _1049_[3], 1'h0 };
assign _1055_[6:1] = 6'h00;
assign { _1056_[6], _1056_[4], _1056_[2] } = { _0929_[6], _0929_[4], _0929_[2] };
assign { _1057_[6], _1057_[4:0] } = { 2'h0, _1057_[5], _1057_[5], 1'h0, _1057_[5] };
assign { _1065_[6:3], _1065_[1:0] } = { 4'h0, _1065_[2], _1065_[2] };
assign { _1069_[6], _1069_[4:0] } = { 2'h0, _1069_[5], _1069_[5], _1069_[5], 1'h0 };
assign { _1071_[6], _1071_[4:0] } = { 2'h0, _1071_[5], 1'h0, _1071_[5], _1071_[5] };
assign { _1074_[6:5], _1074_[1:0] } = { _0935_[6:5], _0935_[1:0] };
assign _1075_[6:1] = 6'h00;
assign _1090_[0] = _0940_[0];
assign _1112_[1] = 1'h0;
assign _1114_[1] = 1'h0;
assign _1116_[1] = 1'h0;
assign _1121_[1] = _0953_[1];
assign _1122_[0] = 1'h0;
assign _1274_[0] = _0336_;
assign _1275_[0] = _0041_;
assign alu_multicycle_o = 1'h0;
assign alu_multicycle_o_t0 = 1'h0;
assign bt_a_mux_sel_o = 2'h2;
assign bt_a_mux_sel_o_t0 = 2'h0;
assign bt_b_mux_sel_o = 3'h0;
assign bt_b_mux_sel_o_t0 = 3'h0;
assign imm_b_type_o = { instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[7], instr_rdata_i[30:25], instr_rdata_i[11:8], 1'h0 };
assign imm_b_type_o_t0 = { instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[7], instr_rdata_i_t0[30:25], instr_rdata_i_t0[11:8], 1'h0 };
assign imm_i_type_o = { instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31:20] };
assign imm_i_type_o_t0 = { instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31:20] };
assign imm_j_type_o = { instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[19:12], instr_rdata_i[20], instr_rdata_i[30:21], 1'h0 };
assign imm_j_type_o_t0 = { instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[19:12], instr_rdata_i_t0[20], instr_rdata_i_t0[30:21], 1'h0 };
assign imm_s_type_o = { instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31], instr_rdata_i[31:25], instr_rdata_i[11:7] };
assign imm_s_type_o_t0 = { instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31], instr_rdata_i_t0[31:25], instr_rdata_i_t0[11:7] };
assign imm_u_type_o = { instr_rdata_i[31:12], 12'h000 };
assign imm_u_type_o_t0 = { instr_rdata_i_t0[31:12], 12'h000 };
assign rf_raddr_a_o = instr_rdata_i[19:15];
assign rf_raddr_a_o_t0 = instr_rdata_i_t0[19:15];
assign rf_raddr_b_o = instr_rdata_i[24:20];
assign rf_raddr_b_o_t0 = instr_rdata_i_t0[24:20];
assign rf_waddr_o = instr_rdata_i[11:7];
assign rf_waddr_o_t0 = instr_rdata_i_t0[11:7];
assign zimm_rs1_type_o = { 27'h0000000, instr_rdata_i[19:15] };
assign zimm_rs1_type_o_t0 = { 27'h0000000, instr_rdata_i_t0[19:15] };
endmodule

module \$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _00_;
wire [31:0] _01_;
wire [31:0] _02_;
wire [31:0] _03_;
wire [31:0] _04_;
wire [31:0] _05_;
wire [31:0] _06_;
wire [31:0] _07_;
wire [31:0] _08_;
/* src = "generated/sv2v_out.v:14871.13-14871.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14875.28-14875.37" */
output [31:0] rd_data_o;
reg [31:0] rd_data_o;
/* cellift = 32'd1 */
output [31:0] rd_data_o_t0;
reg [31:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14876.14-14876.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14872.13-14872.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14873.27-14873.36" */
input [31:0] wr_data_i;
wire [31:0] wr_data_i;
/* cellift = 32'd1 */
input [31:0] wr_data_i_t0;
wire [31:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14874.13-14874.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _00_ = ~ wr_en_i;
assign _08_ = wr_data_i ^ rd_data_o;
assign _04_ = wr_data_i_t0 | rd_data_o_t0;
assign _05_ = _08_ | _04_;
assign _01_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _02_ = { _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_ } & rd_data_o_t0;
assign _03_ = _05_ & { wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0 };
assign _06_ = _01_ | _02_;
assign _07_ = _06_ | _03_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 32'd0;
else rd_data_o_t0 <= _07_;
/* src = "generated/sv2v_out.v:14878.2-14882.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 32'd0;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage (clk_i, rst_ni, boot_addr_i, req_i, instr_req_o, instr_addr_o, instr_gnt_i, instr_rvalid_i, instr_rdata_i, instr_bus_err_i, instr_intg_err_o, ic_tag_req_o, ic_tag_write_o, ic_tag_addr_o, ic_tag_wdata_o, ic_tag_rdata_i, ic_data_req_o, ic_data_write_o, ic_data_addr_o, ic_data_wdata_o, ic_data_rdata_i
, ic_scr_key_valid_i, ic_scr_key_req_o, instr_valid_id_o, instr_new_id_o, instr_rdata_id_o, instr_rdata_alu_id_o, instr_rdata_c_id_o, instr_is_compressed_id_o, instr_bp_taken_o, instr_fetch_err_o, instr_fetch_err_plus2_o, illegal_c_insn_id_o, dummy_instr_id_o, pc_if_o, pc_id_o, pmp_err_if_i, pmp_err_if_plus2_i, instr_valid_clear_i, pc_set_i, pc_mux_i, nt_branch_mispredict_i
, nt_branch_addr_i, exc_pc_mux_i, exc_cause, dummy_instr_en_i, dummy_instr_mask_i, dummy_instr_seed_en_i, dummy_instr_seed_i, icache_enable_i, icache_inval_i, icache_ecc_error_o, branch_target_ex_i, csr_mepc_i, csr_depc_i, csr_mtvec_i, csr_mtvec_init_o, id_in_ready_i, pc_mismatch_alert_o, if_busy_o, pmp_err_if_plus2_i_t0, pmp_err_if_i_t0, pc_set_i_t0
, pc_mux_i_t0, pc_mismatch_alert_o_t0, pc_if_o_t0, pc_id_o_t0, nt_branch_mispredict_i_t0, nt_branch_addr_i_t0, instr_valid_id_o_t0, instr_valid_clear_i_t0, instr_rdata_id_o_t0, instr_rdata_c_id_o_t0, instr_rdata_alu_id_o_t0, instr_new_id_o_t0, instr_is_compressed_id_o_t0, instr_intg_err_o_t0, instr_fetch_err_plus2_o_t0, instr_fetch_err_o_t0, instr_bus_err_i_t0, instr_bp_taken_o_t0, illegal_c_insn_id_o_t0, if_busy_o_t0, icache_inval_i_t0
, icache_enable_i_t0, icache_ecc_error_o_t0, ic_tag_write_o_t0, ic_tag_wdata_o_t0, ic_tag_req_o_t0, ic_tag_rdata_i_t0, ic_tag_addr_o_t0, ic_scr_key_valid_i_t0, ic_scr_key_req_o_t0, ic_data_write_o_t0, ic_data_wdata_o_t0, ic_data_req_o_t0, ic_data_rdata_i_t0, ic_data_addr_o_t0, exc_pc_mux_i_t0, exc_cause_t0, dummy_instr_id_o_t0, csr_mtvec_init_o_t0, csr_mtvec_i_t0, csr_mepc_i_t0, csr_depc_i_t0
, branch_target_ex_i_t0, boot_addr_i_t0, id_in_ready_i_t0, dummy_instr_seed_i_t0, dummy_instr_seed_en_i_t0, dummy_instr_mask_i_t0, dummy_instr_en_i_t0, req_i_t0, instr_rvalid_i_t0, instr_req_o_t0, instr_rdata_i_t0, instr_gnt_i_t0, instr_addr_o_t0);
/* src = "generated/sv2v_out.v:18096.45-18096.84" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18096.45-18096.84" */
wire _001_;
/* src = "generated/sv2v_out.v:18096.44-18096.106" */
wire _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18096.44-18096.106" */
wire _003_;
/* src = "generated/sv2v_out.v:18102.12-18102.36" */
wire _004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18102.12-18102.36" */
wire _005_;
/* src = "generated/sv2v_out.v:18157.29-18157.73" */
wire _006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18157.29-18157.73" */
wire _007_;
/* src = "generated/sv2v_out.v:18157.78-18157.117" */
wire _008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18157.78-18157.117" */
wire _009_;
/* src = "generated/sv2v_out.v:18213.32-18213.81" */
wire _010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18213.32-18213.81" */
wire _011_;
/* src = "generated/sv2v_out.v:18213.31-18213.98" */
wire _012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18213.31-18213.98" */
wire _013_;
wire [31:0] _014_;
wire [31:0] _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire [31:0] _020_;
wire [2:0] _021_;
wire [1:0] _022_;
wire _023_;
wire [1:0] _024_;
wire _025_;
wire _026_;
wire [31:0] _027_;
wire [31:0] _028_;
wire [31:0] _029_;
wire [31:0] _030_;
wire [31:0] _031_;
wire [31:0] _032_;
wire [4:0] _033_;
wire [31:0] _034_;
wire [31:0] _035_;
wire _036_;
wire [4:0] _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire [31:0] _054_;
wire [31:0] _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire [31:0] _104_;
wire [31:0] _105_;
wire [31:0] _106_;
wire [31:0] _107_;
wire [31:0] _108_;
wire [31:0] _109_;
wire [15:0] _110_;
wire [15:0] _111_;
wire [15:0] _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire [31:0] _131_;
wire [31:0] _132_;
wire [31:0] _133_;
wire [31:0] _134_;
wire [31:0] _135_;
wire [31:0] _136_;
wire [31:0] _137_;
wire [31:0] _138_;
wire [31:0] _139_;
wire [31:0] _140_;
wire [31:0] _141_;
wire [31:0] _142_;
wire [31:0] _143_;
wire [31:0] _144_;
wire [31:0] _145_;
wire [31:0] _146_;
wire [31:0] _147_;
wire [31:0] _148_;
wire [2:0] _149_;
wire [31:0] _150_;
wire [31:0] _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire [1:0] _173_;
wire [4:0] _174_;
wire [4:0] _175_;
wire [1:0] _176_;
wire [31:0] _177_;
wire [31:0] _178_;
wire [31:0] _179_;
wire [31:0] _180_;
wire [31:0] _181_;
wire [31:0] _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire [31:0] _189_;
wire [31:0] _190_;
wire [31:0] _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire _206_;
wire _207_;
wire _208_;
wire _209_;
wire _210_;
wire [31:0] _211_;
wire [31:0] _212_;
wire [31:0] _213_;
wire [31:0] _214_;
wire [31:0] _215_;
wire [31:0] _216_;
wire [31:0] _217_;
wire [31:0] _218_;
wire [15:0] _219_;
wire [15:0] _220_;
wire [15:0] _221_;
wire [15:0] _222_;
wire _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire _230_;
wire _231_;
wire _232_;
wire _233_;
wire _234_;
wire _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire [31:0] _241_;
wire [31:0] _242_;
wire [31:0] _243_;
wire [31:0] _244_;
wire [31:0] _245_;
wire [31:0] _246_;
wire [31:0] _247_;
wire [31:0] _248_;
wire [31:0] _249_;
wire [31:0] _250_;
wire [31:0] _251_;
wire [31:0] _252_;
wire [31:0] _253_;
wire [31:0] _254_;
wire [31:0] _255_;
wire [31:0] _256_;
wire [31:0] _257_;
wire [31:0] _258_;
wire [31:0] _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire [4:0] _267_;
wire [31:0] _268_;
wire [31:0] _269_;
wire [31:0] _270_;
wire [31:0] _271_;
wire [31:0] _272_;
wire [31:0] _273_;
wire _274_;
wire _275_;
/* cellift = 32'd1 */
wire _276_;
wire _277_;
/* cellift = 32'd1 */
wire _278_;
wire [31:0] _279_;
wire _280_;
wire [31:0] _281_;
wire [31:0] _282_;
wire [15:0] _283_;
wire _284_;
wire _285_;
wire _286_;
wire _287_;
wire [31:0] _288_;
wire [31:0] _289_;
wire [31:0] _290_;
wire [31:0] _291_;
wire [31:0] _292_;
wire [31:0] _293_;
wire [31:0] _294_;
wire [31:0] _295_;
wire _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire [31:0] _304_;
wire [31:0] _305_;
wire [31:0] _306_;
/* cellift = 32'd1 */
wire [31:0] _307_;
wire [31:0] _308_;
/* cellift = 32'd1 */
wire [31:0] _309_;
wire [31:0] _310_;
/* cellift = 32'd1 */
wire [31:0] _311_;
wire [31:0] _312_;
/* cellift = 32'd1 */
wire [31:0] _313_;
wire [31:0] _314_;
/* cellift = 32'd1 */
wire [31:0] _315_;
/* src = "generated/sv2v_out.v:17981.29-17981.45" */
wire _316_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17981.29-17981.45" */
wire _317_;
/* src = "generated/sv2v_out.v:18224.53-18224.88" */
wire _318_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18224.53-18224.88" */
wire _319_;
/* src = "generated/sv2v_out.v:18096.64-18096.84" */
wire _320_;
/* src = "generated/sv2v_out.v:18157.97-18157.117" */
wire _321_;
/* src = "generated/sv2v_out.v:18213.85-18213.98" */
wire _322_;
/* src = "generated/sv2v_out.v:18098.31-18098.113" */
wire _323_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18098.31-18098.113" */
wire _324_;
/* src = "generated/sv2v_out.v:18213.33-18213.66" */
wire _325_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18213.33-18213.66" */
wire _326_;
wire _327_;
/* cellift = 32'd1 */
wire _328_;
wire _329_;
/* cellift = 32'd1 */
wire _330_;
wire _331_;
/* cellift = 32'd1 */
wire _332_;
wire _333_;
/* cellift = 32'd1 */
wire _334_;
wire _335_;
wire _336_;
/* cellift = 32'd1 */
wire _337_;
wire _338_;
/* cellift = 32'd1 */
wire _339_;
/* src = "generated/sv2v_out.v:18219.45-18219.85" */
wire [31:0] _340_;
/* src = "generated/sv2v_out.v:17852.20-17852.31" */
input [31:0] boot_addr_i;
wire [31:0] boot_addr_i;
/* cellift = 32'd1 */
input [31:0] boot_addr_i_t0;
wire [31:0] boot_addr_i_t0;
/* src = "generated/sv2v_out.v:17902.20-17902.38" */
input [31:0] branch_target_ex_i;
wire [31:0] branch_target_ex_i;
/* cellift = 32'd1 */
input [31:0] branch_target_ex_i_t0;
wire [31:0] branch_target_ex_i_t0;
/* src = "generated/sv2v_out.v:17850.13-17850.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:17904.20-17904.30" */
input [31:0] csr_depc_i;
wire [31:0] csr_depc_i;
/* cellift = 32'd1 */
input [31:0] csr_depc_i_t0;
wire [31:0] csr_depc_i_t0;
/* src = "generated/sv2v_out.v:17903.20-17903.30" */
input [31:0] csr_mepc_i;
wire [31:0] csr_mepc_i;
/* cellift = 32'd1 */
input [31:0] csr_mepc_i_t0;
wire [31:0] csr_mepc_i_t0;
/* src = "generated/sv2v_out.v:17905.20-17905.31" */
input [31:0] csr_mtvec_i;
wire [31:0] csr_mtvec_i;
/* cellift = 32'd1 */
input [31:0] csr_mtvec_i_t0;
wire [31:0] csr_mtvec_i_t0;
/* src = "generated/sv2v_out.v:17906.14-17906.30" */
output csr_mtvec_init_o;
wire csr_mtvec_init_o;
/* cellift = 32'd1 */
output csr_mtvec_init_o_t0;
wire csr_mtvec_init_o_t0;
/* src = "generated/sv2v_out.v:17895.13-17895.29" */
input dummy_instr_en_i;
wire dummy_instr_en_i;
/* cellift = 32'd1 */
input dummy_instr_en_i_t0;
wire dummy_instr_en_i_t0;
/* src = "generated/sv2v_out.v:17883.13-17883.29" */
output dummy_instr_id_o;
reg dummy_instr_id_o;
/* cellift = 32'd1 */
output dummy_instr_id_o_t0;
reg dummy_instr_id_o_t0;
/* src = "generated/sv2v_out.v:17896.19-17896.37" */
input [2:0] dummy_instr_mask_i;
wire [2:0] dummy_instr_mask_i;
/* cellift = 32'd1 */
input [2:0] dummy_instr_mask_i_t0;
wire [2:0] dummy_instr_mask_i_t0;
/* src = "generated/sv2v_out.v:17897.13-17897.34" */
input dummy_instr_seed_en_i;
wire dummy_instr_seed_en_i;
/* cellift = 32'd1 */
input dummy_instr_seed_en_i_t0;
wire dummy_instr_seed_en_i_t0;
/* src = "generated/sv2v_out.v:17898.20-17898.38" */
input [31:0] dummy_instr_seed_i;
wire [31:0] dummy_instr_seed_i;
/* cellift = 32'd1 */
input [31:0] dummy_instr_seed_i_t0;
wire [31:0] dummy_instr_seed_i_t0;
/* src = "generated/sv2v_out.v:17894.19-17894.28" */
input [6:0] exc_cause;
wire [6:0] exc_cause;
/* cellift = 32'd1 */
input [6:0] exc_cause_t0;
wire [6:0] exc_cause_t0;
/* src = "generated/sv2v_out.v:17939.13-17939.19" */
wire [31:0] exc_pc;
/* src = "generated/sv2v_out.v:17893.19-17893.31" */
input [1:0] exc_pc_mux_i;
wire [1:0] exc_pc_mux_i;
/* cellift = 32'd1 */
input [1:0] exc_pc_mux_i_t0;
wire [1:0] exc_pc_mux_i_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17939.13-17939.19" */
wire [31:0] exc_pc_t0;
/* src = "generated/sv2v_out.v:17918.13-17918.25" */
/* unused_bits = "0" */
wire [31:0] fetch_addr_n;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17918.13-17918.25" */
/* unused_bits = "0" */
wire [31:0] fetch_addr_n_t0;
/* src = "generated/sv2v_out.v:17927.7-17927.16" */
wire fetch_err;
/* src = "generated/sv2v_out.v:17928.7-17928.22" */
wire fetch_err_plus2;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17928.7-17928.22" */
wire fetch_err_plus2_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17927.7-17927.16" */
wire fetch_err_t0;
/* src = "generated/sv2v_out.v:17925.14-17925.25" */
wire [31:0] fetch_rdata;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17925.14-17925.25" */
wire [31:0] fetch_rdata_t0;
/* src = "generated/sv2v_out.v:17924.7-17924.18" */
wire fetch_ready;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17924.7-17924.18" */
wire fetch_ready_t0;
/* src = "generated/sv2v_out.v:17923.7-17923.18" */
wire fetch_valid;
/* src = "generated/sv2v_out.v:17922.7-17922.22" */
wire fetch_valid_raw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17922.7-17922.22" */
wire fetch_valid_raw_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17923.7-17923.18" */
wire fetch_valid_t0;
/* src = "generated/sv2v_out.v:17984.15-17984.22" */
wire [1:0] \g_mem_ecc.ecc_err ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17984.15-17984.22" */
wire [1:0] \g_mem_ecc.ecc_err_t0 ;
/* src = "generated/sv2v_out.v:17985.30-17985.45" */
wire [38:0] \g_mem_ecc.instr_rdata_buf ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17985.30-17985.45" */
wire [38:0] \g_mem_ecc.instr_rdata_buf_t0 ;
/* src = "generated/sv2v_out.v:18209.16-18209.36" */
wire [31:0] \g_secure_pc.prev_instr_addr_incr ;
/* src = "generated/sv2v_out.v:18210.16-18210.40" */
wire [31:0] \g_secure_pc.prev_instr_addr_incr_buf ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18210.16-18210.40" */
wire [31:0] \g_secure_pc.prev_instr_addr_incr_buf_t0 ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18209.16-18209.36" */
wire [31:0] \g_secure_pc.prev_instr_addr_incr_t0 ;
/* src = "generated/sv2v_out.v:18212.9-18212.25" */
wire \g_secure_pc.prev_instr_seq_d ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18212.9-18212.25" */
wire \g_secure_pc.prev_instr_seq_d_t0 ;
/* src = "generated/sv2v_out.v:18211.8-18211.24" */
reg \g_secure_pc.prev_instr_seq_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18211.8-18211.24" */
reg \g_secure_pc.prev_instr_seq_q_t0 ;
/* src = "generated/sv2v_out.v:18111.16-18111.32" */
wire [31:0] \gen_dummy_instr.dummy_instr_data ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18111.16-18111.32" */
wire [31:0] \gen_dummy_instr.dummy_instr_data_t0 ;
/* src = "generated/sv2v_out.v:18110.9-18110.27" */
wire \gen_dummy_instr.insert_dummy_instr ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18110.9-18110.27" */
wire \gen_dummy_instr.insert_dummy_instr_t0 ;
/* src = "generated/sv2v_out.v:17868.42-17868.56" */
output [7:0] ic_data_addr_o;
wire [7:0] ic_data_addr_o;
/* cellift = 32'd1 */
output [7:0] ic_data_addr_o_t0;
wire [7:0] ic_data_addr_o_t0;
/* src = "generated/sv2v_out.v:17870.58-17870.73" */
input [127:0] ic_data_rdata_i;
wire [127:0] ic_data_rdata_i;
/* cellift = 32'd1 */
input [127:0] ic_data_rdata_i_t0;
wire [127:0] ic_data_rdata_i_t0;
/* src = "generated/sv2v_out.v:17866.20-17866.33" */
output [1:0] ic_data_req_o;
wire [1:0] ic_data_req_o;
/* cellift = 32'd1 */
output [1:0] ic_data_req_o_t0;
wire [1:0] ic_data_req_o_t0;
/* src = "generated/sv2v_out.v:17869.34-17869.49" */
output [63:0] ic_data_wdata_o;
wire [63:0] ic_data_wdata_o;
/* cellift = 32'd1 */
output [63:0] ic_data_wdata_o_t0;
wire [63:0] ic_data_wdata_o_t0;
/* src = "generated/sv2v_out.v:17867.14-17867.29" */
output ic_data_write_o;
wire ic_data_write_o;
/* cellift = 32'd1 */
output ic_data_write_o_t0;
wire ic_data_write_o_t0;
/* src = "generated/sv2v_out.v:17872.14-17872.30" */
output ic_scr_key_req_o;
wire ic_scr_key_req_o;
/* cellift = 32'd1 */
output ic_scr_key_req_o_t0;
wire ic_scr_key_req_o_t0;
/* src = "generated/sv2v_out.v:17871.13-17871.31" */
input ic_scr_key_valid_i;
wire ic_scr_key_valid_i;
/* cellift = 32'd1 */
input ic_scr_key_valid_i_t0;
wire ic_scr_key_valid_i_t0;
/* src = "generated/sv2v_out.v:17863.42-17863.55" */
output [7:0] ic_tag_addr_o;
wire [7:0] ic_tag_addr_o;
/* cellift = 32'd1 */
output [7:0] ic_tag_addr_o_t0;
wire [7:0] ic_tag_addr_o_t0;
/* src = "generated/sv2v_out.v:17865.57-17865.71" */
input [43:0] ic_tag_rdata_i;
wire [43:0] ic_tag_rdata_i;
/* cellift = 32'd1 */
input [43:0] ic_tag_rdata_i_t0;
wire [43:0] ic_tag_rdata_i_t0;
/* src = "generated/sv2v_out.v:17861.20-17861.32" */
output [1:0] ic_tag_req_o;
wire [1:0] ic_tag_req_o;
/* cellift = 32'd1 */
output [1:0] ic_tag_req_o_t0;
wire [1:0] ic_tag_req_o_t0;
/* src = "generated/sv2v_out.v:17864.33-17864.47" */
output [21:0] ic_tag_wdata_o;
wire [21:0] ic_tag_wdata_o;
/* cellift = 32'd1 */
output [21:0] ic_tag_wdata_o_t0;
wire [21:0] ic_tag_wdata_o_t0;
/* src = "generated/sv2v_out.v:17862.14-17862.28" */
output ic_tag_write_o;
wire ic_tag_write_o;
/* cellift = 32'd1 */
output ic_tag_write_o_t0;
wire ic_tag_write_o_t0;
/* src = "generated/sv2v_out.v:17901.14-17901.32" */
output icache_ecc_error_o;
wire icache_ecc_error_o;
/* cellift = 32'd1 */
output icache_ecc_error_o_t0;
wire icache_ecc_error_o_t0;
/* src = "generated/sv2v_out.v:17899.13-17899.28" */
input icache_enable_i;
wire icache_enable_i;
/* cellift = 32'd1 */
input icache_enable_i_t0;
wire icache_enable_i_t0;
/* src = "generated/sv2v_out.v:17900.13-17900.27" */
input icache_inval_i;
wire icache_inval_i;
/* cellift = 32'd1 */
input icache_inval_i_t0;
wire icache_inval_i_t0;
/* src = "generated/sv2v_out.v:17907.13-17907.26" */
input id_in_ready_i;
wire id_in_ready_i;
/* cellift = 32'd1 */
input id_in_ready_i_t0;
wire id_in_ready_i_t0;
/* src = "generated/sv2v_out.v:17909.14-17909.23" */
output if_busy_o;
wire if_busy_o;
/* cellift = 32'd1 */
output if_busy_o_t0;
wire if_busy_o_t0;
/* src = "generated/sv2v_out.v:17940.7-17940.24" */
wire if_id_pipe_reg_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17940.7-17940.24" */
wire if_id_pipe_reg_we_t0;
/* src = "generated/sv2v_out.v:17937.7-17937.19" */
wire if_instr_err;
/* src = "generated/sv2v_out.v:17938.7-17938.25" */
wire if_instr_err_plus2;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17938.7-17938.25" */
wire if_instr_err_plus2_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17937.7-17937.19" */
wire if_instr_err_t0;
/* src = "generated/sv2v_out.v:17936.7-17936.23" */
wire if_instr_pmp_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17936.7-17936.23" */
wire if_instr_pmp_err_t0;
/* src = "generated/sv2v_out.v:17930.7-17930.21" */
wire illegal_c_insn;
/* src = "generated/sv2v_out.v:17882.13-17882.32" */
output illegal_c_insn_id_o;
reg illegal_c_insn_id_o;
/* cellift = 32'd1 */
output illegal_c_insn_id_o_t0;
reg illegal_c_insn_id_o_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17930.7-17930.21" */
wire illegal_c_insn_t0;
/* src = "generated/sv2v_out.v:17944.7-17944.26" */
wire illegal_c_instr_out;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17944.7-17944.26" */
wire illegal_c_instr_out_t0;
/* src = "generated/sv2v_out.v:17855.21-17855.33" */
output [31:0] instr_addr_o;
wire [31:0] instr_addr_o;
/* cellift = 32'd1 */
output [31:0] instr_addr_o_t0;
wire [31:0] instr_addr_o_t0;
/* src = "generated/sv2v_out.v:17879.14-17879.30" */
output instr_bp_taken_o;
wire instr_bp_taken_o;
/* cellift = 32'd1 */
output instr_bp_taken_o_t0;
wire instr_bp_taken_o_t0;
/* src = "generated/sv2v_out.v:17859.13-17859.28" */
input instr_bus_err_i;
wire instr_bus_err_i;
/* cellift = 32'd1 */
input instr_bus_err_i_t0;
wire instr_bus_err_i_t0;
/* src = "generated/sv2v_out.v:17929.14-17929.32" */
wire [31:0] instr_decompressed;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17929.14-17929.32" */
wire [31:0] instr_decompressed_t0;
/* src = "generated/sv2v_out.v:17914.7-17914.16" */
wire instr_err;
/* src = "generated/sv2v_out.v:17945.7-17945.20" */
wire instr_err_out;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17945.7-17945.20" */
wire instr_err_out_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17914.7-17914.16" */
wire instr_err_t0;
/* src = "generated/sv2v_out.v:17880.13-17880.30" */
output instr_fetch_err_o;
reg instr_fetch_err_o;
/* cellift = 32'd1 */
output instr_fetch_err_o_t0;
reg instr_fetch_err_o_t0;
/* src = "generated/sv2v_out.v:17881.13-17881.36" */
output instr_fetch_err_plus2_o;
reg instr_fetch_err_plus2_o;
/* cellift = 32'd1 */
output instr_fetch_err_plus2_o_t0;
reg instr_fetch_err_plus2_o_t0;
/* src = "generated/sv2v_out.v:17856.13-17856.24" */
input instr_gnt_i;
wire instr_gnt_i;
/* cellift = 32'd1 */
input instr_gnt_i_t0;
wire instr_gnt_i_t0;
/* src = "generated/sv2v_out.v:17915.7-17915.21" */
wire instr_intg_err;
/* src = "generated/sv2v_out.v:17860.14-17860.30" */
output instr_intg_err_o;
wire instr_intg_err_o;
/* cellift = 32'd1 */
output instr_intg_err_o_t0;
wire instr_intg_err_o_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17915.7-17915.21" */
wire instr_intg_err_t0;
/* src = "generated/sv2v_out.v:17931.7-17931.26" */
wire instr_is_compressed;
/* src = "generated/sv2v_out.v:17878.13-17878.37" */
output instr_is_compressed_id_o;
reg instr_is_compressed_id_o;
/* cellift = 32'd1 */
output instr_is_compressed_id_o_t0;
reg instr_is_compressed_id_o_t0;
/* src = "generated/sv2v_out.v:17943.7-17943.30" */
wire instr_is_compressed_out;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17943.7-17943.30" */
wire instr_is_compressed_out_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17931.7-17931.26" */
wire instr_is_compressed_t0;
/* src = "generated/sv2v_out.v:17874.14-17874.28" */
output instr_new_id_o;
reg instr_new_id_o;
/* cellift = 32'd1 */
output instr_new_id_o_t0;
reg instr_new_id_o_t0;
/* src = "generated/sv2v_out.v:17942.14-17942.23" */
wire [31:0] instr_out;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17942.14-17942.23" */
wire [31:0] instr_out_t0;
/* src = "generated/sv2v_out.v:17876.20-17876.40" */
output [31:0] instr_rdata_alu_id_o;
reg [31:0] instr_rdata_alu_id_o;
/* cellift = 32'd1 */
output [31:0] instr_rdata_alu_id_o_t0;
reg [31:0] instr_rdata_alu_id_o_t0;
/* src = "generated/sv2v_out.v:17877.20-17877.38" */
output [15:0] instr_rdata_c_id_o;
reg [15:0] instr_rdata_c_id_o;
/* cellift = 32'd1 */
output [15:0] instr_rdata_c_id_o_t0;
reg [15:0] instr_rdata_c_id_o_t0;
/* src = "generated/sv2v_out.v:17858.34-17858.47" */
input [38:0] instr_rdata_i;
wire [38:0] instr_rdata_i;
/* cellift = 32'd1 */
input [38:0] instr_rdata_i_t0;
wire [38:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:17875.20-17875.36" */
output [31:0] instr_rdata_id_o;
wire [31:0] instr_rdata_id_o;
/* cellift = 32'd1 */
output [31:0] instr_rdata_id_o_t0;
wire [31:0] instr_rdata_id_o_t0;
/* src = "generated/sv2v_out.v:17854.14-17854.25" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:17857.13-17857.27" */
input instr_rvalid_i;
wire instr_rvalid_i;
/* cellift = 32'd1 */
input instr_rvalid_i_t0;
wire instr_rvalid_i_t0;
/* src = "generated/sv2v_out.v:17888.13-17888.32" */
input instr_valid_clear_i;
wire instr_valid_clear_i;
/* cellift = 32'd1 */
input instr_valid_clear_i_t0;
wire instr_valid_clear_i_t0;
/* src = "generated/sv2v_out.v:17910.7-17910.23" */
wire instr_valid_id_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17910.7-17910.23" */
wire instr_valid_id_d_t0;
/* src = "generated/sv2v_out.v:17873.14-17873.30" */
output instr_valid_id_o;
reg instr_valid_id_o;
/* cellift = 32'd1 */
output instr_valid_id_o_t0;
reg instr_valid_id_o_t0;
/* src = "generated/sv2v_out.v:17948.12-17948.19" */
wire [4:0] irq_vec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17948.12-17948.19" */
wire [4:0] irq_vec_t0;
/* src = "generated/sv2v_out.v:17892.20-17892.36" */
input [31:0] nt_branch_addr_i;
wire [31:0] nt_branch_addr_i;
/* cellift = 32'd1 */
input [31:0] nt_branch_addr_i_t0;
wire [31:0] nt_branch_addr_i_t0;
/* src = "generated/sv2v_out.v:17891.13-17891.35" */
input nt_branch_mispredict_i;
wire nt_branch_mispredict_i;
/* cellift = 32'd1 */
input nt_branch_mispredict_i_t0;
wire nt_branch_mispredict_i_t0;
/* src = "generated/sv2v_out.v:17885.20-17885.27" */
output [31:0] pc_id_o;
reg [31:0] pc_id_o;
/* cellift = 32'd1 */
output [31:0] pc_id_o_t0;
reg [31:0] pc_id_o_t0;
/* src = "generated/sv2v_out.v:17884.21-17884.28" */
output [31:0] pc_if_o;
wire [31:0] pc_if_o;
/* cellift = 32'd1 */
output [31:0] pc_if_o_t0;
wire [31:0] pc_if_o_t0;
/* src = "generated/sv2v_out.v:17908.14-17908.33" */
output pc_mismatch_alert_o;
wire pc_mismatch_alert_o;
/* cellift = 32'd1 */
output pc_mismatch_alert_o_t0;
wire pc_mismatch_alert_o_t0;
/* src = "generated/sv2v_out.v:17890.19-17890.27" */
input [2:0] pc_mux_i;
wire [2:0] pc_mux_i;
/* cellift = 32'd1 */
input [2:0] pc_mux_i_t0;
wire [2:0] pc_mux_i_t0;
/* src = "generated/sv2v_out.v:17889.13-17889.21" */
input pc_set_i;
wire pc_set_i;
/* cellift = 32'd1 */
input pc_set_i_t0;
wire pc_set_i_t0;
/* src = "generated/sv2v_out.v:17886.13-17886.25" */
input pmp_err_if_i;
wire pmp_err_if_i;
/* cellift = 32'd1 */
input pmp_err_if_i_t0;
wire pmp_err_if_i_t0;
/* src = "generated/sv2v_out.v:17887.13-17887.31" */
input pmp_err_if_plus2_i;
wire pmp_err_if_plus2_i;
/* cellift = 32'd1 */
input pmp_err_if_plus2_i_t0;
wire pmp_err_if_plus2_i_t0;
/* src = "generated/sv2v_out.v:17921.14-17921.27" */
wire [31:0] prefetch_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17921.14-17921.27" */
wire [31:0] prefetch_addr_t0;
/* src = "generated/sv2v_out.v:17920.7-17920.22" */
wire prefetch_branch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17920.7-17920.22" */
wire prefetch_branch_t0;
/* src = "generated/sv2v_out.v:17853.13-17853.18" */
input req_i;
wire req_i;
/* cellift = 32'd1 */
input req_i_t0;
wire req_i_t0;
/* src = "generated/sv2v_out.v:17851.13-17851.19" */
input rst_ni;
wire rst_ni;
assign \g_secure_pc.prev_instr_addr_incr  = pc_id_o + /* src = "generated/sv2v_out.v:18219.34-18219.86" */ _340_;
assign csr_mtvec_init_o = _316_ & /* src = "generated/sv2v_out.v:17981.28-17981.57" */ pc_set_i;
assign instr_intg_err_o = instr_intg_err & /* src = "generated/sv2v_out.v:18001.28-18001.59" */ instr_rvalid_i;
assign fetch_valid = fetch_valid_raw & /* src = "generated/sv2v_out.v:18004.23-18004.64" */ _050_;
assign _000_ = pc_if_o[1] & /* src = "generated/sv2v_out.v:18098.33-18098.72" */ _320_;
assign _002_ = _000_ & /* src = "generated/sv2v_out.v:18098.32-18098.94" */ pmp_err_if_plus2_i;
assign if_instr_err_plus2 = _323_ & /* src = "generated/sv2v_out.v:18098.30-18098.130" */ _042_;
assign _004_ = fetch_valid & /* src = "generated/sv2v_out.v:18102.12-18102.36" */ _043_;
assign _006_ = if_id_pipe_reg_we & /* src = "generated/sv2v_out.v:18157.29-18157.73" */ _041_;
assign _008_ = instr_valid_id_o & /* src = "generated/sv2v_out.v:18157.78-18157.117" */ _321_;
assign if_id_pipe_reg_we = fetch_valid & /* src = "generated/sv2v_out.v:18158.26-18158.56" */ id_in_ready_i;
assign _010_ = _325_ & /* src = "generated/sv2v_out.v:18213.32-18213.81" */ _041_;
assign _012_ = _010_ & /* src = "generated/sv2v_out.v:18213.31-18213.98" */ _322_;
assign \g_secure_pc.prev_instr_seq_d  = _012_ & /* src = "generated/sv2v_out.v:18213.30-18213.120" */ _036_;
assign pc_mismatch_alert_o = \g_secure_pc.prev_instr_seq_q  & /* src = "generated/sv2v_out.v:18224.33-18224.89" */ _318_;
assign fetch_ready = id_in_ready_i & /* src = "generated/sv2v_out.v:18305.25-18305.59" */ _036_;
assign _014_ = ~ pc_id_o_t0;
assign _015_ = ~ { 29'h00000000, instr_is_compressed_id_o_t0, instr_is_compressed_id_o_t0, 1'h0 };
assign _054_ = pc_id_o & _014_;
assign _055_ = _340_ & _015_;
assign _304_ = _054_ + _055_;
assign _189_ = pc_id_o | pc_id_o_t0;
assign _190_ = _340_ | { 29'h00000000, instr_is_compressed_id_o_t0, instr_is_compressed_id_o_t0, 1'h0 };
assign _305_ = _189_ + _190_;
assign _279_ = _304_ ^ _305_;
assign _191_ = _279_ | pc_id_o_t0;
assign \g_secure_pc.prev_instr_addr_incr_t0  = _191_ | { 29'h00000000, instr_is_compressed_id_o_t0, instr_is_compressed_id_o_t0, 1'h0 };
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME \g_secure_pc.prev_instr_seq_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_secure_pc.prev_instr_seq_q_t0  <= 1'h0;
else \g_secure_pc.prev_instr_seq_q_t0  <= \g_secure_pc.prev_instr_seq_d_t0 ;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_valid_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_valid_id_o_t0 <= 1'h0;
else instr_valid_id_o_t0 <= instr_valid_id_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_new_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_new_id_o_t0 <= 1'h0;
else instr_new_id_o_t0 <= if_id_pipe_reg_we_t0;
assign _016_ = ~ if_id_pipe_reg_we;
assign _280_ = \gen_dummy_instr.insert_dummy_instr  ^ dummy_instr_id_o;
assign _281_ = pc_if_o ^ pc_id_o;
assign _282_ = instr_out ^ instr_rdata_alu_id_o;
assign _283_ = fetch_rdata[15:0] ^ instr_rdata_c_id_o;
assign _284_ = instr_is_compressed_out ^ instr_is_compressed_id_o;
assign _285_ = instr_err_out ^ instr_fetch_err_o;
assign _286_ = if_instr_err_plus2 ^ instr_fetch_err_plus2_o;
assign _287_ = illegal_c_instr_out ^ illegal_c_insn_id_o;
assign _207_ = \gen_dummy_instr.insert_dummy_instr_t0  | dummy_instr_id_o_t0;
assign _211_ = pc_if_o_t0 | pc_id_o_t0;
assign _215_ = instr_out_t0 | instr_rdata_alu_id_o_t0;
assign _219_ = fetch_rdata_t0[15:0] | instr_rdata_c_id_o_t0;
assign _223_ = instr_is_compressed_out_t0 | instr_is_compressed_id_o_t0;
assign _227_ = instr_err_out_t0 | instr_fetch_err_o_t0;
assign _231_ = if_instr_err_plus2_t0 | instr_fetch_err_plus2_o_t0;
assign _235_ = illegal_c_instr_out_t0 | illegal_c_insn_id_o_t0;
assign _208_ = _280_ | _207_;
assign _212_ = _281_ | _211_;
assign _216_ = _282_ | _215_;
assign _220_ = _283_ | _219_;
assign _224_ = _284_ | _223_;
assign _228_ = _285_ | _227_;
assign _232_ = _286_ | _231_;
assign _236_ = _287_ | _235_;
assign _101_ = if_id_pipe_reg_we & \gen_dummy_instr.insert_dummy_instr_t0 ;
assign _104_ = { if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we } & pc_if_o_t0;
assign _107_ = { if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we } & instr_out_t0;
assign _110_ = { if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we, if_id_pipe_reg_we } & fetch_rdata_t0[15:0];
assign _113_ = if_id_pipe_reg_we & instr_is_compressed_out_t0;
assign _116_ = if_id_pipe_reg_we & instr_err_out_t0;
assign _119_ = if_id_pipe_reg_we & if_instr_err_plus2_t0;
assign _122_ = if_id_pipe_reg_we & illegal_c_instr_out_t0;
assign _102_ = _016_ & dummy_instr_id_o_t0;
assign _105_ = { _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_ } & pc_id_o_t0;
assign _108_ = { _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_ } & instr_rdata_alu_id_o_t0;
assign _111_ = { _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_, _016_ } & instr_rdata_c_id_o_t0;
assign _114_ = _016_ & instr_is_compressed_id_o_t0;
assign _117_ = _016_ & instr_fetch_err_o_t0;
assign _120_ = _016_ & instr_fetch_err_plus2_o_t0;
assign _123_ = _016_ & illegal_c_insn_id_o_t0;
assign _103_ = _208_ & if_id_pipe_reg_we_t0;
assign _106_ = _212_ & { if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0 };
assign _109_ = _216_ & { if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0 };
assign _112_ = _220_ & { if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0, if_id_pipe_reg_we_t0 };
assign _115_ = _224_ & if_id_pipe_reg_we_t0;
assign _118_ = _228_ & if_id_pipe_reg_we_t0;
assign _121_ = _232_ & if_id_pipe_reg_we_t0;
assign _124_ = _236_ & if_id_pipe_reg_we_t0;
assign _209_ = _101_ | _102_;
assign _213_ = _104_ | _105_;
assign _217_ = _107_ | _108_;
assign _221_ = _110_ | _111_;
assign _225_ = _113_ | _114_;
assign _229_ = _116_ | _117_;
assign _233_ = _119_ | _120_;
assign _237_ = _122_ | _123_;
assign _210_ = _209_ | _103_;
assign _214_ = _213_ | _106_;
assign _218_ = _217_ | _109_;
assign _222_ = _221_ | _112_;
assign _226_ = _225_ | _115_;
assign _230_ = _229_ | _118_;
assign _234_ = _233_ | _121_;
assign _238_ = _237_ | _124_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME dummy_instr_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_instr_id_o_t0 <= 1'h0;
else dummy_instr_id_o_t0 <= _210_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME pc_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) pc_id_o_t0 <= 32'd0;
else pc_id_o_t0 <= _214_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_rdata_alu_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_rdata_alu_id_o_t0 <= 32'd0;
else instr_rdata_alu_id_o_t0 <= _218_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_rdata_c_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_rdata_c_id_o_t0 <= 16'h0000;
else instr_rdata_c_id_o_t0 <= _222_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_is_compressed_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_is_compressed_id_o_t0 <= 1'h0;
else instr_is_compressed_id_o_t0 <= _226_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_fetch_err_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_fetch_err_o_t0 <= 1'h0;
else instr_fetch_err_o_t0 <= _230_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_fetch_err_plus2_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_fetch_err_plus2_o_t0 <= 1'h0;
else instr_fetch_err_plus2_o_t0 <= _234_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME illegal_c_insn_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) illegal_c_insn_id_o_t0 <= 1'h0;
else illegal_c_insn_id_o_t0 <= _238_;
assign _056_ = _317_ & pc_set_i;
assign _059_ = instr_intg_err_t0 & instr_rvalid_i;
assign _062_ = fetch_valid_raw_t0 & _050_;
assign _065_ = pc_if_o_t0[1] & _320_;
assign _068_ = _001_ & pmp_err_if_plus2_i;
assign _071_ = _324_ & _042_;
assign _074_ = fetch_valid_t0 & _043_;
assign _077_ = if_id_pipe_reg_we_t0 & _041_;
assign _080_ = instr_valid_id_o_t0 & _321_;
assign _083_ = fetch_valid_t0 & id_in_ready_i;
assign _086_ = _326_ & _041_;
assign _089_ = _011_ & _322_;
assign _092_ = _013_ & _036_;
assign _095_ = \g_secure_pc.prev_instr_seq_q_t0  & _318_;
assign _098_ = id_in_ready_i_t0 & _036_;
assign _057_ = pc_set_i_t0 & _316_;
assign _060_ = instr_rvalid_i_t0 & instr_intg_err;
assign _063_ = nt_branch_mispredict_i_t0 & fetch_valid_raw;
assign _066_ = instr_is_compressed_t0 & pc_if_o[1];
assign _069_ = pmp_err_if_plus2_i_t0 & _000_;
assign _072_ = pmp_err_if_i_t0 & _323_;
assign _075_ = fetch_err_t0 & fetch_valid;
assign _078_ = pc_set_i_t0 & if_id_pipe_reg_we;
assign _081_ = instr_valid_clear_i_t0 & instr_valid_id_o;
assign _084_ = id_in_ready_i_t0 & fetch_valid;
assign _087_ = pc_set_i_t0 & _325_;
assign _090_ = if_instr_err_t0 & _010_;
assign _093_ = \gen_dummy_instr.insert_dummy_instr_t0  & _012_;
assign _096_ = _319_ & \g_secure_pc.prev_instr_seq_q ;
assign _099_ = \gen_dummy_instr.insert_dummy_instr_t0  & id_in_ready_i;
assign _058_ = _317_ & pc_set_i_t0;
assign _061_ = instr_intg_err_t0 & instr_rvalid_i_t0;
assign _064_ = fetch_valid_raw_t0 & nt_branch_mispredict_i_t0;
assign _067_ = pc_if_o_t0[1] & instr_is_compressed_t0;
assign _070_ = _001_ & pmp_err_if_plus2_i_t0;
assign _073_ = _324_ & pmp_err_if_i_t0;
assign _076_ = fetch_valid_t0 & fetch_err_t0;
assign _079_ = if_id_pipe_reg_we_t0 & pc_set_i_t0;
assign _082_ = instr_valid_id_o_t0 & instr_valid_clear_i_t0;
assign _085_ = fetch_valid_t0 & id_in_ready_i_t0;
assign _088_ = _326_ & pc_set_i_t0;
assign _091_ = _011_ & if_instr_err_t0;
assign _094_ = _013_ & \gen_dummy_instr.insert_dummy_instr_t0 ;
assign _097_ = \g_secure_pc.prev_instr_seq_q_t0  & _319_;
assign _100_ = id_in_ready_i_t0 & \gen_dummy_instr.insert_dummy_instr_t0 ;
assign _192_ = _056_ | _057_;
assign _193_ = _059_ | _060_;
assign _194_ = _062_ | _063_;
assign _195_ = _065_ | _066_;
assign _196_ = _068_ | _069_;
assign _197_ = _071_ | _072_;
assign _198_ = _074_ | _075_;
assign _199_ = _077_ | _078_;
assign _200_ = _080_ | _081_;
assign _201_ = _083_ | _084_;
assign _202_ = _086_ | _087_;
assign _203_ = _089_ | _090_;
assign _204_ = _092_ | _093_;
assign _205_ = _095_ | _096_;
assign _206_ = _098_ | _099_;
assign csr_mtvec_init_o_t0 = _192_ | _058_;
assign instr_intg_err_o_t0 = _193_ | _061_;
assign fetch_valid_t0 = _194_ | _064_;
assign _001_ = _195_ | _067_;
assign _003_ = _196_ | _070_;
assign if_instr_err_plus2_t0 = _197_ | _073_;
assign _005_ = _198_ | _076_;
assign _007_ = _199_ | _079_;
assign _009_ = _200_ | _082_;
assign if_id_pipe_reg_we_t0 = _201_ | _085_;
assign _011_ = _202_ | _088_;
assign _013_ = _203_ | _091_;
assign \g_secure_pc.prev_instr_seq_d_t0  = _204_ | _094_;
assign pc_mismatch_alert_o_t0 = _205_ | _097_;
assign fetch_ready_t0 = _206_ | _100_;
assign _017_ = | { pc_if_o_t0, \g_secure_pc.prev_instr_addr_incr_buf_t0  };
assign _018_ = | pc_mux_i_t0;
assign _019_ = | exc_pc_mux_i_t0;
assign _259_ = pc_if_o_t0 | \g_secure_pc.prev_instr_addr_incr_buf_t0 ;
assign _020_ = ~ _259_;
assign _021_ = ~ pc_mux_i_t0;
assign _022_ = ~ exc_pc_mux_i_t0;
assign _150_ = pc_if_o & _020_;
assign _149_ = pc_mux_i & _021_;
assign _173_ = exc_pc_mux_i & _022_;
assign _151_ = \g_secure_pc.prev_instr_addr_incr_buf  & _020_;
assign _296_ = _150_ == _151_;
assign _297_ = _149_ == { _021_[2], 2'h0 };
assign _298_ = _149_ == { 1'h0, _021_[1:0] };
assign _299_ = _149_ == { 1'h0, _021_[1], 1'h0 };
assign _300_ = _149_ == { 2'h0, _021_[0] };
assign _301_ = _173_ == _022_;
assign _302_ = _173_ == { _022_[1], 1'h0 };
assign _303_ = _173_ == { 1'h0, _022_[0] };
assign _319_ = _296_ & _017_;
assign _328_ = _297_ & _018_;
assign _330_ = _298_ & _018_;
assign _332_ = _299_ & _018_;
assign _334_ = _300_ & _018_;
assign _313_[3] = _301_ & _019_;
assign _337_ = _302_ & _019_;
assign _339_ = _303_ & _019_;
/* src = "generated/sv2v_out.v:18132.4-18136.45" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME dummy_instr_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) dummy_instr_id_o <= 1'h0;
else if (if_id_pipe_reg_we) dummy_instr_id_o <= \gen_dummy_instr.insert_dummy_instr ;
/* src = "generated/sv2v_out.v:18173.4-18193.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME pc_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) pc_id_o <= 32'd0;
else if (if_id_pipe_reg_we) pc_id_o <= pc_if_o;
/* src = "generated/sv2v_out.v:18173.4-18193.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_rdata_alu_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_rdata_alu_id_o <= 32'd0;
else if (if_id_pipe_reg_we) instr_rdata_alu_id_o <= instr_out;
/* src = "generated/sv2v_out.v:18173.4-18193.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_rdata_c_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_rdata_c_id_o <= 16'h0000;
else if (if_id_pipe_reg_we) instr_rdata_c_id_o <= fetch_rdata[15:0];
/* src = "generated/sv2v_out.v:18173.4-18193.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_is_compressed_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_is_compressed_id_o <= 1'h0;
else if (if_id_pipe_reg_we) instr_is_compressed_id_o <= instr_is_compressed_out;
/* src = "generated/sv2v_out.v:18173.4-18193.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_fetch_err_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_fetch_err_o <= 1'h0;
else if (if_id_pipe_reg_we) instr_fetch_err_o <= instr_err_out;
/* src = "generated/sv2v_out.v:18173.4-18193.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_fetch_err_plus2_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_fetch_err_plus2_o <= 1'h0;
else if (if_id_pipe_reg_we) instr_fetch_err_plus2_o <= if_instr_err_plus2;
/* src = "generated/sv2v_out.v:18173.4-18193.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME illegal_c_insn_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) illegal_c_insn_id_o <= 1'h0;
else if (if_id_pipe_reg_we) illegal_c_insn_id_o <= illegal_c_instr_out;
assign _023_ = | \g_mem_ecc.ecc_err_t0 ;
assign _024_ = ~ \g_mem_ecc.ecc_err_t0 ;
assign _176_ = \g_mem_ecc.ecc_err  & _024_;
assign _025_ = ! _149_;
assign _026_ = ! _176_;
assign _317_ = _025_ & _018_;
assign instr_intg_err_t0 = _026_ & _023_;
assign _027_ = ~ { _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_ };
assign _028_ = ~ { _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_ };
assign _029_ = ~ { _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_ };
assign _030_ = ~ { _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_ };
assign _031_ = ~ { _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_ };
assign _032_ = ~ { _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_ };
assign _033_ = ~ { exc_cause[6], exc_cause[6], exc_cause[6], exc_cause[6], exc_cause[6] };
assign _034_ = ~ { pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i };
assign _035_ = ~ { \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr  };
assign _036_ = ~ \gen_dummy_instr.insert_dummy_instr ;
assign _241_ = { _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_ } | _027_;
assign _244_ = { _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_ } | _028_;
assign _247_ = { _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_ } | _029_;
assign _250_ = { _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_ } | _030_;
assign _253_ = { _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_ } | _031_;
assign _256_ = { _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_ } | _032_;
assign _267_ = { exc_cause_t0[6], exc_cause_t0[6], exc_cause_t0[6], exc_cause_t0[6], exc_cause_t0[6] } | _033_;
assign _268_ = { pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0 } | _034_;
assign _271_ = { \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0  } | _035_;
assign _274_ = \gen_dummy_instr.insert_dummy_instr_t0  | _036_;
assign _242_ = { _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_ } | { _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_, _327_ };
assign _245_ = { _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_ } | { _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_, _333_ };
assign _248_ = { _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_ } | { _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_, _331_ };
assign _251_ = { _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_ } | { _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_, _275_ };
assign _254_ = { _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_ } | { _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_, _338_ };
assign _257_ = { _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_ } | { _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_, _277_ };
assign _269_ = { pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0 } | { pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i, pc_set_i };
assign _272_ = { \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0  } | { \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr , \gen_dummy_instr.insert_dummy_instr  };
assign _131_ = csr_mepc_i_t0 & _241_;
assign _134_ = { boot_addr_i_t0[31:8], 8'h00 } & _244_;
assign _137_ = _309_ & _247_;
assign _140_ = _311_ & _250_;
assign _143_ = { csr_mtvec_i_t0[31:8], 8'h00 } & _253_;
assign _146_ = _315_ & _256_;
assign _174_ = exc_cause_t0[4:0] & _267_;
assign _177_ = nt_branch_addr_i_t0 & _268_;
assign _180_ = instr_decompressed_t0 & _271_;
assign _183_ = instr_is_compressed_t0 & _274_;
assign _185_ = illegal_c_insn_t0 & _274_;
assign _187_ = if_instr_err_t0 & _274_;
assign _132_ = csr_depc_i_t0 & _242_;
assign _135_ = branch_target_ex_i_t0 & _245_;
assign _138_ = exc_pc_t0 & _248_;
assign _141_ = _307_ & _251_;
assign _144_ = { csr_mtvec_i_t0[31:8], 1'h0, irq_vec_t0, 2'h0 } & _254_;
assign _147_ = { 28'h0000000, _313_[3], 3'h0 } & _257_;
assign _178_ = { fetch_addr_n_t0[31:1], 1'h0 } & _269_;
assign _181_ = \gen_dummy_instr.dummy_instr_data_t0  & _272_;
assign _243_ = _131_ | _132_;
assign _246_ = _134_ | _135_;
assign _249_ = _137_ | _138_;
assign _252_ = _140_ | _141_;
assign _255_ = _143_ | _144_;
assign _258_ = _146_ | _147_;
assign _270_ = _177_ | _178_;
assign _273_ = _180_ | _181_;
assign _288_ = csr_mepc_i ^ csr_depc_i;
assign _289_ = { boot_addr_i[31:8], 8'h80 } ^ branch_target_ex_i;
assign _290_ = _308_ ^ exc_pc;
assign _291_ = _310_ ^ _306_;
assign _292_ = { csr_mtvec_i[31:8], 8'h00 } ^ { csr_mtvec_i[31:8], 1'h0, irq_vec, 2'h0 };
assign _293_ = _314_ ^ _312_;
assign _294_ = nt_branch_addr_i ^ { fetch_addr_n[31:1], 1'h0 };
assign _295_ = instr_decompressed ^ \gen_dummy_instr.dummy_instr_data ;
assign _133_ = { _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_, _328_ } & _288_;
assign _136_ = { _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_, _334_ } & _289_;
assign _139_ = { _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_, _332_ } & _290_;
assign _142_ = { _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_, _276_ } & _291_;
assign _145_ = { _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_, _339_ } & _292_;
assign _148_ = { _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_, _278_ } & _293_;
assign _175_ = { exc_cause_t0[6], exc_cause_t0[6], exc_cause_t0[6], exc_cause_t0[6], exc_cause_t0[6] } & _037_;
assign _179_ = { pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0, pc_set_i_t0 } & _294_;
assign _182_ = { \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0 , \gen_dummy_instr.insert_dummy_instr_t0  } & _295_;
assign _184_ = \gen_dummy_instr.insert_dummy_instr_t0  & instr_is_compressed;
assign _186_ = \gen_dummy_instr.insert_dummy_instr_t0  & illegal_c_insn;
assign _188_ = \gen_dummy_instr.insert_dummy_instr_t0  & if_instr_err;
assign _307_ = _133_ | _243_;
assign _309_ = _136_ | _246_;
assign _311_ = _139_ | _249_;
assign fetch_addr_n_t0 = _142_ | _252_;
assign _315_ = _145_ | _255_;
assign exc_pc_t0 = _148_ | _258_;
assign irq_vec_t0 = _175_ | _174_;
assign prefetch_addr_t0 = _179_ | _270_;
assign instr_out_t0 = _182_ | _273_;
assign instr_is_compressed_out_t0 = _184_ | _183_;
assign illegal_c_instr_out_t0 = _186_ | _185_;
assign instr_err_out_t0 = _188_ | _187_;
assign _037_ = ~ exc_cause[4:0];
assign _038_ = ~ _329_;
assign _039_ = ~ _336_;
assign _040_ = ~ instr_intg_err;
assign _041_ = ~ pc_set_i;
assign _042_ = ~ pmp_err_if_i;
assign _043_ = ~ fetch_err;
assign _044_ = ~ _002_;
assign _045_ = ~ _006_;
assign _046_ = ~ \g_secure_pc.prev_instr_seq_q ;
assign _047_ = ~ _327_;
assign _048_ = ~ _335_;
assign _049_ = ~ instr_bus_err_i;
assign _050_ = ~ nt_branch_mispredict_i;
assign _051_ = ~ if_instr_pmp_err;
assign _052_ = ~ fetch_err_plus2;
assign _053_ = ~ _008_;
assign _125_ = _330_ & _047_;
assign _128_ = _337_ & _048_;
assign _152_ = instr_intg_err_t0 & _049_;
assign _155_ = pc_set_i_t0 & _050_;
assign _158_ = pmp_err_if_i_t0 & _044_;
assign _161_ = fetch_err_t0 & _051_;
assign _164_ = _003_ & _052_;
assign _167_ = _007_ & _053_;
assign _170_ = \g_secure_pc.prev_instr_seq_q_t0  & _016_;
assign _126_ = _328_ & _038_;
assign _129_ = _313_[3] & _039_;
assign _153_ = instr_bus_err_i_t0 & _040_;
assign _156_ = nt_branch_mispredict_i_t0 & _041_;
assign _159_ = _003_ & _042_;
assign _162_ = if_instr_pmp_err_t0 & _043_;
assign _165_ = fetch_err_plus2_t0 & _044_;
assign _168_ = _009_ & _045_;
assign _171_ = if_id_pipe_reg_we_t0 & _046_;
assign _127_ = _330_ & _328_;
assign _130_ = _337_ & _313_[3];
assign _154_ = instr_intg_err_t0 & instr_bus_err_i_t0;
assign _157_ = pc_set_i_t0 & nt_branch_mispredict_i_t0;
assign _160_ = pmp_err_if_i_t0 & _003_;
assign _163_ = fetch_err_t0 & if_instr_pmp_err_t0;
assign _166_ = _003_ & fetch_err_plus2_t0;
assign _169_ = _007_ & _009_;
assign _172_ = \g_secure_pc.prev_instr_seq_q_t0  & if_id_pipe_reg_we_t0;
assign _239_ = _125_ | _126_;
assign _240_ = _128_ | _129_;
assign _260_ = _152_ | _153_;
assign _261_ = _155_ | _156_;
assign _262_ = _158_ | _159_;
assign _263_ = _161_ | _162_;
assign _264_ = _164_ | _165_;
assign _265_ = _167_ | _168_;
assign _266_ = _170_ | _171_;
assign _276_ = _239_ | _127_;
assign _278_ = _240_ | _130_;
assign instr_err_t0 = _260_ | _154_;
assign prefetch_branch_t0 = _261_ | _157_;
assign if_instr_pmp_err_t0 = _262_ | _160_;
assign if_instr_err_t0 = _263_ | _163_;
assign _324_ = _264_ | _166_;
assign instr_valid_id_d_t0 = _265_ | _169_;
assign _326_ = _266_ | _172_;
assign _275_ = _329_ | _327_;
assign _277_ = _336_ | _335_;
assign _306_ = _327_ ? csr_depc_i : csr_mepc_i;
assign _308_ = _333_ ? branch_target_ex_i : { boot_addr_i[31:8], 8'h80 };
assign _310_ = _331_ ? exc_pc : _308_;
assign fetch_addr_n = _275_ ? _306_ : _310_;
assign _312_ = _335_ ? 32'd437323784 : 32'd437323776;
assign _314_ = _338_ ? { csr_mtvec_i[31:8], 1'h0, irq_vec, 2'h0 } : { csr_mtvec_i[31:8], 8'h00 };
assign exc_pc = _277_ ? _312_ : _314_;
assign _316_ = ! /* src = "generated/sv2v_out.v:17981.29-17981.45" */ pc_mux_i;
assign _318_ = pc_if_o != /* src = "generated/sv2v_out.v:18224.53-18224.88" */ \g_secure_pc.prev_instr_addr_incr_buf ;
assign _320_ = ~ /* src = "generated/sv2v_out.v:18098.52-18098.72" */ instr_is_compressed;
assign _321_ = ~ /* src = "generated/sv2v_out.v:18157.97-18157.117" */ instr_valid_clear_i;
assign _322_ = ~ /* src = "generated/sv2v_out.v:18213.85-18213.98" */ if_instr_err;
assign instr_err = instr_intg_err | /* src = "generated/sv2v_out.v:18000.21-18000.53" */ instr_bus_err_i;
assign prefetch_branch = pc_set_i | /* src = "generated/sv2v_out.v:18002.27-18002.62" */ nt_branch_mispredict_i;
assign if_instr_pmp_err = pmp_err_if_i | /* src = "generated/sv2v_out.v:18096.28-18096.107" */ _002_;
assign if_instr_err = fetch_err | /* src = "generated/sv2v_out.v:18097.24-18097.59" */ if_instr_pmp_err;
assign _323_ = _002_ | /* src = "generated/sv2v_out.v:18098.31-18098.113" */ fetch_err_plus2;
assign instr_valid_id_d = _006_ | /* src = "generated/sv2v_out.v:18157.28-18157.118" */ _008_;
assign _325_ = \g_secure_pc.prev_instr_seq_q  | /* src = "generated/sv2v_out.v:18213.33-18213.66" */ if_id_pipe_reg_we;
/* src = "generated/sv2v_out.v:18214.4-18218.43" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME \g_secure_pc.prev_instr_seq_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_secure_pc.prev_instr_seq_q  <= 1'h0;
else \g_secure_pc.prev_instr_seq_q  <= \g_secure_pc.prev_instr_seq_d ;
/* src = "generated/sv2v_out.v:18159.2-18167.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_valid_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_valid_id_o <= 1'h0;
else instr_valid_id_o <= instr_valid_id_d;
/* src = "generated/sv2v_out.v:18159.2-18167.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$8b70aa1c3f3184a39244ef702f2b1543a1aeacb2\ibex_if_stage  */
/* PC_TAINT_INFO STATE_NAME instr_new_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_new_id_o <= 1'h0;
else instr_new_id_o <= if_id_pipe_reg_we;
assign _327_ = pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17971.3-17979.10" */ 3'h4;
assign _329_ = pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17971.3-17979.10" */ 3'h3;
assign _331_ = pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17971.3-17979.10" */ 3'h2;
assign _333_ = pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17971.3-17979.10" */ 3'h1;
assign _335_ = exc_pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17961.3-17967.10" */ 2'h3;
assign _336_ = exc_pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17961.3-17967.10" */ 2'h2;
assign _338_ = exc_pc_mux_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17961.3-17967.10" */ 2'h1;
assign irq_vec = exc_cause[6] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17959.7-17959.19|generated/sv2v_out.v:17959.3-17960.43" */ 5'h1f : exc_cause[4:0];
assign instr_intg_err = | /* src = "generated/sv2v_out.v:17994.28-17994.36" */ \g_mem_ecc.ecc_err ;
assign prefetch_addr = pc_set_i ? /* src = "generated/sv2v_out.v:18003.26-18003.84" */ { fetch_addr_n[31:1], 1'h0 } : nt_branch_addr_i;
assign instr_out = \gen_dummy_instr.insert_dummy_instr  ? /* src = "generated/sv2v_out.v:18127.24-18127.82" */ \gen_dummy_instr.dummy_instr_data  : instr_decompressed;
assign instr_is_compressed_out = \gen_dummy_instr.insert_dummy_instr  ? /* src = "generated/sv2v_out.v:18128.38-18128.85" */ 1'h0 : instr_is_compressed;
assign illegal_c_instr_out = \gen_dummy_instr.insert_dummy_instr  ? /* src = "generated/sv2v_out.v:18129.34-18129.76" */ 1'h0 : illegal_c_insn;
assign instr_err_out = \gen_dummy_instr.insert_dummy_instr  ? /* src = "generated/sv2v_out.v:18130.28-18130.68" */ 1'h0 : if_instr_err;
assign _340_ = instr_is_compressed_id_o ? /* src = "generated/sv2v_out.v:18219.45-18219.85" */ 32'd2 : 32'd4;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18099.26-18107.3" */
ibex_compressed_decoder compressed_decoder_i (
.clk_i(clk_i),
.illegal_instr_o(illegal_c_insn),
.illegal_instr_o_t0(illegal_c_insn_t0),
.instr_i(fetch_rdata),
.instr_i_t0(fetch_rdata_t0),
.instr_o(instr_decompressed),
.instr_o_t0(instr_decompressed_t0),
.is_compressed_o(instr_is_compressed),
.is_compressed_o_t0(instr_is_compressed_t0),
.rst_ni(rst_ni),
.valid_i(_004_),
.valid_i_t0(_005_)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:17990.30-17993.5" */
prim_secded_inv_39_32_dec \g_mem_ecc.u_instr_intg_dec  (
.data_i(\g_mem_ecc.instr_rdata_buf ),
.data_i_t0(\g_mem_ecc.instr_rdata_buf_t0 ),
.err_o(\g_mem_ecc.ecc_err ),
.err_o_t0(\g_mem_ecc.ecc_err_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:17986.37-17989.5" */
\$paramod\prim_buf\Width=32'00000000000000000000000000100111  \g_mem_ecc.u_prim_buf_instr_rdata  (
.in_i(instr_rdata_i),
.in_i_t0(instr_rdata_i_t0),
.out_o(\g_mem_ecc.instr_rdata_buf ),
.out_o_t0(\g_mem_ecc.instr_rdata_buf_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18220.27-18223.5" */
\$paramod\prim_buf\Width=s32'00000000000000000000000000100000  \g_secure_pc.u_prev_instr_addr_incr_buf  (
.in_i(\g_secure_pc.prev_instr_addr_incr ),
.in_i_t0(\g_secure_pc.prev_instr_addr_incr_t0 ),
.out_o(\g_secure_pc.prev_instr_addr_incr_buf ),
.out_o_t0(\g_secure_pc.prev_instr_addr_incr_buf_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18115.6-18126.5" */
\$paramod$501c60d7519704ee720c78ef16ad88cf05835059\ibex_dummy_instr  \gen_dummy_instr.dummy_instr_i  (
.clk_i(clk_i),
.dummy_instr_data_o(\gen_dummy_instr.dummy_instr_data ),
.dummy_instr_data_o_t0(\gen_dummy_instr.dummy_instr_data_t0 ),
.dummy_instr_en_i(dummy_instr_en_i),
.dummy_instr_en_i_t0(dummy_instr_en_i_t0),
.dummy_instr_mask_i(dummy_instr_mask_i),
.dummy_instr_mask_i_t0(dummy_instr_mask_i_t0),
.dummy_instr_seed_en_i(dummy_instr_seed_en_i),
.dummy_instr_seed_en_i_t0(dummy_instr_seed_en_i_t0),
.dummy_instr_seed_i(dummy_instr_seed_i),
.dummy_instr_seed_i_t0(dummy_instr_seed_i_t0),
.fetch_valid_i(fetch_valid),
.fetch_valid_i_t0(fetch_valid_t0),
.id_in_ready_i(id_in_ready_i),
.id_in_ready_i_t0(id_in_ready_i_t0),
.insert_dummy_instr_o(\gen_dummy_instr.insert_dummy_instr ),
.insert_dummy_instr_o_t0(\gen_dummy_instr.insert_dummy_instr_t0 ),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18050.48-18069.5" */
\$paramod\ibex_prefetch_buffer\ResetAll=1'1  \gen_prefetch_buffer.prefetch_buffer_i  (
.addr_i(prefetch_addr),
.addr_i_t0(prefetch_addr_t0),
.addr_o(pc_if_o),
.addr_o_t0(pc_if_o_t0),
.branch_i(prefetch_branch),
.branch_i_t0(prefetch_branch_t0),
.busy_o(if_busy_o),
.busy_o_t0(if_busy_o_t0),
.clk_i(clk_i),
.err_o(fetch_err),
.err_o_t0(fetch_err_t0),
.err_plus2_o(fetch_err_plus2),
.err_plus2_o_t0(fetch_err_plus2_t0),
.instr_addr_o(instr_addr_o),
.instr_addr_o_t0(instr_addr_o_t0),
.instr_err_i(instr_err),
.instr_err_i_t0(instr_err_t0),
.instr_gnt_i(instr_gnt_i),
.instr_gnt_i_t0(instr_gnt_i_t0),
.instr_rdata_i(instr_rdata_i[31:0]),
.instr_rdata_i_t0(instr_rdata_i_t0[31:0]),
.instr_req_o(instr_req_o),
.instr_req_o_t0(instr_req_o_t0),
.instr_rvalid_i(instr_rvalid_i),
.instr_rvalid_i_t0(instr_rvalid_i_t0),
.rdata_o(fetch_rdata),
.rdata_o_t0(fetch_rdata_t0),
.ready_i(fetch_ready),
.ready_i_t0(fetch_ready_t0),
.req_i(req_i),
.req_i_t0(req_i_t0),
.rst_ni(rst_ni),
.valid_o(fetch_valid_raw),
.valid_o_t0(fetch_valid_raw_t0)
);
assign { _313_[31:4], _313_[2:0] } = 31'h00000000;
assign ic_data_addr_o = 8'h00;
assign ic_data_addr_o_t0 = 8'h00;
assign ic_data_req_o = 2'h0;
assign ic_data_req_o_t0 = 2'h0;
assign ic_data_wdata_o = 64'h0000000000000000;
assign ic_data_wdata_o_t0 = 64'h0000000000000000;
assign ic_data_write_o = 1'h0;
assign ic_data_write_o_t0 = 1'h0;
assign ic_scr_key_req_o = 1'h0;
assign ic_scr_key_req_o_t0 = 1'h0;
assign ic_tag_addr_o = 8'h00;
assign ic_tag_addr_o_t0 = 8'h00;
assign ic_tag_req_o = 2'h0;
assign ic_tag_req_o_t0 = 2'h0;
assign ic_tag_wdata_o = 22'h000000;
assign ic_tag_wdata_o_t0 = 22'h000000;
assign ic_tag_write_o = 1'h0;
assign ic_tag_write_o_t0 = 1'h0;
assign icache_ecc_error_o = 1'h0;
assign icache_ecc_error_o_t0 = 1'h0;
assign instr_bp_taken_o = 1'h0;
assign instr_bp_taken_o_t0 = 1'h0;
assign instr_rdata_id_o = instr_rdata_alu_id_o;
assign instr_rdata_id_o_t0 = instr_rdata_alu_id_o_t0;
endmodule

module \$paramod$916c47de983e2a42946808797a4a11650abb788f\prim_onehot_check (clk_i, rst_ni, oh_i, addr_i, en_i, err_o, addr_i_t0, en_i_t0, err_o_t0, oh_i_t0);
wire _0000_;
wire _0001_;
wire _0002_;
wire _0003_;
wire _0004_;
wire _0005_;
wire _0006_;
wire _0007_;
wire _0008_;
wire _0009_;
wire _0010_;
wire _0011_;
wire _0012_;
wire _0013_;
wire _0014_;
wire _0015_;
wire _0016_;
wire _0017_;
wire _0018_;
wire _0019_;
wire _0020_;
wire _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire _0026_;
wire _0027_;
wire _0028_;
wire _0029_;
wire _0030_;
wire _0031_;
wire _0032_;
wire _0033_;
wire _0034_;
wire _0035_;
wire _0036_;
wire _0037_;
wire _0038_;
wire _0039_;
wire _0040_;
wire _0041_;
wire _0042_;
wire _0043_;
wire _0044_;
wire _0045_;
wire _0046_;
wire _0047_;
wire _0048_;
wire _0049_;
wire _0050_;
wire _0051_;
wire _0052_;
wire _0053_;
wire _0054_;
wire _0055_;
wire _0056_;
wire _0057_;
wire _0058_;
wire _0059_;
wire _0060_;
wire _0061_;
wire _0062_;
wire _0063_;
wire _0064_;
wire _0065_;
wire _0066_;
wire _0067_;
wire _0068_;
wire _0069_;
wire _0070_;
wire _0071_;
wire _0072_;
wire _0073_;
wire _0074_;
wire _0075_;
wire _0076_;
wire _0077_;
wire _0078_;
wire _0079_;
wire _0080_;
wire _0081_;
wire _0082_;
wire _0083_;
wire _0084_;
wire _0085_;
wire _0086_;
wire _0087_;
wire _0088_;
wire _0089_;
wire _0090_;
wire _0091_;
wire _0092_;
wire _0093_;
wire _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire _0109_;
wire _0110_;
wire _0111_;
wire _0112_;
wire _0113_;
wire _0114_;
wire _0115_;
wire _0116_;
wire _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire _0139_;
wire _0140_;
wire _0141_;
wire _0142_;
wire _0143_;
wire _0144_;
wire _0145_;
wire _0146_;
wire _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
wire _0152_;
wire _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire _0186_;
wire _0187_;
wire _0188_;
wire _0189_;
wire _0190_;
wire _0191_;
wire _0192_;
wire _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire _0199_;
wire _0200_;
wire _0201_;
wire _0202_;
wire _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
wire _0221_;
wire _0222_;
wire _0223_;
wire _0224_;
wire _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire _0241_;
wire _0242_;
wire _0243_;
wire _0244_;
wire _0245_;
wire _0246_;
wire _0247_;
wire _0248_;
wire _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire _0271_;
wire _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire _0276_;
wire _0277_;
wire _0278_;
wire _0279_;
wire _0280_;
wire _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire _0285_;
wire _0286_;
wire _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire _0294_;
wire _0295_;
wire _0296_;
wire _0297_;
wire _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire _0324_;
wire _0325_;
wire _0326_;
wire _0327_;
wire _0328_;
wire _0329_;
wire _0330_;
wire _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire _0335_;
wire _0336_;
wire _0337_;
wire _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire _0344_;
wire _0345_;
wire _0346_;
wire _0347_;
wire _0348_;
wire _0349_;
wire _0350_;
wire _0351_;
wire _0352_;
wire _0353_;
wire _0354_;
wire _0355_;
wire _0356_;
wire _0357_;
wire _0358_;
wire _0359_;
wire _0360_;
wire _0361_;
wire _0362_;
wire _0363_;
wire _0364_;
wire _0365_;
wire _0366_;
wire _0367_;
wire _0368_;
wire _0369_;
wire _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire _0376_;
wire _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire _0382_;
wire _0383_;
wire _0384_;
wire _0385_;
wire _0386_;
wire _0387_;
wire _0388_;
wire _0389_;
wire _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire _0398_;
wire _0399_;
wire _0400_;
wire _0401_;
wire _0402_;
wire _0403_;
wire _0404_;
wire _0405_;
wire _0406_;
wire _0407_;
wire _0408_;
wire _0409_;
wire _0410_;
wire _0411_;
wire _0412_;
wire _0413_;
wire _0414_;
wire _0415_;
wire _0416_;
wire _0417_;
wire _0418_;
wire _0419_;
wire _0420_;
wire _0421_;
wire _0422_;
wire _0423_;
wire _0424_;
wire _0425_;
wire _0426_;
wire _0427_;
wire _0428_;
wire _0429_;
wire _0430_;
wire _0431_;
wire _0432_;
wire _0433_;
wire _0434_;
wire _0435_;
wire _0436_;
wire _0437_;
wire _0438_;
wire _0439_;
wire _0440_;
wire _0441_;
wire _0442_;
wire _0443_;
wire _0444_;
wire _0445_;
wire _0446_;
wire _0447_;
wire _0448_;
wire _0449_;
wire _0450_;
wire _0451_;
wire _0452_;
wire _0453_;
wire _0454_;
wire _0455_;
wire _0456_;
wire _0457_;
wire _0458_;
wire _0459_;
wire _0460_;
wire _0461_;
wire _0462_;
wire _0463_;
wire _0464_;
wire _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire _0469_;
wire _0470_;
wire _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire _0477_;
wire _0478_;
wire _0479_;
wire _0480_;
wire _0481_;
wire _0482_;
wire _0483_;
wire _0484_;
wire _0485_;
wire _0486_;
wire _0487_;
wire _0488_;
wire _0489_;
wire _0490_;
wire _0491_;
wire _0492_;
wire _0493_;
wire _0494_;
wire _0495_;
wire _0496_;
wire _0497_;
wire _0498_;
wire _0499_;
wire _0500_;
wire _0501_;
wire _0502_;
wire _0503_;
wire _0504_;
wire _0505_;
wire _0506_;
wire _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0517_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
wire _0525_;
wire _0526_;
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire _0534_;
wire _0535_;
wire _0536_;
wire _0537_;
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0542_;
wire _0543_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire _0560_;
wire _0561_;
wire _0562_;
wire _0563_;
wire _0564_;
wire _0565_;
wire _0566_;
wire _0567_;
wire _0568_;
wire _0569_;
wire _0570_;
wire _0571_;
wire _0572_;
wire _0573_;
wire _0574_;
wire _0575_;
wire _0576_;
wire _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire _0596_;
wire _0597_;
wire _0598_;
wire _0599_;
wire _0600_;
wire _0601_;
wire _0602_;
wire _0603_;
wire _0604_;
wire _0605_;
wire _0606_;
wire _0607_;
wire _0608_;
wire _0609_;
wire _0610_;
wire _0611_;
wire _0612_;
wire _0613_;
wire _0614_;
wire _0615_;
wire _0616_;
wire _0617_;
wire _0618_;
wire _0619_;
wire _0620_;
wire _0621_;
wire _0622_;
wire _0623_;
wire _0624_;
wire _0625_;
wire _0626_;
wire _0627_;
wire _0628_;
wire _0629_;
wire _0630_;
wire _0631_;
wire _0632_;
wire _0633_;
wire _0634_;
wire _0635_;
wire _0636_;
wire _0637_;
wire _0638_;
wire _0639_;
wire _0640_;
wire _0641_;
wire _0642_;
wire _0643_;
wire _0644_;
wire _0645_;
wire _0646_;
wire _0647_;
wire _0648_;
wire _0649_;
wire _0650_;
wire _0651_;
wire _0652_;
wire _0653_;
wire _0654_;
wire _0655_;
wire _0656_;
wire _0657_;
wire _0658_;
wire _0659_;
wire _0660_;
wire _0661_;
wire _0662_;
wire _0663_;
wire _0664_;
wire _0665_;
wire _0666_;
wire _0667_;
wire _0668_;
wire _0669_;
wire _0670_;
wire _0671_;
wire _0672_;
wire _0673_;
wire _0674_;
wire _0675_;
wire _0676_;
wire _0677_;
wire _0678_;
wire _0679_;
wire _0680_;
wire _0681_;
wire _0682_;
wire _0683_;
wire _0684_;
wire _0685_;
wire _0686_;
wire _0687_;
wire _0688_;
wire _0689_;
wire _0690_;
wire _0691_;
wire _0692_;
wire _0693_;
wire _0694_;
wire _0695_;
wire _0696_;
wire _0697_;
wire _0698_;
wire _0699_;
wire _0700_;
wire _0701_;
wire _0702_;
wire _0703_;
wire _0704_;
wire _0705_;
wire _0706_;
wire _0707_;
wire _0708_;
wire _0709_;
wire _0710_;
wire _0711_;
wire _0712_;
wire _0713_;
wire _0714_;
wire _0715_;
wire _0716_;
wire _0717_;
wire _0718_;
wire _0719_;
wire _0720_;
wire _0721_;
wire _0722_;
wire _0723_;
wire _0724_;
wire _0725_;
wire _0726_;
wire _0727_;
wire _0728_;
wire _0729_;
wire _0730_;
wire _0731_;
wire _0732_;
wire _0733_;
wire _0734_;
wire _0735_;
wire _0736_;
wire _0737_;
wire _0738_;
wire _0739_;
wire _0740_;
wire _0741_;
wire _0742_;
wire _0743_;
wire _0744_;
wire _0745_;
wire _0746_;
wire _0747_;
wire _0748_;
wire _0749_;
wire _0750_;
wire _0751_;
wire _0752_;
wire _0753_;
wire _0754_;
wire _0755_;
wire _0756_;
wire _0757_;
wire _0758_;
wire _0759_;
wire _0760_;
wire _0761_;
wire _0762_;
wire _0763_;
wire _0764_;
wire _0765_;
wire _0766_;
wire _0767_;
wire _0768_;
wire _0769_;
wire _0770_;
wire _0771_;
wire _0772_;
wire _0773_;
wire _0774_;
wire _0775_;
wire _0776_;
wire _0777_;
wire _0778_;
wire _0779_;
wire _0780_;
wire _0781_;
wire _0782_;
wire _0783_;
wire _0784_;
wire _0785_;
wire _0786_;
wire _0787_;
wire _0788_;
wire _0789_;
wire _0790_;
wire _0791_;
wire _0792_;
wire _0793_;
wire _0794_;
wire _0795_;
wire _0796_;
wire _0797_;
wire _0798_;
wire _0799_;
wire _0800_;
wire _0801_;
wire _0802_;
wire _0803_;
wire _0804_;
wire _0805_;
wire _0806_;
wire _0807_;
wire _0808_;
wire _0809_;
wire _0810_;
wire _0811_;
wire _0812_;
wire _0813_;
wire _0814_;
wire _0815_;
wire _0816_;
wire _0817_;
wire _0818_;
wire _0819_;
wire _0820_;
wire _0821_;
wire _0822_;
wire _0823_;
wire _0824_;
wire _0825_;
wire _0826_;
wire _0827_;
wire _0828_;
wire _0829_;
wire _0830_;
wire _0831_;
wire _0832_;
wire _0833_;
wire _0834_;
wire _0835_;
wire _0836_;
wire _0837_;
wire _0838_;
wire _0839_;
wire _0840_;
wire _0841_;
wire _0842_;
wire _0843_;
wire _0844_;
wire _0845_;
wire _0846_;
wire _0847_;
wire _0848_;
wire _0849_;
wire _0850_;
wire _0851_;
wire _0852_;
wire _0853_;
wire _0854_;
wire _0855_;
wire _0856_;
wire _0857_;
wire _0858_;
wire _0859_;
wire _0860_;
wire _0861_;
wire _0862_;
wire _0863_;
wire _0864_;
wire _0865_;
wire _0866_;
wire _0867_;
wire _0868_;
wire _0869_;
wire _0870_;
wire _0871_;
wire _0872_;
wire _0873_;
wire _0874_;
wire _0875_;
wire _0876_;
wire _0877_;
wire _0878_;
wire _0879_;
wire _0880_;
wire _0881_;
wire _0882_;
wire _0883_;
wire _0884_;
wire _0885_;
wire _0886_;
wire _0887_;
wire _0888_;
wire _0889_;
wire _0890_;
wire _0891_;
wire _0892_;
wire _0893_;
wire _0894_;
wire _0895_;
wire _0896_;
wire _0897_;
wire _0898_;
wire _0899_;
wire _0900_;
wire _0901_;
wire _0902_;
wire _0903_;
wire _0904_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0905_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0906_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0907_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0908_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0909_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0910_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0911_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0912_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0913_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0914_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0915_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0916_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0917_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0918_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0919_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0920_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0921_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0922_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0923_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0924_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0925_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0926_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0927_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0928_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0929_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0930_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0931_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0932_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0933_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0934_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0935_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0936_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0937_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0938_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0939_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0940_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0941_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0942_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0943_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0944_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0945_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0946_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0947_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0948_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0949_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0950_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0951_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0952_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0953_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0954_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0955_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0956_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0957_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0958_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0959_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0960_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0961_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0962_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0963_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0964_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0965_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0966_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0967_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0968_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0969_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0970_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0971_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0972_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0973_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0974_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0975_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0976_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0977_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0978_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0979_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0980_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0981_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0982_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0983_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0984_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0985_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0986_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0987_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0988_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0989_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0990_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0991_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0992_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0993_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0994_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0995_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0996_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0997_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _0998_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _0999_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _1000_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _1001_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _1002_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _1003_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _1004_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _1005_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _1006_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _1007_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _1008_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _1009_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _1010_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _1011_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _1012_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _1013_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _1014_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _1015_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _1016_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _1017_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _1018_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _1019_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _1020_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _1021_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _1022_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _1023_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _1024_;
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _1025_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.29-26484.77" */
wire _1026_;
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _1027_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26484.83-26484.130" */
wire _1028_;
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1029_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1030_;
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1031_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1032_;
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1033_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1034_;
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1035_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1036_;
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1037_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1038_;
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1039_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1040_;
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1041_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1042_;
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1043_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1044_;
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1045_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1046_;
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1047_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1048_;
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1049_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1050_;
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1051_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1052_;
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1053_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1054_;
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1055_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1056_;
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1057_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.30-26485.56" */
wire _1058_;
/* src = "generated/sv2v_out.v:26484.29-26484.61" */
wire _1059_;
/* src = "generated/sv2v_out.v:26484.29-26484.61" */
wire _1060_;
/* src = "generated/sv2v_out.v:26484.29-26484.61" */
wire _1061_;
/* src = "generated/sv2v_out.v:26484.29-26484.61" */
wire _1062_;
/* src = "generated/sv2v_out.v:26484.29-26484.61" */
wire _1063_;
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1064_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1065_;
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1066_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1067_;
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1068_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1069_;
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1070_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1071_;
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1072_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1073_;
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1074_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1075_;
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1076_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1077_;
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1078_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1079_;
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1080_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1081_;
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1082_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1083_;
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1084_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1085_;
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1086_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1087_;
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1088_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1089_;
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1090_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1091_;
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1092_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26485.29-26485.73" */
wire _1093_;
/* src = "generated/sv2v_out.v:26493.18-26493.39" */
wire _1094_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26493.18-26493.39" */
wire _1095_;
/* src = "generated/sv2v_out.v:26491.7-26491.15" */
wire addr_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26491.7-26491.15" */
wire addr_err_t0;
/* src = "generated/sv2v_out.v:26454.31-26454.37" */
input [4:0] addr_i;
wire [4:0] addr_i;
/* cellift = 32'd1 */
input [4:0] addr_i_t0;
wire [4:0] addr_i_t0;
/* src = "generated/sv2v_out.v:26459.38-26459.46" */
wire [62:0] and_tree;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26459.38-26459.46" */
wire [62:0] and_tree_t0;
/* src = "generated/sv2v_out.v:26451.8-26451.13" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:26455.13-26455.17" */
input en_i;
wire en_i;
/* cellift = 32'd1 */
input en_i_t0;
wire en_i_t0;
/* src = "generated/sv2v_out.v:26490.7-26490.17" */
wire enable_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26490.7-26490.17" */
wire enable_err_t0;
/* src = "generated/sv2v_out.v:26456.14-26456.19" */
output err_o;
wire err_o;
/* cellift = 32'd1 */
output err_o_t0;
wire err_o_t0;
/* src = "generated/sv2v_out.v:26460.38-26460.46" */
wire [62:0] err_tree;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26460.38-26460.46" */
wire [62:0] err_tree_t0;
/* src = "generated/sv2v_out.v:26492.7-26492.14" */
wire oh0_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26492.7-26492.14" */
wire oh0_err_t0;
/* src = "generated/sv2v_out.v:26453.33-26453.37" */
input [31:0] oh_i;
wire [31:0] oh_i;
/* cellift = 32'd1 */
input [31:0] oh_i_t0;
wire [31:0] oh_i_t0;
/* src = "generated/sv2v_out.v:26458.38-26458.45" */
wire [62:0] or_tree;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:26458.38-26458.45" */
wire [62:0] or_tree_t0;
/* src = "generated/sv2v_out.v:26452.8-26452.14" */
input rst_ni;
wire rst_ni;
assign _0188_ = addr_i_t0[1] & and_tree[17];
assign _0191_ = addr_i_t0[1] & and_tree[18];
assign _0194_ = addr_i_t0[1] & and_tree[19];
assign _0197_ = addr_i_t0[1] & and_tree[20];
assign _0200_ = addr_i_t0[1] & and_tree[21];
assign _0203_ = addr_i_t0[1] & and_tree[22];
assign _0206_ = addr_i_t0[1] & and_tree[23];
assign _0209_ = addr_i_t0[1] & and_tree[24];
assign _0212_ = addr_i_t0[1] & and_tree[25];
assign _0215_ = addr_i_t0[1] & and_tree[26];
assign _0218_ = addr_i_t0[1] & and_tree[27];
assign _0221_ = addr_i_t0[1] & and_tree[28];
assign _0224_ = addr_i_t0[1] & and_tree[29];
assign _0227_ = addr_i_t0[1] & and_tree[30];
assign _0230_ = addr_i_t0[0] & oh_i[0];
assign _0233_ = addr_i_t0[0] & oh_i[1];
assign _0236_ = addr_i_t0[0] & oh_i[2];
assign _0239_ = addr_i_t0[0] & oh_i[3];
assign _0242_ = addr_i_t0[0] & oh_i[4];
assign _0245_ = addr_i_t0[0] & oh_i[5];
assign _0248_ = addr_i_t0[0] & oh_i[6];
assign _0251_ = addr_i_t0[0] & oh_i[7];
assign _0254_ = addr_i_t0[0] & oh_i[8];
assign _0257_ = addr_i_t0[0] & oh_i[9];
assign _0260_ = addr_i_t0[0] & oh_i[10];
assign _0263_ = addr_i_t0[0] & oh_i[11];
assign _0266_ = addr_i_t0[0] & oh_i[12];
assign _0269_ = addr_i_t0[0] & oh_i[13];
assign _0272_ = addr_i_t0[0] & oh_i[14];
assign _0275_ = addr_i_t0[0] & oh_i[15];
assign _0278_ = addr_i_t0[0] & oh_i[16];
assign _0281_ = addr_i_t0[0] & oh_i[17];
assign _0284_ = addr_i_t0[0] & oh_i[18];
assign _0287_ = addr_i_t0[0] & oh_i[19];
assign _0290_ = addr_i_t0[0] & oh_i[20];
assign _0293_ = addr_i_t0[0] & oh_i[21];
assign _0296_ = addr_i_t0[0] & oh_i[22];
assign _0299_ = addr_i_t0[0] & oh_i[23];
assign _0302_ = addr_i_t0[0] & oh_i[24];
assign _0305_ = addr_i_t0[0] & oh_i[25];
assign _0308_ = addr_i_t0[0] & oh_i[26];
assign _0311_ = addr_i_t0[0] & oh_i[27];
assign _0314_ = addr_i_t0[0] & oh_i[28];
assign _0317_ = addr_i_t0[0] & oh_i[29];
assign _0320_ = addr_i_t0[0] & oh_i[30];
assign _0323_ = addr_i_t0[0] & oh_i[31];
assign _0326_ = addr_i_t0[4] & and_tree[1];
assign _0329_ = addr_i_t0[4] & and_tree[2];
assign _0332_ = addr_i_t0[3] & and_tree[3];
assign _0335_ = addr_i_t0[3] & and_tree[4];
assign _0338_ = addr_i_t0[3] & and_tree[5];
assign _0341_ = addr_i_t0[3] & and_tree[6];
assign _0344_ = addr_i_t0[2] & and_tree[7];
assign _0347_ = addr_i_t0[2] & and_tree[8];
assign _0350_ = addr_i_t0[2] & and_tree[9];
assign _0353_ = addr_i_t0[2] & and_tree[10];
assign _0356_ = addr_i_t0[2] & and_tree[11];
assign _0359_ = addr_i_t0[2] & and_tree[12];
assign _0362_ = addr_i_t0[2] & and_tree[13];
assign _0365_ = addr_i_t0[2] & and_tree[14];
assign _0368_ = addr_i_t0[1] & and_tree[15];
assign _0371_ = addr_i_t0[1] & and_tree[16];
assign _0374_ = or_tree_t0[17] & or_tree[18];
assign _0377_ = or_tree_t0[19] & or_tree[20];
assign _0380_ = or_tree_t0[21] & or_tree[22];
assign _0383_ = or_tree_t0[23] & or_tree[24];
assign _0386_ = or_tree_t0[25] & or_tree[26];
assign _0389_ = or_tree_t0[27] & or_tree[28];
assign _0392_ = or_tree_t0[29] & or_tree[30];
assign _0395_ = oh_i_t0[0] & oh_i[1];
assign _0398_ = oh_i_t0[2] & oh_i[3];
assign _0401_ = oh_i_t0[4] & oh_i[5];
assign _0404_ = oh_i_t0[6] & oh_i[7];
assign _0407_ = oh_i_t0[8] & oh_i[9];
assign _0410_ = oh_i_t0[10] & oh_i[11];
assign _0413_ = oh_i_t0[12] & oh_i[13];
assign _0416_ = oh_i_t0[14] & oh_i[15];
assign _0419_ = oh_i_t0[16] & oh_i[17];
assign _0422_ = oh_i_t0[18] & oh_i[19];
assign _0425_ = oh_i_t0[20] & oh_i[21];
assign _0428_ = oh_i_t0[22] & oh_i[23];
assign _0431_ = oh_i_t0[24] & oh_i[25];
assign _0434_ = oh_i_t0[26] & oh_i[27];
assign _0437_ = oh_i_t0[28] & oh_i[29];
assign _0440_ = oh_i_t0[30] & oh_i[31];
assign _0443_ = or_tree_t0[1] & or_tree[2];
assign _0446_ = or_tree_t0[3] & or_tree[4];
assign _0449_ = or_tree_t0[5] & or_tree[6];
assign _0452_ = or_tree_t0[7] & or_tree[8];
assign _0455_ = or_tree_t0[9] & or_tree[10];
assign _0458_ = or_tree_t0[11] & or_tree[12];
assign _0461_ = or_tree_t0[13] & or_tree[14];
assign _0464_ = or_tree_t0[15] & or_tree[16];
assign _0189_ = and_tree_t0[17] & _1059_;
assign _0192_ = and_tree_t0[18] & addr_i[1];
assign _0195_ = and_tree_t0[19] & _1059_;
assign _0198_ = and_tree_t0[20] & addr_i[1];
assign _0201_ = and_tree_t0[21] & _1059_;
assign _0204_ = and_tree_t0[22] & addr_i[1];
assign _0207_ = and_tree_t0[23] & _1059_;
assign _0210_ = and_tree_t0[24] & addr_i[1];
assign _0213_ = and_tree_t0[25] & _1059_;
assign _0216_ = and_tree_t0[26] & addr_i[1];
assign _0219_ = and_tree_t0[27] & _1059_;
assign _0222_ = and_tree_t0[28] & addr_i[1];
assign _0225_ = and_tree_t0[29] & _1059_;
assign _0228_ = and_tree_t0[30] & addr_i[1];
assign _0231_ = oh_i_t0[0] & _1060_;
assign _0234_ = oh_i_t0[1] & addr_i[0];
assign _0237_ = oh_i_t0[2] & _1060_;
assign _0240_ = oh_i_t0[3] & addr_i[0];
assign _0243_ = oh_i_t0[4] & _1060_;
assign _0246_ = oh_i_t0[5] & addr_i[0];
assign _0249_ = oh_i_t0[6] & _1060_;
assign _0252_ = oh_i_t0[7] & addr_i[0];
assign _0255_ = oh_i_t0[8] & _1060_;
assign _0258_ = oh_i_t0[9] & addr_i[0];
assign _0261_ = oh_i_t0[10] & _1060_;
assign _0264_ = oh_i_t0[11] & addr_i[0];
assign _0267_ = oh_i_t0[12] & _1060_;
assign _0270_ = oh_i_t0[13] & addr_i[0];
assign _0273_ = oh_i_t0[14] & _1060_;
assign _0276_ = oh_i_t0[15] & addr_i[0];
assign _0279_ = oh_i_t0[16] & _1060_;
assign _0282_ = oh_i_t0[17] & addr_i[0];
assign _0285_ = oh_i_t0[18] & _1060_;
assign _0288_ = oh_i_t0[19] & addr_i[0];
assign _0291_ = oh_i_t0[20] & _1060_;
assign _0294_ = oh_i_t0[21] & addr_i[0];
assign _0297_ = oh_i_t0[22] & _1060_;
assign _0300_ = oh_i_t0[23] & addr_i[0];
assign _0303_ = oh_i_t0[24] & _1060_;
assign _0306_ = oh_i_t0[25] & addr_i[0];
assign _0309_ = oh_i_t0[26] & _1060_;
assign _0312_ = oh_i_t0[27] & addr_i[0];
assign _0315_ = oh_i_t0[28] & _1060_;
assign _0318_ = oh_i_t0[29] & addr_i[0];
assign _0321_ = oh_i_t0[30] & _1060_;
assign _0324_ = oh_i_t0[31] & addr_i[0];
assign _0327_ = and_tree_t0[1] & _1061_;
assign _0330_ = and_tree_t0[2] & addr_i[4];
assign _0333_ = and_tree_t0[3] & _1062_;
assign _0336_ = and_tree_t0[4] & addr_i[3];
assign _0339_ = and_tree_t0[5] & _1062_;
assign _0342_ = and_tree_t0[6] & addr_i[3];
assign _0345_ = and_tree_t0[7] & _1063_;
assign _0348_ = and_tree_t0[8] & addr_i[2];
assign _0351_ = and_tree_t0[9] & _1063_;
assign _0354_ = and_tree_t0[10] & addr_i[2];
assign _0357_ = and_tree_t0[11] & _1063_;
assign _0360_ = and_tree_t0[12] & addr_i[2];
assign _0363_ = and_tree_t0[13] & _1063_;
assign _0366_ = and_tree_t0[14] & addr_i[2];
assign _0369_ = and_tree_t0[15] & _1059_;
assign _0372_ = and_tree_t0[16] & addr_i[1];
assign _0375_ = or_tree_t0[18] & or_tree[17];
assign _0378_ = or_tree_t0[20] & or_tree[19];
assign _0381_ = or_tree_t0[22] & or_tree[21];
assign _0384_ = or_tree_t0[24] & or_tree[23];
assign _0387_ = or_tree_t0[26] & or_tree[25];
assign _0390_ = or_tree_t0[28] & or_tree[27];
assign _0393_ = or_tree_t0[30] & or_tree[29];
assign _0396_ = oh_i_t0[1] & oh_i[0];
assign _0399_ = oh_i_t0[3] & oh_i[2];
assign _0402_ = oh_i_t0[5] & oh_i[4];
assign _0405_ = oh_i_t0[7] & oh_i[6];
assign _0408_ = oh_i_t0[9] & oh_i[8];
assign _0411_ = oh_i_t0[11] & oh_i[10];
assign _0414_ = oh_i_t0[13] & oh_i[12];
assign _0417_ = oh_i_t0[15] & oh_i[14];
assign _0420_ = oh_i_t0[17] & oh_i[16];
assign _0423_ = oh_i_t0[19] & oh_i[18];
assign _0426_ = oh_i_t0[21] & oh_i[20];
assign _0429_ = oh_i_t0[23] & oh_i[22];
assign _0432_ = oh_i_t0[25] & oh_i[24];
assign _0435_ = oh_i_t0[27] & oh_i[26];
assign _0438_ = oh_i_t0[29] & oh_i[28];
assign _0441_ = oh_i_t0[31] & oh_i[30];
assign _0444_ = or_tree_t0[2] & or_tree[1];
assign _0447_ = or_tree_t0[4] & or_tree[3];
assign _0450_ = or_tree_t0[6] & or_tree[5];
assign _0453_ = or_tree_t0[8] & or_tree[7];
assign _0456_ = or_tree_t0[10] & or_tree[9];
assign _0459_ = or_tree_t0[12] & or_tree[11];
assign _0462_ = or_tree_t0[14] & or_tree[13];
assign _0465_ = or_tree_t0[16] & or_tree[15];
assign _0190_ = addr_i_t0[1] & and_tree_t0[17];
assign _0193_ = addr_i_t0[1] & and_tree_t0[18];
assign _0196_ = addr_i_t0[1] & and_tree_t0[19];
assign _0199_ = addr_i_t0[1] & and_tree_t0[20];
assign _0202_ = addr_i_t0[1] & and_tree_t0[21];
assign _0205_ = addr_i_t0[1] & and_tree_t0[22];
assign _0208_ = addr_i_t0[1] & and_tree_t0[23];
assign _0211_ = addr_i_t0[1] & and_tree_t0[24];
assign _0214_ = addr_i_t0[1] & and_tree_t0[25];
assign _0217_ = addr_i_t0[1] & and_tree_t0[26];
assign _0220_ = addr_i_t0[1] & and_tree_t0[27];
assign _0223_ = addr_i_t0[1] & and_tree_t0[28];
assign _0226_ = addr_i_t0[1] & and_tree_t0[29];
assign _0229_ = addr_i_t0[1] & and_tree_t0[30];
assign _0232_ = addr_i_t0[0] & oh_i_t0[0];
assign _0235_ = addr_i_t0[0] & oh_i_t0[1];
assign _0238_ = addr_i_t0[0] & oh_i_t0[2];
assign _0241_ = addr_i_t0[0] & oh_i_t0[3];
assign _0244_ = addr_i_t0[0] & oh_i_t0[4];
assign _0247_ = addr_i_t0[0] & oh_i_t0[5];
assign _0250_ = addr_i_t0[0] & oh_i_t0[6];
assign _0253_ = addr_i_t0[0] & oh_i_t0[7];
assign _0256_ = addr_i_t0[0] & oh_i_t0[8];
assign _0259_ = addr_i_t0[0] & oh_i_t0[9];
assign _0262_ = addr_i_t0[0] & oh_i_t0[10];
assign _0265_ = addr_i_t0[0] & oh_i_t0[11];
assign _0268_ = addr_i_t0[0] & oh_i_t0[12];
assign _0271_ = addr_i_t0[0] & oh_i_t0[13];
assign _0274_ = addr_i_t0[0] & oh_i_t0[14];
assign _0277_ = addr_i_t0[0] & oh_i_t0[15];
assign _0280_ = addr_i_t0[0] & oh_i_t0[16];
assign _0283_ = addr_i_t0[0] & oh_i_t0[17];
assign _0286_ = addr_i_t0[0] & oh_i_t0[18];
assign _0289_ = addr_i_t0[0] & oh_i_t0[19];
assign _0292_ = addr_i_t0[0] & oh_i_t0[20];
assign _0295_ = addr_i_t0[0] & oh_i_t0[21];
assign _0298_ = addr_i_t0[0] & oh_i_t0[22];
assign _0301_ = addr_i_t0[0] & oh_i_t0[23];
assign _0304_ = addr_i_t0[0] & oh_i_t0[24];
assign _0307_ = addr_i_t0[0] & oh_i_t0[25];
assign _0310_ = addr_i_t0[0] & oh_i_t0[26];
assign _0313_ = addr_i_t0[0] & oh_i_t0[27];
assign _0316_ = addr_i_t0[0] & oh_i_t0[28];
assign _0319_ = addr_i_t0[0] & oh_i_t0[29];
assign _0322_ = addr_i_t0[0] & oh_i_t0[30];
assign _0325_ = addr_i_t0[0] & oh_i_t0[31];
assign _0328_ = addr_i_t0[4] & and_tree_t0[1];
assign _0331_ = addr_i_t0[4] & and_tree_t0[2];
assign _0334_ = addr_i_t0[3] & and_tree_t0[3];
assign _0337_ = addr_i_t0[3] & and_tree_t0[4];
assign _0340_ = addr_i_t0[3] & and_tree_t0[5];
assign _0343_ = addr_i_t0[3] & and_tree_t0[6];
assign _0346_ = addr_i_t0[2] & and_tree_t0[7];
assign _0349_ = addr_i_t0[2] & and_tree_t0[8];
assign _0352_ = addr_i_t0[2] & and_tree_t0[9];
assign _0355_ = addr_i_t0[2] & and_tree_t0[10];
assign _0358_ = addr_i_t0[2] & and_tree_t0[11];
assign _0361_ = addr_i_t0[2] & and_tree_t0[12];
assign _0364_ = addr_i_t0[2] & and_tree_t0[13];
assign _0367_ = addr_i_t0[2] & and_tree_t0[14];
assign _0370_ = addr_i_t0[1] & and_tree_t0[15];
assign _0373_ = addr_i_t0[1] & and_tree_t0[16];
assign _0376_ = or_tree_t0[17] & or_tree_t0[18];
assign _0379_ = or_tree_t0[19] & or_tree_t0[20];
assign _0382_ = or_tree_t0[21] & or_tree_t0[22];
assign _0385_ = or_tree_t0[23] & or_tree_t0[24];
assign _0388_ = or_tree_t0[25] & or_tree_t0[26];
assign _0391_ = or_tree_t0[27] & or_tree_t0[28];
assign _0394_ = or_tree_t0[29] & or_tree_t0[30];
assign _0397_ = oh_i_t0[0] & oh_i_t0[1];
assign _0400_ = oh_i_t0[2] & oh_i_t0[3];
assign _0403_ = oh_i_t0[4] & oh_i_t0[5];
assign _0406_ = oh_i_t0[6] & oh_i_t0[7];
assign _0409_ = oh_i_t0[8] & oh_i_t0[9];
assign _0412_ = oh_i_t0[10] & oh_i_t0[11];
assign _0415_ = oh_i_t0[12] & oh_i_t0[13];
assign _0418_ = oh_i_t0[14] & oh_i_t0[15];
assign _0421_ = oh_i_t0[16] & oh_i_t0[17];
assign _0424_ = oh_i_t0[18] & oh_i_t0[19];
assign _0427_ = oh_i_t0[20] & oh_i_t0[21];
assign _0430_ = oh_i_t0[22] & oh_i_t0[23];
assign _0433_ = oh_i_t0[24] & oh_i_t0[25];
assign _0436_ = oh_i_t0[26] & oh_i_t0[27];
assign _0439_ = oh_i_t0[28] & oh_i_t0[29];
assign _0442_ = oh_i_t0[30] & oh_i_t0[31];
assign _0445_ = or_tree_t0[1] & or_tree_t0[2];
assign _0448_ = or_tree_t0[3] & or_tree_t0[4];
assign _0451_ = or_tree_t0[5] & or_tree_t0[6];
assign _0454_ = or_tree_t0[7] & or_tree_t0[8];
assign _0457_ = or_tree_t0[9] & or_tree_t0[10];
assign _0460_ = or_tree_t0[11] & or_tree_t0[12];
assign _0463_ = or_tree_t0[13] & or_tree_t0[14];
assign _0466_ = or_tree_t0[15] & or_tree_t0[16];
assign _0718_ = _0188_ | _0189_;
assign _0719_ = _0191_ | _0192_;
assign _0720_ = _0194_ | _0195_;
assign _0721_ = _0197_ | _0198_;
assign _0722_ = _0200_ | _0201_;
assign _0723_ = _0203_ | _0204_;
assign _0724_ = _0206_ | _0207_;
assign _0725_ = _0209_ | _0210_;
assign _0726_ = _0212_ | _0213_;
assign _0727_ = _0215_ | _0216_;
assign _0728_ = _0218_ | _0219_;
assign _0729_ = _0221_ | _0222_;
assign _0730_ = _0224_ | _0225_;
assign _0731_ = _0227_ | _0228_;
assign _0732_ = _0230_ | _0231_;
assign _0733_ = _0233_ | _0234_;
assign _0734_ = _0236_ | _0237_;
assign _0735_ = _0239_ | _0240_;
assign _0736_ = _0242_ | _0243_;
assign _0737_ = _0245_ | _0246_;
assign _0738_ = _0248_ | _0249_;
assign _0739_ = _0251_ | _0252_;
assign _0740_ = _0254_ | _0255_;
assign _0741_ = _0257_ | _0258_;
assign _0742_ = _0260_ | _0261_;
assign _0743_ = _0263_ | _0264_;
assign _0744_ = _0266_ | _0267_;
assign _0745_ = _0269_ | _0270_;
assign _0746_ = _0272_ | _0273_;
assign _0747_ = _0275_ | _0276_;
assign _0748_ = _0278_ | _0279_;
assign _0749_ = _0281_ | _0282_;
assign _0750_ = _0284_ | _0285_;
assign _0751_ = _0287_ | _0288_;
assign _0752_ = _0290_ | _0291_;
assign _0753_ = _0293_ | _0294_;
assign _0754_ = _0296_ | _0297_;
assign _0755_ = _0299_ | _0300_;
assign _0756_ = _0302_ | _0303_;
assign _0757_ = _0305_ | _0306_;
assign _0758_ = _0308_ | _0309_;
assign _0759_ = _0311_ | _0312_;
assign _0760_ = _0314_ | _0315_;
assign _0761_ = _0317_ | _0318_;
assign _0762_ = _0320_ | _0321_;
assign _0763_ = _0323_ | _0324_;
assign _0764_ = _0326_ | _0327_;
assign _0765_ = _0329_ | _0330_;
assign _0766_ = _0332_ | _0333_;
assign _0767_ = _0335_ | _0336_;
assign _0768_ = _0338_ | _0339_;
assign _0769_ = _0341_ | _0342_;
assign _0770_ = _0344_ | _0345_;
assign _0771_ = _0347_ | _0348_;
assign _0772_ = _0350_ | _0351_;
assign _0773_ = _0353_ | _0354_;
assign _0774_ = _0356_ | _0357_;
assign _0775_ = _0359_ | _0360_;
assign _0776_ = _0362_ | _0363_;
assign _0777_ = _0365_ | _0366_;
assign _0778_ = _0368_ | _0369_;
assign _0779_ = _0371_ | _0372_;
assign _0780_ = _0374_ | _0375_;
assign _0781_ = _0377_ | _0378_;
assign _0782_ = _0380_ | _0381_;
assign _0783_ = _0383_ | _0384_;
assign _0784_ = _0386_ | _0387_;
assign _0785_ = _0389_ | _0390_;
assign _0786_ = _0392_ | _0393_;
assign _0787_ = _0395_ | _0396_;
assign _0788_ = _0398_ | _0399_;
assign _0789_ = _0401_ | _0402_;
assign _0790_ = _0404_ | _0405_;
assign _0791_ = _0407_ | _0408_;
assign _0792_ = _0410_ | _0411_;
assign _0793_ = _0413_ | _0414_;
assign _0794_ = _0416_ | _0417_;
assign _0795_ = _0419_ | _0420_;
assign _0796_ = _0422_ | _0423_;
assign _0797_ = _0425_ | _0426_;
assign _0798_ = _0428_ | _0429_;
assign _0799_ = _0431_ | _0432_;
assign _0800_ = _0434_ | _0435_;
assign _0801_ = _0437_ | _0438_;
assign _0802_ = _0440_ | _0441_;
assign _0803_ = _0443_ | _0444_;
assign _0804_ = _0446_ | _0447_;
assign _0805_ = _0449_ | _0450_;
assign _0806_ = _0452_ | _0453_;
assign _0807_ = _0455_ | _0456_;
assign _0808_ = _0458_ | _0459_;
assign _0809_ = _0461_ | _0462_;
assign _0810_ = _0464_ | _0465_;
assign _0906_ = _0718_ | _0190_;
assign _0908_ = _0719_ | _0193_;
assign _0910_ = _0720_ | _0196_;
assign _0912_ = _0721_ | _0199_;
assign _0914_ = _0722_ | _0202_;
assign _0916_ = _0723_ | _0205_;
assign _0918_ = _0724_ | _0208_;
assign _0920_ = _0725_ | _0211_;
assign _0922_ = _0726_ | _0214_;
assign _0924_ = _0727_ | _0217_;
assign _0926_ = _0728_ | _0220_;
assign _0928_ = _0729_ | _0223_;
assign _0930_ = _0730_ | _0226_;
assign _0932_ = _0731_ | _0229_;
assign _0934_ = _0732_ | _0232_;
assign _0936_ = _0733_ | _0235_;
assign _0938_ = _0734_ | _0238_;
assign _0940_ = _0735_ | _0241_;
assign _0942_ = _0736_ | _0244_;
assign _0944_ = _0737_ | _0247_;
assign _0946_ = _0738_ | _0250_;
assign _0948_ = _0739_ | _0253_;
assign _0950_ = _0740_ | _0256_;
assign _0952_ = _0741_ | _0259_;
assign _0954_ = _0742_ | _0262_;
assign _0956_ = _0743_ | _0265_;
assign _0958_ = _0744_ | _0268_;
assign _0960_ = _0745_ | _0271_;
assign _0962_ = _0746_ | _0274_;
assign _0964_ = _0747_ | _0277_;
assign _0966_ = _0748_ | _0280_;
assign _0968_ = _0749_ | _0283_;
assign _0970_ = _0750_ | _0286_;
assign _0972_ = _0751_ | _0289_;
assign _0974_ = _0752_ | _0292_;
assign _0976_ = _0753_ | _0295_;
assign _0978_ = _0754_ | _0298_;
assign _0980_ = _0755_ | _0301_;
assign _0982_ = _0756_ | _0304_;
assign _0984_ = _0757_ | _0307_;
assign _0986_ = _0758_ | _0310_;
assign _0988_ = _0759_ | _0313_;
assign _0990_ = _0760_ | _0316_;
assign _0992_ = _0761_ | _0319_;
assign _0994_ = _0762_ | _0322_;
assign _0996_ = _0763_ | _0325_;
assign _0998_ = _0764_ | _0328_;
assign _1000_ = _0765_ | _0331_;
assign _1002_ = _0766_ | _0334_;
assign _1004_ = _0767_ | _0337_;
assign _1006_ = _0768_ | _0340_;
assign _1008_ = _0769_ | _0343_;
assign _1010_ = _0770_ | _0346_;
assign _1012_ = _0771_ | _0349_;
assign _1014_ = _0772_ | _0352_;
assign _1016_ = _0773_ | _0355_;
assign _1018_ = _0774_ | _0358_;
assign _1020_ = _0775_ | _0361_;
assign _1022_ = _0776_ | _0364_;
assign _1024_ = _0777_ | _0367_;
assign _1026_ = _0778_ | _0370_;
assign _1028_ = _0779_ | _0373_;
assign _1030_ = _0780_ | _0376_;
assign _1032_ = _0781_ | _0379_;
assign _1034_ = _0782_ | _0382_;
assign _1036_ = _0783_ | _0385_;
assign _1038_ = _0784_ | _0388_;
assign _1040_ = _0785_ | _0391_;
assign _1042_ = _0786_ | _0394_;
assign err_tree_t0[15] = _0787_ | _0397_;
assign err_tree_t0[16] = _0788_ | _0400_;
assign err_tree_t0[17] = _0789_ | _0403_;
assign err_tree_t0[18] = _0790_ | _0406_;
assign err_tree_t0[19] = _0791_ | _0409_;
assign err_tree_t0[20] = _0792_ | _0412_;
assign err_tree_t0[21] = _0793_ | _0415_;
assign err_tree_t0[22] = _0794_ | _0418_;
assign err_tree_t0[23] = _0795_ | _0421_;
assign err_tree_t0[24] = _0796_ | _0424_;
assign err_tree_t0[25] = _0797_ | _0427_;
assign err_tree_t0[26] = _0798_ | _0430_;
assign err_tree_t0[27] = _0799_ | _0433_;
assign err_tree_t0[28] = _0800_ | _0436_;
assign err_tree_t0[29] = _0801_ | _0439_;
assign err_tree_t0[30] = _0802_ | _0442_;
assign _1044_ = _0803_ | _0445_;
assign _1046_ = _0804_ | _0448_;
assign _1048_ = _0805_ | _0451_;
assign _1050_ = _0806_ | _0454_;
assign _1052_ = _0807_ | _0457_;
assign _1054_ = _0808_ | _0460_;
assign _1056_ = _0809_ | _0463_;
assign _1058_ = _0810_ | _0466_;
assign _0000_ = ~ or_tree[19];
assign _0001_ = ~ or_tree[21];
assign _0002_ = ~ or_tree[23];
assign _0003_ = ~ or_tree[25];
assign _0004_ = ~ or_tree[27];
assign _0005_ = ~ or_tree[29];
assign _0006_ = ~ oh_i[0];
assign _0007_ = ~ oh_i[2];
assign _0008_ = ~ oh_i[4];
assign _0009_ = ~ oh_i[6];
assign _0010_ = ~ oh_i[8];
assign _0011_ = ~ oh_i[10];
assign _0012_ = ~ oh_i[12];
assign _0013_ = ~ oh_i[14];
assign _0014_ = ~ oh_i[16];
assign _0015_ = ~ oh_i[18];
assign _0016_ = ~ oh_i[20];
assign _0017_ = ~ oh_i[22];
assign _0018_ = ~ oh_i[24];
assign _0019_ = ~ oh_i[26];
assign _0020_ = ~ oh_i[28];
assign _0021_ = ~ oh_i[30];
assign _0022_ = ~ or_tree[1];
assign _0023_ = ~ or_tree[3];
assign _0024_ = ~ or_tree[5];
assign _0025_ = ~ or_tree[7];
assign _0026_ = ~ or_tree[9];
assign _0027_ = ~ or_tree[11];
assign _0028_ = ~ or_tree[13];
assign _0029_ = ~ or_tree[15];
assign _0030_ = ~ or_tree[17];
assign _0031_ = ~ _0905_;
assign _0032_ = ~ _0909_;
assign _0033_ = ~ _0913_;
assign _0034_ = ~ _0917_;
assign _0035_ = ~ _0921_;
assign _0036_ = ~ _0925_;
assign _0037_ = ~ _0929_;
assign _0038_ = ~ _0933_;
assign _0039_ = ~ _0937_;
assign _0040_ = ~ _0941_;
assign _0041_ = ~ _0945_;
assign _0042_ = ~ _0949_;
assign _0043_ = ~ _0953_;
assign _0044_ = ~ _0957_;
assign _0045_ = ~ _0961_;
assign _0046_ = ~ _0965_;
assign _0047_ = ~ _0969_;
assign _0048_ = ~ _0973_;
assign _0049_ = ~ _0977_;
assign _0050_ = ~ _0981_;
assign _0051_ = ~ _0985_;
assign _0052_ = ~ _0989_;
assign _0053_ = ~ _0993_;
assign _0054_ = ~ _0997_;
assign _0055_ = ~ _1001_;
assign _0056_ = ~ _1005_;
assign _0057_ = ~ _1009_;
assign _0058_ = ~ _1013_;
assign _0059_ = ~ _1017_;
assign _0060_ = ~ _1021_;
assign _0061_ = ~ _1025_;
assign _0062_ = ~ _1029_;
assign _0063_ = ~ _1064_;
assign _0064_ = ~ _1031_;
assign _0065_ = ~ _1066_;
assign _0066_ = ~ _1033_;
assign _0067_ = ~ _1068_;
assign _0068_ = ~ _1035_;
assign _0069_ = ~ _1070_;
assign _0070_ = ~ _1037_;
assign _0071_ = ~ _1072_;
assign _0072_ = ~ _1039_;
assign _0073_ = ~ _1074_;
assign _0074_ = ~ _1041_;
assign _0075_ = ~ _1076_;
assign _0076_ = ~ _1043_;
assign _0077_ = ~ _1078_;
assign _0078_ = ~ _1045_;
assign _0079_ = ~ _1080_;
assign _0080_ = ~ _1047_;
assign _0081_ = ~ _1082_;
assign _0082_ = ~ _1049_;
assign _0083_ = ~ _1084_;
assign _0084_ = ~ _1051_;
assign _0085_ = ~ _1086_;
assign _0086_ = ~ _1053_;
assign _0087_ = ~ _1088_;
assign _0088_ = ~ _1055_;
assign _0089_ = ~ _1090_;
assign _0090_ = ~ _1057_;
assign _0091_ = ~ _1092_;
assign _0092_ = ~ oh0_err;
assign _0093_ = ~ _1094_;
assign _0094_ = ~ or_tree[20];
assign _0095_ = ~ or_tree[22];
assign _0096_ = ~ or_tree[24];
assign _0097_ = ~ or_tree[26];
assign _0098_ = ~ or_tree[28];
assign _0099_ = ~ or_tree[30];
assign _0100_ = ~ oh_i[1];
assign _0101_ = ~ oh_i[3];
assign _0102_ = ~ oh_i[5];
assign _0103_ = ~ oh_i[7];
assign _0104_ = ~ oh_i[9];
assign _0105_ = ~ oh_i[11];
assign _0106_ = ~ oh_i[13];
assign _0107_ = ~ oh_i[15];
assign _0108_ = ~ oh_i[17];
assign _0109_ = ~ oh_i[19];
assign _0110_ = ~ oh_i[21];
assign _0111_ = ~ oh_i[23];
assign _0112_ = ~ oh_i[25];
assign _0113_ = ~ oh_i[27];
assign _0114_ = ~ oh_i[29];
assign _0115_ = ~ oh_i[31];
assign _0116_ = ~ or_tree[2];
assign _0117_ = ~ or_tree[4];
assign _0118_ = ~ or_tree[6];
assign _0119_ = ~ or_tree[8];
assign _0120_ = ~ or_tree[10];
assign _0121_ = ~ or_tree[12];
assign _0122_ = ~ or_tree[14];
assign _0123_ = ~ or_tree[16];
assign _0124_ = ~ or_tree[18];
assign _0125_ = ~ _0907_;
assign _0126_ = ~ _0911_;
assign _0127_ = ~ _0915_;
assign _0128_ = ~ _0919_;
assign _0129_ = ~ _0923_;
assign _0130_ = ~ _0927_;
assign _0131_ = ~ _0931_;
assign _0132_ = ~ _0935_;
assign _0133_ = ~ _0939_;
assign _0134_ = ~ _0943_;
assign _0135_ = ~ _0947_;
assign _0136_ = ~ _0951_;
assign _0137_ = ~ _0955_;
assign _0138_ = ~ _0959_;
assign _0139_ = ~ _0963_;
assign _0140_ = ~ _0967_;
assign _0141_ = ~ _0971_;
assign _0142_ = ~ _0975_;
assign _0143_ = ~ _0979_;
assign _0144_ = ~ _0983_;
assign _0145_ = ~ _0987_;
assign _0146_ = ~ _0991_;
assign _0147_ = ~ _0995_;
assign _0148_ = ~ _0999_;
assign _0149_ = ~ _1003_;
assign _0150_ = ~ _1007_;
assign _0151_ = ~ _1011_;
assign _0152_ = ~ _1015_;
assign _0153_ = ~ _1019_;
assign _0154_ = ~ _1023_;
assign _0155_ = ~ _1027_;
assign _0156_ = ~ err_tree[17];
assign _0157_ = ~ err_tree[18];
assign _0158_ = ~ err_tree[19];
assign _0159_ = ~ err_tree[20];
assign _0160_ = ~ err_tree[21];
assign _0161_ = ~ err_tree[22];
assign _0162_ = ~ err_tree[23];
assign _0163_ = ~ err_tree[24];
assign _0164_ = ~ err_tree[25];
assign _0165_ = ~ err_tree[26];
assign _0166_ = ~ err_tree[27];
assign _0167_ = ~ err_tree[28];
assign _0168_ = ~ err_tree[29];
assign _0169_ = ~ err_tree[30];
assign _0170_ = ~ err_tree[1];
assign _0171_ = ~ err_tree[2];
assign _0172_ = ~ err_tree[3];
assign _0173_ = ~ err_tree[4];
assign _0174_ = ~ err_tree[5];
assign _0175_ = ~ err_tree[6];
assign _0176_ = ~ err_tree[7];
assign _0177_ = ~ err_tree[8];
assign _0178_ = ~ err_tree[9];
assign _0179_ = ~ err_tree[10];
assign _0180_ = ~ err_tree[11];
assign _0181_ = ~ err_tree[12];
assign _0182_ = ~ err_tree[13];
assign _0183_ = ~ err_tree[14];
assign _0184_ = ~ err_tree[15];
assign _0185_ = ~ err_tree[16];
assign _0186_ = ~ enable_err;
assign _0187_ = ~ addr_err;
assign _0467_ = or_tree_t0[19] & _0094_;
assign _0469_ = or_tree_t0[21] & _0095_;
assign _0471_ = or_tree_t0[23] & _0096_;
assign _0473_ = or_tree_t0[25] & _0097_;
assign _0475_ = or_tree_t0[27] & _0098_;
assign _0477_ = or_tree_t0[29] & _0099_;
assign _0479_ = oh_i_t0[0] & _0100_;
assign _0481_ = oh_i_t0[2] & _0101_;
assign _0483_ = oh_i_t0[4] & _0102_;
assign _0485_ = oh_i_t0[6] & _0103_;
assign _0487_ = oh_i_t0[8] & _0104_;
assign _0489_ = oh_i_t0[10] & _0105_;
assign _0491_ = oh_i_t0[12] & _0106_;
assign _0493_ = oh_i_t0[14] & _0107_;
assign _0495_ = oh_i_t0[16] & _0108_;
assign _0497_ = oh_i_t0[18] & _0109_;
assign _0499_ = oh_i_t0[20] & _0110_;
assign _0501_ = oh_i_t0[22] & _0111_;
assign _0503_ = oh_i_t0[24] & _0112_;
assign _0505_ = oh_i_t0[26] & _0113_;
assign _0507_ = oh_i_t0[28] & _0114_;
assign _0509_ = oh_i_t0[30] & _0115_;
assign _0511_ = or_tree_t0[1] & _0116_;
assign _0513_ = or_tree_t0[3] & _0117_;
assign _0515_ = or_tree_t0[5] & _0118_;
assign _0517_ = or_tree_t0[7] & _0119_;
assign _0519_ = or_tree_t0[9] & _0120_;
assign _0521_ = or_tree_t0[11] & _0121_;
assign _0523_ = or_tree_t0[13] & _0122_;
assign _0525_ = or_tree_t0[15] & _0123_;
assign _0527_ = or_tree_t0[17] & _0124_;
assign _0529_ = _0906_ & _0125_;
assign _0532_ = _0910_ & _0126_;
assign _0535_ = _0914_ & _0127_;
assign _0538_ = _0918_ & _0128_;
assign _0541_ = _0922_ & _0129_;
assign _0544_ = _0926_ & _0130_;
assign _0547_ = _0930_ & _0131_;
assign _0550_ = _0934_ & _0132_;
assign _0553_ = _0938_ & _0133_;
assign _0556_ = _0942_ & _0134_;
assign _0559_ = _0946_ & _0135_;
assign _0562_ = _0950_ & _0136_;
assign _0565_ = _0954_ & _0137_;
assign _0568_ = _0958_ & _0138_;
assign _0571_ = _0962_ & _0139_;
assign _0574_ = _0966_ & _0140_;
assign _0577_ = _0970_ & _0141_;
assign _0580_ = _0974_ & _0142_;
assign _0583_ = _0978_ & _0143_;
assign _0586_ = _0982_ & _0144_;
assign _0589_ = _0986_ & _0145_;
assign _0592_ = _0990_ & _0146_;
assign _0595_ = _0994_ & _0147_;
assign _0598_ = _0998_ & _0148_;
assign _0601_ = _1002_ & _0149_;
assign _0604_ = _1006_ & _0150_;
assign _0607_ = _1010_ & _0151_;
assign _0610_ = _1014_ & _0152_;
assign _0613_ = _1018_ & _0153_;
assign _0616_ = _1022_ & _0154_;
assign _0619_ = _1026_ & _0155_;
assign _0622_ = _1030_ & _0156_;
assign _0625_ = _1065_ & _0157_;
assign _0628_ = _1032_ & _0158_;
assign _0631_ = _1067_ & _0159_;
assign _0634_ = _1034_ & _0160_;
assign _0637_ = _1069_ & _0161_;
assign _0640_ = _1036_ & _0162_;
assign _0643_ = _1071_ & _0163_;
assign _0646_ = _1038_ & _0164_;
assign _0649_ = _1073_ & _0165_;
assign _0652_ = _1040_ & _0166_;
assign _0655_ = _1075_ & _0167_;
assign _0658_ = _1042_ & _0168_;
assign _0661_ = _1077_ & _0169_;
assign _0664_ = _1044_ & _0170_;
assign _0667_ = _1079_ & _0171_;
assign _0670_ = _1046_ & _0172_;
assign _0673_ = _1081_ & _0173_;
assign _0676_ = _1048_ & _0174_;
assign _0679_ = _1083_ & _0175_;
assign _0682_ = _1050_ & _0176_;
assign _0685_ = _1085_ & _0177_;
assign _0688_ = _1052_ & _0178_;
assign _0691_ = _1087_ & _0179_;
assign _0694_ = _1054_ & _0180_;
assign _0697_ = _1089_ & _0181_;
assign _0700_ = _1056_ & _0182_;
assign _0703_ = _1091_ & _0183_;
assign _0706_ = _1058_ & _0184_;
assign _0709_ = _1093_ & _0185_;
assign _0712_ = oh0_err_t0 & _0186_;
assign _0715_ = _1095_ & _0187_;
assign _0468_ = or_tree_t0[20] & _0000_;
assign _0470_ = or_tree_t0[22] & _0001_;
assign _0472_ = or_tree_t0[24] & _0002_;
assign _0474_ = or_tree_t0[26] & _0003_;
assign _0476_ = or_tree_t0[28] & _0004_;
assign _0478_ = or_tree_t0[30] & _0005_;
assign _0480_ = oh_i_t0[1] & _0006_;
assign _0482_ = oh_i_t0[3] & _0007_;
assign _0484_ = oh_i_t0[5] & _0008_;
assign _0486_ = oh_i_t0[7] & _0009_;
assign _0488_ = oh_i_t0[9] & _0010_;
assign _0490_ = oh_i_t0[11] & _0011_;
assign _0492_ = oh_i_t0[13] & _0012_;
assign _0494_ = oh_i_t0[15] & _0013_;
assign _0496_ = oh_i_t0[17] & _0014_;
assign _0498_ = oh_i_t0[19] & _0015_;
assign _0500_ = oh_i_t0[21] & _0016_;
assign _0502_ = oh_i_t0[23] & _0017_;
assign _0504_ = oh_i_t0[25] & _0018_;
assign _0506_ = oh_i_t0[27] & _0019_;
assign _0508_ = oh_i_t0[29] & _0020_;
assign _0510_ = oh_i_t0[31] & _0021_;
assign _0512_ = or_tree_t0[2] & _0022_;
assign _0514_ = or_tree_t0[4] & _0023_;
assign _0516_ = or_tree_t0[6] & _0024_;
assign _0518_ = or_tree_t0[8] & _0025_;
assign _0520_ = or_tree_t0[10] & _0026_;
assign _0522_ = or_tree_t0[12] & _0027_;
assign _0524_ = or_tree_t0[14] & _0028_;
assign _0526_ = or_tree_t0[16] & _0029_;
assign _0528_ = or_tree_t0[18] & _0030_;
assign _0530_ = _0908_ & _0031_;
assign _0533_ = _0912_ & _0032_;
assign _0536_ = _0916_ & _0033_;
assign _0539_ = _0920_ & _0034_;
assign _0542_ = _0924_ & _0035_;
assign _0545_ = _0928_ & _0036_;
assign _0548_ = _0932_ & _0037_;
assign _0551_ = _0936_ & _0038_;
assign _0554_ = _0940_ & _0039_;
assign _0557_ = _0944_ & _0040_;
assign _0560_ = _0948_ & _0041_;
assign _0563_ = _0952_ & _0042_;
assign _0566_ = _0956_ & _0043_;
assign _0569_ = _0960_ & _0044_;
assign _0572_ = _0964_ & _0045_;
assign _0575_ = _0968_ & _0046_;
assign _0578_ = _0972_ & _0047_;
assign _0581_ = _0976_ & _0048_;
assign _0584_ = _0980_ & _0049_;
assign _0587_ = _0984_ & _0050_;
assign _0590_ = _0988_ & _0051_;
assign _0593_ = _0992_ & _0052_;
assign _0596_ = _0996_ & _0053_;
assign _0599_ = _1000_ & _0054_;
assign _0602_ = _1004_ & _0055_;
assign _0605_ = _1008_ & _0056_;
assign _0608_ = _1012_ & _0057_;
assign _0611_ = _1016_ & _0058_;
assign _0614_ = _1020_ & _0059_;
assign _0617_ = _1024_ & _0060_;
assign _0620_ = _1028_ & _0061_;
assign _0623_ = err_tree_t0[17] & _0062_;
assign _0626_ = err_tree_t0[18] & _0063_;
assign _0629_ = err_tree_t0[19] & _0064_;
assign _0632_ = err_tree_t0[20] & _0065_;
assign _0635_ = err_tree_t0[21] & _0066_;
assign _0638_ = err_tree_t0[22] & _0067_;
assign _0641_ = err_tree_t0[23] & _0068_;
assign _0644_ = err_tree_t0[24] & _0069_;
assign _0647_ = err_tree_t0[25] & _0070_;
assign _0650_ = err_tree_t0[26] & _0071_;
assign _0653_ = err_tree_t0[27] & _0072_;
assign _0656_ = err_tree_t0[28] & _0073_;
assign _0659_ = err_tree_t0[29] & _0074_;
assign _0662_ = err_tree_t0[30] & _0075_;
assign _0665_ = err_tree_t0[1] & _0076_;
assign _0668_ = err_tree_t0[2] & _0077_;
assign _0671_ = err_tree_t0[3] & _0078_;
assign _0674_ = err_tree_t0[4] & _0079_;
assign _0677_ = err_tree_t0[5] & _0080_;
assign _0680_ = err_tree_t0[6] & _0081_;
assign _0683_ = err_tree_t0[7] & _0082_;
assign _0686_ = err_tree_t0[8] & _0083_;
assign _0689_ = err_tree_t0[9] & _0084_;
assign _0692_ = err_tree_t0[10] & _0085_;
assign _0695_ = err_tree_t0[11] & _0086_;
assign _0698_ = err_tree_t0[12] & _0087_;
assign _0701_ = err_tree_t0[13] & _0088_;
assign _0704_ = err_tree_t0[14] & _0089_;
assign _0707_ = err_tree_t0[15] & _0090_;
assign _0710_ = err_tree_t0[16] & _0091_;
assign _0713_ = enable_err_t0 & _0092_;
assign _0716_ = addr_err_t0 & _0093_;
assign _0531_ = _0906_ & _0908_;
assign _0534_ = _0910_ & _0912_;
assign _0537_ = _0914_ & _0916_;
assign _0540_ = _0918_ & _0920_;
assign _0543_ = _0922_ & _0924_;
assign _0546_ = _0926_ & _0928_;
assign _0549_ = _0930_ & _0932_;
assign _0552_ = _0934_ & _0936_;
assign _0555_ = _0938_ & _0940_;
assign _0558_ = _0942_ & _0944_;
assign _0561_ = _0946_ & _0948_;
assign _0564_ = _0950_ & _0952_;
assign _0567_ = _0954_ & _0956_;
assign _0570_ = _0958_ & _0960_;
assign _0573_ = _0962_ & _0964_;
assign _0576_ = _0966_ & _0968_;
assign _0579_ = _0970_ & _0972_;
assign _0582_ = _0974_ & _0976_;
assign _0585_ = _0978_ & _0980_;
assign _0588_ = _0982_ & _0984_;
assign _0591_ = _0986_ & _0988_;
assign _0594_ = _0990_ & _0992_;
assign _0597_ = _0994_ & _0996_;
assign _0600_ = _0998_ & _1000_;
assign _0603_ = _1002_ & _1004_;
assign _0606_ = _1006_ & _1008_;
assign _0609_ = _1010_ & _1012_;
assign _0612_ = _1014_ & _1016_;
assign _0615_ = _1018_ & _1020_;
assign _0618_ = _1022_ & _1024_;
assign _0621_ = _1026_ & _1028_;
assign _0624_ = _1030_ & err_tree_t0[17];
assign _0627_ = _1065_ & err_tree_t0[18];
assign _0630_ = _1032_ & err_tree_t0[19];
assign _0633_ = _1067_ & err_tree_t0[20];
assign _0636_ = _1034_ & err_tree_t0[21];
assign _0639_ = _1069_ & err_tree_t0[22];
assign _0642_ = _1036_ & err_tree_t0[23];
assign _0645_ = _1071_ & err_tree_t0[24];
assign _0648_ = _1038_ & err_tree_t0[25];
assign _0651_ = _1073_ & err_tree_t0[26];
assign _0654_ = _1040_ & err_tree_t0[27];
assign _0657_ = _1075_ & err_tree_t0[28];
assign _0660_ = _1042_ & err_tree_t0[29];
assign _0663_ = _1077_ & err_tree_t0[30];
assign _0666_ = _1044_ & err_tree_t0[1];
assign _0669_ = _1079_ & err_tree_t0[2];
assign _0672_ = _1046_ & err_tree_t0[3];
assign _0675_ = _1081_ & err_tree_t0[4];
assign _0678_ = _1048_ & err_tree_t0[5];
assign _0681_ = _1083_ & err_tree_t0[6];
assign _0684_ = _1050_ & err_tree_t0[7];
assign _0687_ = _1085_ & err_tree_t0[8];
assign _0690_ = _1052_ & err_tree_t0[9];
assign _0693_ = _1087_ & err_tree_t0[10];
assign _0696_ = _1054_ & err_tree_t0[11];
assign _0699_ = _1089_ & err_tree_t0[12];
assign _0702_ = _1056_ & err_tree_t0[13];
assign _0705_ = _1091_ & err_tree_t0[14];
assign _0708_ = _1058_ & err_tree_t0[15];
assign _0711_ = _1093_ & err_tree_t0[16];
assign _0714_ = oh0_err_t0 & enable_err_t0;
assign _0717_ = _1095_ & addr_err_t0;
assign _0811_ = _0467_ | _0468_;
assign _0812_ = _0469_ | _0470_;
assign _0813_ = _0471_ | _0472_;
assign _0814_ = _0473_ | _0474_;
assign _0815_ = _0475_ | _0476_;
assign _0816_ = _0477_ | _0478_;
assign _0817_ = _0479_ | _0480_;
assign _0818_ = _0481_ | _0482_;
assign _0819_ = _0483_ | _0484_;
assign _0820_ = _0485_ | _0486_;
assign _0821_ = _0487_ | _0488_;
assign _0822_ = _0489_ | _0490_;
assign _0823_ = _0491_ | _0492_;
assign _0824_ = _0493_ | _0494_;
assign _0825_ = _0495_ | _0496_;
assign _0826_ = _0497_ | _0498_;
assign _0827_ = _0499_ | _0500_;
assign _0828_ = _0501_ | _0502_;
assign _0829_ = _0503_ | _0504_;
assign _0830_ = _0505_ | _0506_;
assign _0831_ = _0507_ | _0508_;
assign _0832_ = _0509_ | _0510_;
assign _0833_ = _0511_ | _0512_;
assign _0834_ = _0513_ | _0514_;
assign _0835_ = _0515_ | _0516_;
assign _0836_ = _0517_ | _0518_;
assign _0837_ = _0519_ | _0520_;
assign _0838_ = _0521_ | _0522_;
assign _0839_ = _0523_ | _0524_;
assign _0840_ = _0525_ | _0526_;
assign _0841_ = _0527_ | _0528_;
assign _0842_ = _0529_ | _0530_;
assign _0843_ = _0532_ | _0533_;
assign _0844_ = _0535_ | _0536_;
assign _0845_ = _0538_ | _0539_;
assign _0846_ = _0541_ | _0542_;
assign _0847_ = _0544_ | _0545_;
assign _0848_ = _0547_ | _0548_;
assign _0849_ = _0550_ | _0551_;
assign _0850_ = _0553_ | _0554_;
assign _0851_ = _0556_ | _0557_;
assign _0852_ = _0559_ | _0560_;
assign _0853_ = _0562_ | _0563_;
assign _0854_ = _0565_ | _0566_;
assign _0855_ = _0568_ | _0569_;
assign _0856_ = _0571_ | _0572_;
assign _0857_ = _0574_ | _0575_;
assign _0858_ = _0577_ | _0578_;
assign _0859_ = _0580_ | _0581_;
assign _0860_ = _0583_ | _0584_;
assign _0861_ = _0586_ | _0587_;
assign _0862_ = _0589_ | _0590_;
assign _0863_ = _0592_ | _0593_;
assign _0864_ = _0595_ | _0596_;
assign _0865_ = _0598_ | _0599_;
assign _0866_ = _0601_ | _0602_;
assign _0867_ = _0604_ | _0605_;
assign _0868_ = _0607_ | _0608_;
assign _0869_ = _0610_ | _0611_;
assign _0870_ = _0613_ | _0614_;
assign _0871_ = _0616_ | _0617_;
assign _0872_ = _0619_ | _0620_;
assign _0873_ = _0622_ | _0623_;
assign _0874_ = _0625_ | _0626_;
assign _0875_ = _0628_ | _0629_;
assign _0876_ = _0631_ | _0632_;
assign _0877_ = _0634_ | _0635_;
assign _0878_ = _0637_ | _0638_;
assign _0879_ = _0640_ | _0641_;
assign _0880_ = _0643_ | _0644_;
assign _0881_ = _0646_ | _0647_;
assign _0882_ = _0649_ | _0650_;
assign _0883_ = _0652_ | _0653_;
assign _0884_ = _0655_ | _0656_;
assign _0885_ = _0658_ | _0659_;
assign _0886_ = _0661_ | _0662_;
assign _0887_ = _0664_ | _0665_;
assign _0888_ = _0667_ | _0668_;
assign _0889_ = _0670_ | _0671_;
assign _0890_ = _0673_ | _0674_;
assign _0891_ = _0676_ | _0677_;
assign _0892_ = _0679_ | _0680_;
assign _0893_ = _0682_ | _0683_;
assign _0894_ = _0685_ | _0686_;
assign _0895_ = _0688_ | _0689_;
assign _0896_ = _0691_ | _0692_;
assign _0897_ = _0694_ | _0695_;
assign _0898_ = _0697_ | _0698_;
assign _0899_ = _0700_ | _0701_;
assign _0900_ = _0703_ | _0704_;
assign _0901_ = _0706_ | _0707_;
assign _0902_ = _0709_ | _0710_;
assign _0903_ = _0712_ | _0713_;
assign _0904_ = _0715_ | _0716_;
assign or_tree_t0[9] = _0811_ | _0379_;
assign or_tree_t0[10] = _0812_ | _0382_;
assign or_tree_t0[11] = _0813_ | _0385_;
assign or_tree_t0[12] = _0814_ | _0388_;
assign or_tree_t0[13] = _0815_ | _0391_;
assign or_tree_t0[14] = _0816_ | _0394_;
assign or_tree_t0[15] = _0817_ | _0397_;
assign or_tree_t0[16] = _0818_ | _0400_;
assign or_tree_t0[17] = _0819_ | _0403_;
assign or_tree_t0[18] = _0820_ | _0406_;
assign or_tree_t0[19] = _0821_ | _0409_;
assign or_tree_t0[20] = _0822_ | _0412_;
assign or_tree_t0[21] = _0823_ | _0415_;
assign or_tree_t0[22] = _0824_ | _0418_;
assign or_tree_t0[23] = _0825_ | _0421_;
assign or_tree_t0[24] = _0826_ | _0424_;
assign or_tree_t0[25] = _0827_ | _0427_;
assign or_tree_t0[26] = _0828_ | _0430_;
assign or_tree_t0[27] = _0829_ | _0433_;
assign or_tree_t0[28] = _0830_ | _0436_;
assign or_tree_t0[29] = _0831_ | _0439_;
assign or_tree_t0[30] = _0832_ | _0442_;
assign or_tree_t0[0] = _0833_ | _0445_;
assign or_tree_t0[1] = _0834_ | _0448_;
assign or_tree_t0[2] = _0835_ | _0451_;
assign or_tree_t0[3] = _0836_ | _0454_;
assign or_tree_t0[4] = _0837_ | _0457_;
assign or_tree_t0[5] = _0838_ | _0460_;
assign or_tree_t0[6] = _0839_ | _0463_;
assign or_tree_t0[7] = _0840_ | _0466_;
assign or_tree_t0[8] = _0841_ | _0376_;
assign and_tree_t0[8] = _0842_ | _0531_;
assign and_tree_t0[9] = _0843_ | _0534_;
assign and_tree_t0[10] = _0844_ | _0537_;
assign and_tree_t0[11] = _0845_ | _0540_;
assign and_tree_t0[12] = _0846_ | _0543_;
assign and_tree_t0[13] = _0847_ | _0546_;
assign and_tree_t0[14] = _0848_ | _0549_;
assign and_tree_t0[15] = _0849_ | _0552_;
assign and_tree_t0[16] = _0850_ | _0555_;
assign and_tree_t0[17] = _0851_ | _0558_;
assign and_tree_t0[18] = _0852_ | _0561_;
assign and_tree_t0[19] = _0853_ | _0564_;
assign and_tree_t0[20] = _0854_ | _0567_;
assign and_tree_t0[21] = _0855_ | _0570_;
assign and_tree_t0[22] = _0856_ | _0573_;
assign and_tree_t0[23] = _0857_ | _0576_;
assign and_tree_t0[24] = _0858_ | _0579_;
assign and_tree_t0[25] = _0859_ | _0582_;
assign and_tree_t0[26] = _0860_ | _0585_;
assign and_tree_t0[27] = _0861_ | _0588_;
assign and_tree_t0[28] = _0862_ | _0591_;
assign and_tree_t0[29] = _0863_ | _0594_;
assign and_tree_t0[30] = _0864_ | _0597_;
assign and_tree_t0[0] = _0865_ | _0600_;
assign and_tree_t0[1] = _0866_ | _0603_;
assign and_tree_t0[2] = _0867_ | _0606_;
assign and_tree_t0[3] = _0868_ | _0609_;
assign and_tree_t0[4] = _0869_ | _0612_;
assign and_tree_t0[5] = _0870_ | _0615_;
assign and_tree_t0[6] = _0871_ | _0618_;
assign and_tree_t0[7] = _0872_ | _0621_;
assign _1065_ = _0873_ | _0624_;
assign err_tree_t0[8] = _0874_ | _0627_;
assign _1067_ = _0875_ | _0630_;
assign err_tree_t0[9] = _0876_ | _0633_;
assign _1069_ = _0877_ | _0636_;
assign err_tree_t0[10] = _0878_ | _0639_;
assign _1071_ = _0879_ | _0642_;
assign err_tree_t0[11] = _0880_ | _0645_;
assign _1073_ = _0881_ | _0648_;
assign err_tree_t0[12] = _0882_ | _0651_;
assign _1075_ = _0883_ | _0654_;
assign err_tree_t0[13] = _0884_ | _0657_;
assign _1077_ = _0885_ | _0660_;
assign err_tree_t0[14] = _0886_ | _0663_;
assign _1079_ = _0887_ | _0666_;
assign oh0_err_t0 = _0888_ | _0669_;
assign _1081_ = _0889_ | _0672_;
assign err_tree_t0[1] = _0890_ | _0675_;
assign _1083_ = _0891_ | _0678_;
assign err_tree_t0[2] = _0892_ | _0681_;
assign _1085_ = _0893_ | _0684_;
assign err_tree_t0[3] = _0894_ | _0687_;
assign _1087_ = _0895_ | _0690_;
assign err_tree_t0[4] = _0896_ | _0693_;
assign _1089_ = _0897_ | _0696_;
assign err_tree_t0[5] = _0898_ | _0699_;
assign _1091_ = _0899_ | _0702_;
assign err_tree_t0[6] = _0900_ | _0705_;
assign _1093_ = _0901_ | _0708_;
assign err_tree_t0[7] = _0902_ | _0711_;
assign _1095_ = _0903_ | _0714_;
assign err_o_t0 = _0904_ | _0717_;
assign enable_err_t0 = or_tree_t0[0] | en_i_t0;
assign addr_err_t0 = or_tree_t0[0] | and_tree_t0[0];
assign _0905_ = _1059_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ and_tree[17];
assign _0907_ = addr_i[1] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ and_tree[18];
assign _0909_ = _1059_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ and_tree[19];
assign _0911_ = addr_i[1] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ and_tree[20];
assign _0913_ = _1059_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ and_tree[21];
assign _0915_ = addr_i[1] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ and_tree[22];
assign _0917_ = _1059_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ and_tree[23];
assign _0919_ = addr_i[1] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ and_tree[24];
assign _0921_ = _1059_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ and_tree[25];
assign _0923_ = addr_i[1] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ and_tree[26];
assign _0925_ = _1059_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ and_tree[27];
assign _0927_ = addr_i[1] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ and_tree[28];
assign _0929_ = _1059_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ and_tree[29];
assign _0931_ = addr_i[1] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ and_tree[30];
assign _0933_ = _1060_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ oh_i[0];
assign _0935_ = addr_i[0] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ oh_i[1];
assign _0937_ = _1060_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ oh_i[2];
assign _0939_ = addr_i[0] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ oh_i[3];
assign _0941_ = _1060_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ oh_i[4];
assign _0943_ = addr_i[0] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ oh_i[5];
assign _0945_ = _1060_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ oh_i[6];
assign _0947_ = addr_i[0] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ oh_i[7];
assign _0949_ = _1060_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ oh_i[8];
assign _0951_ = addr_i[0] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ oh_i[9];
assign _0953_ = _1060_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ oh_i[10];
assign _0955_ = addr_i[0] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ oh_i[11];
assign _0957_ = _1060_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ oh_i[12];
assign _0959_ = addr_i[0] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ oh_i[13];
assign _0961_ = _1060_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ oh_i[14];
assign _0963_ = addr_i[0] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ oh_i[15];
assign _0965_ = _1060_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ oh_i[16];
assign _0967_ = addr_i[0] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ oh_i[17];
assign _0969_ = _1060_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ oh_i[18];
assign _0971_ = addr_i[0] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ oh_i[19];
assign _0973_ = _1060_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ oh_i[20];
assign _0975_ = addr_i[0] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ oh_i[21];
assign _0977_ = _1060_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ oh_i[22];
assign _0979_ = addr_i[0] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ oh_i[23];
assign _0981_ = _1060_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ oh_i[24];
assign _0983_ = addr_i[0] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ oh_i[25];
assign _0985_ = _1060_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ oh_i[26];
assign _0987_ = addr_i[0] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ oh_i[27];
assign _0989_ = _1060_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ oh_i[28];
assign _0991_ = addr_i[0] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ oh_i[29];
assign _0993_ = _1060_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ oh_i[30];
assign _0995_ = addr_i[0] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ oh_i[31];
assign _0997_ = _1061_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ and_tree[1];
assign _0999_ = addr_i[4] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ and_tree[2];
assign _1001_ = _1062_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ and_tree[3];
assign _1003_ = addr_i[3] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ and_tree[4];
assign _1005_ = _1062_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ and_tree[5];
assign _1007_ = addr_i[3] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ and_tree[6];
assign _1009_ = _1063_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ and_tree[7];
assign _1011_ = addr_i[2] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ and_tree[8];
assign _1013_ = _1063_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ and_tree[9];
assign _1015_ = addr_i[2] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ and_tree[10];
assign _1017_ = _1063_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ and_tree[11];
assign _1019_ = addr_i[2] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ and_tree[12];
assign _1021_ = _1063_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ and_tree[13];
assign _1023_ = addr_i[2] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ and_tree[14];
assign _1025_ = _1059_ && /* src = "generated/sv2v_out.v:26484.29-26484.77" */ and_tree[15];
assign _1027_ = addr_i[1] && /* src = "generated/sv2v_out.v:26484.83-26484.130" */ and_tree[16];
assign _1029_ = or_tree[17] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ or_tree[18];
assign _1031_ = or_tree[19] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ or_tree[20];
assign _1033_ = or_tree[21] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ or_tree[22];
assign _1035_ = or_tree[23] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ or_tree[24];
assign _1037_ = or_tree[25] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ or_tree[26];
assign _1039_ = or_tree[27] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ or_tree[28];
assign _1041_ = or_tree[29] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ or_tree[30];
assign err_tree[15] = oh_i[0] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ oh_i[1];
assign err_tree[16] = oh_i[2] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ oh_i[3];
assign err_tree[17] = oh_i[4] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ oh_i[5];
assign err_tree[18] = oh_i[6] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ oh_i[7];
assign err_tree[19] = oh_i[8] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ oh_i[9];
assign err_tree[20] = oh_i[10] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ oh_i[11];
assign err_tree[21] = oh_i[12] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ oh_i[13];
assign err_tree[22] = oh_i[14] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ oh_i[15];
assign err_tree[23] = oh_i[16] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ oh_i[17];
assign err_tree[24] = oh_i[18] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ oh_i[19];
assign err_tree[25] = oh_i[20] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ oh_i[21];
assign err_tree[26] = oh_i[22] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ oh_i[23];
assign err_tree[27] = oh_i[24] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ oh_i[25];
assign err_tree[28] = oh_i[26] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ oh_i[27];
assign err_tree[29] = oh_i[28] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ oh_i[29];
assign err_tree[30] = oh_i[30] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ oh_i[31];
assign _1043_ = or_tree[1] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ or_tree[2];
assign _1045_ = or_tree[3] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ or_tree[4];
assign _1047_ = or_tree[5] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ or_tree[6];
assign _1049_ = or_tree[7] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ or_tree[8];
assign _1051_ = or_tree[9] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ or_tree[10];
assign _1053_ = or_tree[11] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ or_tree[12];
assign _1055_ = or_tree[13] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ or_tree[14];
assign _1057_ = or_tree[15] && /* src = "generated/sv2v_out.v:26485.30-26485.56" */ or_tree[16];
assign _1059_ = ! /* src = "generated/sv2v_out.v:26484.29-26484.61" */ addr_i[1];
assign _1060_ = ! /* src = "generated/sv2v_out.v:26484.29-26484.61" */ addr_i[0];
assign _1061_ = ! /* src = "generated/sv2v_out.v:26484.29-26484.61" */ addr_i[4];
assign _1062_ = ! /* src = "generated/sv2v_out.v:26484.29-26484.61" */ addr_i[3];
assign _1063_ = ! /* src = "generated/sv2v_out.v:26484.29-26484.61" */ addr_i[2];
assign or_tree[9] = or_tree[19] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ or_tree[20];
assign or_tree[10] = or_tree[21] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ or_tree[22];
assign or_tree[11] = or_tree[23] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ or_tree[24];
assign or_tree[12] = or_tree[25] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ or_tree[26];
assign or_tree[13] = or_tree[27] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ or_tree[28];
assign or_tree[14] = or_tree[29] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ or_tree[30];
assign or_tree[15] = oh_i[0] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ oh_i[1];
assign or_tree[16] = oh_i[2] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ oh_i[3];
assign or_tree[17] = oh_i[4] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ oh_i[5];
assign or_tree[18] = oh_i[6] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ oh_i[7];
assign or_tree[19] = oh_i[8] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ oh_i[9];
assign or_tree[20] = oh_i[10] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ oh_i[11];
assign or_tree[21] = oh_i[12] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ oh_i[13];
assign or_tree[22] = oh_i[14] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ oh_i[15];
assign or_tree[23] = oh_i[16] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ oh_i[17];
assign or_tree[24] = oh_i[18] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ oh_i[19];
assign or_tree[25] = oh_i[20] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ oh_i[21];
assign or_tree[26] = oh_i[22] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ oh_i[23];
assign or_tree[27] = oh_i[24] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ oh_i[25];
assign or_tree[28] = oh_i[26] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ oh_i[27];
assign or_tree[29] = oh_i[28] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ oh_i[29];
assign or_tree[30] = oh_i[30] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ oh_i[31];
assign or_tree[0] = or_tree[1] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ or_tree[2];
assign or_tree[1] = or_tree[3] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ or_tree[4];
assign or_tree[2] = or_tree[5] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ or_tree[6];
assign or_tree[3] = or_tree[7] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ or_tree[8];
assign or_tree[4] = or_tree[9] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ or_tree[10];
assign or_tree[5] = or_tree[11] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ or_tree[12];
assign or_tree[6] = or_tree[13] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ or_tree[14];
assign or_tree[7] = or_tree[15] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ or_tree[16];
assign or_tree[8] = or_tree[17] || /* src = "generated/sv2v_out.v:26483.27-26483.53" */ or_tree[18];
assign and_tree[8] = _0905_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0907_;
assign and_tree[9] = _0909_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0911_;
assign and_tree[10] = _0913_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0915_;
assign and_tree[11] = _0917_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0919_;
assign and_tree[12] = _0921_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0923_;
assign and_tree[13] = _0925_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0927_;
assign and_tree[14] = _0929_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0931_;
assign and_tree[15] = _0933_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0935_;
assign and_tree[16] = _0937_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0939_;
assign and_tree[17] = _0941_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0943_;
assign and_tree[18] = _0945_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0947_;
assign and_tree[19] = _0949_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0951_;
assign and_tree[20] = _0953_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0955_;
assign and_tree[21] = _0957_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0959_;
assign and_tree[22] = _0961_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0963_;
assign and_tree[23] = _0965_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0967_;
assign and_tree[24] = _0969_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0971_;
assign and_tree[25] = _0973_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0975_;
assign and_tree[26] = _0977_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0979_;
assign and_tree[27] = _0981_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0983_;
assign and_tree[28] = _0985_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0987_;
assign and_tree[29] = _0989_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0991_;
assign and_tree[30] = _0993_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0995_;
assign and_tree[0] = _0997_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _0999_;
assign and_tree[1] = _1001_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _1003_;
assign and_tree[2] = _1005_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _1007_;
assign and_tree[3] = _1009_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _1011_;
assign and_tree[4] = _1013_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _1015_;
assign and_tree[5] = _1017_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _1019_;
assign and_tree[6] = _1021_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _1023_;
assign and_tree[7] = _1025_ || /* src = "generated/sv2v_out.v:26484.28-26484.131" */ _1027_;
assign _1064_ = _1029_ || /* src = "generated/sv2v_out.v:26485.29-26485.73" */ err_tree[17];
assign err_tree[8] = _1064_ || /* src = "generated/sv2v_out.v:26485.28-26485.90" */ err_tree[18];
assign _1066_ = _1031_ || /* src = "generated/sv2v_out.v:26485.29-26485.73" */ err_tree[19];
assign err_tree[9] = _1066_ || /* src = "generated/sv2v_out.v:26485.28-26485.90" */ err_tree[20];
assign _1068_ = _1033_ || /* src = "generated/sv2v_out.v:26485.29-26485.73" */ err_tree[21];
assign err_tree[10] = _1068_ || /* src = "generated/sv2v_out.v:26485.28-26485.90" */ err_tree[22];
assign _1070_ = _1035_ || /* src = "generated/sv2v_out.v:26485.29-26485.73" */ err_tree[23];
assign err_tree[11] = _1070_ || /* src = "generated/sv2v_out.v:26485.28-26485.90" */ err_tree[24];
assign _1072_ = _1037_ || /* src = "generated/sv2v_out.v:26485.29-26485.73" */ err_tree[25];
assign err_tree[12] = _1072_ || /* src = "generated/sv2v_out.v:26485.28-26485.90" */ err_tree[26];
assign _1074_ = _1039_ || /* src = "generated/sv2v_out.v:26485.29-26485.73" */ err_tree[27];
assign err_tree[13] = _1074_ || /* src = "generated/sv2v_out.v:26485.28-26485.90" */ err_tree[28];
assign _1076_ = _1041_ || /* src = "generated/sv2v_out.v:26485.29-26485.73" */ err_tree[29];
assign err_tree[14] = _1076_ || /* src = "generated/sv2v_out.v:26485.28-26485.90" */ err_tree[30];
assign _1078_ = _1043_ || /* src = "generated/sv2v_out.v:26485.29-26485.73" */ err_tree[1];
assign oh0_err = _1078_ || /* src = "generated/sv2v_out.v:26485.28-26485.90" */ err_tree[2];
assign _1080_ = _1045_ || /* src = "generated/sv2v_out.v:26485.29-26485.73" */ err_tree[3];
assign err_tree[1] = _1080_ || /* src = "generated/sv2v_out.v:26485.28-26485.90" */ err_tree[4];
assign _1082_ = _1047_ || /* src = "generated/sv2v_out.v:26485.29-26485.73" */ err_tree[5];
assign err_tree[2] = _1082_ || /* src = "generated/sv2v_out.v:26485.28-26485.90" */ err_tree[6];
assign _1084_ = _1049_ || /* src = "generated/sv2v_out.v:26485.29-26485.73" */ err_tree[7];
assign err_tree[3] = _1084_ || /* src = "generated/sv2v_out.v:26485.28-26485.90" */ err_tree[8];
assign _1086_ = _1051_ || /* src = "generated/sv2v_out.v:26485.29-26485.73" */ err_tree[9];
assign err_tree[4] = _1086_ || /* src = "generated/sv2v_out.v:26485.28-26485.90" */ err_tree[10];
assign _1088_ = _1053_ || /* src = "generated/sv2v_out.v:26485.29-26485.73" */ err_tree[11];
assign err_tree[5] = _1088_ || /* src = "generated/sv2v_out.v:26485.28-26485.90" */ err_tree[12];
assign _1090_ = _1055_ || /* src = "generated/sv2v_out.v:26485.29-26485.73" */ err_tree[13];
assign err_tree[6] = _1090_ || /* src = "generated/sv2v_out.v:26485.28-26485.90" */ err_tree[14];
assign _1092_ = _1057_ || /* src = "generated/sv2v_out.v:26485.29-26485.73" */ err_tree[15];
assign err_tree[7] = _1092_ || /* src = "generated/sv2v_out.v:26485.28-26485.90" */ err_tree[16];
assign _1094_ = oh0_err || /* src = "generated/sv2v_out.v:26493.18-26493.39" */ enable_err;
assign err_o = _1094_ || /* src = "generated/sv2v_out.v:26493.17-26493.52" */ addr_err;
assign enable_err = or_tree[0] ^ /* src = "generated/sv2v_out.v:26498.25-26498.42" */ en_i;
assign addr_err = or_tree[0] ^ /* src = "generated/sv2v_out.v:26510.22-26510.46" */ and_tree[0];
assign and_tree[62:31] = oh_i;
assign and_tree_t0[62:31] = oh_i_t0;
assign { err_tree[62:31], err_tree[0] } = { 32'h00000000, oh0_err };
assign { err_tree_t0[62:31], err_tree_t0[0] } = { 32'h00000000, oh0_err_t0 };
assign or_tree[62:31] = oh_i;
assign or_tree_t0[62:31] = oh_i_t0;
endmodule

module \$paramod$9a435d8f6db004a67362aa9a56f32ea481a74dbe\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _00_;
wire [31:0] _01_;
wire [31:0] _02_;
wire [31:0] _03_;
wire [31:0] _04_;
wire [31:0] _05_;
wire [31:0] _06_;
wire [31:0] _07_;
wire [31:0] _08_;
/* src = "generated/sv2v_out.v:14871.13-14871.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14875.28-14875.37" */
output [31:0] rd_data_o;
reg [31:0] rd_data_o;
/* cellift = 32'd1 */
output [31:0] rd_data_o_t0;
reg [31:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14876.14-14876.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14872.13-14872.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14873.27-14873.36" */
input [31:0] wr_data_i;
wire [31:0] wr_data_i;
/* cellift = 32'd1 */
input [31:0] wr_data_i_t0;
wire [31:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14874.13-14874.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _00_ = ~ wr_en_i;
assign _08_ = wr_data_i ^ rd_data_o;
assign _04_ = wr_data_i_t0 | rd_data_o_t0;
assign _05_ = _08_ | _04_;
assign _01_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _02_ = { _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_ } & rd_data_o_t0;
assign _03_ = _05_ & { wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0 };
assign _06_ = _01_ | _02_;
assign _07_ = _06_ | _03_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$9a435d8f6db004a67362aa9a56f32ea481a74dbe\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 32'd0;
else rd_data_o_t0 <= _07_;
/* src = "generated/sv2v_out.v:14878.2-14882.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$9a435d8f6db004a67362aa9a56f32ea481a74dbe\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 32'd1073741827;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$a088b13b9337f1e1fba58a671f47d7c7701ffa49\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _00_;
wire [7:0] _01_;
wire [7:0] _02_;
wire [7:0] _03_;
wire [7:0] _04_;
wire [7:0] _05_;
wire [7:0] _06_;
wire [7:0] _07_;
wire [7:0] _08_;
/* src = "generated/sv2v_out.v:14871.13-14871.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14875.28-14875.37" */
output [7:0] rd_data_o;
reg [7:0] rd_data_o;
/* cellift = 32'd1 */
output [7:0] rd_data_o_t0;
reg [7:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14876.14-14876.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14872.13-14872.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14873.27-14873.36" */
input [7:0] wr_data_i;
wire [7:0] wr_data_i;
/* cellift = 32'd1 */
input [7:0] wr_data_i_t0;
wire [7:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14874.13-14874.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _00_ = ~ wr_en_i;
assign _08_ = wr_data_i ^ rd_data_o;
assign _04_ = wr_data_i_t0 | rd_data_o_t0;
assign _05_ = _08_ | _04_;
assign _01_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _02_ = { _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_ } & rd_data_o_t0;
assign _03_ = _05_ & { wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0 };
assign _06_ = _01_ | _02_;
assign _07_ = _06_ | _03_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a088b13b9337f1e1fba58a671f47d7c7701ffa49\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 8'h00;
else rd_data_o_t0 <= _07_;
/* src = "generated/sv2v_out.v:14878.2-14882.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a088b13b9337f1e1fba58a671f47d7c7701ffa49\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 8'h00;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$a308247794889ee6093207090edbf289adef8be1\ibex_ex_block (clk_i, rst_ni, alu_operator_i, alu_operand_a_i, alu_operand_b_i, alu_instr_first_cycle_i, bt_a_operand_i, bt_b_operand_i, multdiv_operator_i, mult_en_i, div_en_i, mult_sel_i, div_sel_i, multdiv_signed_mode_i, multdiv_operand_a_i, multdiv_operand_b_i, multdiv_ready_id_i, data_ind_timing_i, imd_val_we_o, imd_val_d_o, imd_val_q_i
, alu_adder_result_ex_o, result_ex_o, branch_target_o, branch_decision_o, ex_valid_o, data_ind_timing_i_t0, div_en_i_t0, div_sel_i_t0, imd_val_d_o_t0, imd_val_q_i_t0, imd_val_we_o_t0, mult_en_i_t0, mult_sel_i_t0, multdiv_ready_id_i_t0, multdiv_operand_a_i_t0, multdiv_operand_b_i_t0, alu_adder_result_ex_o_t0, alu_instr_first_cycle_i_t0, alu_operand_a_i_t0, alu_operand_b_i_t0, alu_operator_i_t0
, branch_decision_o_t0, branch_target_o_t0, bt_a_operand_i_t0, bt_b_operand_i_t0, ex_valid_o_t0, multdiv_operator_i_t0, multdiv_signed_mode_i_t0, result_ex_o_t0);
wire _000_;
wire [1:0] _001_;
wire _002_;
wire [33:0] _003_;
wire [1:0] _004_;
wire [31:0] _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire [1:0] _012_;
wire [33:0] _013_;
wire [33:0] _014_;
wire [33:0] _015_;
wire [33:0] _016_;
wire [33:0] _017_;
wire [33:0] _018_;
wire [1:0] _019_;
wire [1:0] _020_;
wire [1:0] _021_;
wire [31:0] _022_;
wire [31:0] _023_;
wire [31:0] _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire [33:0] _029_;
wire [33:0] _030_;
wire [33:0] _031_;
wire [33:0] _032_;
wire [1:0] _033_;
wire [1:0] _034_;
wire [1:0] _035_;
wire [31:0] _036_;
wire [31:0] _037_;
wire [31:0] _038_;
wire _039_;
wire _040_;
wire _041_;
wire [33:0] _042_;
wire [33:0] _043_;
wire [1:0] _044_;
wire [31:0] _045_;
wire _046_;
/* src = "generated/sv2v_out.v:16057.53-16057.71" */
wire _047_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16057.53-16057.71" */
wire _048_;
/* src = "generated/sv2v_out.v:16057.55-16057.70" */
wire _049_;
/* src = "generated/sv2v_out.v:15937.21-15937.42" */
output [31:0] alu_adder_result_ex_o;
wire [31:0] alu_adder_result_ex_o;
/* cellift = 32'd1 */
output [31:0] alu_adder_result_ex_o_t0;
wire [31:0] alu_adder_result_ex_o_t0;
/* src = "generated/sv2v_out.v:15946.14-15946.34" */
wire [33:0] alu_adder_result_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15946.14-15946.34" */
wire [33:0] alu_adder_result_ext_t0;
/* src = "generated/sv2v_out.v:15952.14-15952.27" */
wire [63:0] alu_imd_val_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15952.14-15952.27" */
wire [63:0] alu_imd_val_d_t0;
/* src = "generated/sv2v_out.v:15953.13-15953.27" */
wire [1:0] alu_imd_val_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15953.13-15953.27" */
wire [1:0] alu_imd_val_we_t0;
/* src = "generated/sv2v_out.v:15921.13-15921.36" */
input alu_instr_first_cycle_i;
wire alu_instr_first_cycle_i;
/* cellift = 32'd1 */
input alu_instr_first_cycle_i_t0;
wire alu_instr_first_cycle_i_t0;
/* src = "generated/sv2v_out.v:15948.7-15948.26" */
wire alu_is_equal_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15948.7-15948.26" */
wire alu_is_equal_result_t0;
/* src = "generated/sv2v_out.v:15919.20-15919.35" */
input [31:0] alu_operand_a_i;
wire [31:0] alu_operand_a_i;
/* cellift = 32'd1 */
input [31:0] alu_operand_a_i_t0;
wire [31:0] alu_operand_a_i_t0;
/* src = "generated/sv2v_out.v:15920.20-15920.35" */
input [31:0] alu_operand_b_i;
wire [31:0] alu_operand_b_i;
/* cellift = 32'd1 */
input [31:0] alu_operand_b_i_t0;
wire [31:0] alu_operand_b_i_t0;
/* src = "generated/sv2v_out.v:15918.19-15918.33" */
input [6:0] alu_operator_i;
wire [6:0] alu_operator_i;
/* cellift = 32'd1 */
input [6:0] alu_operator_i_t0;
wire [6:0] alu_operator_i_t0;
/* src = "generated/sv2v_out.v:15942.14-15942.24" */
wire [31:0] alu_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15942.14-15942.24" */
wire [31:0] alu_result_t0;
/* src = "generated/sv2v_out.v:15940.14-15940.31" */
output branch_decision_o;
wire branch_decision_o;
/* cellift = 32'd1 */
output branch_decision_o_t0;
wire branch_decision_o_t0;
/* src = "generated/sv2v_out.v:15939.21-15939.36" */
output [31:0] branch_target_o;
wire [31:0] branch_target_o;
/* cellift = 32'd1 */
output [31:0] branch_target_o_t0;
wire [31:0] branch_target_o_t0;
/* src = "generated/sv2v_out.v:15922.20-15922.34" */
input [31:0] bt_a_operand_i;
wire [31:0] bt_a_operand_i;
/* cellift = 32'd1 */
input [31:0] bt_a_operand_i_t0;
wire [31:0] bt_a_operand_i_t0;
/* src = "generated/sv2v_out.v:15923.20-15923.34" */
input [31:0] bt_b_operand_i;
wire [31:0] bt_b_operand_i;
/* cellift = 32'd1 */
input [31:0] bt_b_operand_i_t0;
wire [31:0] bt_b_operand_i_t0;
/* src = "generated/sv2v_out.v:15916.13-15916.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:15933.13-15933.30" */
input data_ind_timing_i;
wire data_ind_timing_i;
/* cellift = 32'd1 */
input data_ind_timing_i_t0;
wire data_ind_timing_i_t0;
/* src = "generated/sv2v_out.v:15926.13-15926.21" */
input div_en_i;
wire div_en_i;
/* cellift = 32'd1 */
input div_en_i_t0;
wire div_en_i_t0;
/* src = "generated/sv2v_out.v:15928.13-15928.22" */
input div_sel_i;
wire div_sel_i;
/* cellift = 32'd1 */
input div_sel_i_t0;
wire div_sel_i_t0;
/* src = "generated/sv2v_out.v:15941.14-15941.24" */
output ex_valid_o;
wire ex_valid_o;
/* cellift = 32'd1 */
output ex_valid_o_t0;
wire ex_valid_o_t0;
/* src = "generated/sv2v_out.v:15935.21-15935.32" */
output [67:0] imd_val_d_o;
wire [67:0] imd_val_d_o;
/* cellift = 32'd1 */
output [67:0] imd_val_d_o_t0;
wire [67:0] imd_val_d_o_t0;
/* src = "generated/sv2v_out.v:15936.20-15936.31" */
input [67:0] imd_val_q_i;
wire [67:0] imd_val_q_i;
/* cellift = 32'd1 */
input [67:0] imd_val_q_i_t0;
wire [67:0] imd_val_q_i_t0;
/* src = "generated/sv2v_out.v:15934.20-15934.32" */
output [1:0] imd_val_we_o;
wire [1:0] imd_val_we_o;
/* cellift = 32'd1 */
output [1:0] imd_val_we_o_t0;
wire [1:0] imd_val_we_o_t0;
/* src = "generated/sv2v_out.v:15925.13-15925.22" */
input mult_en_i;
wire mult_en_i;
/* cellift = 32'd1 */
input mult_en_i_t0;
wire mult_en_i_t0;
/* src = "generated/sv2v_out.v:15927.13-15927.23" */
input mult_sel_i;
wire mult_sel_i;
/* cellift = 32'd1 */
input mult_sel_i_t0;
wire mult_sel_i_t0;
/* src = "generated/sv2v_out.v:15945.14-15945.35" */
wire [32:0] multdiv_alu_operand_a;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15945.14-15945.35" */
wire [32:0] multdiv_alu_operand_a_t0;
/* src = "generated/sv2v_out.v:15944.14-15944.35" */
wire [32:0] multdiv_alu_operand_b;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15944.14-15944.35" */
wire [32:0] multdiv_alu_operand_b_t0;
/* src = "generated/sv2v_out.v:15954.14-15954.31" */
wire [67:0] multdiv_imd_val_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15954.14-15954.31" */
wire [67:0] multdiv_imd_val_d_t0;
/* src = "generated/sv2v_out.v:15955.13-15955.31" */
wire [1:0] multdiv_imd_val_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15955.13-15955.31" */
wire [1:0] multdiv_imd_val_we_t0;
/* src = "generated/sv2v_out.v:15930.20-15930.39" */
input [31:0] multdiv_operand_a_i;
wire [31:0] multdiv_operand_a_i;
/* cellift = 32'd1 */
input [31:0] multdiv_operand_a_i_t0;
wire [31:0] multdiv_operand_a_i_t0;
/* src = "generated/sv2v_out.v:15931.20-15931.39" */
input [31:0] multdiv_operand_b_i;
wire [31:0] multdiv_operand_b_i;
/* cellift = 32'd1 */
input [31:0] multdiv_operand_b_i_t0;
wire [31:0] multdiv_operand_b_i_t0;
/* src = "generated/sv2v_out.v:15924.19-15924.37" */
input [1:0] multdiv_operator_i;
wire [1:0] multdiv_operator_i;
/* cellift = 32'd1 */
input [1:0] multdiv_operator_i_t0;
wire [1:0] multdiv_operator_i_t0;
/* src = "generated/sv2v_out.v:15932.13-15932.31" */
input multdiv_ready_id_i;
wire multdiv_ready_id_i;
/* cellift = 32'd1 */
input multdiv_ready_id_i_t0;
wire multdiv_ready_id_i_t0;
/* src = "generated/sv2v_out.v:15943.14-15943.28" */
wire [31:0] multdiv_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15943.14-15943.28" */
wire [31:0] multdiv_result_t0;
/* src = "generated/sv2v_out.v:15950.7-15950.18" */
wire multdiv_sel;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15950.7-15950.18" */
wire multdiv_sel_t0;
/* src = "generated/sv2v_out.v:15929.19-15929.40" */
input [1:0] multdiv_signed_mode_i;
wire [1:0] multdiv_signed_mode_i;
/* cellift = 32'd1 */
input [1:0] multdiv_signed_mode_i_t0;
wire [1:0] multdiv_signed_mode_i_t0;
/* src = "generated/sv2v_out.v:15949.7-15949.20" */
wire multdiv_valid;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:15949.7-15949.20" */
wire multdiv_valid_t0;
/* src = "generated/sv2v_out.v:15938.21-15938.32" */
output [31:0] result_ex_o;
wire [31:0] result_ex_o;
/* cellift = 32'd1 */
output [31:0] result_ex_o_t0;
wire [31:0] result_ex_o_t0;
/* src = "generated/sv2v_out.v:15917.13-15917.19" */
input rst_ni;
wire rst_ni;
assign _000_ = | alu_imd_val_we_t0;
assign _001_ = ~ alu_imd_val_we_t0;
assign _012_ = alu_imd_val_we & _001_;
assign _002_ = ! _012_;
assign _048_ = _002_ & _000_;
assign _003_ = ~ { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel };
assign _004_ = ~ { multdiv_sel, multdiv_sel };
assign _005_ = ~ { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel };
assign _006_ = ~ multdiv_sel;
assign _029_ = { multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0 } | _003_;
assign _033_ = { multdiv_sel_t0, multdiv_sel_t0 } | _004_;
assign _036_ = { multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0 } | _005_;
assign _039_ = multdiv_sel_t0 | _006_;
assign _030_ = { multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0 } | { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel };
assign _034_ = { multdiv_sel_t0, multdiv_sel_t0 } | { multdiv_sel, multdiv_sel };
assign _037_ = { multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0 } | { multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel, multdiv_sel };
assign _040_ = multdiv_sel_t0 | multdiv_sel;
assign _013_ = { 2'h0, alu_imd_val_d_t0[63:32] } & _029_;
assign _016_ = { 2'h0, alu_imd_val_d_t0[31:0] } & _029_;
assign _019_ = alu_imd_val_we_t0 & _033_;
assign _022_ = alu_result_t0 & _036_;
assign _025_ = _048_ & _039_;
assign _014_ = multdiv_imd_val_d_t0[67:34] & _030_;
assign _017_ = multdiv_imd_val_d_t0[33:0] & _030_;
assign _020_ = multdiv_imd_val_we_t0 & _034_;
assign _023_ = multdiv_result_t0 & _037_;
assign _026_ = multdiv_valid_t0 & _040_;
assign _031_ = _013_ | _014_;
assign _032_ = _016_ | _017_;
assign _035_ = _019_ | _020_;
assign _038_ = _022_ | _023_;
assign _041_ = _025_ | _026_;
assign _042_ = { 2'h0, alu_imd_val_d[63:32] } ^ multdiv_imd_val_d[67:34];
assign _043_ = { 2'h0, alu_imd_val_d[31:0] } ^ multdiv_imd_val_d[33:0];
assign _044_ = alu_imd_val_we ^ multdiv_imd_val_we;
assign _045_ = alu_result ^ multdiv_result;
assign _046_ = _047_ ^ multdiv_valid;
assign _015_ = { multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0 } & _042_;
assign _018_ = { multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0 } & _043_;
assign _021_ = { multdiv_sel_t0, multdiv_sel_t0 } & _044_;
assign _024_ = { multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0, multdiv_sel_t0 } & _045_;
assign _027_ = multdiv_sel_t0 & _046_;
assign imd_val_d_o_t0[67:34] = _015_ | _031_;
assign imd_val_d_o_t0[33:0] = _018_ | _032_;
assign imd_val_we_o_t0 = _021_ | _035_;
assign result_ex_o_t0 = _024_ | _038_;
assign ex_valid_o_t0 = _027_ | _041_;
assign _007_ = ~ mult_sel_i;
assign _008_ = ~ div_sel_i;
assign _009_ = mult_sel_i_t0 & _008_;
assign _010_ = div_sel_i_t0 & _007_;
assign _011_ = mult_sel_i_t0 & div_sel_i_t0;
assign _028_ = _009_ | _010_;
assign multdiv_sel_t0 = _028_ | _011_;
assign _047_ = ~ /* src = "generated/sv2v_out.v:16057.53-16057.71" */ _049_;
assign multdiv_sel = mult_sel_i | /* src = "generated/sv2v_out.v:15958.25-15958.47" */ div_sel_i;
assign _049_ = | /* src = "generated/sv2v_out.v:16057.55-16057.70" */ alu_imd_val_we;
assign imd_val_d_o[67:34] = multdiv_sel ? /* src = "generated/sv2v_out.v:15964.32-15964.104" */ multdiv_imd_val_d[67:34] : { 2'h0, alu_imd_val_d[63:32] };
assign imd_val_d_o[33:0] = multdiv_sel ? /* src = "generated/sv2v_out.v:15965.31-15965.101" */ multdiv_imd_val_d[33:0] : { 2'h0, alu_imd_val_d[31:0] };
assign imd_val_we_o = multdiv_sel ? /* src = "generated/sv2v_out.v:15966.25-15966.74" */ multdiv_imd_val_we : alu_imd_val_we;
assign result_ex_o = multdiv_sel ? /* src = "generated/sv2v_out.v:15968.24-15968.65" */ multdiv_result : alu_result;
assign ex_valid_o = multdiv_sel ? /* src = "generated/sv2v_out.v:16057.23-16057.71" */ multdiv_valid : _047_;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:15986.28-16002.3" */
\$paramod\ibex_alu\RV32B=s32'00000000000000000000000000000000  alu_i (
.adder_result_ext_o(alu_adder_result_ext),
.adder_result_ext_o_t0(alu_adder_result_ext_t0),
.adder_result_o(alu_adder_result_ex_o),
.adder_result_o_t0(alu_adder_result_ex_o_t0),
.comparison_result_o(branch_decision_o),
.comparison_result_o_t0(branch_decision_o_t0),
.imd_val_d_o(alu_imd_val_d),
.imd_val_d_o_t0(alu_imd_val_d_t0),
.imd_val_q_i({ imd_val_q_i[65:34], imd_val_q_i[31:0] }),
.imd_val_q_i_t0({ imd_val_q_i_t0[65:34], imd_val_q_i_t0[31:0] }),
.imd_val_we_o(alu_imd_val_we),
.imd_val_we_o_t0(alu_imd_val_we_t0),
.instr_first_cycle_i(alu_instr_first_cycle_i),
.instr_first_cycle_i_t0(alu_instr_first_cycle_i_t0),
.is_equal_result_o(alu_is_equal_result),
.is_equal_result_o_t0(alu_is_equal_result_t0),
.multdiv_operand_a_i(multdiv_alu_operand_a),
.multdiv_operand_a_i_t0(multdiv_alu_operand_a_t0),
.multdiv_operand_b_i(multdiv_alu_operand_b),
.multdiv_operand_b_i_t0(multdiv_alu_operand_b_t0),
.multdiv_sel_i(multdiv_sel),
.multdiv_sel_i_t0(multdiv_sel_t0),
.operand_a_i(alu_operand_a_i),
.operand_a_i_t0(alu_operand_a_i_t0),
.operand_b_i(alu_operand_b_i),
.operand_b_i_t0(alu_operand_b_i_t0),
.operator_i(alu_operator_i),
.operator_i_t0(alu_operator_i_t0),
.result_o(alu_result),
.result_o_t0(alu_result_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:16005.22-16028.5" */
ibex_multdiv_slow \gen_multdiv_slow.multdiv_i  (
.alu_adder_ext_i(alu_adder_result_ext),
.alu_adder_ext_i_t0(alu_adder_result_ext_t0),
.alu_adder_i(alu_adder_result_ex_o),
.alu_adder_i_t0(alu_adder_result_ex_o_t0),
.alu_operand_a_o(multdiv_alu_operand_a),
.alu_operand_a_o_t0(multdiv_alu_operand_a_t0),
.alu_operand_b_o(multdiv_alu_operand_b),
.alu_operand_b_o_t0(multdiv_alu_operand_b_t0),
.clk_i(clk_i),
.data_ind_timing_i(data_ind_timing_i),
.data_ind_timing_i_t0(data_ind_timing_i_t0),
.div_en_i(div_en_i),
.div_en_i_t0(div_en_i_t0),
.div_sel_i(div_sel_i),
.div_sel_i_t0(div_sel_i_t0),
.equal_to_zero_i(alu_is_equal_result),
.equal_to_zero_i_t0(alu_is_equal_result_t0),
.imd_val_d_o(multdiv_imd_val_d),
.imd_val_d_o_t0(multdiv_imd_val_d_t0),
.imd_val_q_i(imd_val_q_i),
.imd_val_q_i_t0(imd_val_q_i_t0),
.imd_val_we_o(multdiv_imd_val_we),
.imd_val_we_o_t0(multdiv_imd_val_we_t0),
.mult_en_i(mult_en_i),
.mult_en_i_t0(mult_en_i_t0),
.mult_sel_i(mult_sel_i),
.mult_sel_i_t0(mult_sel_i_t0),
.multdiv_ready_id_i(multdiv_ready_id_i),
.multdiv_ready_id_i_t0(multdiv_ready_id_i_t0),
.multdiv_result_o(multdiv_result),
.multdiv_result_o_t0(multdiv_result_t0),
.op_a_i(multdiv_operand_a_i),
.op_a_i_t0(multdiv_operand_a_i_t0),
.op_b_i(multdiv_operand_b_i),
.op_b_i_t0(multdiv_operand_b_i_t0),
.operator_i(multdiv_operator_i),
.operator_i_t0(multdiv_operator_i_t0),
.rst_ni(rst_ni),
.signed_mode_i(multdiv_signed_mode_i),
.signed_mode_i_t0(multdiv_signed_mode_i_t0),
.valid_o(multdiv_valid),
.valid_o_t0(multdiv_valid_t0)
);
assign branch_target_o = alu_adder_result_ex_o;
assign branch_target_o_t0 = alu_adder_result_ex_o_t0;
endmodule

module \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff (clk_i, rst_ni, test_en_i, dummy_instr_id_i, dummy_instr_wb_i, raddr_a_i, rdata_a_o, raddr_b_i, rdata_b_o, waddr_a_i, wdata_a_i, we_a_i, err_o, test_en_i_t0, err_o_t0, dummy_instr_id_i_t0, dummy_instr_wb_i_t0, raddr_a_i_t0, raddr_b_i_t0, rdata_a_o_t0, rdata_b_o_t0
, waddr_a_i_t0, wdata_a_i_t0, we_a_i_t0);
wire _0000_;
wire _0001_;
wire _0002_;
wire _0003_;
wire _0004_;
wire _0005_;
wire _0006_;
wire _0007_;
wire _0008_;
wire _0009_;
wire _0010_;
wire _0011_;
wire _0012_;
wire _0013_;
wire _0014_;
wire _0015_;
wire _0016_;
wire _0017_;
wire _0018_;
wire _0019_;
wire _0020_;
wire _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire _0026_;
wire _0027_;
wire _0028_;
wire _0029_;
wire _0030_;
wire _0031_;
wire _0032_;
wire _0033_;
wire _0034_;
wire [4:0] _0035_;
wire [4:0] _0036_;
wire [4:0] _0037_;
wire _0038_;
wire _0039_;
wire _0040_;
wire _0041_;
wire _0042_;
wire _0043_;
wire _0044_;
wire _0045_;
wire _0046_;
wire _0047_;
wire _0048_;
wire _0049_;
wire _0050_;
wire _0051_;
wire [2:0] _0052_;
wire [2:0] _0053_;
wire [5:0] _0054_;
wire [2:0] _0055_;
wire [2:0] _0056_;
wire [5:0] _0057_;
wire [11:0] _0058_;
wire [2:0] _0059_;
wire [2:0] _0060_;
wire [5:0] _0061_;
wire [2:0] _0062_;
wire [2:0] _0063_;
wire [5:0] _0064_;
wire [11:0] _0065_;
wire _0066_;
wire _0067_;
wire _0068_;
wire _0069_;
wire _0070_;
wire _0071_;
wire _0072_;
wire _0073_;
wire _0074_;
wire _0075_;
wire _0076_;
wire _0077_;
wire _0078_;
wire _0079_;
wire _0080_;
wire [38:0] _0081_;
wire [38:0] _0082_;
wire [38:0] _0083_;
wire [38:0] _0084_;
wire [38:0] _0085_;
wire [38:0] _0086_;
wire [38:0] _0087_;
wire [38:0] _0088_;
wire [38:0] _0089_;
wire [38:0] _0090_;
wire [38:0] _0091_;
wire [38:0] _0092_;
wire [38:0] _0093_;
wire [38:0] _0094_;
wire [38:0] _0095_;
wire [38:0] _0096_;
wire [38:0] _0097_;
wire [38:0] _0098_;
wire [38:0] _0099_;
wire [38:0] _0100_;
wire [38:0] _0101_;
wire [38:0] _0102_;
wire [38:0] _0103_;
wire [38:0] _0104_;
wire [38:0] _0105_;
wire [38:0] _0106_;
wire [38:0] _0107_;
wire [38:0] _0108_;
wire [38:0] _0109_;
wire [38:0] _0110_;
wire [38:0] _0111_;
wire [38:0] _0112_;
wire [38:0] _0113_;
wire [38:0] _0114_;
wire [38:0] _0115_;
wire [38:0] _0116_;
wire [38:0] _0117_;
wire [38:0] _0118_;
wire [38:0] _0119_;
wire [38:0] _0120_;
wire [38:0] _0121_;
wire [38:0] _0122_;
wire [38:0] _0123_;
wire [38:0] _0124_;
wire [38:0] _0125_;
wire [38:0] _0126_;
wire [38:0] _0127_;
wire [38:0] _0128_;
wire [38:0] _0129_;
wire [38:0] _0130_;
wire [38:0] _0131_;
wire [38:0] _0132_;
wire [38:0] _0133_;
wire [38:0] _0134_;
wire [38:0] _0135_;
wire [38:0] _0136_;
wire [38:0] _0137_;
wire [38:0] _0138_;
wire [38:0] _0139_;
wire [38:0] _0140_;
wire [38:0] _0141_;
wire [38:0] _0142_;
wire [2:0] _0143_;
wire _0144_;
wire _0145_;
wire _0146_;
wire _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
wire _0152_;
wire _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
/* cellift = 32'd1 */
wire _0177_;
wire _0178_;
/* cellift = 32'd1 */
wire _0179_;
wire _0180_;
/* cellift = 32'd1 */
wire _0181_;
wire _0182_;
/* cellift = 32'd1 */
wire _0183_;
wire _0184_;
/* cellift = 32'd1 */
wire _0185_;
wire _0186_;
/* cellift = 32'd1 */
wire _0187_;
wire _0188_;
/* cellift = 32'd1 */
wire _0189_;
wire _0190_;
/* cellift = 32'd1 */
wire _0191_;
wire _0192_;
/* cellift = 32'd1 */
wire _0193_;
wire _0194_;
/* cellift = 32'd1 */
wire _0195_;
wire _0196_;
/* cellift = 32'd1 */
wire _0197_;
wire _0198_;
/* cellift = 32'd1 */
wire _0199_;
wire _0200_;
/* cellift = 32'd1 */
wire _0201_;
wire _0202_;
/* cellift = 32'd1 */
wire _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire [38:0] _0207_;
wire [38:0] _0208_;
wire [38:0] _0209_;
wire [38:0] _0210_;
wire [38:0] _0211_;
wire [38:0] _0212_;
wire [38:0] _0213_;
wire [38:0] _0214_;
wire [38:0] _0215_;
wire [38:0] _0216_;
wire [38:0] _0217_;
wire [38:0] _0218_;
wire [38:0] _0219_;
wire [38:0] _0220_;
wire [38:0] _0221_;
wire [38:0] _0222_;
wire [38:0] _0223_;
wire [38:0] _0224_;
wire [38:0] _0225_;
wire [38:0] _0226_;
wire [38:0] _0227_;
wire [38:0] _0228_;
wire [38:0] _0229_;
wire [38:0] _0230_;
wire [38:0] _0231_;
wire [38:0] _0232_;
wire [38:0] _0233_;
wire [38:0] _0234_;
wire [38:0] _0235_;
wire [38:0] _0236_;
wire [38:0] _0237_;
wire [38:0] _0238_;
wire [38:0] _0239_;
wire [38:0] _0240_;
wire [38:0] _0241_;
wire [38:0] _0242_;
wire [38:0] _0243_;
wire [38:0] _0244_;
wire [38:0] _0245_;
wire [38:0] _0246_;
wire [38:0] _0247_;
wire [38:0] _0248_;
wire [38:0] _0249_;
wire [38:0] _0250_;
wire [38:0] _0251_;
wire [38:0] _0252_;
wire [38:0] _0253_;
wire [38:0] _0254_;
wire [38:0] _0255_;
wire [38:0] _0256_;
wire [38:0] _0257_;
wire [38:0] _0258_;
wire [38:0] _0259_;
wire [38:0] _0260_;
wire [38:0] _0261_;
wire [38:0] _0262_;
wire [38:0] _0263_;
wire [38:0] _0264_;
wire [38:0] _0265_;
wire [38:0] _0266_;
wire [38:0] _0267_;
wire [38:0] _0268_;
wire [38:0] _0269_;
wire [38:0] _0270_;
wire [38:0] _0271_;
wire [38:0] _0272_;
wire [38:0] _0273_;
wire [38:0] _0274_;
wire [38:0] _0275_;
wire [38:0] _0276_;
wire [38:0] _0277_;
wire [38:0] _0278_;
wire [38:0] _0279_;
wire [38:0] _0280_;
wire [38:0] _0281_;
wire [38:0] _0282_;
wire [38:0] _0283_;
wire [38:0] _0284_;
wire [38:0] _0285_;
wire [38:0] _0286_;
wire [38:0] _0287_;
wire [38:0] _0288_;
wire [38:0] _0289_;
wire [38:0] _0290_;
wire [38:0] _0291_;
wire [38:0] _0292_;
wire [38:0] _0293_;
wire [38:0] _0294_;
wire [38:0] _0295_;
wire [38:0] _0296_;
wire [38:0] _0297_;
wire [38:0] _0298_;
wire [38:0] _0299_;
wire [38:0] _0300_;
wire [38:0] _0301_;
wire [38:0] _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire _0324_;
wire _0325_;
wire _0326_;
wire _0327_;
wire _0328_;
wire _0329_;
wire _0330_;
wire _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire _0335_;
wire _0336_;
wire _0337_;
wire _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire _0344_;
wire _0345_;
wire _0346_;
wire _0347_;
wire _0348_;
wire _0349_;
wire _0350_;
wire [2:0] _0351_;
wire [2:0] _0352_;
wire [5:0] _0353_;
wire [2:0] _0354_;
wire [2:0] _0355_;
wire [5:0] _0356_;
wire [11:0] _0357_;
wire [2:0] _0358_;
wire [2:0] _0359_;
wire [5:0] _0360_;
wire [2:0] _0361_;
wire [2:0] _0362_;
wire [5:0] _0363_;
wire [11:0] _0364_;
wire [38:0] _0365_;
wire [38:0] _0366_;
wire [38:0] _0367_;
wire [38:0] _0368_;
wire [38:0] _0369_;
wire [38:0] _0370_;
wire [38:0] _0371_;
wire [38:0] _0372_;
wire [38:0] _0373_;
wire [38:0] _0374_;
wire [38:0] _0375_;
wire [38:0] _0376_;
wire [38:0] _0377_;
wire [38:0] _0378_;
wire [38:0] _0379_;
wire [38:0] _0380_;
wire [38:0] _0381_;
wire [38:0] _0382_;
wire [38:0] _0383_;
wire [38:0] _0384_;
wire [38:0] _0385_;
wire [38:0] _0386_;
wire [38:0] _0387_;
wire [38:0] _0388_;
wire [38:0] _0389_;
wire [38:0] _0390_;
wire [38:0] _0391_;
wire [38:0] _0392_;
wire [38:0] _0393_;
wire [38:0] _0394_;
wire [38:0] _0395_;
wire [38:0] _0396_;
wire [38:0] _0397_;
wire [38:0] _0398_;
wire [38:0] _0399_;
wire [38:0] _0400_;
wire [38:0] _0401_;
wire [38:0] _0402_;
wire [38:0] _0403_;
wire [38:0] _0404_;
wire [38:0] _0405_;
wire [38:0] _0406_;
wire [38:0] _0407_;
wire [38:0] _0408_;
wire [38:0] _0409_;
wire [38:0] _0410_;
wire [38:0] _0411_;
wire [38:0] _0412_;
wire [38:0] _0413_;
wire [38:0] _0414_;
wire [38:0] _0415_;
wire [38:0] _0416_;
wire [38:0] _0417_;
wire [38:0] _0418_;
wire [38:0] _0419_;
wire [38:0] _0420_;
wire [38:0] _0421_;
wire [38:0] _0422_;
wire [38:0] _0423_;
wire [38:0] _0424_;
wire [38:0] _0425_;
wire [38:0] _0426_;
wire [38:0] _0427_;
wire [38:0] _0428_;
wire [38:0] _0429_;
wire [38:0] _0430_;
wire [38:0] _0431_;
wire [38:0] _0432_;
wire [38:0] _0433_;
wire [38:0] _0434_;
wire [38:0] _0435_;
wire [38:0] _0436_;
wire [38:0] _0437_;
wire [38:0] _0438_;
wire [38:0] _0439_;
wire [38:0] _0440_;
wire [38:0] _0441_;
wire [38:0] _0442_;
wire [38:0] _0443_;
wire [38:0] _0444_;
wire [38:0] _0445_;
wire [38:0] _0446_;
wire [38:0] _0447_;
wire [38:0] _0448_;
wire [38:0] _0449_;
wire [38:0] _0450_;
wire [38:0] _0451_;
wire [38:0] _0452_;
wire [38:0] _0453_;
wire [38:0] _0454_;
wire [38:0] _0455_;
wire [38:0] _0456_;
wire [38:0] _0457_;
wire [38:0] _0458_;
wire [38:0] _0459_;
wire [38:0] _0460_;
wire [38:0] _0461_;
wire [38:0] _0462_;
wire [38:0] _0463_;
wire [38:0] _0464_;
wire [38:0] _0465_;
wire [38:0] _0466_;
wire [38:0] _0467_;
wire [38:0] _0468_;
wire [38:0] _0469_;
wire [38:0] _0470_;
wire [38:0] _0471_;
wire [38:0] _0472_;
wire [38:0] _0473_;
wire [38:0] _0474_;
wire [38:0] _0475_;
wire [38:0] _0476_;
wire [38:0] _0477_;
wire [38:0] _0478_;
wire [38:0] _0479_;
wire [38:0] _0480_;
wire [38:0] _0481_;
wire [38:0] _0482_;
wire [38:0] _0483_;
wire [38:0] _0484_;
wire [38:0] _0485_;
wire [38:0] _0486_;
wire [38:0] _0487_;
wire [38:0] _0488_;
wire [38:0] _0489_;
wire [38:0] _0490_;
wire [38:0] _0491_;
wire [38:0] _0492_;
wire [38:0] _0493_;
wire [38:0] _0494_;
wire [38:0] _0495_;
wire [38:0] _0496_;
wire [38:0] _0497_;
wire [38:0] _0498_;
wire [38:0] _0499_;
wire [38:0] _0500_;
wire [38:0] _0501_;
wire [38:0] _0502_;
wire [38:0] _0503_;
wire [38:0] _0504_;
wire [38:0] _0505_;
wire [38:0] _0506_;
wire [38:0] _0507_;
wire [38:0] _0508_;
wire [38:0] _0509_;
wire [38:0] _0510_;
wire [38:0] _0511_;
wire [38:0] _0512_;
wire [38:0] _0513_;
wire [38:0] _0514_;
wire [38:0] _0515_;
wire [38:0] _0516_;
wire [38:0] _0517_;
wire [38:0] _0518_;
wire [38:0] _0519_;
wire [38:0] _0520_;
wire [38:0] _0521_;
wire [38:0] _0522_;
wire [38:0] _0523_;
wire [38:0] _0524_;
wire [38:0] _0525_;
wire [38:0] _0526_;
wire [38:0] _0527_;
wire [38:0] _0528_;
wire [38:0] _0529_;
wire [38:0] _0530_;
wire [38:0] _0531_;
wire [38:0] _0532_;
wire [38:0] _0533_;
wire [38:0] _0534_;
wire [38:0] _0535_;
wire [38:0] _0536_;
wire [38:0] _0537_;
wire [38:0] _0538_;
wire [38:0] _0539_;
wire [38:0] _0540_;
wire [38:0] _0541_;
wire [38:0] _0542_;
wire [38:0] _0543_;
wire [38:0] _0544_;
wire [38:0] _0545_;
wire [38:0] _0546_;
wire [38:0] _0547_;
wire [38:0] _0548_;
wire [38:0] _0549_;
wire [38:0] _0550_;
wire [4:0] _0551_;
wire [4:0] _0552_;
wire [4:0] _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire _0560_;
wire _0561_;
wire _0562_;
wire _0563_;
wire _0564_;
wire _0565_;
wire _0566_;
wire _0567_;
wire _0568_;
wire _0569_;
wire _0570_;
wire _0571_;
wire _0572_;
wire _0573_;
wire _0574_;
wire _0575_;
wire _0576_;
wire _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire _0596_;
wire _0597_;
wire _0598_;
wire _0599_;
wire _0600_;
wire _0601_;
wire _0602_;
wire _0603_;
wire _0604_;
wire _0605_;
wire _0606_;
wire _0607_;
wire _0608_;
wire _0609_;
wire _0610_;
wire _0611_;
wire _0612_;
wire _0613_;
wire _0614_;
wire _0615_;
wire _0616_;
wire _0617_;
wire [38:0] _0618_;
wire [38:0] _0619_;
wire _0620_;
wire [38:0] _0621_;
wire [38:0] _0622_;
wire [38:0] _0623_;
wire [38:0] _0624_;
wire [38:0] _0625_;
wire [38:0] _0626_;
wire [38:0] _0627_;
wire [38:0] _0628_;
wire [38:0] _0629_;
wire [38:0] _0630_;
wire [38:0] _0631_;
wire [38:0] _0632_;
wire [38:0] _0633_;
wire [38:0] _0634_;
wire [38:0] _0635_;
wire [38:0] _0636_;
wire [38:0] _0637_;
wire [38:0] _0638_;
wire [38:0] _0639_;
wire [38:0] _0640_;
wire [38:0] _0641_;
wire [38:0] _0642_;
wire [38:0] _0643_;
wire [38:0] _0644_;
wire [38:0] _0645_;
wire [38:0] _0646_;
wire [38:0] _0647_;
wire [38:0] _0648_;
wire [38:0] _0649_;
wire [38:0] _0650_;
wire [38:0] _0651_;
wire [38:0] _0652_;
wire [38:0] _0653_;
wire [38:0] _0654_;
wire [38:0] _0655_;
wire [38:0] _0656_;
wire [38:0] _0657_;
wire [38:0] _0658_;
wire [38:0] _0659_;
wire [38:0] _0660_;
wire [38:0] _0661_;
wire [38:0] _0662_;
wire [38:0] _0663_;
wire [38:0] _0664_;
wire [38:0] _0665_;
wire [38:0] _0666_;
wire [38:0] _0667_;
wire [38:0] _0668_;
wire [38:0] _0669_;
wire [38:0] _0670_;
wire [38:0] _0671_;
wire [38:0] _0672_;
wire [38:0] _0673_;
wire [38:0] _0674_;
wire [38:0] _0675_;
wire [38:0] _0676_;
wire [38:0] _0677_;
wire [38:0] _0678_;
wire [38:0] _0679_;
wire [38:0] _0680_;
wire [38:0] _0681_;
wire [38:0] _0682_;
wire [38:0] _0683_;
wire [38:0] _0684_;
wire [38:0] _0685_;
wire [38:0] _0686_;
wire [38:0] _0687_;
wire [38:0] _0688_;
wire [38:0] _0689_;
wire [38:0] _0690_;
wire [38:0] _0691_;
wire [38:0] _0692_;
wire [38:0] _0693_;
wire [38:0] _0694_;
wire [38:0] _0695_;
wire [38:0] _0696_;
wire [38:0] _0697_;
wire [38:0] _0698_;
wire [38:0] _0699_;
wire [38:0] _0700_;
wire [38:0] _0701_;
wire [38:0] _0702_;
wire [38:0] _0703_;
wire [38:0] _0704_;
wire [38:0] _0705_;
wire [38:0] _0706_;
wire [38:0] _0707_;
wire [38:0] _0708_;
wire [38:0] _0709_;
wire [38:0] _0710_;
wire [38:0] _0711_;
wire [38:0] _0712_;
wire [38:0] _0713_;
wire [38:0] _0714_;
wire [38:0] _0715_;
wire [38:0] _0716_;
wire [38:0] _0717_;
wire [38:0] _0718_;
wire [38:0] _0719_;
wire [38:0] _0720_;
wire [38:0] _0721_;
wire [38:0] _0722_;
wire [38:0] _0723_;
wire [38:0] _0724_;
wire [38:0] _0725_;
wire [38:0] _0726_;
wire [38:0] _0727_;
wire [38:0] _0728_;
wire [38:0] _0729_;
wire [38:0] _0730_;
wire [38:0] _0731_;
wire [38:0] _0732_;
wire [38:0] _0733_;
wire [38:0] _0734_;
wire [38:0] _0735_;
wire [38:0] _0736_;
wire [38:0] _0737_;
wire [38:0] _0738_;
wire [38:0] _0739_;
wire [38:0] _0740_;
wire [38:0] _0741_;
wire [38:0] _0742_;
wire [38:0] _0743_;
wire [38:0] _0744_;
wire [38:0] _0745_;
wire [38:0] _0746_;
wire [38:0] _0747_;
wire [38:0] _0748_;
wire _0749_;
wire _0750_;
wire _0751_;
wire _0752_;
wire _0753_;
wire _0754_;
wire _0755_;
wire _0756_;
wire _0757_;
wire _0758_;
wire _0759_;
wire _0760_;
wire _0761_;
wire _0762_;
wire _0763_;
wire _0764_;
wire [38:0] _0765_;
wire [38:0] _0766_;
wire [38:0] _0767_;
wire [38:0] _0768_;
wire [38:0] _0769_;
wire [38:0] _0770_;
wire [38:0] _0771_;
wire [38:0] _0772_;
wire [38:0] _0773_;
wire [38:0] _0774_;
wire [38:0] _0775_;
wire [38:0] _0776_;
wire [38:0] _0777_;
wire [38:0] _0778_;
wire [38:0] _0779_;
wire [38:0] _0780_;
wire [38:0] _0781_;
wire [38:0] _0782_;
wire [38:0] _0783_;
wire [38:0] _0784_;
wire [38:0] _0785_;
wire [38:0] _0786_;
wire [38:0] _0787_;
wire [38:0] _0788_;
wire [38:0] _0789_;
wire [38:0] _0790_;
wire [38:0] _0791_;
wire [38:0] _0792_;
wire [38:0] _0793_;
wire [38:0] _0794_;
wire [38:0] _0795_;
wire [38:0] _0796_;
wire [38:0] _0797_;
wire [38:0] _0798_;
wire [38:0] _0799_;
wire [38:0] _0800_;
wire [38:0] _0801_;
wire [38:0] _0802_;
wire [38:0] _0803_;
wire [38:0] _0804_;
wire [38:0] _0805_;
wire [38:0] _0806_;
wire [38:0] _0807_;
wire [38:0] _0808_;
wire [38:0] _0809_;
wire [38:0] _0810_;
wire [38:0] _0811_;
wire [38:0] _0812_;
wire [38:0] _0813_;
wire [38:0] _0814_;
wire [38:0] _0815_;
wire [38:0] _0816_;
wire [38:0] _0817_;
wire [38:0] _0818_;
wire [38:0] _0819_;
wire [38:0] _0820_;
wire [38:0] _0821_;
wire [38:0] _0822_;
wire [38:0] _0823_;
wire [38:0] _0824_;
wire [38:0] _0825_;
wire [38:0] _0826_;
wire [38:0] _0827_;
wire [38:0] _0828_;
wire [38:0] _0829_;
wire [38:0] _0830_;
wire [38:0] _0831_;
wire [38:0] _0832_;
wire [38:0] _0833_;
wire [38:0] _0834_;
wire [38:0] _0835_;
wire [38:0] _0836_;
wire [38:0] _0837_;
wire [38:0] _0838_;
wire [38:0] _0839_;
wire [38:0] _0840_;
wire [38:0] _0841_;
wire [38:0] _0842_;
wire [38:0] _0843_;
wire [38:0] _0844_;
wire [38:0] _0845_;
wire [38:0] _0846_;
wire [38:0] _0847_;
wire [38:0] _0848_;
wire [38:0] _0849_;
wire [38:0] _0850_;
wire [38:0] _0851_;
wire [38:0] _0852_;
wire [38:0] _0853_;
wire [38:0] _0854_;
wire [38:0] _0855_;
wire [38:0] _0856_;
wire [38:0] _0857_;
wire [38:0] _0858_;
wire [38:0] _0859_;
wire [38:0] _0860_;
wire [38:0] _0861_;
wire [38:0] _0862_;
wire [38:0] _0863_;
wire [38:0] _0864_;
wire [38:0] _0865_;
wire [38:0] _0866_;
wire [38:0] _0867_;
wire [38:0] _0868_;
wire [38:0] _0869_;
wire [38:0] _0870_;
wire [38:0] _0871_;
wire [38:0] _0872_;
wire [38:0] _0873_;
wire [38:0] _0874_;
wire [38:0] _0875_;
wire [38:0] _0876_;
wire [38:0] _0877_;
wire [38:0] _0878_;
wire [38:0] _0879_;
wire [38:0] _0880_;
wire [38:0] _0881_;
wire [38:0] _0882_;
wire [38:0] _0883_;
wire [38:0] _0884_;
wire [38:0] _0885_;
wire [38:0] _0886_;
wire [38:0] _0887_;
wire [38:0] _0888_;
wire [38:0] _0889_;
wire [38:0] _0890_;
wire [38:0] _0891_;
wire [38:0] _0892_;
wire [38:0] _0893_;
wire [38:0] _0894_;
wire [38:0] _0895_;
wire [38:0] _0896_;
wire [38:0] _0897_;
wire [38:0] _0898_;
wire [38:0] _0899_;
wire [38:0] _0900_;
wire [38:0] _0901_;
wire [38:0] _0902_;
wire [38:0] _0903_;
wire [38:0] _0904_;
wire [38:0] _0905_;
wire [38:0] _0906_;
wire [38:0] _0907_;
wire [38:0] _0908_;
wire [38:0] _0909_;
wire [38:0] _0910_;
wire [38:0] _0911_;
wire [38:0] _0912_;
wire [38:0] _0913_;
wire [38:0] _0914_;
wire [38:0] _0915_;
wire [38:0] _0916_;
wire [38:0] _0917_;
wire [38:0] _0918_;
wire [38:0] _0919_;
wire [38:0] _0920_;
wire [38:0] _0921_;
wire [38:0] _0922_;
wire [38:0] _0923_;
wire [38:0] _0924_;
wire [38:0] _0925_;
wire [38:0] _0926_;
wire [38:0] _0927_;
wire [38:0] _0928_;
wire [38:0] _0929_;
wire [38:0] _0930_;
wire [38:0] _0931_;
wire [38:0] _0932_;
wire [38:0] _0933_;
wire [38:0] _0934_;
wire [38:0] _0935_;
wire [38:0] _0936_;
wire [38:0] _0937_;
wire [38:0] _0938_;
wire [38:0] _0939_;
wire [38:0] _0940_;
wire [38:0] _0941_;
wire [38:0] _0942_;
wire [38:0] _0943_;
wire [38:0] _0944_;
wire [38:0] _0945_;
wire [38:0] _0946_;
wire [38:0] _0947_;
wire [38:0] _0948_;
wire [38:0] _0949_;
wire [38:0] _0950_;
wire _0951_;
wire _0952_;
wire _0953_;
wire _0954_;
wire _0955_;
wire _0956_;
wire _0957_;
wire _0958_;
wire _0959_;
wire _0960_;
wire _0961_;
wire _0962_;
wire _0963_;
wire _0964_;
wire _0965_;
wire _0966_;
wire _0967_;
wire _0968_;
wire _0969_;
wire _0970_;
wire _0971_;
wire _0972_;
wire _0973_;
wire _0974_;
wire _0975_;
wire _0976_;
wire _0977_;
wire _0978_;
wire _0979_;
wire _0980_;
wire _0981_;
wire _0982_;
wire [38:0] _0983_;
wire _0984_;
/* cellift = 32'd1 */
wire _0985_;
wire _0986_;
/* cellift = 32'd1 */
wire _0987_;
wire _0988_;
/* cellift = 32'd1 */
wire _0989_;
wire _0990_;
/* cellift = 32'd1 */
wire _0991_;
wire _0992_;
/* cellift = 32'd1 */
wire _0993_;
wire _0994_;
/* cellift = 32'd1 */
wire _0995_;
wire _0996_;
/* cellift = 32'd1 */
wire _0997_;
wire _0998_;
/* cellift = 32'd1 */
wire _0999_;
wire _1000_;
/* cellift = 32'd1 */
wire _1001_;
wire _1002_;
/* cellift = 32'd1 */
wire _1003_;
wire _1004_;
/* cellift = 32'd1 */
wire _1005_;
wire _1006_;
/* cellift = 32'd1 */
wire _1007_;
wire _1008_;
/* cellift = 32'd1 */
wire _1009_;
wire _1010_;
/* cellift = 32'd1 */
wire _1011_;
wire _1012_;
/* cellift = 32'd1 */
wire _1013_;
wire _1014_;
/* cellift = 32'd1 */
wire _1015_;
wire [38:0] _1016_;
wire [38:0] _1017_;
wire [38:0] _1018_;
wire [38:0] _1019_;
wire [38:0] _1020_;
wire [38:0] _1021_;
wire [38:0] _1022_;
wire [38:0] _1023_;
wire [38:0] _1024_;
wire [38:0] _1025_;
wire [38:0] _1026_;
wire [38:0] _1027_;
wire [38:0] _1028_;
wire [38:0] _1029_;
wire [38:0] _1030_;
wire [38:0] _1031_;
wire [38:0] _1032_;
wire [38:0] _1033_;
wire [38:0] _1034_;
wire [38:0] _1035_;
wire [38:0] _1036_;
wire [38:0] _1037_;
wire [38:0] _1038_;
wire [38:0] _1039_;
wire [38:0] _1040_;
wire [38:0] _1041_;
wire [38:0] _1042_;
wire [38:0] _1043_;
wire [38:0] _1044_;
wire [38:0] _1045_;
wire [38:0] _1046_;
wire [38:0] _1047_;
wire [38:0] _1048_;
wire [38:0] _1049_;
wire [38:0] _1050_;
wire [38:0] _1051_;
wire [38:0] _1052_;
wire [38:0] _1053_;
wire [38:0] _1054_;
wire [38:0] _1055_;
wire [38:0] _1056_;
wire [38:0] _1057_;
wire [38:0] _1058_;
wire [38:0] _1059_;
wire [38:0] _1060_;
wire [38:0] _1061_;
wire [38:0] _1062_;
wire [38:0] _1063_;
wire [38:0] _1064_;
wire [38:0] _1065_;
wire [38:0] _1066_;
wire [38:0] _1067_;
wire [38:0] _1068_;
wire [38:0] _1069_;
wire [38:0] _1070_;
wire [38:0] _1071_;
wire [38:0] _1072_;
wire [38:0] _1073_;
wire [38:0] _1074_;
wire [38:0] _1075_;
wire [38:0] _1076_;
wire [38:0] _1077_;
wire [38:0] _1078_;
wire [38:0] _1079_;
wire [38:0] _1080_;
wire [38:0] _1081_;
wire [38:0] _1082_;
wire [38:0] _1083_;
wire [38:0] _1084_;
wire [38:0] _1085_;
wire [38:0] _1086_;
wire [38:0] _1087_;
wire [38:0] _1088_;
wire [38:0] _1089_;
wire [38:0] _1090_;
wire [38:0] _1091_;
wire [38:0] _1092_;
wire [38:0] _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire _1122_;
wire _1123_;
wire _1124_;
wire _1125_;
wire _1126_;
wire _1127_;
wire _1128_;
wire _1129_;
wire _1130_;
wire _1131_;
wire _1132_;
wire _1133_;
wire _1134_;
wire _1135_;
wire _1136_;
wire _1137_;
wire _1138_;
wire _1139_;
wire _1140_;
wire _1141_;
wire _1142_;
wire _1143_;
wire _1144_;
wire _1145_;
wire _1146_;
wire _1147_;
wire _1148_;
wire _1149_;
wire _1150_;
wire _1151_;
wire _1152_;
wire _1153_;
wire _1154_;
wire _1155_;
wire _1156_;
wire _1157_;
wire _1158_;
wire _1159_;
wire _1160_;
wire _1161_;
wire _1162_;
wire _1163_;
wire _1164_;
wire _1165_;
wire _1166_;
wire _1167_;
wire _1168_;
wire _1169_;
wire _1170_;
wire _1171_;
wire _1172_;
wire _1173_;
wire _1174_;
wire _1175_;
wire _1176_;
wire _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire _1181_;
wire _1182_;
wire _1183_;
wire _1184_;
wire _1185_;
wire _1186_;
wire [38:0] _1187_;
/* cellift = 32'd1 */
wire [38:0] _1188_;
wire [38:0] _1189_;
/* cellift = 32'd1 */
wire [38:0] _1190_;
wire [38:0] _1191_;
/* cellift = 32'd1 */
wire [38:0] _1192_;
wire [38:0] _1193_;
/* cellift = 32'd1 */
wire [38:0] _1194_;
wire [38:0] _1195_;
/* cellift = 32'd1 */
wire [38:0] _1196_;
wire [38:0] _1197_;
/* cellift = 32'd1 */
wire [38:0] _1198_;
wire [38:0] _1199_;
/* cellift = 32'd1 */
wire [38:0] _1200_;
wire [38:0] _1201_;
/* cellift = 32'd1 */
wire [38:0] _1202_;
wire [38:0] _1203_;
/* cellift = 32'd1 */
wire [38:0] _1204_;
wire [38:0] _1205_;
/* cellift = 32'd1 */
wire [38:0] _1206_;
wire [38:0] _1207_;
/* cellift = 32'd1 */
wire [38:0] _1208_;
wire [38:0] _1209_;
/* cellift = 32'd1 */
wire [38:0] _1210_;
wire [38:0] _1211_;
/* cellift = 32'd1 */
wire [38:0] _1212_;
wire [38:0] _1213_;
/* cellift = 32'd1 */
wire [38:0] _1214_;
wire [38:0] _1215_;
/* cellift = 32'd1 */
wire [38:0] _1216_;
wire [38:0] _1217_;
/* cellift = 32'd1 */
wire [38:0] _1218_;
wire [38:0] _1219_;
/* cellift = 32'd1 */
wire [38:0] _1220_;
wire [38:0] _1221_;
/* cellift = 32'd1 */
wire [38:0] _1222_;
wire [38:0] _1223_;
/* cellift = 32'd1 */
wire [38:0] _1224_;
wire [38:0] _1225_;
/* cellift = 32'd1 */
wire [38:0] _1226_;
wire [38:0] _1227_;
/* cellift = 32'd1 */
wire [38:0] _1228_;
wire [38:0] _1229_;
/* cellift = 32'd1 */
wire [38:0] _1230_;
wire [38:0] _1231_;
/* cellift = 32'd1 */
wire [38:0] _1232_;
wire [38:0] _1233_;
/* cellift = 32'd1 */
wire [38:0] _1234_;
wire [38:0] _1235_;
/* cellift = 32'd1 */
wire [38:0] _1236_;
wire [38:0] _1237_;
/* cellift = 32'd1 */
wire [38:0] _1238_;
wire [38:0] _1239_;
/* cellift = 32'd1 */
wire [38:0] _1240_;
wire [38:0] _1241_;
/* cellift = 32'd1 */
wire [38:0] _1242_;
wire [38:0] _1243_;
/* cellift = 32'd1 */
wire [38:0] _1244_;
wire [38:0] _1245_;
/* cellift = 32'd1 */
wire [38:0] _1246_;
wire [38:0] _1247_;
/* cellift = 32'd1 */
wire [38:0] _1248_;
wire [38:0] _1249_;
/* cellift = 32'd1 */
wire [38:0] _1250_;
wire [38:0] _1251_;
/* cellift = 32'd1 */
wire [38:0] _1252_;
wire [38:0] _1253_;
/* cellift = 32'd1 */
wire [38:0] _1254_;
wire [38:0] _1255_;
/* cellift = 32'd1 */
wire [38:0] _1256_;
wire [38:0] _1257_;
/* cellift = 32'd1 */
wire [38:0] _1258_;
wire [38:0] _1259_;
/* cellift = 32'd1 */
wire [38:0] _1260_;
wire [38:0] _1261_;
/* cellift = 32'd1 */
wire [38:0] _1262_;
wire [38:0] _1263_;
/* cellift = 32'd1 */
wire [38:0] _1264_;
wire [38:0] _1265_;
/* cellift = 32'd1 */
wire [38:0] _1266_;
wire [38:0] _1267_;
/* cellift = 32'd1 */
wire [38:0] _1268_;
wire [38:0] _1269_;
/* cellift = 32'd1 */
wire [38:0] _1270_;
wire [38:0] _1271_;
/* cellift = 32'd1 */
wire [38:0] _1272_;
wire [38:0] _1273_;
/* cellift = 32'd1 */
wire [38:0] _1274_;
wire [38:0] _1275_;
/* cellift = 32'd1 */
wire [38:0] _1276_;
wire [38:0] _1277_;
/* cellift = 32'd1 */
wire [38:0] _1278_;
wire [38:0] _1279_;
/* cellift = 32'd1 */
wire [38:0] _1280_;
wire [38:0] _1281_;
/* cellift = 32'd1 */
wire [38:0] _1282_;
wire [38:0] _1283_;
/* cellift = 32'd1 */
wire [38:0] _1284_;
wire [38:0] _1285_;
/* cellift = 32'd1 */
wire [38:0] _1286_;
wire [38:0] _1287_;
/* cellift = 32'd1 */
wire [38:0] _1288_;
wire [38:0] _1289_;
/* cellift = 32'd1 */
wire [38:0] _1290_;
wire [38:0] _1291_;
/* cellift = 32'd1 */
wire [38:0] _1292_;
wire [38:0] _1293_;
/* cellift = 32'd1 */
wire [38:0] _1294_;
wire [38:0] _1295_;
/* cellift = 32'd1 */
wire [38:0] _1296_;
wire [38:0] _1297_;
/* cellift = 32'd1 */
wire [38:0] _1298_;
wire [38:0] _1299_;
/* cellift = 32'd1 */
wire [38:0] _1300_;
wire [38:0] _1301_;
/* cellift = 32'd1 */
wire [38:0] _1302_;
wire [38:0] _1303_;
/* cellift = 32'd1 */
wire [38:0] _1304_;
wire [38:0] _1305_;
/* cellift = 32'd1 */
wire [38:0] _1306_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1307_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1308_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1309_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1310_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1311_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1312_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1313_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1314_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1315_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1316_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1317_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1318_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1319_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1320_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1321_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1322_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1323_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1324_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1325_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1326_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1327_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1328_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1329_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1330_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1331_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1332_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1333_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1334_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1335_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1336_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1337_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1338_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1339_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1340_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1341_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1342_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1343_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1344_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1345_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1346_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1347_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1348_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1349_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1350_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1351_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1352_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1353_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1354_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1355_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1356_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1357_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1358_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1359_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1360_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1361_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1362_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1363_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1364_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1365_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1366_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1367_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1368_;
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1369_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20074.20-20074.47" */
wire _1370_;
wire _1371_;
/* cellift = 32'd1 */
wire _1372_;
wire _1373_;
/* cellift = 32'd1 */
wire _1374_;
wire _1375_;
/* cellift = 32'd1 */
wire _1376_;
wire _1377_;
/* cellift = 32'd1 */
wire _1378_;
wire _1379_;
/* cellift = 32'd1 */
wire _1380_;
wire _1381_;
/* cellift = 32'd1 */
wire _1382_;
wire _1383_;
/* cellift = 32'd1 */
wire _1384_;
wire _1385_;
/* cellift = 32'd1 */
wire _1386_;
wire _1387_;
/* cellift = 32'd1 */
wire _1388_;
wire _1389_;
/* cellift = 32'd1 */
wire _1390_;
wire _1391_;
/* cellift = 32'd1 */
wire _1392_;
wire _1393_;
/* cellift = 32'd1 */
wire _1394_;
wire _1395_;
/* cellift = 32'd1 */
wire _1396_;
wire _1397_;
/* cellift = 32'd1 */
wire _1398_;
wire _1399_;
/* cellift = 32'd1 */
wire _1400_;
wire _1401_;
/* cellift = 32'd1 */
wire _1402_;
wire _1403_;
/* cellift = 32'd1 */
wire _1404_;
wire _1405_;
/* cellift = 32'd1 */
wire _1406_;
wire _1407_;
/* cellift = 32'd1 */
wire _1408_;
wire _1409_;
/* cellift = 32'd1 */
wire _1410_;
wire _1411_;
/* cellift = 32'd1 */
wire _1412_;
wire _1413_;
/* cellift = 32'd1 */
wire _1414_;
wire _1415_;
/* cellift = 32'd1 */
wire _1416_;
wire _1417_;
/* cellift = 32'd1 */
wire _1418_;
wire _1419_;
/* cellift = 32'd1 */
wire _1420_;
wire _1421_;
/* cellift = 32'd1 */
wire _1422_;
wire _1423_;
/* cellift = 32'd1 */
wire _1424_;
wire _1425_;
/* cellift = 32'd1 */
wire _1426_;
wire _1427_;
/* cellift = 32'd1 */
wire _1428_;
wire _1429_;
/* cellift = 32'd1 */
wire _1430_;
wire _1431_;
/* cellift = 32'd1 */
wire _1432_;
wire _1433_;
/* cellift = 32'd1 */
wire _1434_;
wire _1435_;
/* cellift = 32'd1 */
wire _1436_;
wire _1437_;
/* cellift = 32'd1 */
wire _1438_;
wire _1439_;
/* cellift = 32'd1 */
wire _1440_;
wire _1441_;
/* cellift = 32'd1 */
wire _1442_;
wire _1443_;
/* cellift = 32'd1 */
wire _1444_;
wire _1445_;
/* cellift = 32'd1 */
wire _1446_;
wire _1447_;
/* cellift = 32'd1 */
wire _1448_;
wire _1449_;
/* cellift = 32'd1 */
wire _1450_;
wire _1451_;
/* cellift = 32'd1 */
wire _1452_;
wire _1453_;
/* cellift = 32'd1 */
wire _1454_;
wire _1455_;
/* cellift = 32'd1 */
wire _1456_;
wire _1457_;
/* cellift = 32'd1 */
wire _1458_;
wire _1459_;
/* cellift = 32'd1 */
wire _1460_;
wire _1461_;
/* cellift = 32'd1 */
wire _1462_;
wire _1463_;
/* cellift = 32'd1 */
wire _1464_;
wire _1465_;
/* cellift = 32'd1 */
wire _1466_;
wire _1467_;
/* cellift = 32'd1 */
wire _1468_;
wire _1469_;
/* cellift = 32'd1 */
wire _1470_;
wire _1471_;
/* cellift = 32'd1 */
wire _1472_;
wire _1473_;
/* cellift = 32'd1 */
wire _1474_;
wire _1475_;
/* cellift = 32'd1 */
wire _1476_;
wire _1477_;
/* cellift = 32'd1 */
wire _1478_;
wire _1479_;
/* cellift = 32'd1 */
wire _1480_;
wire _1481_;
/* cellift = 32'd1 */
wire _1482_;
wire _1483_;
/* cellift = 32'd1 */
wire _1484_;
wire _1485_;
/* cellift = 32'd1 */
wire _1486_;
wire _1487_;
/* cellift = 32'd1 */
wire _1488_;
wire _1489_;
/* cellift = 32'd1 */
wire _1490_;
wire _1491_;
/* cellift = 32'd1 */
wire _1492_;
wire _1493_;
/* cellift = 32'd1 */
wire _1494_;
/* src = "generated/sv2v_out.v:20049.13-20049.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:20052.13-20052.29" */
input dummy_instr_id_i;
wire dummy_instr_id_i;
/* cellift = 32'd1 */
input dummy_instr_id_i_t0;
wire dummy_instr_id_i_t0;
/* src = "generated/sv2v_out.v:20053.13-20053.29" */
input dummy_instr_wb_i;
wire dummy_instr_wb_i;
/* cellift = 32'd1 */
input dummy_instr_wb_i_t0;
wire dummy_instr_wb_i_t0;
/* src = "generated/sv2v_out.v:20061.14-20061.19" */
output err_o;
wire err_o;
/* cellift = 32'd1 */
output err_o_t0;
wire err_o_t0;
/* src = "generated/sv2v_out.v:20116.26-20116.33" */
reg [38:0] \g_dummy_r0.rf_r0_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20116.26-20116.33" */
reg [38:0] \g_dummy_r0.rf_r0_q_t0 ;
/* src = "generated/sv2v_out.v:20115.9-20115.20" */
wire \g_dummy_r0.we_r0_dummy ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20115.9-20115.20" */
wire \g_dummy_r0.we_r0_dummy_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[10].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[10].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[11].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[11].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[12].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[12].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[13].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[13].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[14].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[14].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[15].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[15].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[16].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[16].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[17].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[17].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[18].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[18].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[19].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[19].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[1].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[1].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[20].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[20].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[21].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[21].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[22].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[22].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[23].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[23].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[24].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[24].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[25].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[25].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[26].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[26].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[27].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[27].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[28].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[28].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[29].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[29].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[2].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[2].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[30].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[30].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[31].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[31].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[3].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[3].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[4].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[4].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[5].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[5].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[6].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[6].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[7].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[7].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[8].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[8].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[9].rf_reg_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20106.26-20106.34" */
reg [38:0] \g_rf_flops[9].rf_reg_q_t0 ;
/* src = "generated/sv2v_out.v:20079.27-20079.39" */
wire [31:0] \gen_wren_check.we_a_dec_buf ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20079.27-20079.39" */
wire [31:0] \gen_wren_check.we_a_dec_buf_t0 ;
/* src = "generated/sv2v_out.v:20054.19-20054.28" */
input [4:0] raddr_a_i;
wire [4:0] raddr_a_i;
/* cellift = 32'd1 */
input [4:0] raddr_a_i_t0;
wire [4:0] raddr_a_i_t0;
/* src = "generated/sv2v_out.v:20056.19-20056.28" */
input [4:0] raddr_b_i;
wire [4:0] raddr_b_i;
/* cellift = 32'd1 */
input [4:0] raddr_b_i_t0;
wire [4:0] raddr_b_i_t0;
/* src = "generated/sv2v_out.v:20055.32-20055.41" */
output [38:0] rdata_a_o;
wire [38:0] rdata_a_o;
/* cellift = 32'd1 */
output [38:0] rdata_a_o_t0;
wire [38:0] rdata_a_o_t0;
/* src = "generated/sv2v_out.v:20057.32-20057.41" */
output [38:0] rdata_b_o;
wire [38:0] rdata_b_o;
/* cellift = 32'd1 */
output [38:0] rdata_b_o_t0;
wire [38:0] rdata_b_o_t0;
/* src = "generated/sv2v_out.v:20064.25-20064.31" */
wire [38:0] \rf_reg[0] ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20064.25-20064.31" */
wire [38:0] \rf_reg[0]_t0 ;
/* src = "generated/sv2v_out.v:20050.13-20050.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:20051.13-20051.22" */
input test_en_i;
wire test_en_i;
/* cellift = 32'd1 */
input test_en_i_t0;
wire test_en_i_t0;
/* src = "generated/sv2v_out.v:20058.19-20058.28" */
input [4:0] waddr_a_i;
wire [4:0] waddr_a_i;
/* cellift = 32'd1 */
input [4:0] waddr_a_i_t0;
wire [4:0] waddr_a_i_t0;
/* src = "generated/sv2v_out.v:20059.31-20059.40" */
input [38:0] wdata_a_i;
wire [38:0] wdata_a_i;
/* cellift = 32'd1 */
input [38:0] wdata_a_i_t0;
wire [38:0] wdata_a_i_t0;
/* src = "generated/sv2v_out.v:20065.24-20065.32" */
wire [31:0] we_a_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20065.24-20065.32" */
wire [31:0] we_a_dec_t0;
/* src = "generated/sv2v_out.v:20060.13-20060.19" */
input we_a_i;
wire we_a_i;
/* cellift = 32'd1 */
input we_a_i_t0;
wire we_a_i_t0;
assign \g_dummy_r0.we_r0_dummy  = we_a_i & /* src = "generated/sv2v_out.v:20117.25-20117.50" */ dummy_instr_wb_i;
assign _0000_ = ~ we_a_dec[31];
assign _0001_ = ~ we_a_dec[30];
assign _0002_ = ~ we_a_dec[29];
assign _0003_ = ~ we_a_dec[28];
assign _0004_ = ~ we_a_dec[27];
assign _0005_ = ~ we_a_dec[26];
assign _0006_ = ~ we_a_dec[25];
assign _0007_ = ~ we_a_dec[24];
assign _0008_ = ~ we_a_dec[23];
assign _0009_ = ~ we_a_dec[22];
assign _0010_ = ~ we_a_dec[21];
assign _0011_ = ~ we_a_dec[20];
assign _0012_ = ~ we_a_dec[19];
assign _0013_ = ~ we_a_dec[18];
assign _0014_ = ~ we_a_dec[17];
assign _0015_ = ~ we_a_dec[16];
assign _0016_ = ~ we_a_dec[15];
assign _0017_ = ~ we_a_dec[14];
assign _0018_ = ~ we_a_dec[13];
assign _0019_ = ~ we_a_dec[12];
assign _0020_ = ~ we_a_dec[11];
assign _0021_ = ~ we_a_dec[10];
assign _0022_ = ~ we_a_dec[9];
assign _0023_ = ~ we_a_dec[8];
assign _0024_ = ~ we_a_dec[7];
assign _0025_ = ~ we_a_dec[6];
assign _0026_ = ~ we_a_dec[5];
assign _0027_ = ~ we_a_dec[4];
assign _0028_ = ~ we_a_dec[3];
assign _0029_ = ~ we_a_dec[2];
assign _0030_ = ~ we_a_dec[1];
assign _0031_ = ~ \g_dummy_r0.we_r0_dummy ;
assign _1016_ = wdata_a_i ^ \g_rf_flops[31].rf_reg_q ;
assign _1017_ = wdata_a_i ^ \g_rf_flops[30].rf_reg_q ;
assign _1018_ = wdata_a_i ^ \g_rf_flops[29].rf_reg_q ;
assign _1019_ = wdata_a_i ^ \g_rf_flops[28].rf_reg_q ;
assign _1020_ = wdata_a_i ^ \g_rf_flops[27].rf_reg_q ;
assign _1021_ = wdata_a_i ^ \g_rf_flops[26].rf_reg_q ;
assign _1022_ = wdata_a_i ^ \g_rf_flops[25].rf_reg_q ;
assign _1023_ = wdata_a_i ^ \g_rf_flops[24].rf_reg_q ;
assign _1024_ = wdata_a_i ^ \g_rf_flops[23].rf_reg_q ;
assign _1025_ = wdata_a_i ^ \g_rf_flops[22].rf_reg_q ;
assign _1026_ = wdata_a_i ^ \g_rf_flops[21].rf_reg_q ;
assign _1027_ = wdata_a_i ^ \g_rf_flops[20].rf_reg_q ;
assign _1028_ = wdata_a_i ^ \g_rf_flops[19].rf_reg_q ;
assign _1029_ = wdata_a_i ^ \g_rf_flops[18].rf_reg_q ;
assign _1030_ = wdata_a_i ^ \g_rf_flops[17].rf_reg_q ;
assign _1031_ = wdata_a_i ^ \g_rf_flops[16].rf_reg_q ;
assign _1032_ = wdata_a_i ^ \g_rf_flops[15].rf_reg_q ;
assign _1033_ = wdata_a_i ^ \g_rf_flops[14].rf_reg_q ;
assign _1034_ = wdata_a_i ^ \g_rf_flops[13].rf_reg_q ;
assign _1035_ = wdata_a_i ^ \g_rf_flops[12].rf_reg_q ;
assign _1036_ = wdata_a_i ^ \g_rf_flops[11].rf_reg_q ;
assign _1037_ = wdata_a_i ^ \g_rf_flops[10].rf_reg_q ;
assign _1038_ = wdata_a_i ^ \g_rf_flops[9].rf_reg_q ;
assign _1039_ = wdata_a_i ^ \g_rf_flops[8].rf_reg_q ;
assign _1040_ = wdata_a_i ^ \g_rf_flops[7].rf_reg_q ;
assign _1041_ = wdata_a_i ^ \g_rf_flops[6].rf_reg_q ;
assign _1042_ = wdata_a_i ^ \g_rf_flops[5].rf_reg_q ;
assign _1043_ = wdata_a_i ^ \g_rf_flops[4].rf_reg_q ;
assign _1044_ = wdata_a_i ^ \g_rf_flops[3].rf_reg_q ;
assign _1045_ = wdata_a_i ^ \g_rf_flops[2].rf_reg_q ;
assign _1046_ = wdata_a_i ^ \g_rf_flops[1].rf_reg_q ;
assign _1047_ = wdata_a_i ^ \g_dummy_r0.rf_r0_q ;
assign _0621_ = wdata_a_i_t0 | \g_rf_flops[31].rf_reg_q_t0 ;
assign _0625_ = wdata_a_i_t0 | \g_rf_flops[30].rf_reg_q_t0 ;
assign _0629_ = wdata_a_i_t0 | \g_rf_flops[29].rf_reg_q_t0 ;
assign _0633_ = wdata_a_i_t0 | \g_rf_flops[28].rf_reg_q_t0 ;
assign _0637_ = wdata_a_i_t0 | \g_rf_flops[27].rf_reg_q_t0 ;
assign _0641_ = wdata_a_i_t0 | \g_rf_flops[26].rf_reg_q_t0 ;
assign _0645_ = wdata_a_i_t0 | \g_rf_flops[25].rf_reg_q_t0 ;
assign _0649_ = wdata_a_i_t0 | \g_rf_flops[24].rf_reg_q_t0 ;
assign _0653_ = wdata_a_i_t0 | \g_rf_flops[23].rf_reg_q_t0 ;
assign _0657_ = wdata_a_i_t0 | \g_rf_flops[22].rf_reg_q_t0 ;
assign _0661_ = wdata_a_i_t0 | \g_rf_flops[21].rf_reg_q_t0 ;
assign _0665_ = wdata_a_i_t0 | \g_rf_flops[20].rf_reg_q_t0 ;
assign _0669_ = wdata_a_i_t0 | \g_rf_flops[19].rf_reg_q_t0 ;
assign _0673_ = wdata_a_i_t0 | \g_rf_flops[18].rf_reg_q_t0 ;
assign _0677_ = wdata_a_i_t0 | \g_rf_flops[17].rf_reg_q_t0 ;
assign _0681_ = wdata_a_i_t0 | \g_rf_flops[16].rf_reg_q_t0 ;
assign _0685_ = wdata_a_i_t0 | \g_rf_flops[15].rf_reg_q_t0 ;
assign _0689_ = wdata_a_i_t0 | \g_rf_flops[14].rf_reg_q_t0 ;
assign _0693_ = wdata_a_i_t0 | \g_rf_flops[13].rf_reg_q_t0 ;
assign _0697_ = wdata_a_i_t0 | \g_rf_flops[12].rf_reg_q_t0 ;
assign _0701_ = wdata_a_i_t0 | \g_rf_flops[11].rf_reg_q_t0 ;
assign _0705_ = wdata_a_i_t0 | \g_rf_flops[10].rf_reg_q_t0 ;
assign _0709_ = wdata_a_i_t0 | \g_rf_flops[9].rf_reg_q_t0 ;
assign _0713_ = wdata_a_i_t0 | \g_rf_flops[8].rf_reg_q_t0 ;
assign _0717_ = wdata_a_i_t0 | \g_rf_flops[7].rf_reg_q_t0 ;
assign _0721_ = wdata_a_i_t0 | \g_rf_flops[6].rf_reg_q_t0 ;
assign _0725_ = wdata_a_i_t0 | \g_rf_flops[5].rf_reg_q_t0 ;
assign _0729_ = wdata_a_i_t0 | \g_rf_flops[4].rf_reg_q_t0 ;
assign _0733_ = wdata_a_i_t0 | \g_rf_flops[3].rf_reg_q_t0 ;
assign _0737_ = wdata_a_i_t0 | \g_rf_flops[2].rf_reg_q_t0 ;
assign _0741_ = wdata_a_i_t0 | \g_rf_flops[1].rf_reg_q_t0 ;
assign _0745_ = wdata_a_i_t0 | \g_dummy_r0.rf_r0_q_t0 ;
assign _0622_ = _1016_ | _0621_;
assign _0626_ = _1017_ | _0625_;
assign _0630_ = _1018_ | _0629_;
assign _0634_ = _1019_ | _0633_;
assign _0638_ = _1020_ | _0637_;
assign _0642_ = _1021_ | _0641_;
assign _0646_ = _1022_ | _0645_;
assign _0650_ = _1023_ | _0649_;
assign _0654_ = _1024_ | _0653_;
assign _0658_ = _1025_ | _0657_;
assign _0662_ = _1026_ | _0661_;
assign _0666_ = _1027_ | _0665_;
assign _0670_ = _1028_ | _0669_;
assign _0674_ = _1029_ | _0673_;
assign _0678_ = _1030_ | _0677_;
assign _0682_ = _1031_ | _0681_;
assign _0686_ = _1032_ | _0685_;
assign _0690_ = _1033_ | _0689_;
assign _0694_ = _1034_ | _0693_;
assign _0698_ = _1035_ | _0697_;
assign _0702_ = _1036_ | _0701_;
assign _0706_ = _1037_ | _0705_;
assign _0710_ = _1038_ | _0709_;
assign _0714_ = _1039_ | _0713_;
assign _0718_ = _1040_ | _0717_;
assign _0722_ = _1041_ | _0721_;
assign _0726_ = _1042_ | _0725_;
assign _0730_ = _1043_ | _0729_;
assign _0734_ = _1044_ | _0733_;
assign _0738_ = _1045_ | _0737_;
assign _0742_ = _1046_ | _0741_;
assign _0746_ = _1047_ | _0745_;
assign _0207_ = { we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31], we_a_dec[31] } & wdata_a_i_t0;
assign _0210_ = { we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30], we_a_dec[30] } & wdata_a_i_t0;
assign _0213_ = { we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29], we_a_dec[29] } & wdata_a_i_t0;
assign _0216_ = { we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28], we_a_dec[28] } & wdata_a_i_t0;
assign _0219_ = { we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27], we_a_dec[27] } & wdata_a_i_t0;
assign _0222_ = { we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26], we_a_dec[26] } & wdata_a_i_t0;
assign _0225_ = { we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25], we_a_dec[25] } & wdata_a_i_t0;
assign _0228_ = { we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24], we_a_dec[24] } & wdata_a_i_t0;
assign _0231_ = { we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23], we_a_dec[23] } & wdata_a_i_t0;
assign _0234_ = { we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22], we_a_dec[22] } & wdata_a_i_t0;
assign _0237_ = { we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21], we_a_dec[21] } & wdata_a_i_t0;
assign _0240_ = { we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20], we_a_dec[20] } & wdata_a_i_t0;
assign _0243_ = { we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19], we_a_dec[19] } & wdata_a_i_t0;
assign _0246_ = { we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18], we_a_dec[18] } & wdata_a_i_t0;
assign _0249_ = { we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17], we_a_dec[17] } & wdata_a_i_t0;
assign _0252_ = { we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16], we_a_dec[16] } & wdata_a_i_t0;
assign _0255_ = { we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15], we_a_dec[15] } & wdata_a_i_t0;
assign _0258_ = { we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14], we_a_dec[14] } & wdata_a_i_t0;
assign _0261_ = { we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13], we_a_dec[13] } & wdata_a_i_t0;
assign _0264_ = { we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12], we_a_dec[12] } & wdata_a_i_t0;
assign _0267_ = { we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11], we_a_dec[11] } & wdata_a_i_t0;
assign _0270_ = { we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10], we_a_dec[10] } & wdata_a_i_t0;
assign _0273_ = { we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9], we_a_dec[9] } & wdata_a_i_t0;
assign _0276_ = { we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8], we_a_dec[8] } & wdata_a_i_t0;
assign _0279_ = { we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7], we_a_dec[7] } & wdata_a_i_t0;
assign _0282_ = { we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6], we_a_dec[6] } & wdata_a_i_t0;
assign _0285_ = { we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5], we_a_dec[5] } & wdata_a_i_t0;
assign _0288_ = { we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4], we_a_dec[4] } & wdata_a_i_t0;
assign _0291_ = { we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3], we_a_dec[3] } & wdata_a_i_t0;
assign _0294_ = { we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2], we_a_dec[2] } & wdata_a_i_t0;
assign _0297_ = { we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1], we_a_dec[1] } & wdata_a_i_t0;
assign _0300_ = { \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy , \g_dummy_r0.we_r0_dummy  } & wdata_a_i_t0;
assign _0208_ = { _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_, _0000_ } & \g_rf_flops[31].rf_reg_q_t0 ;
assign _0211_ = { _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_, _0001_ } & \g_rf_flops[30].rf_reg_q_t0 ;
assign _0214_ = { _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_, _0002_ } & \g_rf_flops[29].rf_reg_q_t0 ;
assign _0217_ = { _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_, _0003_ } & \g_rf_flops[28].rf_reg_q_t0 ;
assign _0220_ = { _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_ } & \g_rf_flops[27].rf_reg_q_t0 ;
assign _0223_ = { _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_, _0005_ } & \g_rf_flops[26].rf_reg_q_t0 ;
assign _0226_ = { _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_, _0006_ } & \g_rf_flops[25].rf_reg_q_t0 ;
assign _0229_ = { _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_, _0007_ } & \g_rf_flops[24].rf_reg_q_t0 ;
assign _0232_ = { _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_, _0008_ } & \g_rf_flops[23].rf_reg_q_t0 ;
assign _0235_ = { _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_, _0009_ } & \g_rf_flops[22].rf_reg_q_t0 ;
assign _0238_ = { _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_, _0010_ } & \g_rf_flops[21].rf_reg_q_t0 ;
assign _0241_ = { _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_, _0011_ } & \g_rf_flops[20].rf_reg_q_t0 ;
assign _0244_ = { _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_, _0012_ } & \g_rf_flops[19].rf_reg_q_t0 ;
assign _0247_ = { _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_, _0013_ } & \g_rf_flops[18].rf_reg_q_t0 ;
assign _0250_ = { _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_, _0014_ } & \g_rf_flops[17].rf_reg_q_t0 ;
assign _0253_ = { _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_, _0015_ } & \g_rf_flops[16].rf_reg_q_t0 ;
assign _0256_ = { _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_, _0016_ } & \g_rf_flops[15].rf_reg_q_t0 ;
assign _0259_ = { _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_, _0017_ } & \g_rf_flops[14].rf_reg_q_t0 ;
assign _0262_ = { _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_, _0018_ } & \g_rf_flops[13].rf_reg_q_t0 ;
assign _0265_ = { _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_, _0019_ } & \g_rf_flops[12].rf_reg_q_t0 ;
assign _0268_ = { _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_, _0020_ } & \g_rf_flops[11].rf_reg_q_t0 ;
assign _0271_ = { _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_, _0021_ } & \g_rf_flops[10].rf_reg_q_t0 ;
assign _0274_ = { _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_, _0022_ } & \g_rf_flops[9].rf_reg_q_t0 ;
assign _0277_ = { _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_, _0023_ } & \g_rf_flops[8].rf_reg_q_t0 ;
assign _0280_ = { _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_, _0024_ } & \g_rf_flops[7].rf_reg_q_t0 ;
assign _0283_ = { _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_, _0025_ } & \g_rf_flops[6].rf_reg_q_t0 ;
assign _0286_ = { _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_, _0026_ } & \g_rf_flops[5].rf_reg_q_t0 ;
assign _0289_ = { _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_, _0027_ } & \g_rf_flops[4].rf_reg_q_t0 ;
assign _0292_ = { _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_ } & \g_rf_flops[3].rf_reg_q_t0 ;
assign _0295_ = { _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_, _0029_ } & \g_rf_flops[2].rf_reg_q_t0 ;
assign _0298_ = { _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_, _0030_ } & \g_rf_flops[1].rf_reg_q_t0 ;
assign _0301_ = { _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_, _0031_ } & \g_dummy_r0.rf_r0_q_t0 ;
assign _0209_ = _0622_ & { we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31], we_a_dec_t0[31] };
assign _0212_ = _0626_ & { we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30], we_a_dec_t0[30] };
assign _0215_ = _0630_ & { we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29], we_a_dec_t0[29] };
assign _0218_ = _0634_ & { we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28], we_a_dec_t0[28] };
assign _0221_ = _0638_ & { we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27], we_a_dec_t0[27] };
assign _0224_ = _0642_ & { we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26], we_a_dec_t0[26] };
assign _0227_ = _0646_ & { we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25], we_a_dec_t0[25] };
assign _0230_ = _0650_ & { we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24], we_a_dec_t0[24] };
assign _0233_ = _0654_ & { we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23], we_a_dec_t0[23] };
assign _0236_ = _0658_ & { we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22], we_a_dec_t0[22] };
assign _0239_ = _0662_ & { we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21], we_a_dec_t0[21] };
assign _0242_ = _0666_ & { we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20], we_a_dec_t0[20] };
assign _0245_ = _0670_ & { we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19], we_a_dec_t0[19] };
assign _0248_ = _0674_ & { we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18], we_a_dec_t0[18] };
assign _0251_ = _0678_ & { we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17], we_a_dec_t0[17] };
assign _0254_ = _0682_ & { we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16], we_a_dec_t0[16] };
assign _0257_ = _0686_ & { we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15], we_a_dec_t0[15] };
assign _0260_ = _0690_ & { we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14], we_a_dec_t0[14] };
assign _0263_ = _0694_ & { we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13], we_a_dec_t0[13] };
assign _0266_ = _0698_ & { we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12], we_a_dec_t0[12] };
assign _0269_ = _0702_ & { we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11], we_a_dec_t0[11] };
assign _0272_ = _0706_ & { we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10], we_a_dec_t0[10] };
assign _0275_ = _0710_ & { we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9], we_a_dec_t0[9] };
assign _0278_ = _0714_ & { we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8], we_a_dec_t0[8] };
assign _0281_ = _0718_ & { we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7], we_a_dec_t0[7] };
assign _0284_ = _0722_ & { we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6], we_a_dec_t0[6] };
assign _0287_ = _0726_ & { we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5], we_a_dec_t0[5] };
assign _0290_ = _0730_ & { we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4], we_a_dec_t0[4] };
assign _0293_ = _0734_ & { we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3], we_a_dec_t0[3] };
assign _0296_ = _0738_ & { we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2], we_a_dec_t0[2] };
assign _0299_ = _0742_ & { we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1], we_a_dec_t0[1] };
assign _0302_ = _0746_ & { \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0 , \g_dummy_r0.we_r0_dummy_t0  };
assign _0623_ = _0207_ | _0208_;
assign _0627_ = _0210_ | _0211_;
assign _0631_ = _0213_ | _0214_;
assign _0635_ = _0216_ | _0217_;
assign _0639_ = _0219_ | _0220_;
assign _0643_ = _0222_ | _0223_;
assign _0647_ = _0225_ | _0226_;
assign _0651_ = _0228_ | _0229_;
assign _0655_ = _0231_ | _0232_;
assign _0659_ = _0234_ | _0235_;
assign _0663_ = _0237_ | _0238_;
assign _0667_ = _0240_ | _0241_;
assign _0671_ = _0243_ | _0244_;
assign _0675_ = _0246_ | _0247_;
assign _0679_ = _0249_ | _0250_;
assign _0683_ = _0252_ | _0253_;
assign _0687_ = _0255_ | _0256_;
assign _0691_ = _0258_ | _0259_;
assign _0695_ = _0261_ | _0262_;
assign _0699_ = _0264_ | _0265_;
assign _0703_ = _0267_ | _0268_;
assign _0707_ = _0270_ | _0271_;
assign _0711_ = _0273_ | _0274_;
assign _0715_ = _0276_ | _0277_;
assign _0719_ = _0279_ | _0280_;
assign _0723_ = _0282_ | _0283_;
assign _0727_ = _0285_ | _0286_;
assign _0731_ = _0288_ | _0289_;
assign _0735_ = _0291_ | _0292_;
assign _0739_ = _0294_ | _0295_;
assign _0743_ = _0297_ | _0298_;
assign _0747_ = _0300_ | _0301_;
assign _0624_ = _0623_ | _0209_;
assign _0628_ = _0627_ | _0212_;
assign _0632_ = _0631_ | _0215_;
assign _0636_ = _0635_ | _0218_;
assign _0640_ = _0639_ | _0221_;
assign _0644_ = _0643_ | _0224_;
assign _0648_ = _0647_ | _0227_;
assign _0652_ = _0651_ | _0230_;
assign _0656_ = _0655_ | _0233_;
assign _0660_ = _0659_ | _0236_;
assign _0664_ = _0663_ | _0239_;
assign _0668_ = _0667_ | _0242_;
assign _0672_ = _0671_ | _0245_;
assign _0676_ = _0675_ | _0248_;
assign _0680_ = _0679_ | _0251_;
assign _0684_ = _0683_ | _0254_;
assign _0688_ = _0687_ | _0257_;
assign _0692_ = _0691_ | _0260_;
assign _0696_ = _0695_ | _0263_;
assign _0700_ = _0699_ | _0266_;
assign _0704_ = _0703_ | _0269_;
assign _0708_ = _0707_ | _0272_;
assign _0712_ = _0711_ | _0275_;
assign _0716_ = _0715_ | _0278_;
assign _0720_ = _0719_ | _0281_;
assign _0724_ = _0723_ | _0284_;
assign _0728_ = _0727_ | _0287_;
assign _0732_ = _0731_ | _0290_;
assign _0736_ = _0735_ | _0293_;
assign _0740_ = _0739_ | _0296_;
assign _0744_ = _0743_ | _0299_;
assign _0748_ = _0747_ | _0302_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[31].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[31].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[31].rf_reg_q_t0  <= _0624_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[30].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[30].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[30].rf_reg_q_t0  <= _0628_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[29].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[29].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[29].rf_reg_q_t0  <= _0632_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[28].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[28].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[28].rf_reg_q_t0  <= _0636_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[27].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[27].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[27].rf_reg_q_t0  <= _0640_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[26].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[26].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[26].rf_reg_q_t0  <= _0644_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[25].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[25].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[25].rf_reg_q_t0  <= _0648_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[24].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[24].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[24].rf_reg_q_t0  <= _0652_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[23].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[23].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[23].rf_reg_q_t0  <= _0656_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[22].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[22].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[22].rf_reg_q_t0  <= _0660_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[21].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[21].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[21].rf_reg_q_t0  <= _0664_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[20].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[20].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[20].rf_reg_q_t0  <= _0668_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[19].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[19].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[19].rf_reg_q_t0  <= _0672_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[18].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[18].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[18].rf_reg_q_t0  <= _0676_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[17].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[17].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[17].rf_reg_q_t0  <= _0680_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[16].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[16].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[16].rf_reg_q_t0  <= _0684_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[15].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[15].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[15].rf_reg_q_t0  <= _0688_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[14].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[14].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[14].rf_reg_q_t0  <= _0692_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[13].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[13].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[13].rf_reg_q_t0  <= _0696_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[12].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[12].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[12].rf_reg_q_t0  <= _0700_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[11].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[11].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[11].rf_reg_q_t0  <= _0704_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[10].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[10].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[10].rf_reg_q_t0  <= _0708_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[9].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[9].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[9].rf_reg_q_t0  <= _0712_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[8].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[8].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[8].rf_reg_q_t0  <= _0716_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[7].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[7].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[7].rf_reg_q_t0  <= _0720_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[6].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[6].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[6].rf_reg_q_t0  <= _0724_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[5].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[5].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[5].rf_reg_q_t0  <= _0728_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[4].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[4].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[4].rf_reg_q_t0  <= _0732_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[3].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[3].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[3].rf_reg_q_t0  <= _0736_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[2].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[2].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[2].rf_reg_q_t0  <= _0740_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[1].rf_reg_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[1].rf_reg_q_t0  <= 39'h0000000000;
else \g_rf_flops[1].rf_reg_q_t0  <= _0744_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_dummy_r0.rf_r0_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_dummy_r0.rf_r0_q_t0  <= 39'h0000000000;
else \g_dummy_r0.rf_r0_q_t0  <= _0748_;
assign _0204_ = we_a_i_t0 & dummy_instr_wb_i;
assign _0205_ = dummy_instr_wb_i_t0 & we_a_i;
assign _0206_ = we_a_i_t0 & dummy_instr_wb_i_t0;
assign _0620_ = _0204_ | _0205_;
assign \g_dummy_r0.we_r0_dummy_t0  = _0620_ | _0206_;
assign _0033_ = | raddr_b_i_t0;
assign _0034_ = | raddr_a_i_t0;
assign _0035_ = ~ waddr_a_i_t0;
assign _0036_ = ~ raddr_b_i_t0;
assign _0037_ = ~ raddr_a_i_t0;
assign _0551_ = waddr_a_i & _0035_;
assign _0552_ = raddr_b_i & _0036_;
assign _0553_ = raddr_a_i & _0037_;
assign _1094_ = _0551_ == { 4'h0, _0035_[0] };
assign _1095_ = _0551_ == { 3'h0, _0035_[1], 1'h0 };
assign _1096_ = _0551_ == { 3'h0, _0035_[1:0] };
assign _1097_ = _0551_ == { 2'h0, _0035_[2], 2'h0 };
assign _1098_ = _0551_ == { 2'h0, _0035_[2], 1'h0, _0035_[0] };
assign _1099_ = _0551_ == { 2'h0, _0035_[2:1], 1'h0 };
assign _1100_ = _0551_ == { 2'h0, _0035_[2:0] };
assign _1101_ = _0551_ == { 1'h0, _0035_[3], 3'h0 };
assign _1102_ = _0551_ == { 1'h0, _0035_[3], 2'h0, _0035_[0] };
assign _1103_ = _0551_ == { 1'h0, _0035_[3], 1'h0, _0035_[1], 1'h0 };
assign _1104_ = _0551_ == { 1'h0, _0035_[3], 1'h0, _0035_[1:0] };
assign _1105_ = _0551_ == { 1'h0, _0035_[3:2], 2'h0 };
assign _1106_ = _0551_ == { 1'h0, _0035_[3:2], 1'h0, _0035_[0] };
assign _1107_ = _0551_ == { 1'h0, _0035_[3:1], 1'h0 };
assign _1108_ = _0551_ == { 1'h0, _0035_[3:0] };
assign _1109_ = _0551_ == { _0035_[4], 4'h0 };
assign _1110_ = _0551_ == { _0035_[4], 3'h0, _0035_[0] };
assign _1111_ = _0551_ == { _0035_[4], 2'h0, _0035_[1], 1'h0 };
assign _1112_ = _0551_ == { _0035_[4], 2'h0, _0035_[1:0] };
assign _1113_ = _0551_ == { _0035_[4], 1'h0, _0035_[2], 2'h0 };
assign _1114_ = _0551_ == { _0035_[4], 1'h0, _0035_[2], 1'h0, _0035_[0] };
assign _1115_ = _0551_ == { _0035_[4], 1'h0, _0035_[2:1], 1'h0 };
assign _1116_ = _0551_ == { _0035_[4], 1'h0, _0035_[2:0] };
assign _1117_ = _0551_ == { _0035_[4:3], 3'h0 };
assign _1118_ = _0551_ == { _0035_[4:3], 2'h0, _0035_[0] };
assign _1119_ = _0551_ == { _0035_[4:3], 1'h0, _0035_[1], 1'h0 };
assign _1120_ = _0551_ == { _0035_[4:3], 1'h0, _0035_[1:0] };
assign _1121_ = _0551_ == { _0035_[4:2], 2'h0 };
assign _1122_ = _0551_ == { _0035_[4:2], 1'h0, _0035_[0] };
assign _1123_ = _0551_ == { _0035_[4:1], 1'h0 };
assign _1124_ = _0551_ == _0035_;
assign _1125_ = _0552_ == _0036_;
assign _1126_ = _0552_ == { _0036_[4:1], 1'h0 };
assign _1127_ = _0552_ == { _0036_[4:2], 1'h0, _0036_[0] };
assign _1128_ = _0552_ == { _0036_[4:2], 2'h0 };
assign _1129_ = _0552_ == { _0036_[4:3], 1'h0, _0036_[1:0] };
assign _1130_ = _0552_ == { _0036_[4:3], 1'h0, _0036_[1], 1'h0 };
assign _1131_ = _0552_ == { _0036_[4:3], 2'h0, _0036_[0] };
assign _1132_ = _0552_ == { _0036_[4:3], 3'h0 };
assign _1133_ = _0552_ == { _0036_[4], 1'h0, _0036_[2:0] };
assign _1134_ = _0552_ == { _0036_[4], 1'h0, _0036_[2:1], 1'h0 };
assign _1135_ = _0552_ == { _0036_[4], 1'h0, _0036_[2], 1'h0, _0036_[0] };
assign _1136_ = _0552_ == { _0036_[4], 1'h0, _0036_[2], 2'h0 };
assign _1137_ = _0552_ == { _0036_[4], 2'h0, _0036_[1:0] };
assign _1138_ = _0552_ == { _0036_[4], 2'h0, _0036_[1], 1'h0 };
assign _1139_ = _0552_ == { _0036_[4], 3'h0, _0036_[0] };
assign _1140_ = _0552_ == { _0036_[4], 4'h0 };
assign _1141_ = _0552_ == { 1'h0, _0036_[3:0] };
assign _1142_ = _0552_ == { 1'h0, _0036_[3:1], 1'h0 };
assign _1143_ = _0552_ == { 1'h0, _0036_[3:2], 1'h0, _0036_[0] };
assign _1144_ = _0552_ == { 1'h0, _0036_[3:2], 2'h0 };
assign _1145_ = _0552_ == { 1'h0, _0036_[3], 1'h0, _0036_[1:0] };
assign _1146_ = _0552_ == { 1'h0, _0036_[3], 1'h0, _0036_[1], 1'h0 };
assign _1147_ = _0552_ == { 1'h0, _0036_[3], 2'h0, _0036_[0] };
assign _1148_ = _0552_ == { 1'h0, _0036_[3], 3'h0 };
assign _1149_ = _0552_ == { 2'h0, _0036_[2:0] };
assign _1150_ = _0552_ == { 2'h0, _0036_[2:1], 1'h0 };
assign _1151_ = _0552_ == { 2'h0, _0036_[2], 1'h0, _0036_[0] };
assign _1152_ = _0552_ == { 2'h0, _0036_[2], 2'h0 };
assign _1153_ = _0552_ == { 3'h0, _0036_[1:0] };
assign _1154_ = _0552_ == { 3'h0, _0036_[1], 1'h0 };
assign _1155_ = _0552_ == { 4'h0, _0036_[0] };
assign _1156_ = _0553_ == _0037_;
assign _1157_ = _0553_ == { _0037_[4:1], 1'h0 };
assign _1158_ = _0553_ == { _0037_[4:2], 1'h0, _0037_[0] };
assign _1159_ = _0553_ == { _0037_[4:2], 2'h0 };
assign _1160_ = _0553_ == { _0037_[4:3], 1'h0, _0037_[1:0] };
assign _1161_ = _0553_ == { _0037_[4:3], 1'h0, _0037_[1], 1'h0 };
assign _1162_ = _0553_ == { _0037_[4:3], 2'h0, _0037_[0] };
assign _1163_ = _0553_ == { _0037_[4:3], 3'h0 };
assign _1164_ = _0553_ == { _0037_[4], 1'h0, _0037_[2:0] };
assign _1165_ = _0553_ == { _0037_[4], 1'h0, _0037_[2:1], 1'h0 };
assign _1166_ = _0553_ == { _0037_[4], 1'h0, _0037_[2], 1'h0, _0037_[0] };
assign _1167_ = _0553_ == { _0037_[4], 1'h0, _0037_[2], 2'h0 };
assign _1168_ = _0553_ == { _0037_[4], 2'h0, _0037_[1:0] };
assign _1169_ = _0553_ == { _0037_[4], 2'h0, _0037_[1], 1'h0 };
assign _1170_ = _0553_ == { _0037_[4], 3'h0, _0037_[0] };
assign _1171_ = _0553_ == { _0037_[4], 4'h0 };
assign _1172_ = _0553_ == { 1'h0, _0037_[3:0] };
assign _1173_ = _0553_ == { 1'h0, _0037_[3:1], 1'h0 };
assign _1174_ = _0553_ == { 1'h0, _0037_[3:2], 1'h0, _0037_[0] };
assign _1175_ = _0553_ == { 1'h0, _0037_[3:2], 2'h0 };
assign _1176_ = _0553_ == { 1'h0, _0037_[3], 1'h0, _0037_[1:0] };
assign _1177_ = _0553_ == { 1'h0, _0037_[3], 1'h0, _0037_[1], 1'h0 };
assign _1178_ = _0553_ == { 1'h0, _0037_[3], 2'h0, _0037_[0] };
assign _1179_ = _0553_ == { 1'h0, _0037_[3], 3'h0 };
assign _1180_ = _0553_ == { 2'h0, _0037_[2:0] };
assign _1181_ = _0553_ == { 2'h0, _0037_[2:1], 1'h0 };
assign _1182_ = _0553_ == { 2'h0, _0037_[2], 1'h0, _0037_[0] };
assign _1183_ = _0553_ == { 2'h0, _0037_[2], 2'h0 };
assign _1184_ = _0553_ == { 3'h0, _0037_[1:0] };
assign _1185_ = _0553_ == { 3'h0, _0037_[1], 1'h0 };
assign _1186_ = _0553_ == { 4'h0, _0037_[0] };
assign _1310_ = _1094_ & _0032_;
assign _1312_ = _1095_ & _0032_;
assign _1314_ = _1096_ & _0032_;
assign _1316_ = _1097_ & _0032_;
assign _1318_ = _1098_ & _0032_;
assign _1320_ = _1099_ & _0032_;
assign _1322_ = _1100_ & _0032_;
assign _1324_ = _1101_ & _0032_;
assign _1326_ = _1102_ & _0032_;
assign _1328_ = _1103_ & _0032_;
assign _1330_ = _1104_ & _0032_;
assign _1332_ = _1105_ & _0032_;
assign _1334_ = _1106_ & _0032_;
assign _1336_ = _1107_ & _0032_;
assign _1338_ = _1108_ & _0032_;
assign _1340_ = _1109_ & _0032_;
assign _1342_ = _1110_ & _0032_;
assign _1344_ = _1111_ & _0032_;
assign _1346_ = _1112_ & _0032_;
assign _1348_ = _1113_ & _0032_;
assign _1350_ = _1114_ & _0032_;
assign _1352_ = _1115_ & _0032_;
assign _1354_ = _1116_ & _0032_;
assign _1356_ = _1117_ & _0032_;
assign _1358_ = _1118_ & _0032_;
assign _1360_ = _1119_ & _0032_;
assign _1362_ = _1120_ & _0032_;
assign _1364_ = _1121_ & _0032_;
assign _1366_ = _1122_ & _0032_;
assign _1368_ = _1123_ & _0032_;
assign _1370_ = _1124_ & _0032_;
assign _1372_ = _1125_ & _0033_;
assign _1374_ = _1126_ & _0033_;
assign _1376_ = _1127_ & _0033_;
assign _1378_ = _1128_ & _0033_;
assign _1380_ = _1129_ & _0033_;
assign _1382_ = _1130_ & _0033_;
assign _1384_ = _1131_ & _0033_;
assign _1386_ = _1132_ & _0033_;
assign _1388_ = _1133_ & _0033_;
assign _1390_ = _1134_ & _0033_;
assign _1392_ = _1135_ & _0033_;
assign _1394_ = _1136_ & _0033_;
assign _1396_ = _1137_ & _0033_;
assign _1398_ = _1138_ & _0033_;
assign _1400_ = _1139_ & _0033_;
assign _1402_ = _1140_ & _0033_;
assign _1404_ = _1141_ & _0033_;
assign _1406_ = _1142_ & _0033_;
assign _1408_ = _1143_ & _0033_;
assign _1410_ = _1144_ & _0033_;
assign _1412_ = _1145_ & _0033_;
assign _1414_ = _1146_ & _0033_;
assign _1416_ = _1147_ & _0033_;
assign _1418_ = _1148_ & _0033_;
assign _1420_ = _1149_ & _0033_;
assign _1422_ = _1150_ & _0033_;
assign _1424_ = _1151_ & _0033_;
assign _1426_ = _1152_ & _0033_;
assign _1428_ = _1153_ & _0033_;
assign _1430_ = _1154_ & _0033_;
assign _1432_ = _1155_ & _0033_;
assign _1434_ = _1156_ & _0034_;
assign _1436_ = _1157_ & _0034_;
assign _1438_ = _1158_ & _0034_;
assign _1440_ = _1159_ & _0034_;
assign _1442_ = _1160_ & _0034_;
assign _1444_ = _1161_ & _0034_;
assign _1446_ = _1162_ & _0034_;
assign _1448_ = _1163_ & _0034_;
assign _1450_ = _1164_ & _0034_;
assign _1452_ = _1165_ & _0034_;
assign _1454_ = _1166_ & _0034_;
assign _1456_ = _1167_ & _0034_;
assign _1458_ = _1168_ & _0034_;
assign _1460_ = _1169_ & _0034_;
assign _1462_ = _1170_ & _0034_;
assign _1464_ = _1171_ & _0034_;
assign _1466_ = _1172_ & _0034_;
assign _1468_ = _1173_ & _0034_;
assign _1470_ = _1174_ & _0034_;
assign _1472_ = _1175_ & _0034_;
assign _1474_ = _1176_ & _0034_;
assign _1476_ = _1177_ & _0034_;
assign _1478_ = _1178_ & _0034_;
assign _1480_ = _1179_ & _0034_;
assign _1482_ = _1180_ & _0034_;
assign _1484_ = _1181_ & _0034_;
assign _1486_ = _1182_ & _0034_;
assign _1488_ = _1183_ & _0034_;
assign _1490_ = _1184_ & _0034_;
assign _1492_ = _1185_ & _0034_;
assign _1494_ = _1186_ & _0034_;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[31].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[31].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[31]) \g_rf_flops[31].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[30].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[30].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[30]) \g_rf_flops[30].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[29].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[29].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[29]) \g_rf_flops[29].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[28].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[28].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[28]) \g_rf_flops[28].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[27].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[27].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[27]) \g_rf_flops[27].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[26].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[26].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[26]) \g_rf_flops[26].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[25].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[25].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[25]) \g_rf_flops[25].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[24].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[24].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[24]) \g_rf_flops[24].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[23].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[23].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[23]) \g_rf_flops[23].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[22].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[22].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[22]) \g_rf_flops[22].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[21].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[21].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[21]) \g_rf_flops[21].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[20].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[20].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[20]) \g_rf_flops[20].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[19].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[19].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[19]) \g_rf_flops[19].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[18].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[18].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[18]) \g_rf_flops[18].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[17].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[17].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[17]) \g_rf_flops[17].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[16].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[16].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[16]) \g_rf_flops[16].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[15].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[15].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[15]) \g_rf_flops[15].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[14].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[14].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[14]) \g_rf_flops[14].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[13].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[13].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[13]) \g_rf_flops[13].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[12].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[12].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[12]) \g_rf_flops[12].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[11].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[11].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[11]) \g_rf_flops[11].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[10].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[10].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[10]) \g_rf_flops[10].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[9].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[9].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[9]) \g_rf_flops[9].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[8].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[8].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[8]) \g_rf_flops[8].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[7].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[7].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[7]) \g_rf_flops[7].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[6].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[6].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[6]) \g_rf_flops[6].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[5].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[5].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[5]) \g_rf_flops[5].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[4].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[4].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[4]) \g_rf_flops[4].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[3].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[3].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[3]) \g_rf_flops[3].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[2].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[2].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[2]) \g_rf_flops[2].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20107.4-20111.28" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_rf_flops[1].rf_reg_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_rf_flops[1].rf_reg_q  <= 39'h2a00000000;
else if (we_a_dec[1]) \g_rf_flops[1].rf_reg_q  <= wdata_a_i;
/* src = "generated/sv2v_out.v:20118.4-20122.27" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  */
/* PC_TAINT_INFO STATE_NAME \g_dummy_r0.rf_r0_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_dummy_r0.rf_r0_q  <= 39'h2a00000000;
else if (\g_dummy_r0.we_r0_dummy ) \g_dummy_r0.rf_r0_q  <= wdata_a_i;
assign _0038_ = | { _1378_, _1376_, _0985_ };
assign _0039_ = | { _1394_, _1392_, _0989_ };
assign _0040_ = | { _1386_, _1384_, _1378_, _1376_, _0987_, _0985_ };
assign _0041_ = | { _1410_, _1408_, _0993_ };
assign _0042_ = | { _1426_, _1424_, _0997_ };
assign _0043_ = | { _1418_, _1416_, _1410_, _1408_, _0995_, _0993_ };
assign _0044_ = | { _1400_, _1402_, _1386_, _1384_, _1394_, _1392_, _1378_, _1376_, _0991_, _0989_, _0987_, _0985_ };
assign _0045_ = | { _1438_, _1440_, _1001_ };
assign _0046_ = | { _1456_, _1454_, _1005_ };
assign _0047_ = | { _1448_, _1446_, _1438_, _1440_, _1003_, _1001_ };
assign _0048_ = | { _1472_, _1470_, _1009_ };
assign _0049_ = | { _1488_, _1486_, _1013_ };
assign _0050_ = | { _1480_, _1478_, _1472_, _1470_, _1011_, _1009_ };
assign _0051_ = | { _1464_, _1462_, _1448_, _1446_, _1456_, _1454_, _1438_, _1440_, _1007_, _1005_, _1003_, _1001_ };
assign _0032_ = | waddr_a_i_t0;
assign _0052_ = ~ { _0985_, _1378_, _1376_ };
assign _0053_ = ~ { _0989_, _1394_, _1392_ };
assign _0054_ = ~ { _0985_, _0987_, _1386_, _1384_, _1378_, _1376_ };
assign _0055_ = ~ { _0993_, _1410_, _1408_ };
assign _0056_ = ~ { _0997_, _1426_, _1424_ };
assign _0057_ = ~ { _0993_, _0995_, _1418_, _1416_, _1410_, _1408_ };
assign _0058_ = ~ { _0985_, _0987_, _0989_, _0991_, _1400_, _1402_, _1394_, _1392_, _1386_, _1384_, _1378_, _1376_ };
assign _0059_ = ~ { _1001_, _1438_, _1440_ };
assign _0060_ = ~ { _1005_, _1456_, _1454_ };
assign _0061_ = ~ { _1001_, _1003_, _1448_, _1446_, _1438_, _1440_ };
assign _0062_ = ~ { _1009_, _1472_, _1470_ };
assign _0063_ = ~ { _1013_, _1488_, _1486_ };
assign _0064_ = ~ { _1009_, _1011_, _1480_, _1478_, _1472_, _1470_ };
assign _0065_ = ~ { _1001_, _1003_, _1005_, _1007_, _1464_, _1462_, _1456_, _1454_, _1448_, _1446_, _1438_, _1440_ };
assign _0351_ = { _0984_, _1377_, _1375_ } & _0052_;
assign _0352_ = { _0988_, _1393_, _1391_ } & _0053_;
assign _0353_ = { _0984_, _0986_, _1385_, _1383_, _1377_, _1375_ } & _0054_;
assign _0354_ = { _0992_, _1409_, _1407_ } & _0055_;
assign _0355_ = { _0996_, _1425_, _1423_ } & _0056_;
assign _0356_ = { _0992_, _0994_, _1417_, _1415_, _1409_, _1407_ } & _0057_;
assign _0357_ = { _0984_, _0986_, _0988_, _0990_, _1399_, _1401_, _1393_, _1391_, _1385_, _1383_, _1377_, _1375_ } & _0058_;
assign _0358_ = { _1000_, _1437_, _1439_ } & _0059_;
assign _0359_ = { _1004_, _1455_, _1453_ } & _0060_;
assign _0360_ = { _1000_, _1002_, _1447_, _1445_, _1437_, _1439_ } & _0061_;
assign _0361_ = { _1008_, _1471_, _1469_ } & _0062_;
assign _0362_ = { _1012_, _1487_, _1485_ } & _0063_;
assign _0363_ = { _1008_, _1010_, _1479_, _1477_, _1471_, _1469_ } & _0064_;
assign _0364_ = { _1000_, _1002_, _1004_, _1006_, _1463_, _1461_, _1455_, _1453_, _1447_, _1445_, _1437_, _1439_ } & _0065_;
assign _0066_ = ! _0351_;
assign _0067_ = ! _0352_;
assign _0068_ = ! _0353_;
assign _0069_ = ! _0354_;
assign _0070_ = ! _0355_;
assign _0071_ = ! _0356_;
assign _0072_ = ! _0357_;
assign _0073_ = ! _0358_;
assign _0074_ = ! _0359_;
assign _0075_ = ! _0360_;
assign _0076_ = ! _0361_;
assign _0077_ = ! _0362_;
assign _0078_ = ! _0363_;
assign _0079_ = ! _0364_;
assign _0080_ = ! _0551_;
assign _0177_ = _0066_ & _0038_;
assign _0179_ = _0067_ & _0039_;
assign _0181_ = _0068_ & _0040_;
assign _0183_ = _0069_ & _0041_;
assign _0185_ = _0070_ & _0042_;
assign _0187_ = _0071_ & _0043_;
assign _0189_ = _0072_ & _0044_;
assign _0191_ = _0073_ & _0045_;
assign _0193_ = _0074_ & _0046_;
assign _0195_ = _0075_ & _0047_;
assign _0197_ = _0076_ & _0048_;
assign _0199_ = _0077_ & _0049_;
assign _0201_ = _0078_ & _0050_;
assign _0203_ = _0079_ & _0051_;
assign _1308_ = _0080_ & _0032_;
assign _0081_ = ~ { _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_ };
assign _0082_ = ~ { _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_ };
assign _0083_ = ~ { _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_ };
assign _0084_ = ~ { _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_ };
assign _0085_ = ~ { _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_ };
assign _0086_ = ~ { _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_ };
assign _0087_ = ~ { _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_ };
assign _0088_ = ~ { _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_ };
assign _0089_ = ~ { _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_ };
assign _0090_ = ~ { _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_ };
assign _0091_ = ~ { _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_ };
assign _0092_ = ~ { _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_ };
assign _0093_ = ~ { _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_ };
assign _0094_ = ~ { _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_ };
assign _0095_ = ~ { _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_ };
assign _0096_ = ~ { _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_ };
assign _0097_ = ~ { _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_ };
assign _0098_ = ~ { _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_ };
assign _0099_ = ~ { _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_ };
assign _0100_ = ~ { _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_ };
assign _0101_ = ~ { _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_ };
assign _0102_ = ~ { _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_ };
assign _0103_ = ~ { _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_ };
assign _0104_ = ~ { _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_ };
assign _0105_ = ~ { _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_ };
assign _0106_ = ~ { _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_ };
assign _0107_ = ~ { _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_ };
assign _0108_ = ~ { _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_ };
assign _0109_ = ~ { _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_ };
assign _0110_ = ~ { _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_ };
assign _0111_ = ~ { _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_ };
assign _0112_ = ~ { _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_ };
assign _0113_ = ~ { _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_ };
assign _0114_ = ~ { _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_ };
assign _0115_ = ~ { _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_ };
assign _0116_ = ~ { _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_ };
assign _0117_ = ~ { _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_ };
assign _0118_ = ~ { _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_ };
assign _0119_ = ~ { _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_ };
assign _0120_ = ~ { _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_ };
assign _0121_ = ~ { _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_ };
assign _0122_ = ~ { _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_ };
assign _0123_ = ~ { _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_ };
assign _0124_ = ~ { _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_ };
assign _0125_ = ~ { _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_ };
assign _0126_ = ~ { _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_ };
assign _0127_ = ~ { _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_ };
assign _0128_ = ~ { _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_ };
assign _0129_ = ~ { _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_ };
assign _0130_ = ~ { _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_ };
assign _0131_ = ~ { _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_ };
assign _0132_ = ~ { _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_ };
assign _0133_ = ~ { _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_ };
assign _0134_ = ~ { _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_ };
assign _0135_ = ~ { _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_ };
assign _0136_ = ~ { _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_ };
assign _0137_ = ~ { _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_ };
assign _0138_ = ~ { _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_ };
assign _0139_ = ~ { _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_ };
assign _0140_ = ~ { _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_ };
assign _0141_ = ~ { _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_ };
assign _0142_ = ~ { _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_ };
assign _0765_ = { _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_ } | _0081_;
assign _0768_ = { _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_ } | _0082_;
assign _0771_ = { _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_ } | _0083_;
assign _0774_ = { _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_ } | _0084_;
assign _0777_ = { _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_ } | _0085_;
assign _0780_ = { _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_ } | _0086_;
assign _0783_ = { _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_ } | _0087_;
assign _0786_ = { _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_ } | _0088_;
assign _0789_ = { _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_ } | _0089_;
assign _0792_ = { _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_ } | _0090_;
assign _0795_ = { _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_ } | _0091_;
assign _0798_ = { _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_ } | _0092_;
assign _0801_ = { _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_ } | _0093_;
assign _0804_ = { _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_ } | _0094_;
assign _0807_ = { _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_ } | _0095_;
assign _0810_ = { _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_ } | _0096_;
assign _0813_ = { _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_ } | _0097_;
assign _0816_ = { _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_ } | _0098_;
assign _0819_ = { _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_ } | _0099_;
assign _0822_ = { _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_ } | _0100_;
assign _0825_ = { _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_ } | _0101_;
assign _0828_ = { _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_ } | _0102_;
assign _0831_ = { _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_ } | _0103_;
assign _0834_ = { _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_ } | _0104_;
assign _0837_ = { _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_ } | _0105_;
assign _0840_ = { _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_ } | _0106_;
assign _0843_ = { _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_ } | _0107_;
assign _0846_ = { _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_ } | _0108_;
assign _0849_ = { _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_ } | _0109_;
assign _0852_ = { _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_ } | _0110_;
assign _0855_ = { _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_ } | _0111_;
assign _0858_ = { _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_ } | _0112_;
assign _0861_ = { _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_ } | _0113_;
assign _0864_ = { _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_ } | _0114_;
assign _0867_ = { _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_ } | _0115_;
assign _0870_ = { _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_ } | _0116_;
assign _0873_ = { _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_ } | _0117_;
assign _0876_ = { _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_ } | _0118_;
assign _0879_ = { _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_ } | _0119_;
assign _0882_ = { _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_ } | _0120_;
assign _0885_ = { _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_ } | _0121_;
assign _0888_ = { _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_ } | _0122_;
assign _0891_ = { _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_ } | _0123_;
assign _0894_ = { _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_ } | _0124_;
assign _0897_ = { _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_ } | _0125_;
assign _0900_ = { _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_ } | _0126_;
assign _0903_ = { _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_ } | _0127_;
assign _0906_ = { _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_ } | _0128_;
assign _0909_ = { _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_ } | _0129_;
assign _0912_ = { _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_ } | _0130_;
assign _0915_ = { _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_ } | _0131_;
assign _0918_ = { _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_ } | _0132_;
assign _0921_ = { _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_ } | _0133_;
assign _0924_ = { _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_ } | _0134_;
assign _0927_ = { _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_ } | _0135_;
assign _0930_ = { _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_ } | _0136_;
assign _0933_ = { _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_ } | _0137_;
assign _0936_ = { _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_ } | _0138_;
assign _0939_ = { _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_ } | _0139_;
assign _0942_ = { _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_ } | _0140_;
assign _0945_ = { _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_ } | _0141_;
assign _0948_ = { _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_ } | _0142_;
assign _0766_ = { _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_ } | { _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_, _1371_ };
assign _0769_ = { _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_ } | { _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_, _1375_ };
assign _0772_ = { _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_ } | { _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_, _0984_ };
assign _0775_ = { _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_ } | { _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_ };
assign _0778_ = { _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_ } | { _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_, _1383_ };
assign _0781_ = { _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_ } | { _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_, _0986_ };
assign _0784_ = { _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_ } | { _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_, _0176_ };
assign _0787_ = { _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_ } | { _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_, _1387_ };
assign _0790_ = { _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_ } | { _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_, _1391_ };
assign _0793_ = { _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_ } | { _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_, _0988_ };
assign _0796_ = { _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_ } | { _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_, _1395_ };
assign _0799_ = { _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_ } | { _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_, _1399_ };
assign _0802_ = { _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_ } | { _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_, _0990_ };
assign _0805_ = { _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_ } | { _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_, _0178_ };
assign _0808_ = { _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_ } | { _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_ };
assign _0811_ = { _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_ } | { _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_, _1403_ };
assign _0814_ = { _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_ } | { _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_, _1407_ };
assign _0817_ = { _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_ } | { _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_, _0992_ };
assign _0820_ = { _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_ } | { _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_, _1411_ };
assign _0823_ = { _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_ } | { _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_, _1415_ };
assign _0826_ = { _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_ } | { _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_, _0994_ };
assign _0829_ = { _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_ } | { _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_, _0182_ };
assign _0832_ = { _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_ } | { _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_, _1419_ };
assign _0835_ = { _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_ } | { _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_, _1423_ };
assign _0838_ = { _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_ } | { _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_, _0996_ };
assign _0841_ = { _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_ } | { _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_, _1427_ };
assign _0844_ = { _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_ } | { _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_, _1431_ };
assign _0847_ = { _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_ } | { _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_, _0998_ };
assign _0850_ = { _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_ } | { _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_, _0184_ };
assign _0853_ = { _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_ } | { _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_ };
assign _0856_ = { _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_ } | { _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_, _0188_ };
assign _0859_ = { _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_ } | { _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_ };
assign _0862_ = { _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_ } | { _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_, _1437_ };
assign _0865_ = { _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_ } | { _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_, _1000_ };
assign _0868_ = { _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_ } | { _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_, _1441_ };
assign _0871_ = { _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_ } | { _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_, _1445_ };
assign _0874_ = { _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_ } | { _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_, _1002_ };
assign _0877_ = { _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_ } | { _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_, _0190_ };
assign _0880_ = { _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_ } | { _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_, _1449_ };
assign _0883_ = { _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_ } | { _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_, _1453_ };
assign _0886_ = { _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_ } | { _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_, _1004_ };
assign _0889_ = { _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_ } | { _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_, _1457_ };
assign _0892_ = { _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_ } | { _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_, _1461_ };
assign _0895_ = { _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_ } | { _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_, _1006_ };
assign _0898_ = { _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_ } | { _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_, _0192_ };
assign _0901_ = { _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_ } | { _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_, _0194_ };
assign _0904_ = { _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_ } | { _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_, _1465_ };
assign _0907_ = { _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_ } | { _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_, _1469_ };
assign _0910_ = { _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_ } | { _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_, _1008_ };
assign _0913_ = { _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_ } | { _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_, _1473_ };
assign _0916_ = { _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_ } | { _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_, _1477_ };
assign _0919_ = { _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_ } | { _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_, _1010_ };
assign _0922_ = { _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_ } | { _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_, _0196_ };
assign _0925_ = { _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_ } | { _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_, _1481_ };
assign _0928_ = { _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_ } | { _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_, _1485_ };
assign _0931_ = { _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_ } | { _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_, _1012_ };
assign _0934_ = { _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_ } | { _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_, _1489_ };
assign _0937_ = { _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_ } | { _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_, _1493_ };
assign _0940_ = { _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_ } | { _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_, _1014_ };
assign _0943_ = { _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_ } | { _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_ };
assign _0946_ = { _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_ } | { _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_ };
assign _0949_ = { _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_ } | { _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_, _0202_ };
assign _0951_ = _1308_ | _1307_;
assign _0952_ = _1310_ | _1309_;
assign _0953_ = _1312_ | _1311_;
assign _0954_ = _1314_ | _1313_;
assign _0955_ = _1316_ | _1315_;
assign _0956_ = _1318_ | _1317_;
assign _0957_ = _1320_ | _1319_;
assign _0958_ = _1322_ | _1321_;
assign _0959_ = _1324_ | _1323_;
assign _0960_ = _1326_ | _1325_;
assign _0961_ = _1328_ | _1327_;
assign _0962_ = _1330_ | _1329_;
assign _0963_ = _1332_ | _1331_;
assign _0964_ = _1334_ | _1333_;
assign _0965_ = _1336_ | _1335_;
assign _0966_ = _1338_ | _1337_;
assign _0967_ = _1340_ | _1339_;
assign _0968_ = _1342_ | _1341_;
assign _0969_ = _1344_ | _1343_;
assign _0970_ = _1346_ | _1345_;
assign _0971_ = _1348_ | _1347_;
assign _0972_ = _1350_ | _1349_;
assign _0973_ = _1352_ | _1351_;
assign _0974_ = _1354_ | _1353_;
assign _0975_ = _1356_ | _1355_;
assign _0976_ = _1358_ | _1357_;
assign _0977_ = _1360_ | _1359_;
assign _0978_ = _1362_ | _1361_;
assign _0979_ = _1364_ | _1363_;
assign _0980_ = _1366_ | _1365_;
assign _0981_ = _1368_ | _1367_;
assign _0982_ = _1370_ | _1369_;
assign _0983_ = { dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0 } | { dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i, dummy_instr_id_i };
assign _0365_ = \g_rf_flops[30].rf_reg_q_t0  & _0765_;
assign _0368_ = \g_rf_flops[28].rf_reg_q_t0  & _0768_;
assign _0371_ = _1190_ & _0771_;
assign _0374_ = \g_rf_flops[26].rf_reg_q_t0  & _0774_;
assign _0377_ = \g_rf_flops[24].rf_reg_q_t0  & _0777_;
assign _0380_ = _1196_ & _0780_;
assign _0383_ = _1198_ & _0783_;
assign _0386_ = \g_rf_flops[22].rf_reg_q_t0  & _0786_;
assign _0389_ = \g_rf_flops[20].rf_reg_q_t0  & _0789_;
assign _0392_ = _1204_ & _0792_;
assign _0395_ = \g_rf_flops[18].rf_reg_q_t0  & _0795_;
assign _0398_ = \g_rf_flops[16].rf_reg_q_t0  & _0798_;
assign _0401_ = _1210_ & _0801_;
assign _0404_ = _1212_ & _0804_;
assign _0407_ = _1214_ & _0807_;
assign _0410_ = \g_rf_flops[14].rf_reg_q_t0  & _0810_;
assign _0413_ = \g_rf_flops[12].rf_reg_q_t0  & _0813_;
assign _0416_ = _1220_ & _0816_;
assign _0419_ = \g_rf_flops[10].rf_reg_q_t0  & _0819_;
assign _0422_ = \g_rf_flops[8].rf_reg_q_t0  & _0822_;
assign _0425_ = _1226_ & _0825_;
assign _0428_ = _1228_ & _0828_;
assign _0431_ = \g_rf_flops[6].rf_reg_q_t0  & _0831_;
assign _0434_ = \g_rf_flops[4].rf_reg_q_t0  & _0834_;
assign _0437_ = _1234_ & _0837_;
assign _0440_ = \g_rf_flops[2].rf_reg_q_t0  & _0840_;
assign _0443_ = \rf_reg[0]_t0  & _0843_;
assign _0446_ = _1240_ & _0846_;
assign _0449_ = _1242_ & _0849_;
assign _0452_ = _1244_ & _0852_;
assign _0455_ = _1246_ & _0855_;
assign _0458_ = \g_rf_flops[30].rf_reg_q_t0  & _0858_;
assign _0461_ = \g_rf_flops[28].rf_reg_q_t0  & _0861_;
assign _0464_ = _1250_ & _0864_;
assign _0467_ = \g_rf_flops[26].rf_reg_q_t0  & _0867_;
assign _0470_ = \g_rf_flops[24].rf_reg_q_t0  & _0870_;
assign _0473_ = _1256_ & _0873_;
assign _0476_ = _1258_ & _0876_;
assign _0479_ = \g_rf_flops[22].rf_reg_q_t0  & _0879_;
assign _0482_ = \g_rf_flops[20].rf_reg_q_t0  & _0882_;
assign _0485_ = _1264_ & _0885_;
assign _0488_ = \g_rf_flops[18].rf_reg_q_t0  & _0888_;
assign _0491_ = \g_rf_flops[16].rf_reg_q_t0  & _0891_;
assign _0494_ = _1270_ & _0894_;
assign _0497_ = _1272_ & _0897_;
assign _0500_ = _1274_ & _0900_;
assign _0503_ = \g_rf_flops[14].rf_reg_q_t0  & _0903_;
assign _0506_ = \g_rf_flops[12].rf_reg_q_t0  & _0906_;
assign _0509_ = _1280_ & _0909_;
assign _0512_ = \g_rf_flops[10].rf_reg_q_t0  & _0912_;
assign _0515_ = \g_rf_flops[8].rf_reg_q_t0  & _0915_;
assign _0518_ = _1286_ & _0918_;
assign _0521_ = _1288_ & _0921_;
assign _0524_ = \g_rf_flops[6].rf_reg_q_t0  & _0924_;
assign _0527_ = \g_rf_flops[4].rf_reg_q_t0  & _0927_;
assign _0530_ = _1294_ & _0930_;
assign _0533_ = \g_rf_flops[2].rf_reg_q_t0  & _0933_;
assign _0536_ = \rf_reg[0]_t0  & _0936_;
assign _0539_ = _1300_ & _0939_;
assign _0542_ = _1302_ & _0942_;
assign _0545_ = _1304_ & _0945_;
assign _0548_ = _1306_ & _0948_;
assign _0366_ = \g_rf_flops[31].rf_reg_q_t0  & _0766_;
assign _0369_ = \g_rf_flops[29].rf_reg_q_t0  & _0769_;
assign _0372_ = _1188_ & _0772_;
assign _0375_ = \g_rf_flops[27].rf_reg_q_t0  & _0775_;
assign _0378_ = \g_rf_flops[25].rf_reg_q_t0  & _0778_;
assign _0381_ = _1194_ & _0781_;
assign _0384_ = _1192_ & _0784_;
assign _0387_ = \g_rf_flops[23].rf_reg_q_t0  & _0787_;
assign _0390_ = \g_rf_flops[21].rf_reg_q_t0  & _0790_;
assign _0393_ = _1202_ & _0793_;
assign _0396_ = \g_rf_flops[19].rf_reg_q_t0  & _0796_;
assign _0399_ = \g_rf_flops[17].rf_reg_q_t0  & _0799_;
assign _0402_ = _1208_ & _0802_;
assign _0405_ = _1206_ & _0805_;
assign _0408_ = _1200_ & _0808_;
assign _0411_ = \g_rf_flops[15].rf_reg_q_t0  & _0811_;
assign _0414_ = \g_rf_flops[13].rf_reg_q_t0  & _0814_;
assign _0417_ = _1218_ & _0817_;
assign _0420_ = \g_rf_flops[11].rf_reg_q_t0  & _0820_;
assign _0423_ = \g_rf_flops[9].rf_reg_q_t0  & _0823_;
assign _0426_ = _1224_ & _0826_;
assign _0429_ = _1222_ & _0829_;
assign _0432_ = \g_rf_flops[7].rf_reg_q_t0  & _0832_;
assign _0435_ = \g_rf_flops[5].rf_reg_q_t0  & _0835_;
assign _0438_ = _1232_ & _0838_;
assign _0441_ = \g_rf_flops[3].rf_reg_q_t0  & _0841_;
assign _0444_ = \g_rf_flops[1].rf_reg_q_t0  & _0844_;
assign _0447_ = _1238_ & _0847_;
assign _0450_ = _1236_ & _0850_;
assign _0453_ = _1230_ & _0853_;
assign _0456_ = _1216_ & _0856_;
assign _0459_ = \g_rf_flops[31].rf_reg_q_t0  & _0859_;
assign _0462_ = \g_rf_flops[29].rf_reg_q_t0  & _0862_;
assign _0465_ = _1248_ & _0865_;
assign _0468_ = \g_rf_flops[27].rf_reg_q_t0  & _0868_;
assign _0471_ = \g_rf_flops[25].rf_reg_q_t0  & _0871_;
assign _0474_ = _1254_ & _0874_;
assign _0477_ = _1252_ & _0877_;
assign _0480_ = \g_rf_flops[23].rf_reg_q_t0  & _0880_;
assign _0483_ = \g_rf_flops[21].rf_reg_q_t0  & _0883_;
assign _0486_ = _1262_ & _0886_;
assign _0489_ = \g_rf_flops[19].rf_reg_q_t0  & _0889_;
assign _0492_ = \g_rf_flops[17].rf_reg_q_t0  & _0892_;
assign _0495_ = _1268_ & _0895_;
assign _0498_ = _1266_ & _0898_;
assign _0501_ = _1260_ & _0901_;
assign _0504_ = \g_rf_flops[15].rf_reg_q_t0  & _0904_;
assign _0507_ = \g_rf_flops[13].rf_reg_q_t0  & _0907_;
assign _0510_ = _1278_ & _0910_;
assign _0513_ = \g_rf_flops[11].rf_reg_q_t0  & _0913_;
assign _0516_ = \g_rf_flops[9].rf_reg_q_t0  & _0916_;
assign _0519_ = _1284_ & _0919_;
assign _0522_ = _1282_ & _0922_;
assign _0525_ = \g_rf_flops[7].rf_reg_q_t0  & _0925_;
assign _0528_ = \g_rf_flops[5].rf_reg_q_t0  & _0928_;
assign _0531_ = _1292_ & _0931_;
assign _0534_ = \g_rf_flops[3].rf_reg_q_t0  & _0934_;
assign _0537_ = \g_rf_flops[1].rf_reg_q_t0  & _0937_;
assign _0540_ = _1298_ & _0940_;
assign _0543_ = _1296_ & _0943_;
assign _0546_ = _1290_ & _0946_;
assign _0549_ = _1276_ & _0949_;
assign _0554_ = we_a_i_t0 & _0951_;
assign _0556_ = we_a_i_t0 & _0952_;
assign _0558_ = we_a_i_t0 & _0953_;
assign _0560_ = we_a_i_t0 & _0954_;
assign _0562_ = we_a_i_t0 & _0955_;
assign _0564_ = we_a_i_t0 & _0956_;
assign _0566_ = we_a_i_t0 & _0957_;
assign _0568_ = we_a_i_t0 & _0958_;
assign _0570_ = we_a_i_t0 & _0959_;
assign _0572_ = we_a_i_t0 & _0960_;
assign _0574_ = we_a_i_t0 & _0961_;
assign _0576_ = we_a_i_t0 & _0962_;
assign _0578_ = we_a_i_t0 & _0963_;
assign _0580_ = we_a_i_t0 & _0964_;
assign _0582_ = we_a_i_t0 & _0965_;
assign _0584_ = we_a_i_t0 & _0966_;
assign _0586_ = we_a_i_t0 & _0967_;
assign _0588_ = we_a_i_t0 & _0968_;
assign _0590_ = we_a_i_t0 & _0969_;
assign _0592_ = we_a_i_t0 & _0970_;
assign _0594_ = we_a_i_t0 & _0971_;
assign _0596_ = we_a_i_t0 & _0972_;
assign _0598_ = we_a_i_t0 & _0973_;
assign _0600_ = we_a_i_t0 & _0974_;
assign _0602_ = we_a_i_t0 & _0975_;
assign _0604_ = we_a_i_t0 & _0976_;
assign _0606_ = we_a_i_t0 & _0977_;
assign _0608_ = we_a_i_t0 & _0978_;
assign _0610_ = we_a_i_t0 & _0979_;
assign _0612_ = we_a_i_t0 & _0980_;
assign _0614_ = we_a_i_t0 & _0981_;
assign _0616_ = we_a_i_t0 & _0982_;
assign _0618_ = \g_dummy_r0.rf_r0_q_t0  & _0983_;
assign _0767_ = _0365_ | _0366_;
assign _0770_ = _0368_ | _0369_;
assign _0773_ = _0371_ | _0372_;
assign _0776_ = _0374_ | _0375_;
assign _0779_ = _0377_ | _0378_;
assign _0782_ = _0380_ | _0381_;
assign _0785_ = _0383_ | _0384_;
assign _0788_ = _0386_ | _0387_;
assign _0791_ = _0389_ | _0390_;
assign _0794_ = _0392_ | _0393_;
assign _0797_ = _0395_ | _0396_;
assign _0800_ = _0398_ | _0399_;
assign _0803_ = _0401_ | _0402_;
assign _0806_ = _0404_ | _0405_;
assign _0809_ = _0407_ | _0408_;
assign _0812_ = _0410_ | _0411_;
assign _0815_ = _0413_ | _0414_;
assign _0818_ = _0416_ | _0417_;
assign _0821_ = _0419_ | _0420_;
assign _0824_ = _0422_ | _0423_;
assign _0827_ = _0425_ | _0426_;
assign _0830_ = _0428_ | _0429_;
assign _0833_ = _0431_ | _0432_;
assign _0836_ = _0434_ | _0435_;
assign _0839_ = _0437_ | _0438_;
assign _0842_ = _0440_ | _0441_;
assign _0845_ = _0443_ | _0444_;
assign _0848_ = _0446_ | _0447_;
assign _0851_ = _0449_ | _0450_;
assign _0854_ = _0452_ | _0453_;
assign _0857_ = _0455_ | _0456_;
assign _0860_ = _0458_ | _0459_;
assign _0863_ = _0461_ | _0462_;
assign _0866_ = _0464_ | _0465_;
assign _0869_ = _0467_ | _0468_;
assign _0872_ = _0470_ | _0471_;
assign _0875_ = _0473_ | _0474_;
assign _0878_ = _0476_ | _0477_;
assign _0881_ = _0479_ | _0480_;
assign _0884_ = _0482_ | _0483_;
assign _0887_ = _0485_ | _0486_;
assign _0890_ = _0488_ | _0489_;
assign _0893_ = _0491_ | _0492_;
assign _0896_ = _0494_ | _0495_;
assign _0899_ = _0497_ | _0498_;
assign _0902_ = _0500_ | _0501_;
assign _0905_ = _0503_ | _0504_;
assign _0908_ = _0506_ | _0507_;
assign _0911_ = _0509_ | _0510_;
assign _0914_ = _0512_ | _0513_;
assign _0917_ = _0515_ | _0516_;
assign _0920_ = _0518_ | _0519_;
assign _0923_ = _0521_ | _0522_;
assign _0926_ = _0524_ | _0525_;
assign _0929_ = _0527_ | _0528_;
assign _0932_ = _0530_ | _0531_;
assign _0935_ = _0533_ | _0534_;
assign _0938_ = _0536_ | _0537_;
assign _0941_ = _0539_ | _0540_;
assign _0944_ = _0542_ | _0543_;
assign _0947_ = _0545_ | _0546_;
assign _0950_ = _0548_ | _0549_;
assign _1048_ = \g_rf_flops[30].rf_reg_q  ^ \g_rf_flops[31].rf_reg_q ;
assign _1049_ = \g_rf_flops[28].rf_reg_q  ^ \g_rf_flops[29].rf_reg_q ;
assign _1050_ = _1189_ ^ _1187_;
assign _1051_ = \g_rf_flops[26].rf_reg_q  ^ \g_rf_flops[27].rf_reg_q ;
assign _1052_ = \g_rf_flops[24].rf_reg_q  ^ \g_rf_flops[25].rf_reg_q ;
assign _1053_ = _1195_ ^ _1193_;
assign _1054_ = _1197_ ^ _1191_;
assign _1055_ = \g_rf_flops[22].rf_reg_q  ^ \g_rf_flops[23].rf_reg_q ;
assign _1056_ = \g_rf_flops[20].rf_reg_q  ^ \g_rf_flops[21].rf_reg_q ;
assign _1057_ = _1203_ ^ _1201_;
assign _1058_ = \g_rf_flops[18].rf_reg_q  ^ \g_rf_flops[19].rf_reg_q ;
assign _1059_ = \g_rf_flops[16].rf_reg_q  ^ \g_rf_flops[17].rf_reg_q ;
assign _1060_ = _1209_ ^ _1207_;
assign _1061_ = _1211_ ^ _1205_;
assign _1062_ = _1213_ ^ _1199_;
assign _1063_ = \g_rf_flops[14].rf_reg_q  ^ \g_rf_flops[15].rf_reg_q ;
assign _1064_ = \g_rf_flops[12].rf_reg_q  ^ \g_rf_flops[13].rf_reg_q ;
assign _1065_ = _1219_ ^ _1217_;
assign _1066_ = \g_rf_flops[10].rf_reg_q  ^ \g_rf_flops[11].rf_reg_q ;
assign _1067_ = \g_rf_flops[8].rf_reg_q  ^ \g_rf_flops[9].rf_reg_q ;
assign _1068_ = _1225_ ^ _1223_;
assign _1069_ = _1227_ ^ _1221_;
assign _1070_ = \g_rf_flops[6].rf_reg_q  ^ \g_rf_flops[7].rf_reg_q ;
assign _1071_ = \g_rf_flops[4].rf_reg_q  ^ \g_rf_flops[5].rf_reg_q ;
assign _1072_ = _1233_ ^ _1231_;
assign _1073_ = \g_rf_flops[2].rf_reg_q  ^ \g_rf_flops[3].rf_reg_q ;
assign _1074_ = \rf_reg[0]  ^ \g_rf_flops[1].rf_reg_q ;
assign _1075_ = _1239_ ^ _1237_;
assign _1076_ = _1241_ ^ _1235_;
assign _1077_ = _1243_ ^ _1229_;
assign _1078_ = _1245_ ^ _1215_;
assign _1079_ = _1249_ ^ _1247_;
assign _1080_ = _1255_ ^ _1253_;
assign _1081_ = _1257_ ^ _1251_;
assign _1082_ = _1263_ ^ _1261_;
assign _1083_ = _1269_ ^ _1267_;
assign _1084_ = _1271_ ^ _1265_;
assign _1085_ = _1273_ ^ _1259_;
assign _1086_ = _1279_ ^ _1277_;
assign _1087_ = _1285_ ^ _1283_;
assign _1088_ = _1287_ ^ _1281_;
assign _1089_ = _1293_ ^ _1291_;
assign _1090_ = _1299_ ^ _1297_;
assign _1091_ = _1301_ ^ _1295_;
assign _1092_ = _1303_ ^ _1289_;
assign _1093_ = _1305_ ^ _1275_;
assign _0367_ = { _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_, _1372_ } & _1048_;
assign _0370_ = { _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_ } & _1049_;
assign _0373_ = { _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_, _0985_ } & _1050_;
assign _0376_ = { _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_ } & _1051_;
assign _0379_ = { _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_, _1384_ } & _1052_;
assign _0382_ = { _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_, _0987_ } & _1053_;
assign _0385_ = { _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_, _0177_ } & _1054_;
assign _0388_ = { _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_, _1388_ } & _1055_;
assign _0391_ = { _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_, _1392_ } & _1056_;
assign _0394_ = { _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_, _0989_ } & _1057_;
assign _0397_ = { _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_, _1396_ } & _1058_;
assign _0400_ = { _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_, _1400_ } & _1059_;
assign _0403_ = { _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_, _0991_ } & _1060_;
assign _0406_ = { _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_ } & _1061_;
assign _0409_ = { _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_, _0181_ } & _1062_;
assign _0412_ = { _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_, _1404_ } & _1063_;
assign _0415_ = { _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_, _1408_ } & _1064_;
assign _0418_ = { _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_, _0993_ } & _1065_;
assign _0421_ = { _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_, _1412_ } & _1066_;
assign _0424_ = { _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_, _1416_ } & _1067_;
assign _0427_ = { _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_, _0995_ } & _1068_;
assign _0430_ = { _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_, _0183_ } & _1069_;
assign _0433_ = { _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_, _1420_ } & _1070_;
assign _0436_ = { _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_, _1424_ } & _1071_;
assign _0439_ = { _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_, _0997_ } & _1072_;
assign _0442_ = { _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_, _1428_ } & _1073_;
assign _0445_ = { _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_, _1432_ } & _1074_;
assign _0448_ = { _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_, _0999_ } & _1075_;
assign _0451_ = { _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_, _0185_ } & _1076_;
assign _0454_ = { _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_ } & _1077_;
assign _0457_ = { _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_, _0189_ } & _1078_;
assign _0460_ = { _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_ } & _1048_;
assign _0463_ = { _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_, _1438_ } & _1049_;
assign _0466_ = { _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_, _1001_ } & _1079_;
assign _0469_ = { _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_, _1442_ } & _1051_;
assign _0472_ = { _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_, _1446_ } & _1052_;
assign _0475_ = { _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_, _1003_ } & _1080_;
assign _0478_ = { _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_, _0191_ } & _1081_;
assign _0481_ = { _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_, _1450_ } & _1055_;
assign _0484_ = { _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_, _1454_ } & _1056_;
assign _0487_ = { _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_, _1005_ } & _1082_;
assign _0490_ = { _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_, _1458_ } & _1058_;
assign _0493_ = { _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_, _1462_ } & _1059_;
assign _0496_ = { _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_, _1007_ } & _1083_;
assign _0499_ = { _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_ } & _1084_;
assign _0502_ = { _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_, _0195_ } & _1085_;
assign _0505_ = { _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_, _1466_ } & _1063_;
assign _0508_ = { _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_, _1470_ } & _1064_;
assign _0511_ = { _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_, _1009_ } & _1086_;
assign _0514_ = { _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_, _1474_ } & _1066_;
assign _0517_ = { _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_, _1478_ } & _1067_;
assign _0520_ = { _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_, _1011_ } & _1087_;
assign _0523_ = { _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_, _0197_ } & _1088_;
assign _0526_ = { _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_, _1482_ } & _1070_;
assign _0529_ = { _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_, _1486_ } & _1071_;
assign _0532_ = { _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_, _1013_ } & _1089_;
assign _0535_ = { _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_, _1490_ } & _1073_;
assign _0538_ = { _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_, _1494_ } & _1074_;
assign _0541_ = { _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_, _1015_ } & _1090_;
assign _0544_ = { _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_ } & _1091_;
assign _0547_ = { _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_ } & _1092_;
assign _0550_ = { _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_, _0203_ } & _1093_;
assign _0555_ = _1308_ & we_a_i;
assign _0557_ = _1310_ & we_a_i;
assign _0559_ = _1312_ & we_a_i;
assign _0561_ = _1314_ & we_a_i;
assign _0563_ = _1316_ & we_a_i;
assign _0565_ = _1318_ & we_a_i;
assign _0567_ = _1320_ & we_a_i;
assign _0569_ = _1322_ & we_a_i;
assign _0571_ = _1324_ & we_a_i;
assign _0573_ = _1326_ & we_a_i;
assign _0575_ = _1328_ & we_a_i;
assign _0577_ = _1330_ & we_a_i;
assign _0579_ = _1332_ & we_a_i;
assign _0581_ = _1334_ & we_a_i;
assign _0583_ = _1336_ & we_a_i;
assign _0585_ = _1338_ & we_a_i;
assign _0587_ = _1340_ & we_a_i;
assign _0589_ = _1342_ & we_a_i;
assign _0591_ = _1344_ & we_a_i;
assign _0593_ = _1346_ & we_a_i;
assign _0595_ = _1348_ & we_a_i;
assign _0597_ = _1350_ & we_a_i;
assign _0599_ = _1352_ & we_a_i;
assign _0601_ = _1354_ & we_a_i;
assign _0603_ = _1356_ & we_a_i;
assign _0605_ = _1358_ & we_a_i;
assign _0607_ = _1360_ & we_a_i;
assign _0609_ = _1362_ & we_a_i;
assign _0611_ = _1364_ & we_a_i;
assign _0613_ = _1366_ & we_a_i;
assign _0615_ = _1368_ & we_a_i;
assign _0617_ = _1370_ & we_a_i;
assign _0619_ = { dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0, dummy_instr_id_i_t0 } & { \g_dummy_r0.rf_r0_q [38], _0143_[2], \g_dummy_r0.rf_r0_q [36], _0143_[1], \g_dummy_r0.rf_r0_q [34], _0143_[0], \g_dummy_r0.rf_r0_q [32:0] };
assign _1188_ = _0367_ | _0767_;
assign _1190_ = _0370_ | _0770_;
assign _1192_ = _0373_ | _0773_;
assign _1194_ = _0376_ | _0776_;
assign _1196_ = _0379_ | _0779_;
assign _1198_ = _0382_ | _0782_;
assign _1200_ = _0385_ | _0785_;
assign _1202_ = _0388_ | _0788_;
assign _1204_ = _0391_ | _0791_;
assign _1206_ = _0394_ | _0794_;
assign _1208_ = _0397_ | _0797_;
assign _1210_ = _0400_ | _0800_;
assign _1212_ = _0403_ | _0803_;
assign _1214_ = _0406_ | _0806_;
assign _1216_ = _0409_ | _0809_;
assign _1218_ = _0412_ | _0812_;
assign _1220_ = _0415_ | _0815_;
assign _1222_ = _0418_ | _0818_;
assign _1224_ = _0421_ | _0821_;
assign _1226_ = _0424_ | _0824_;
assign _1228_ = _0427_ | _0827_;
assign _1230_ = _0430_ | _0830_;
assign _1232_ = _0433_ | _0833_;
assign _1234_ = _0436_ | _0836_;
assign _1236_ = _0439_ | _0839_;
assign _1238_ = _0442_ | _0842_;
assign _1240_ = _0445_ | _0845_;
assign _1242_ = _0448_ | _0848_;
assign _1244_ = _0451_ | _0851_;
assign _1246_ = _0454_ | _0854_;
assign rdata_b_o_t0 = _0457_ | _0857_;
assign _1248_ = _0460_ | _0860_;
assign _1250_ = _0463_ | _0863_;
assign _1252_ = _0466_ | _0866_;
assign _1254_ = _0469_ | _0869_;
assign _1256_ = _0472_ | _0872_;
assign _1258_ = _0475_ | _0875_;
assign _1260_ = _0478_ | _0878_;
assign _1262_ = _0481_ | _0881_;
assign _1264_ = _0484_ | _0884_;
assign _1266_ = _0487_ | _0887_;
assign _1268_ = _0490_ | _0890_;
assign _1270_ = _0493_ | _0893_;
assign _1272_ = _0496_ | _0896_;
assign _1274_ = _0499_ | _0899_;
assign _1276_ = _0502_ | _0902_;
assign _1278_ = _0505_ | _0905_;
assign _1280_ = _0508_ | _0908_;
assign _1282_ = _0511_ | _0911_;
assign _1284_ = _0514_ | _0914_;
assign _1286_ = _0517_ | _0917_;
assign _1288_ = _0520_ | _0920_;
assign _1290_ = _0523_ | _0923_;
assign _1292_ = _0526_ | _0926_;
assign _1294_ = _0529_ | _0929_;
assign _1296_ = _0532_ | _0932_;
assign _1298_ = _0535_ | _0935_;
assign _1300_ = _0538_ | _0938_;
assign _1302_ = _0541_ | _0941_;
assign _1304_ = _0544_ | _0944_;
assign _1306_ = _0547_ | _0947_;
assign rdata_a_o_t0 = _0550_ | _0950_;
assign we_a_dec_t0[0] = _0555_ | _0554_;
assign we_a_dec_t0[1] = _0557_ | _0556_;
assign we_a_dec_t0[2] = _0559_ | _0558_;
assign we_a_dec_t0[3] = _0561_ | _0560_;
assign we_a_dec_t0[4] = _0563_ | _0562_;
assign we_a_dec_t0[5] = _0565_ | _0564_;
assign we_a_dec_t0[6] = _0567_ | _0566_;
assign we_a_dec_t0[7] = _0569_ | _0568_;
assign we_a_dec_t0[8] = _0571_ | _0570_;
assign we_a_dec_t0[9] = _0573_ | _0572_;
assign we_a_dec_t0[10] = _0575_ | _0574_;
assign we_a_dec_t0[11] = _0577_ | _0576_;
assign we_a_dec_t0[12] = _0579_ | _0578_;
assign we_a_dec_t0[13] = _0581_ | _0580_;
assign we_a_dec_t0[14] = _0583_ | _0582_;
assign we_a_dec_t0[15] = _0585_ | _0584_;
assign we_a_dec_t0[16] = _0587_ | _0586_;
assign we_a_dec_t0[17] = _0589_ | _0588_;
assign we_a_dec_t0[18] = _0591_ | _0590_;
assign we_a_dec_t0[19] = _0593_ | _0592_;
assign we_a_dec_t0[20] = _0595_ | _0594_;
assign we_a_dec_t0[21] = _0597_ | _0596_;
assign we_a_dec_t0[22] = _0599_ | _0598_;
assign we_a_dec_t0[23] = _0601_ | _0600_;
assign we_a_dec_t0[24] = _0603_ | _0602_;
assign we_a_dec_t0[25] = _0605_ | _0604_;
assign we_a_dec_t0[26] = _0607_ | _0606_;
assign we_a_dec_t0[27] = _0609_ | _0608_;
assign we_a_dec_t0[28] = _0611_ | _0610_;
assign we_a_dec_t0[29] = _0613_ | _0612_;
assign we_a_dec_t0[30] = _0615_ | _0614_;
assign we_a_dec_t0[31] = _0617_ | _0616_;
assign \rf_reg[0]_t0  = _0619_ | _0618_;
assign _0143_ = ~ { \g_dummy_r0.rf_r0_q [37], \g_dummy_r0.rf_r0_q [35], \g_dummy_r0.rf_r0_q [33] };
assign _0144_ = ~ _1373_;
assign _0145_ = ~ _1381_;
assign _0146_ = ~ _1389_;
assign _0147_ = ~ _1397_;
assign _0148_ = ~ _1405_;
assign _0149_ = ~ _1413_;
assign _0150_ = ~ _1421_;
assign _0151_ = ~ _1429_;
assign _0152_ = ~ _1435_;
assign _0153_ = ~ _1443_;
assign _0154_ = ~ _1451_;
assign _0155_ = ~ _1459_;
assign _0156_ = ~ _1467_;
assign _0157_ = ~ _1475_;
assign _0158_ = ~ _1483_;
assign _0159_ = ~ _1491_;
assign _0160_ = ~ _1371_;
assign _0161_ = ~ _1379_;
assign _0162_ = ~ _1387_;
assign _0163_ = ~ _1395_;
assign _0164_ = ~ _1403_;
assign _0165_ = ~ _1411_;
assign _0166_ = ~ _1419_;
assign _0167_ = ~ _1427_;
assign _0168_ = ~ _1433_;
assign _0169_ = ~ _1441_;
assign _0170_ = ~ _1449_;
assign _0171_ = ~ _1457_;
assign _0172_ = ~ _1465_;
assign _0173_ = ~ _1473_;
assign _0174_ = ~ _1481_;
assign _0175_ = ~ _1489_;
assign _0303_ = _1374_ & _0160_;
assign _0306_ = _1382_ & _0161_;
assign _0309_ = _1390_ & _0162_;
assign _0312_ = _1398_ & _0163_;
assign _0315_ = _1406_ & _0164_;
assign _0318_ = _1414_ & _0165_;
assign _0321_ = _1422_ & _0166_;
assign _0324_ = _1430_ & _0167_;
assign _0327_ = _1436_ & _0168_;
assign _0330_ = _1444_ & _0169_;
assign _0333_ = _1452_ & _0170_;
assign _0336_ = _1460_ & _0171_;
assign _0339_ = _1468_ & _0172_;
assign _0342_ = _1476_ & _0173_;
assign _0345_ = _1484_ & _0174_;
assign _0348_ = _1492_ & _0175_;
assign _0304_ = _1372_ & _0144_;
assign _0307_ = _1380_ & _0145_;
assign _0310_ = _1388_ & _0146_;
assign _0313_ = _1396_ & _0147_;
assign _0316_ = _1404_ & _0148_;
assign _0319_ = _1412_ & _0149_;
assign _0322_ = _1420_ & _0150_;
assign _0325_ = _1428_ & _0151_;
assign _0328_ = _1434_ & _0152_;
assign _0331_ = _1442_ & _0153_;
assign _0334_ = _1450_ & _0154_;
assign _0337_ = _1458_ & _0155_;
assign _0340_ = _1466_ & _0156_;
assign _0343_ = _1474_ & _0157_;
assign _0346_ = _1482_ & _0158_;
assign _0349_ = _1490_ & _0159_;
assign _0305_ = _1374_ & _1372_;
assign _0308_ = _1382_ & _1380_;
assign _0311_ = _1390_ & _1388_;
assign _0314_ = _1398_ & _1396_;
assign _0317_ = _1406_ & _1404_;
assign _0320_ = _1414_ & _1412_;
assign _0323_ = _1422_ & _1420_;
assign _0326_ = _1430_ & _1428_;
assign _0329_ = _1436_ & _1434_;
assign _0332_ = _1444_ & _1442_;
assign _0335_ = _1452_ & _1450_;
assign _0338_ = _1460_ & _1458_;
assign _0341_ = _1468_ & _1466_;
assign _0344_ = _1476_ & _1474_;
assign _0347_ = _1484_ & _1482_;
assign _0350_ = _1492_ & _1490_;
assign _0749_ = _0303_ | _0304_;
assign _0750_ = _0306_ | _0307_;
assign _0751_ = _0309_ | _0310_;
assign _0752_ = _0312_ | _0313_;
assign _0753_ = _0315_ | _0316_;
assign _0754_ = _0318_ | _0319_;
assign _0755_ = _0321_ | _0322_;
assign _0756_ = _0324_ | _0325_;
assign _0757_ = _0327_ | _0328_;
assign _0758_ = _0330_ | _0331_;
assign _0759_ = _0333_ | _0334_;
assign _0760_ = _0336_ | _0337_;
assign _0761_ = _0339_ | _0340_;
assign _0762_ = _0342_ | _0343_;
assign _0763_ = _0345_ | _0346_;
assign _0764_ = _0348_ | _0349_;
assign _0985_ = _0749_ | _0305_;
assign _0987_ = _0750_ | _0308_;
assign _0989_ = _0751_ | _0311_;
assign _0991_ = _0752_ | _0314_;
assign _0993_ = _0753_ | _0317_;
assign _0995_ = _0754_ | _0320_;
assign _0997_ = _0755_ | _0323_;
assign _0999_ = _0756_ | _0326_;
assign _1001_ = _0757_ | _0329_;
assign _1003_ = _0758_ | _0332_;
assign _1005_ = _0759_ | _0335_;
assign _1007_ = _0760_ | _0338_;
assign _1009_ = _0761_ | _0341_;
assign _1011_ = _0762_ | _0344_;
assign _1013_ = _0763_ | _0347_;
assign _1015_ = _0764_ | _0350_;
assign _0984_ = _1373_ | _1371_;
assign _0986_ = _1381_ | _1379_;
assign _0988_ = _1389_ | _1387_;
assign _0990_ = _1397_ | _1395_;
assign _0992_ = _1405_ | _1403_;
assign _0994_ = _1413_ | _1411_;
assign _0996_ = _1421_ | _1419_;
assign _0998_ = _1429_ | _1427_;
assign _1000_ = _1435_ | _1433_;
assign _1002_ = _1443_ | _1441_;
assign _1004_ = _1451_ | _1449_;
assign _1006_ = _1459_ | _1457_;
assign _1008_ = _1467_ | _1465_;
assign _1010_ = _1475_ | _1473_;
assign _1012_ = _1483_ | _1481_;
assign _1014_ = _1491_ | _1489_;
assign _0176_ = | { _0984_, _1377_, _1375_ };
assign _0178_ = | { _0988_, _1393_, _1391_ };
assign _0180_ = | { _0984_, _0986_, _1385_, _1383_, _1377_, _1375_ };
assign _0182_ = | { _0992_, _1409_, _1407_ };
assign _0184_ = | { _0996_, _1425_, _1423_ };
assign _0186_ = | { _0992_, _0994_, _1417_, _1415_, _1409_, _1407_ };
assign _0188_ = | { _0984_, _0986_, _0988_, _0990_, _1399_, _1401_, _1393_, _1391_, _1385_, _1383_, _1377_, _1375_ };
assign _0190_ = | { _1000_, _1437_, _1439_ };
assign _0192_ = | { _1004_, _1455_, _1453_ };
assign _0194_ = | { _1000_, _1002_, _1447_, _1445_, _1437_, _1439_ };
assign _0196_ = | { _1008_, _1471_, _1469_ };
assign _0198_ = | { _1012_, _1487_, _1485_ };
assign _0200_ = | { _1008_, _1010_, _1479_, _1477_, _1471_, _1469_ };
assign _0202_ = | { _1000_, _1002_, _1004_, _1006_, _1463_, _1461_, _1455_, _1453_, _1447_, _1445_, _1437_, _1439_ };
assign _1187_ = _1371_ ? \g_rf_flops[31].rf_reg_q  : \g_rf_flops[30].rf_reg_q ;
assign _1189_ = _1375_ ? \g_rf_flops[29].rf_reg_q  : \g_rf_flops[28].rf_reg_q ;
assign _1191_ = _0984_ ? _1187_ : _1189_;
assign _1193_ = _1379_ ? \g_rf_flops[27].rf_reg_q  : \g_rf_flops[26].rf_reg_q ;
assign _1195_ = _1383_ ? \g_rf_flops[25].rf_reg_q  : \g_rf_flops[24].rf_reg_q ;
assign _1197_ = _0986_ ? _1193_ : _1195_;
assign _1199_ = _0176_ ? _1191_ : _1197_;
assign _1201_ = _1387_ ? \g_rf_flops[23].rf_reg_q  : \g_rf_flops[22].rf_reg_q ;
assign _1203_ = _1391_ ? \g_rf_flops[21].rf_reg_q  : \g_rf_flops[20].rf_reg_q ;
assign _1205_ = _0988_ ? _1201_ : _1203_;
assign _1207_ = _1395_ ? \g_rf_flops[19].rf_reg_q  : \g_rf_flops[18].rf_reg_q ;
assign _1209_ = _1399_ ? \g_rf_flops[17].rf_reg_q  : \g_rf_flops[16].rf_reg_q ;
assign _1211_ = _0990_ ? _1207_ : _1209_;
assign _1213_ = _0178_ ? _1205_ : _1211_;
assign _1215_ = _0180_ ? _1199_ : _1213_;
assign _1217_ = _1403_ ? \g_rf_flops[15].rf_reg_q  : \g_rf_flops[14].rf_reg_q ;
assign _1219_ = _1407_ ? \g_rf_flops[13].rf_reg_q  : \g_rf_flops[12].rf_reg_q ;
assign _1221_ = _0992_ ? _1217_ : _1219_;
assign _1223_ = _1411_ ? \g_rf_flops[11].rf_reg_q  : \g_rf_flops[10].rf_reg_q ;
assign _1225_ = _1415_ ? \g_rf_flops[9].rf_reg_q  : \g_rf_flops[8].rf_reg_q ;
assign _1227_ = _0994_ ? _1223_ : _1225_;
assign _1229_ = _0182_ ? _1221_ : _1227_;
assign _1231_ = _1419_ ? \g_rf_flops[7].rf_reg_q  : \g_rf_flops[6].rf_reg_q ;
assign _1233_ = _1423_ ? \g_rf_flops[5].rf_reg_q  : \g_rf_flops[4].rf_reg_q ;
assign _1235_ = _0996_ ? _1231_ : _1233_;
assign _1237_ = _1427_ ? \g_rf_flops[3].rf_reg_q  : \g_rf_flops[2].rf_reg_q ;
assign _1239_ = _1431_ ? \g_rf_flops[1].rf_reg_q  : \rf_reg[0] ;
assign _1241_ = _0998_ ? _1237_ : _1239_;
assign _1243_ = _0184_ ? _1235_ : _1241_;
assign _1245_ = _0186_ ? _1229_ : _1243_;
assign rdata_b_o = _0188_ ? _1215_ : _1245_;
assign _1247_ = _1433_ ? \g_rf_flops[31].rf_reg_q  : \g_rf_flops[30].rf_reg_q ;
assign _1249_ = _1437_ ? \g_rf_flops[29].rf_reg_q  : \g_rf_flops[28].rf_reg_q ;
assign _1251_ = _1000_ ? _1247_ : _1249_;
assign _1253_ = _1441_ ? \g_rf_flops[27].rf_reg_q  : \g_rf_flops[26].rf_reg_q ;
assign _1255_ = _1445_ ? \g_rf_flops[25].rf_reg_q  : \g_rf_flops[24].rf_reg_q ;
assign _1257_ = _1002_ ? _1253_ : _1255_;
assign _1259_ = _0190_ ? _1251_ : _1257_;
assign _1261_ = _1449_ ? \g_rf_flops[23].rf_reg_q  : \g_rf_flops[22].rf_reg_q ;
assign _1263_ = _1453_ ? \g_rf_flops[21].rf_reg_q  : \g_rf_flops[20].rf_reg_q ;
assign _1265_ = _1004_ ? _1261_ : _1263_;
assign _1267_ = _1457_ ? \g_rf_flops[19].rf_reg_q  : \g_rf_flops[18].rf_reg_q ;
assign _1269_ = _1461_ ? \g_rf_flops[17].rf_reg_q  : \g_rf_flops[16].rf_reg_q ;
assign _1271_ = _1006_ ? _1267_ : _1269_;
assign _1273_ = _0192_ ? _1265_ : _1271_;
assign _1275_ = _0194_ ? _1259_ : _1273_;
assign _1277_ = _1465_ ? \g_rf_flops[15].rf_reg_q  : \g_rf_flops[14].rf_reg_q ;
assign _1279_ = _1469_ ? \g_rf_flops[13].rf_reg_q  : \g_rf_flops[12].rf_reg_q ;
assign _1281_ = _1008_ ? _1277_ : _1279_;
assign _1283_ = _1473_ ? \g_rf_flops[11].rf_reg_q  : \g_rf_flops[10].rf_reg_q ;
assign _1285_ = _1477_ ? \g_rf_flops[9].rf_reg_q  : \g_rf_flops[8].rf_reg_q ;
assign _1287_ = _1010_ ? _1283_ : _1285_;
assign _1289_ = _0196_ ? _1281_ : _1287_;
assign _1291_ = _1481_ ? \g_rf_flops[7].rf_reg_q  : \g_rf_flops[6].rf_reg_q ;
assign _1293_ = _1485_ ? \g_rf_flops[5].rf_reg_q  : \g_rf_flops[4].rf_reg_q ;
assign _1295_ = _1012_ ? _1291_ : _1293_;
assign _1297_ = _1489_ ? \g_rf_flops[3].rf_reg_q  : \g_rf_flops[2].rf_reg_q ;
assign _1299_ = _1493_ ? \g_rf_flops[1].rf_reg_q  : \rf_reg[0] ;
assign _1301_ = _1014_ ? _1297_ : _1299_;
assign _1303_ = _0198_ ? _1295_ : _1301_;
assign _1305_ = _0200_ ? _1289_ : _1303_;
assign rdata_a_o = _0202_ ? _1275_ : _1305_;
assign _1307_ = ! /* src = "generated/sv2v_out.v:20074.20-20074.47" */ waddr_a_i;
assign _1309_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h01;
assign _1311_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h02;
assign _1313_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h03;
assign _1315_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h04;
assign _1317_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h05;
assign _1319_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h06;
assign _1321_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h07;
assign _1323_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h08;
assign _1325_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h09;
assign _1327_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h0a;
assign _1329_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h0b;
assign _1331_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h0c;
assign _1333_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h0d;
assign _1335_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h0e;
assign _1337_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h0f;
assign _1339_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h10;
assign _1341_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h11;
assign _1343_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h12;
assign _1345_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h13;
assign _1347_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h14;
assign _1349_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h15;
assign _1351_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h16;
assign _1353_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h17;
assign _1355_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h18;
assign _1357_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h19;
assign _1359_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h1a;
assign _1361_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h1b;
assign _1363_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h1c;
assign _1365_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h1d;
assign _1367_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h1e;
assign _1369_ = waddr_a_i == /* src = "generated/sv2v_out.v:20074.20-20074.47" */ 5'h1f;
assign _1371_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1f;
assign _1373_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1e;
assign _1375_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1d;
assign _1377_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1c;
assign _1379_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1b;
assign _1381_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1a;
assign _1383_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h19;
assign _1385_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h18;
assign _1387_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h17;
assign _1389_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h16;
assign _1391_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h15;
assign _1393_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h14;
assign _1395_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h13;
assign _1397_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h12;
assign _1399_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h11;
assign _1401_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h10;
assign _1403_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0f;
assign _1405_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0e;
assign _1407_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0d;
assign _1409_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0c;
assign _1411_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0b;
assign _1413_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0a;
assign _1415_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h09;
assign _1417_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h08;
assign _1419_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h07;
assign _1421_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h06;
assign _1423_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h05;
assign _1425_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h04;
assign _1427_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h03;
assign _1429_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h02;
assign _1431_ = raddr_b_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h01;
assign _1433_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1f;
assign _1435_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1e;
assign _1437_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1d;
assign _1439_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1c;
assign _1441_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1b;
assign _1443_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1a;
assign _1445_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h19;
assign _1447_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h18;
assign _1449_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h17;
assign _1451_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h16;
assign _1453_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h15;
assign _1455_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h14;
assign _1457_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h13;
assign _1459_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h12;
assign _1461_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h11;
assign _1463_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h10;
assign _1465_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0f;
assign _1467_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0e;
assign _1469_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0d;
assign _1471_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0c;
assign _1473_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0b;
assign _1475_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0a;
assign _1477_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h09;
assign _1479_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h08;
assign _1481_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h07;
assign _1483_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h06;
assign _1485_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h05;
assign _1487_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h04;
assign _1489_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h03;
assign _1491_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h02;
assign _1493_ = raddr_a_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h01;
assign we_a_dec[0] = _1307_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[1] = _1309_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[2] = _1311_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[3] = _1313_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[4] = _1315_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[5] = _1317_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[6] = _1319_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[7] = _1321_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[8] = _1323_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[9] = _1325_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[10] = _1327_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[11] = _1329_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[12] = _1331_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[13] = _1333_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[14] = _1335_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[15] = _1337_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[16] = _1339_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[17] = _1341_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[18] = _1343_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[19] = _1345_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[20] = _1347_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[21] = _1349_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[22] = _1351_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[23] = _1353_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[24] = _1355_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[25] = _1357_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[26] = _1359_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[27] = _1361_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[28] = _1363_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[29] = _1365_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[30] = _1367_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign we_a_dec[31] = _1369_ ? /* src = "generated/sv2v_out.v:20074.20-20074.63" */ we_a_i : 1'h0;
assign \rf_reg[0]  = dummy_instr_id_i ? /* src = "generated/sv2v_out.v:20123.24-20123.64" */ \g_dummy_r0.rf_r0_q  : 39'h2a00000000;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20080.34-20083.5" */
\$paramod\prim_buf\Width=32'00000000000000000000000000100000  \gen_wren_check.u_prim_buf  (
.in_i(we_a_dec),
.in_i_t0(we_a_dec_t0),
.out_o(\gen_wren_check.we_a_dec_buf ),
.out_o_t0(\gen_wren_check.we_a_dec_buf_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20088.6-20095.5" */
\$paramod$916c47de983e2a42946808797a4a11650abb788f\prim_onehot_check  \gen_wren_check.u_prim_onehot_check  (
.addr_i(waddr_a_i),
.addr_i_t0(waddr_a_i_t0),
.clk_i(clk_i),
.en_i(we_a_i),
.en_i_t0(we_a_i_t0),
.err_o(err_o),
.err_o_t0(err_o_t0),
.oh_i(\gen_wren_check.we_a_dec_buf ),
.oh_i_t0(\gen_wren_check.we_a_dec_buf_t0 ),
.rst_ni(rst_ni)
);
endmodule

module \$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers (clk_i, rst_ni, hart_id_i, priv_mode_id_o, priv_mode_lsu_o, csr_mstatus_tw_o, csr_mtvec_o, csr_mtvec_init_i, boot_addr_i, csr_access_i, csr_addr_i, csr_wdata_i, csr_op_i, csr_op_en_i, csr_rdata_o, irq_software_i, irq_timer_i, irq_external_i, irq_fast_i, nmi_mode_i, irq_pending_o
, irqs_o, csr_mstatus_mie_o, csr_mepc_o, csr_mtval_o, csr_pmp_cfg_o, csr_pmp_addr_o, csr_pmp_mseccfg_o, debug_mode_i, debug_mode_entering_i, debug_cause_i, debug_csr_save_i, csr_depc_o, debug_single_step_o, debug_ebreakm_o, debug_ebreaku_o, trigger_match_o, pc_if_i, pc_id_i, pc_wb_i, data_ind_timing_o, dummy_instr_en_o
, dummy_instr_mask_o, dummy_instr_seed_en_o, dummy_instr_seed_o, icache_enable_o, csr_shadow_err_o, ic_scr_key_valid_i, csr_save_if_i, csr_save_id_i, csr_save_wb_i, csr_restore_mret_i, csr_restore_dret_i, csr_save_cause_i, csr_mcause_i, csr_mtval_i, illegal_csr_insn_o, double_fault_seen_o, instr_ret_i, instr_ret_compressed_i, instr_ret_spec_i, instr_ret_compressed_spec_i, iside_wait_i
, jump_i, branch_i, branch_taken_i, mem_load_i, mem_store_i, dside_wait_i, mul_wait_i, div_wait_i, branch_taken_i_t0, csr_mtval_o_t0, pc_id_i_t0, ic_scr_key_valid_i_t0, boot_addr_i_t0, branch_i_t0, csr_access_i_t0, csr_addr_i_t0, csr_depc_o_t0, csr_mcause_i_t0, csr_mepc_o_t0, csr_mstatus_mie_o_t0, csr_mstatus_tw_o_t0
, csr_mtval_i_t0, csr_mtvec_init_i_t0, csr_mtvec_o_t0, csr_op_en_i_t0, csr_op_i_t0, csr_pmp_addr_o_t0, csr_pmp_cfg_o_t0, csr_pmp_mseccfg_o_t0, csr_rdata_o_t0, csr_restore_dret_i_t0, csr_restore_mret_i_t0, csr_save_cause_i_t0, csr_save_id_i_t0, csr_save_if_i_t0, csr_save_wb_i_t0, csr_shadow_err_o_t0, csr_wdata_i_t0, data_ind_timing_o_t0, debug_cause_i_t0, debug_csr_save_i_t0, debug_ebreakm_o_t0
, debug_ebreaku_o_t0, debug_mode_entering_i_t0, debug_mode_i_t0, debug_single_step_o_t0, div_wait_i_t0, double_fault_seen_o_t0, dside_wait_i_t0, dummy_instr_en_o_t0, dummy_instr_mask_o_t0, dummy_instr_seed_en_o_t0, dummy_instr_seed_o_t0, hart_id_i_t0, icache_enable_o_t0, illegal_csr_insn_o_t0, instr_ret_compressed_i_t0, instr_ret_compressed_spec_i_t0, instr_ret_i_t0, instr_ret_spec_i_t0, irq_external_i_t0, irq_fast_i_t0, irq_pending_o_t0
, irq_software_i_t0, irq_timer_i_t0, irqs_o_t0, iside_wait_i_t0, jump_i_t0, mem_load_i_t0, mem_store_i_t0, mul_wait_i_t0, nmi_mode_i_t0, pc_if_i_t0, pc_wb_i_t0, priv_mode_id_o_t0, priv_mode_lsu_o_t0, trigger_match_o_t0);
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [7:0] _0000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [7:0] _0001_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0003_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0005_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0007_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0009_;
/* src = "generated/sv2v_out.v:13959.2-14089.5" */
wire _0010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13959.2-14089.5" */
wire _0011_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0013_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0015_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [5:0] _0016_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [5:0] _0017_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0018_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0019_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0021_;
/* src = "generated/sv2v_out.v:13959.2-14089.5" */
wire [63:0] _0022_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13959.2-14089.5" */
wire [63:0] _0023_;
/* src = "generated/sv2v_out.v:13959.2-14089.5" */
wire [31:0] _0024_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [7:0] _0025_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [7:0] _0026_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0027_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0028_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0029_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0030_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0031_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0032_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0033_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0034_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0035_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0036_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0037_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0038_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0039_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0040_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0041_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0042_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0043_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0044_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [6:0] _0045_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [6:0] _0046_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0047_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0048_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0049_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0050_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0051_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0052_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0053_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0054_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0055_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0056_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0057_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0058_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0059_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0060_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0061_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0062_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0063_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0064_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [5:0] _0065_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [5:0] _0066_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0067_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0068_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0069_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0070_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0071_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0072_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0073_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0074_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [1:0] _0075_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [1:0] _0076_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0077_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0078_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [6:0] _0079_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [6:0] _0080_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0081_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0082_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0083_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [1:0] _0084_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [1:0] _0085_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0086_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0087_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [1:0] _0088_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [1:0] _0089_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0090_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0091_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0092_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0093_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0094_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0095_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0096_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0097_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [6:0] _0098_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [6:0] _0099_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0100_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0101_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0102_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [31:0] _0103_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0104_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0105_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0106_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0107_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0108_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0109_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [1:0] _0110_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [1:0] _0111_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0112_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0113_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0114_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0115_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0116_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0117_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0118_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [3:0] _0119_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [3:0] _0120_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0121_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0122_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0123_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0124_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [1:0] _0125_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [1:0] _0126_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0127_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0128_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [1:0] _0129_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [1:0] _0130_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0131_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0132_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0133_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0134_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [3:0] _0135_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [3:0] _0136_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0137_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0138_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [2:0] _0139_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [2:0] _0140_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0141_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire _0142_;
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [2:0] _0143_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14094.2-14233.5" */
wire [2:0] _0144_;
/* src = "generated/sv2v_out.v:14245.26-14245.52" */
wire [31:0] _0145_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14245.26-14245.52" */
wire [31:0] _0146_;
/* src = "generated/sv2v_out.v:14250.23-14250.43" */
wire _0147_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14250.23-14250.43" */
wire _0148_;
/* src = "generated/sv2v_out.v:14622.18-14622.57" */
wire _0149_;
/* src = "generated/sv2v_out.v:14634.18-14634.57" */
wire _0150_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14634.18-14634.57" */
wire _0151_;
/* src = "generated/sv2v_out.v:14641.27-14641.63" */
wire _0152_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14641.27-14641.63" */
wire _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire [1:0] _0164_;
wire [1:0] _0165_;
wire [1:0] _0166_;
wire [1:0] _0167_;
wire [1:0] _0168_;
wire [1:0] _0169_;
wire [11:0] _0170_;
wire [4:0] _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire _0186_;
wire _0187_;
wire _0188_;
wire _0189_;
wire _0190_;
wire _0191_;
wire _0192_;
wire _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire [2:0] _0199_;
wire [135:0] _0200_;
wire [3:0] _0201_;
wire [1:0] _0202_;
wire [29:0] _0203_;
wire [64:0] _0204_;
wire [60:0] _0205_;
wire [64:0] _0206_;
wire [2:0] _0207_;
wire [33:0] _0208_;
wire [33:0] _0209_;
wire [90:0] _0210_;
wire [2:0] _0211_;
wire [93:0] _0212_;
wire [30:0] _0213_;
wire [2:0] _0214_;
wire [63:0] _0215_;
wire [30:0] _0216_;
wire [30:0] _0217_;
wire [28:0] _0218_;
wire [19:0] _0219_;
wire [2:0] _0220_;
wire [17:0] _0221_;
wire _0222_;
wire _0223_;
wire _0224_;
wire _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire _0241_;
wire _0242_;
wire _0243_;
wire _0244_;
wire _0245_;
wire _0246_;
wire _0247_;
wire _0248_;
wire _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire [2:0] _0267_;
wire [2:0] _0268_;
wire [2:0] _0269_;
wire [2:0] _0270_;
wire [2:0] _0271_;
wire [2:0] _0272_;
wire [2:0] _0273_;
wire [2:0] _0274_;
wire [2:0] _0275_;
wire [2:0] _0276_;
wire [2:0] _0277_;
wire [2:0] _0278_;
wire [2:0] _0279_;
wire [2:0] _0280_;
wire [2:0] _0281_;
wire [2:0] _0282_;
wire [2:0] _0283_;
wire [2:0] _0284_;
wire [2:0] _0285_;
wire [2:0] _0286_;
wire [2:0] _0287_;
wire [2:0] _0288_;
wire [2:0] _0289_;
wire [2:0] _0290_;
wire [2:0] _0291_;
wire [2:0] _0292_;
wire [2:0] _0293_;
wire [2:0] _0294_;
wire _0295_;
wire _0296_;
wire _0297_;
wire _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire [2:0] _0309_;
wire [2:0] _0310_;
wire [2:0] _0311_;
wire [2:0] _0312_;
wire [8:0] _0313_;
wire [8:0] _0314_;
wire [8:0] _0315_;
wire [8:0] _0316_;
wire [8:0] _0317_;
wire [8:0] _0318_;
wire [8:0] _0319_;
wire [8:0] _0320_;
wire [8:0] _0321_;
wire [8:0] _0322_;
wire [8:0] _0323_;
wire [8:0] _0324_;
wire [8:0] _0325_;
wire [8:0] _0326_;
wire [8:0] _0327_;
wire [63:0] _0328_;
wire [63:0] _0329_;
wire [31:0] _0330_;
wire [31:0] _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire _0335_;
wire [2:0] _0336_;
wire [2:0] _0337_;
wire _0338_;
wire _0339_;
wire [31:0] _0340_;
wire _0341_;
wire [2:0] _0342_;
wire [2:0] _0343_;
wire [2:0] _0344_;
wire _0345_;
wire _0346_;
wire _0347_;
wire _0348_;
wire _0349_;
wire [1:0] _0350_;
wire [6:0] _0351_;
wire [31:0] _0352_;
wire _0353_;
wire [31:0] _0354_;
wire [2:0] _0355_;
wire [1:0] _0356_;
wire [6:0] _0357_;
wire [3:0] _0358_;
wire [31:0] _0359_;
wire [31:0] _0360_;
wire [31:0] _0361_;
wire [31:0] _0362_;
wire [1:0] _0363_;
wire [6:0] _0364_;
wire [6:0] _0365_;
wire [6:0] _0366_;
wire [31:0] _0367_;
wire [31:0] _0368_;
wire [6:0] _0369_;
wire [1:0] _0370_;
wire [3:0] _0371_;
wire [1:0] _0372_;
wire [11:0] _0373_;
wire [1:0] _0374_;
wire [1:0] _0375_;
wire [1:0] _0376_;
wire [7:0] _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire [7:0] _0381_;
wire [31:0] _0382_;
wire [5:0] _0383_;
wire _0384_;
wire [31:0] _0385_;
wire [1:0] _0386_;
wire [63:0] _0387_;
wire [31:0] _0388_;
wire [31:0] _0389_;
wire [31:0] _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire _0398_;
wire _0399_;
wire _0400_;
wire _0401_;
wire _0402_;
wire _0403_;
wire _0404_;
wire _0405_;
wire _0406_;
wire _0407_;
wire [1:0] _0408_;
wire _0409_;
wire _0410_;
wire _0411_;
wire _0412_;
wire _0413_;
wire [31:0] _0414_;
wire _0415_;
wire _0416_;
wire _0417_;
wire _0418_;
wire _0419_;
wire _0420_;
wire [31:0] _0421_;
wire _0422_;
wire _0423_;
wire _0424_;
wire _0425_;
/* cellift = 32'd1 */
wire _0426_;
wire _0427_;
/* cellift = 32'd1 */
wire _0428_;
wire _0429_;
/* cellift = 32'd1 */
wire _0430_;
wire _0431_;
/* cellift = 32'd1 */
wire _0432_;
wire _0433_;
/* cellift = 32'd1 */
wire _0434_;
wire _0435_;
/* cellift = 32'd1 */
wire _0436_;
wire _0437_;
/* cellift = 32'd1 */
wire _0438_;
wire _0439_;
/* cellift = 32'd1 */
wire _0440_;
wire _0441_;
/* cellift = 32'd1 */
wire _0442_;
wire _0443_;
/* cellift = 32'd1 */
wire _0444_;
wire _0445_;
/* cellift = 32'd1 */
wire _0446_;
wire _0447_;
/* cellift = 32'd1 */
wire _0448_;
wire _0449_;
wire _0450_;
wire _0451_;
wire _0452_;
/* cellift = 32'd1 */
wire _0453_;
wire _0454_;
wire _0455_;
wire _0456_;
/* cellift = 32'd1 */
wire _0457_;
wire _0458_;
/* cellift = 32'd1 */
wire _0459_;
wire _0460_;
wire _0461_;
wire _0462_;
wire _0463_;
wire _0464_;
wire _0465_;
wire [31:0] _0466_;
wire [31:0] _0467_;
wire [31:0] _0468_;
wire _0469_;
wire _0470_;
wire _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire [17:0] _0475_;
wire [17:0] _0476_;
wire [17:0] _0477_;
wire _0478_;
wire _0479_;
wire _0480_;
wire _0481_;
wire _0482_;
wire _0483_;
wire _0484_;
wire _0485_;
wire _0486_;
wire [1:0] _0487_;
wire [1:0] _0488_;
wire [1:0] _0489_;
wire [1:0] _0490_;
wire [1:0] _0491_;
wire [1:0] _0492_;
wire [2:0] _0493_;
wire [135:0] _0494_;
wire [3:0] _0495_;
wire [1:0] _0496_;
wire [29:0] _0497_;
wire _0498_;
wire _0499_;
wire _0500_;
wire _0501_;
wire _0502_;
wire _0503_;
wire _0504_;
wire _0505_;
wire _0506_;
wire _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0517_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
wire _0525_;
wire _0526_;
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire [64:0] _0534_;
wire [60:0] _0535_;
wire [64:0] _0536_;
wire [2:0] _0537_;
wire [33:0] _0538_;
wire [33:0] _0539_;
wire [90:0] _0540_;
wire [2:0] _0541_;
wire [93:0] _0542_;
wire [30:0] _0543_;
wire [2:0] _0544_;
wire [63:0] _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire _0560_;
wire _0561_;
wire _0562_;
wire _0563_;
wire _0564_;
wire _0565_;
wire _0566_;
wire _0567_;
wire _0568_;
wire _0569_;
wire _0570_;
wire _0571_;
wire _0572_;
wire _0573_;
wire _0574_;
wire _0575_;
wire _0576_;
wire _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire [2:0] _0595_;
wire [2:0] _0596_;
wire [2:0] _0597_;
wire [2:0] _0598_;
wire [2:0] _0599_;
wire [2:0] _0600_;
wire [2:0] _0601_;
wire [2:0] _0602_;
wire [2:0] _0603_;
wire [2:0] _0604_;
wire [2:0] _0605_;
wire [2:0] _0606_;
wire [2:0] _0607_;
wire [2:0] _0608_;
wire [2:0] _0609_;
wire [2:0] _0610_;
wire [2:0] _0611_;
wire [2:0] _0612_;
wire [2:0] _0613_;
wire [2:0] _0614_;
wire [2:0] _0615_;
wire [2:0] _0616_;
wire [2:0] _0617_;
wire [2:0] _0618_;
wire [2:0] _0619_;
wire [2:0] _0620_;
wire [2:0] _0621_;
wire [2:0] _0622_;
wire [2:0] _0623_;
wire [2:0] _0624_;
wire [2:0] _0625_;
wire [2:0] _0626_;
wire [2:0] _0627_;
wire [2:0] _0628_;
wire [2:0] _0629_;
wire [2:0] _0630_;
wire [2:0] _0631_;
wire [2:0] _0632_;
wire [2:0] _0633_;
wire [2:0] _0634_;
wire [2:0] _0635_;
wire [2:0] _0636_;
wire [2:0] _0637_;
wire [2:0] _0638_;
wire [2:0] _0639_;
wire [2:0] _0640_;
wire [2:0] _0641_;
wire [2:0] _0642_;
wire [2:0] _0643_;
wire [2:0] _0644_;
wire [2:0] _0645_;
wire [2:0] _0646_;
wire [2:0] _0647_;
wire [2:0] _0648_;
wire [2:0] _0649_;
wire [2:0] _0650_;
wire [2:0] _0651_;
wire [2:0] _0652_;
wire [2:0] _0653_;
wire [2:0] _0654_;
wire [2:0] _0655_;
wire [2:0] _0656_;
wire [2:0] _0657_;
wire [2:0] _0658_;
wire [2:0] _0659_;
wire [2:0] _0660_;
wire [2:0] _0661_;
wire [2:0] _0662_;
wire [2:0] _0663_;
wire [2:0] _0664_;
wire [2:0] _0665_;
wire [2:0] _0666_;
wire [2:0] _0667_;
wire [2:0] _0668_;
wire [2:0] _0669_;
wire [2:0] _0670_;
wire [2:0] _0671_;
wire [2:0] _0672_;
wire [2:0] _0673_;
wire [2:0] _0674_;
wire [2:0] _0675_;
wire [2:0] _0676_;
wire [2:0] _0677_;
wire [2:0] _0678_;
wire [2:0] _0679_;
wire [2:0] _0680_;
wire [2:0] _0681_;
wire [2:0] _0682_;
wire [2:0] _0683_;
wire [2:0] _0684_;
wire [2:0] _0685_;
wire [2:0] _0686_;
wire [2:0] _0687_;
wire [2:0] _0688_;
wire [2:0] _0689_;
wire [2:0] _0690_;
wire [2:0] _0691_;
wire [2:0] _0692_;
wire [2:0] _0693_;
wire [2:0] _0694_;
wire [2:0] _0695_;
wire [2:0] _0696_;
wire [2:0] _0697_;
wire [2:0] _0698_;
wire [2:0] _0699_;
wire [2:0] _0700_;
wire [2:0] _0701_;
wire [2:0] _0702_;
wire [2:0] _0703_;
wire [2:0] _0704_;
wire [2:0] _0705_;
wire [2:0] _0706_;
wire [2:0] _0707_;
wire [2:0] _0708_;
wire [2:0] _0709_;
wire [2:0] _0710_;
wire [2:0] _0711_;
wire [2:0] _0712_;
wire [2:0] _0713_;
wire [2:0] _0714_;
wire [2:0] _0715_;
wire [2:0] _0716_;
wire [2:0] _0717_;
wire [2:0] _0718_;
wire [2:0] _0719_;
wire [2:0] _0720_;
wire [2:0] _0721_;
wire [2:0] _0722_;
wire [2:0] _0723_;
wire _0724_;
wire _0725_;
wire _0726_;
wire _0727_;
wire _0728_;
wire _0729_;
wire _0730_;
wire _0731_;
wire _0732_;
wire _0733_;
wire _0734_;
wire _0735_;
wire _0736_;
wire _0737_;
wire _0738_;
wire _0739_;
wire _0740_;
wire _0741_;
wire _0742_;
wire _0743_;
wire _0744_;
wire _0745_;
wire _0746_;
wire _0747_;
wire _0748_;
wire _0749_;
wire _0750_;
wire _0751_;
wire _0752_;
wire _0753_;
wire _0754_;
wire _0755_;
wire _0756_;
wire _0757_;
wire _0758_;
wire _0759_;
wire _0760_;
wire _0761_;
wire _0762_;
wire _0763_;
wire _0764_;
wire _0765_;
wire _0766_;
wire _0767_;
wire _0768_;
wire _0769_;
wire _0770_;
wire _0771_;
wire _0772_;
wire _0773_;
wire _0774_;
wire _0775_;
wire _0776_;
wire _0777_;
wire _0778_;
wire _0779_;
wire _0780_;
wire _0781_;
wire _0782_;
wire _0783_;
wire _0784_;
wire _0785_;
wire _0786_;
wire _0787_;
wire _0788_;
wire _0789_;
wire _0790_;
wire _0791_;
wire _0792_;
wire _0793_;
wire _0794_;
wire _0795_;
wire _0796_;
wire _0797_;
wire _0798_;
wire _0799_;
wire _0800_;
wire _0801_;
wire _0802_;
wire _0803_;
wire _0804_;
wire _0805_;
wire _0806_;
wire _0807_;
wire _0808_;
wire _0809_;
wire _0810_;
wire _0811_;
wire [2:0] _0812_;
wire [2:0] _0813_;
wire [2:0] _0814_;
wire [2:0] _0815_;
wire [2:0] _0816_;
wire [2:0] _0817_;
wire [2:0] _0818_;
wire [2:0] _0819_;
wire [2:0] _0820_;
wire [2:0] _0821_;
wire [2:0] _0822_;
wire [2:0] _0823_;
wire [2:0] _0824_;
wire [2:0] _0825_;
wire [2:0] _0826_;
wire [2:0] _0827_;
wire [2:0] _0828_;
wire [2:0] _0829_;
wire [2:0] _0830_;
wire [2:0] _0831_;
wire [2:0] _0832_;
wire [2:0] _0833_;
wire [2:0] _0834_;
wire [2:0] _0835_;
wire [2:0] _0836_;
wire [2:0] _0837_;
wire [2:0] _0838_;
wire [2:0] _0839_;
wire [2:0] _0840_;
wire [2:0] _0841_;
wire [2:0] _0842_;
wire [2:0] _0843_;
wire [2:0] _0844_;
wire [2:0] _0845_;
wire [2:0] _0846_;
wire [2:0] _0847_;
wire [2:0] _0848_;
wire _0849_;
wire _0850_;
wire _0851_;
wire _0852_;
wire _0853_;
wire _0854_;
wire _0855_;
wire _0856_;
wire _0857_;
wire _0858_;
wire _0859_;
wire _0860_;
wire _0861_;
wire _0862_;
wire _0863_;
wire _0864_;
wire _0865_;
wire _0866_;
wire _0867_;
wire _0868_;
wire _0869_;
wire _0870_;
wire _0871_;
wire _0872_;
wire _0873_;
wire _0874_;
wire _0875_;
wire _0876_;
wire _0877_;
wire _0878_;
wire _0879_;
wire _0880_;
wire _0881_;
wire _0882_;
wire _0883_;
wire _0884_;
wire _0885_;
wire _0886_;
wire _0887_;
wire _0888_;
wire _0889_;
wire _0890_;
wire [8:0] _0891_;
wire [8:0] _0892_;
wire [8:0] _0893_;
wire [8:0] _0894_;
wire [8:0] _0895_;
wire [8:0] _0896_;
wire [8:0] _0897_;
wire [8:0] _0898_;
wire [8:0] _0899_;
wire [8:0] _0900_;
wire [8:0] _0901_;
wire [8:0] _0902_;
wire [8:0] _0903_;
wire [8:0] _0904_;
wire [8:0] _0905_;
wire [8:0] _0906_;
wire [8:0] _0907_;
wire [8:0] _0908_;
wire [8:0] _0909_;
wire [8:0] _0910_;
wire [8:0] _0911_;
wire [8:0] _0912_;
wire [8:0] _0913_;
wire [8:0] _0914_;
wire [8:0] _0915_;
wire [8:0] _0916_;
wire [8:0] _0917_;
wire [8:0] _0918_;
wire [8:0] _0919_;
wire [8:0] _0920_;
wire [8:0] _0921_;
wire [8:0] _0922_;
wire [8:0] _0923_;
wire [8:0] _0924_;
wire [8:0] _0925_;
wire [8:0] _0926_;
wire [8:0] _0927_;
wire [8:0] _0928_;
wire [8:0] _0929_;
wire [8:0] _0930_;
wire [8:0] _0931_;
wire [8:0] _0932_;
wire [8:0] _0933_;
wire [8:0] _0934_;
wire [8:0] _0935_;
wire _0936_;
wire _0937_;
wire _0938_;
wire _0939_;
wire _0940_;
wire _0941_;
wire _0942_;
wire _0943_;
wire _0944_;
wire _0945_;
wire _0946_;
wire _0947_;
wire _0948_;
wire _0949_;
wire _0950_;
wire _0951_;
wire _0952_;
wire _0953_;
wire _0954_;
wire _0955_;
wire _0956_;
wire _0957_;
wire _0958_;
wire _0959_;
wire _0960_;
wire _0961_;
wire _0962_;
wire _0963_;
wire _0964_;
wire _0965_;
wire _0966_;
wire _0967_;
wire _0968_;
wire _0969_;
wire _0970_;
wire _0971_;
wire _0972_;
wire _0973_;
wire _0974_;
wire _0975_;
wire _0976_;
wire _0977_;
wire _0978_;
wire _0979_;
wire _0980_;
wire [63:0] _0981_;
wire [63:0] _0982_;
wire [63:0] _0983_;
wire [63:0] _0984_;
wire [63:0] _0985_;
wire _0986_;
wire _0987_;
wire _0988_;
wire _0989_;
wire _0990_;
wire _0991_;
wire _0992_;
wire _0993_;
wire _0994_;
wire _0995_;
wire _0996_;
wire _0997_;
wire _0998_;
wire _0999_;
wire _1000_;
wire _1001_;
wire _1002_;
wire _1003_;
wire _1004_;
wire _1005_;
wire _1006_;
wire _1007_;
wire _1008_;
wire _1009_;
wire _1010_;
wire _1011_;
wire _1012_;
wire _1013_;
wire _1014_;
wire _1015_;
wire _1016_;
wire _1017_;
wire _1018_;
wire _1019_;
wire _1020_;
wire _1021_;
wire _1022_;
wire _1023_;
wire _1024_;
wire _1025_;
wire _1026_;
wire _1027_;
wire _1028_;
wire _1029_;
wire _1030_;
wire [31:0] _1031_;
wire [31:0] _1032_;
wire [31:0] _1033_;
wire [31:0] _1034_;
wire [31:0] _1035_;
wire [31:0] _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire _1045_;
wire _1046_;
wire _1047_;
wire _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1052_;
wire _1053_;
wire _1054_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire _1061_;
wire _1062_;
wire _1063_;
wire _1064_;
wire _1065_;
wire _1066_;
wire _1067_;
wire _1068_;
wire _1069_;
wire _1070_;
wire _1071_;
wire _1072_;
wire _1073_;
wire _1074_;
wire _1075_;
wire _1076_;
wire _1077_;
wire _1078_;
wire _1079_;
wire _1080_;
wire _1081_;
wire _1082_;
wire _1083_;
wire _1084_;
wire _1085_;
wire _1086_;
wire _1087_;
wire _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire [2:0] _1122_;
wire [2:0] _1123_;
wire [2:0] _1124_;
wire [2:0] _1125_;
wire [2:0] _1126_;
wire [2:0] _1127_;
wire [2:0] _1128_;
wire [2:0] _1129_;
wire [2:0] _1130_;
wire [2:0] _1131_;
wire [2:0] _1132_;
wire [2:0] _1133_;
wire [2:0] _1134_;
wire [2:0] _1135_;
wire [2:0] _1136_;
wire [2:0] _1137_;
wire [2:0] _1138_;
wire [2:0] _1139_;
wire [2:0] _1140_;
wire [2:0] _1141_;
wire [2:0] _1142_;
wire [2:0] _1143_;
wire [2:0] _1144_;
wire [2:0] _1145_;
wire [2:0] _1146_;
wire [2:0] _1147_;
wire [2:0] _1148_;
wire [2:0] _1149_;
wire [2:0] _1150_;
wire [2:0] _1151_;
wire [2:0] _1152_;
wire [2:0] _1153_;
wire [2:0] _1154_;
wire [2:0] _1155_;
wire [2:0] _1156_;
wire [2:0] _1157_;
wire [2:0] _1158_;
wire [2:0] _1159_;
wire [2:0] _1160_;
wire [2:0] _1161_;
wire [2:0] _1162_;
wire [1:0] _1163_;
wire [1:0] _1164_;
wire _1165_;
wire _1166_;
wire _1167_;
wire _1168_;
wire _1169_;
wire _1170_;
wire _1171_;
wire _1172_;
wire _1173_;
wire _1174_;
wire _1175_;
wire _1176_;
wire _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire _1181_;
wire _1182_;
wire _1183_;
wire [1:0] _1184_;
wire [1:0] _1185_;
wire [1:0] _1186_;
wire [31:0] _1187_;
wire _1188_;
wire _1189_;
wire _1190_;
wire _1191_;
wire _1192_;
wire _1193_;
wire _1194_;
wire _1195_;
wire _1196_;
wire _1197_;
wire _1198_;
wire _1199_;
wire [31:0] _1200_;
wire _1201_;
wire _1202_;
wire _1203_;
wire _1204_;
wire _1205_;
wire _1206_;
wire _1207_;
wire _1208_;
wire _1209_;
wire [1:0] _1210_;
wire _1211_;
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire [31:0] _1216_;
wire [31:0] _1217_;
wire [31:0] _1218_;
wire _1219_;
wire _1220_;
wire [1:0] _1221_;
wire [1:0] _1222_;
wire _1223_;
wire _1224_;
wire _1225_;
wire _1226_;
wire [2:0] _1227_;
wire [2:0] _1228_;
wire [2:0] _1229_;
wire [2:0] _1230_;
wire [2:0] _1231_;
wire [2:0] _1232_;
wire [2:0] _1233_;
wire [2:0] _1234_;
wire [2:0] _1235_;
wire _1236_;
wire _1237_;
wire _1238_;
wire _1239_;
wire _1240_;
wire _1241_;
wire _1242_;
wire _1243_;
wire _1244_;
wire _1245_;
wire _1246_;
wire _1247_;
wire _1248_;
wire _1249_;
wire _1250_;
wire _1251_;
wire _1252_;
wire _1253_;
wire _1254_;
wire _1255_;
wire _1256_;
wire _1257_;
wire _1258_;
wire _1259_;
wire _1260_;
wire _1261_;
wire _1262_;
wire _1263_;
wire _1264_;
wire [1:0] _1265_;
wire [1:0] _1266_;
wire [1:0] _1267_;
wire _1268_;
wire _1269_;
wire [6:0] _1270_;
wire [6:0] _1271_;
wire [6:0] _1272_;
wire _1273_;
wire _1274_;
wire [31:0] _1275_;
wire [31:0] _1276_;
wire [31:0] _1277_;
wire _1278_;
wire _1279_;
wire _1280_;
wire _1281_;
wire _1282_;
wire [1:0] _1283_;
wire [1:0] _1284_;
wire [1:0] _1285_;
wire _1286_;
wire _1287_;
wire _1288_;
wire _1289_;
wire _1290_;
wire [31:0] _1291_;
wire [31:0] _1292_;
wire [31:0] _1293_;
wire _1294_;
wire _1295_;
wire _1296_;
wire _1297_;
wire [31:0] _1298_;
wire [31:0] _1299_;
wire [31:0] _1300_;
wire _1301_;
wire _1302_;
wire [2:0] _1303_;
wire [2:0] _1304_;
wire [2:0] _1305_;
wire [1:0] _1306_;
wire [1:0] _1307_;
wire [1:0] _1308_;
wire _1309_;
wire _1310_;
wire _1311_;
wire [1:0] _1312_;
wire [1:0] _1313_;
wire [1:0] _1314_;
wire _1315_;
wire _1316_;
wire _1317_;
wire _1318_;
wire _1319_;
wire [31:0] _1320_;
wire [31:0] _1321_;
wire [31:0] _1322_;
wire _1323_;
wire _1324_;
wire _1325_;
wire [6:0] _1326_;
wire [6:0] _1327_;
wire [6:0] _1328_;
wire _1329_;
wire _1330_;
wire _1331_;
wire [31:0] _1332_;
wire [31:0] _1333_;
wire [31:0] _1334_;
wire _1335_;
wire _1336_;
wire _1337_;
wire [3:0] _1338_;
wire [3:0] _1339_;
wire [3:0] _1340_;
wire _1341_;
wire _1342_;
wire [31:0] _1343_;
wire [31:0] _1344_;
wire [31:0] _1345_;
wire [31:0] _1346_;
wire [31:0] _1347_;
wire [31:0] _1348_;
wire [31:0] _1349_;
wire [31:0] _1350_;
wire [31:0] _1351_;
wire _1352_;
wire _1353_;
wire _1354_;
wire _1355_;
wire _1356_;
wire _1357_;
wire _1358_;
wire _1359_;
wire _1360_;
wire _1361_;
wire _1362_;
wire _1363_;
wire _1364_;
wire _1365_;
wire _1366_;
wire _1367_;
wire _1368_;
wire _1369_;
wire _1370_;
wire _1371_;
wire _1372_;
wire [31:0] _1373_;
wire [31:0] _1374_;
wire [31:0] _1375_;
wire _1376_;
wire _1377_;
wire _1378_;
wire [2:0] _1379_;
wire [2:0] _1380_;
wire [2:0] _1381_;
wire [1:0] _1382_;
wire [1:0] _1383_;
wire [1:0] _1384_;
wire _1385_;
wire _1386_;
wire _1387_;
wire [31:0] _1388_;
wire [31:0] _1389_;
wire [31:0] _1390_;
wire _1391_;
wire _1392_;
wire _1393_;
wire _1394_;
wire _1395_;
wire _1396_;
wire _1397_;
wire _1398_;
wire _1399_;
wire [6:0] _1400_;
wire [6:0] _1401_;
wire [6:0] _1402_;
wire [6:0] _1403_;
wire [6:0] _1404_;
wire [6:0] _1405_;
wire [6:0] _1406_;
wire [6:0] _1407_;
wire [6:0] _1408_;
wire _1409_;
wire _1410_;
wire _1411_;
wire _1412_;
wire _1413_;
wire _1414_;
wire _1415_;
wire _1416_;
wire _1417_;
wire [31:0] _1418_;
wire [31:0] _1419_;
wire [31:0] _1420_;
wire [31:0] _1421_;
wire [31:0] _1422_;
wire [31:0] _1423_;
wire [31:0] _1424_;
wire [31:0] _1425_;
wire [31:0] _1426_;
wire _1427_;
wire _1428_;
wire _1429_;
wire _1430_;
wire _1431_;
wire _1432_;
wire _1433_;
wire _1434_;
wire [6:0] _1435_;
wire [6:0] _1436_;
wire [6:0] _1437_;
wire _1438_;
wire _1439_;
wire [1:0] _1440_;
wire [1:0] _1441_;
wire [1:0] _1442_;
wire [1:0] _1443_;
wire [1:0] _1444_;
wire _1445_;
wire _1446_;
wire [3:0] _1447_;
wire [3:0] _1448_;
wire [1:0] _1449_;
wire [1:0] _1450_;
wire [1:0] _1451_;
wire [1:0] _1452_;
wire [1:0] _1453_;
wire [1:0] _1454_;
wire _1455_;
wire _1456_;
wire _1457_;
wire _1458_;
wire _1459_;
wire [11:0] _1460_;
wire [11:0] _1461_;
wire [1:0] _1462_;
wire [1:0] _1463_;
wire [1:0] _1464_;
wire [1:0] _1465_;
wire [1:0] _1466_;
wire [1:0] _1467_;
wire _1468_;
wire _1469_;
wire _1470_;
wire _1471_;
wire _1472_;
wire _1473_;
wire _1474_;
wire _1475_;
wire _1476_;
wire [1:0] _1477_;
wire [1:0] _1478_;
wire [1:0] _1479_;
wire _1480_;
wire _1481_;
wire [1:0] _1482_;
wire [1:0] _1483_;
wire _1484_;
wire _1485_;
wire [1:0] _1486_;
wire [1:0] _1487_;
wire [30:0] _1488_;
wire [7:0] _1489_;
wire [7:0] _1490_;
wire [7:0] _1491_;
wire [31:0] _1492_;
wire [31:0] _1493_;
wire [31:0] _1494_;
wire [31:0] _1495_;
wire _1496_;
wire _1497_;
wire _1498_;
wire _1499_;
wire _1500_;
wire _1501_;
wire [7:0] _1502_;
wire [7:0] _1503_;
wire [7:0] _1504_;
wire [31:0] _1505_;
wire [31:0] _1506_;
wire [31:0] _1507_;
wire [31:0] _1508_;
wire _1509_;
wire _1510_;
wire _1511_;
wire _1512_;
wire _1513_;
wire _1514_;
wire _1515_;
wire _1516_;
wire _1517_;
wire _1518_;
wire [31:0] _1519_;
wire [31:0] _1520_;
wire [31:0] _1521_;
wire _1522_;
wire _1523_;
wire _1524_;
wire _1525_;
wire _1526_;
wire _1527_;
wire _1528_;
wire _1529_;
wire _1530_;
wire _1531_;
wire _1532_;
wire _1533_;
wire _1534_;
wire _1535_;
wire _1536_;
wire [5:0] _1537_;
wire [5:0] _1538_;
wire [5:0] _1539_;
wire _1540_;
wire _1541_;
wire [30:0] _1542_;
wire [11:0] _1543_;
wire [28:0] _1544_;
wire [4:0] _1545_;
wire [19:0] _1546_;
wire [2:0] _1547_;
wire [17:0] _1548_;
wire [31:0] _1549_;
wire [31:0] _1550_;
wire [31:0] _1551_;
wire [1:0] _1552_;
wire [1:0] _1553_;
wire [1:0] _1554_;
wire [63:0] _1555_;
wire [63:0] _1556_;
wire [63:0] _1557_;
wire _1558_;
/* cellift = 32'd1 */
wire _1559_;
wire _1560_;
/* cellift = 32'd1 */
wire _1561_;
wire _1562_;
/* cellift = 32'd1 */
wire _1563_;
wire _1564_;
/* cellift = 32'd1 */
wire _1565_;
wire _1566_;
/* cellift = 32'd1 */
wire _1567_;
wire _1568_;
/* cellift = 32'd1 */
wire _1569_;
wire _1570_;
/* cellift = 32'd1 */
wire _1571_;
wire _1572_;
/* cellift = 32'd1 */
wire _1573_;
wire _1574_;
/* cellift = 32'd1 */
wire _1575_;
wire _1576_;
/* cellift = 32'd1 */
wire _1577_;
wire _1578_;
/* cellift = 32'd1 */
wire _1579_;
wire _1580_;
wire _1581_;
wire [31:0] _1582_;
wire _1583_;
wire _1584_;
wire [17:0] _1585_;
wire _1586_;
wire _1587_;
wire _1588_;
wire [1:0] _1589_;
wire [1:0] _1590_;
wire [1:0] _1591_;
wire [1:0] _1592_;
wire [1:0] _1593_;
wire [1:0] _1594_;
wire [1:0] _1595_;
wire [1:0] _1596_;
wire _1597_;
wire _1598_;
wire _1599_;
wire _1600_;
wire _1601_;
wire _1602_;
wire _1603_;
wire _1604_;
wire _1605_;
wire _1606_;
wire _1607_;
wire _1608_;
wire _1609_;
wire _1610_;
wire _1611_;
wire _1612_;
wire _1613_;
wire _1614_;
wire _1615_;
wire _1616_;
wire _1617_;
wire _1618_;
wire _1619_;
wire _1620_;
wire _1621_;
wire _1622_;
wire _1623_;
wire _1624_;
wire _1625_;
wire _1626_;
wire _1627_;
wire _1628_;
wire _1629_;
wire _1630_;
wire _1631_;
wire _1632_;
wire _1633_;
wire _1634_;
wire _1635_;
wire _1636_;
wire _1637_;
wire _1638_;
wire _1639_;
wire _1640_;
wire _1641_;
wire _1642_;
wire _1643_;
wire _1644_;
wire _1645_;
wire _1646_;
wire _1647_;
wire _1648_;
wire _1649_;
wire _1650_;
wire _1651_;
wire _1652_;
wire _1653_;
wire _1654_;
wire _1655_;
wire [2:0] _1656_;
wire [2:0] _1657_;
wire [2:0] _1658_;
wire [2:0] _1659_;
wire [2:0] _1660_;
wire [2:0] _1661_;
wire [2:0] _1662_;
wire [2:0] _1663_;
wire [2:0] _1664_;
wire [2:0] _1665_;
wire [2:0] _1666_;
wire [2:0] _1667_;
wire [2:0] _1668_;
wire [2:0] _1669_;
wire [2:0] _1670_;
wire [2:0] _1671_;
wire [2:0] _1672_;
wire [2:0] _1673_;
wire [2:0] _1674_;
wire [2:0] _1675_;
wire [2:0] _1676_;
wire [2:0] _1677_;
wire [2:0] _1678_;
wire [2:0] _1679_;
wire [2:0] _1680_;
wire [2:0] _1681_;
wire [2:0] _1682_;
wire [2:0] _1683_;
wire [2:0] _1684_;
wire [2:0] _1685_;
wire [2:0] _1686_;
wire [2:0] _1687_;
wire [2:0] _1688_;
wire [2:0] _1689_;
wire [2:0] _1690_;
wire [2:0] _1691_;
wire [2:0] _1692_;
wire [2:0] _1693_;
wire [2:0] _1694_;
wire [2:0] _1695_;
wire [2:0] _1696_;
wire [2:0] _1697_;
wire [2:0] _1698_;
wire [2:0] _1699_;
wire [2:0] _1700_;
wire [2:0] _1701_;
wire [2:0] _1702_;
wire [2:0] _1703_;
wire [2:0] _1704_;
wire [2:0] _1705_;
wire [2:0] _1706_;
wire [2:0] _1707_;
wire [2:0] _1708_;
wire [2:0] _1709_;
wire [2:0] _1710_;
wire [2:0] _1711_;
wire [2:0] _1712_;
wire [2:0] _1713_;
wire [2:0] _1714_;
wire [2:0] _1715_;
wire [2:0] _1716_;
wire [2:0] _1717_;
wire [2:0] _1718_;
wire [2:0] _1719_;
wire [2:0] _1720_;
wire [2:0] _1721_;
wire [2:0] _1722_;
wire [2:0] _1723_;
wire [2:0] _1724_;
wire [2:0] _1725_;
wire [2:0] _1726_;
wire [2:0] _1727_;
wire [2:0] _1728_;
wire [2:0] _1729_;
wire [2:0] _1730_;
wire [2:0] _1731_;
wire [2:0] _1732_;
wire [2:0] _1733_;
wire [2:0] _1734_;
wire [2:0] _1735_;
wire [2:0] _1736_;
wire [2:0] _1737_;
wire [2:0] _1738_;
wire [2:0] _1739_;
wire [2:0] _1740_;
wire [2:0] _1741_;
wire [2:0] _1742_;
wire [2:0] _1743_;
wire [2:0] _1744_;
wire [2:0] _1745_;
wire [2:0] _1746_;
wire [2:0] _1747_;
wire [2:0] _1748_;
wire _1749_;
wire _1750_;
wire _1751_;
wire _1752_;
wire _1753_;
wire _1754_;
wire _1755_;
wire _1756_;
wire _1757_;
wire _1758_;
wire _1759_;
wire _1760_;
wire _1761_;
wire _1762_;
wire _1763_;
wire _1764_;
wire _1765_;
wire _1766_;
wire _1767_;
wire _1768_;
wire _1769_;
wire _1770_;
wire _1771_;
wire _1772_;
wire _1773_;
wire _1774_;
wire _1775_;
wire _1776_;
wire _1777_;
wire _1778_;
wire _1779_;
wire _1780_;
wire _1781_;
wire _1782_;
wire _1783_;
wire _1784_;
wire _1785_;
wire _1786_;
wire _1787_;
wire _1788_;
wire _1789_;
wire _1790_;
wire _1791_;
wire _1792_;
wire _1793_;
wire _1794_;
wire _1795_;
wire _1796_;
wire _1797_;
wire _1798_;
wire _1799_;
wire _1800_;
wire [2:0] _1801_;
wire [2:0] _1802_;
wire [2:0] _1803_;
wire [2:0] _1804_;
wire [2:0] _1805_;
wire [2:0] _1806_;
wire [2:0] _1807_;
wire [2:0] _1808_;
wire [2:0] _1809_;
wire [2:0] _1810_;
wire [2:0] _1811_;
wire [2:0] _1812_;
wire [2:0] _1813_;
wire [2:0] _1814_;
wire [2:0] _1815_;
wire [2:0] _1816_;
wire [2:0] _1817_;
wire [2:0] _1818_;
wire [2:0] _1819_;
wire _1820_;
wire _1821_;
wire _1822_;
wire _1823_;
wire _1824_;
wire _1825_;
wire _1826_;
wire _1827_;
wire _1828_;
wire _1829_;
wire _1830_;
wire _1831_;
wire _1832_;
wire [8:0] _1833_;
wire [8:0] _1834_;
wire [8:0] _1835_;
wire [8:0] _1836_;
wire [8:0] _1837_;
wire [8:0] _1838_;
wire [8:0] _1839_;
wire [8:0] _1840_;
wire [8:0] _1841_;
wire [8:0] _1842_;
wire [8:0] _1843_;
wire [8:0] _1844_;
wire [8:0] _1845_;
wire [8:0] _1846_;
wire [8:0] _1847_;
wire [8:0] _1848_;
wire [8:0] _1849_;
wire [8:0] _1850_;
wire [8:0] _1851_;
wire [8:0] _1852_;
wire [8:0] _1853_;
wire [8:0] _1854_;
wire [8:0] _1855_;
wire [8:0] _1856_;
wire [8:0] _1857_;
wire [8:0] _1858_;
wire [8:0] _1859_;
wire [8:0] _1860_;
wire [8:0] _1861_;
wire [8:0] _1862_;
wire [8:0] _1863_;
wire [8:0] _1864_;
wire [8:0] _1865_;
wire [8:0] _1866_;
wire [8:0] _1867_;
wire [8:0] _1868_;
wire [8:0] _1869_;
wire [8:0] _1870_;
wire [8:0] _1871_;
wire [8:0] _1872_;
wire [8:0] _1873_;
wire [8:0] _1874_;
wire _1875_;
wire _1876_;
wire _1877_;
wire _1878_;
wire _1879_;
wire _1880_;
wire _1881_;
wire _1882_;
wire _1883_;
wire _1884_;
wire _1885_;
wire _1886_;
wire _1887_;
wire _1888_;
wire [63:0] _1889_;
wire [63:0] _1890_;
wire [63:0] _1891_;
wire [63:0] _1892_;
wire _1893_;
wire _1894_;
wire _1895_;
wire _1896_;
wire _1897_;
wire _1898_;
wire _1899_;
wire _1900_;
wire _1901_;
wire _1902_;
wire _1903_;
wire _1904_;
wire _1905_;
wire _1906_;
wire [31:0] _1907_;
wire [31:0] _1908_;
wire [31:0] _1909_;
wire [31:0] _1910_;
wire [31:0] _1911_;
wire [31:0] _1912_;
wire _1913_;
wire _1914_;
wire _1915_;
wire _1916_;
wire _1917_;
wire _1918_;
wire _1919_;
wire _1920_;
wire _1921_;
wire _1922_;
wire _1923_;
wire _1924_;
wire _1925_;
wire _1926_;
wire _1927_;
wire _1928_;
wire _1929_;
wire _1930_;
wire _1931_;
wire _1932_;
wire _1933_;
wire _1934_;
wire _1935_;
wire _1936_;
wire _1937_;
wire _1938_;
wire _1939_;
wire _1940_;
wire _1941_;
wire _1942_;
wire _1943_;
wire _1944_;
wire _1945_;
wire _1946_;
wire [2:0] _1947_;
wire [2:0] _1948_;
wire [2:0] _1949_;
wire [2:0] _1950_;
wire [2:0] _1951_;
wire [2:0] _1952_;
wire [2:0] _1953_;
wire [2:0] _1954_;
wire [2:0] _1955_;
wire [2:0] _1956_;
wire [2:0] _1957_;
wire [2:0] _1958_;
wire [2:0] _1959_;
wire [2:0] _1960_;
wire [2:0] _1961_;
wire [2:0] _1962_;
wire [2:0] _1963_;
wire _1964_;
wire _1965_;
wire _1966_;
wire _1967_;
wire _1968_;
wire _1969_;
wire _1970_;
wire _1971_;
wire _1972_;
wire [31:0] _1973_;
wire _1974_;
wire _1975_;
wire _1976_;
wire _1977_;
wire [31:0] _1978_;
wire _1979_;
wire _1980_;
wire _1981_;
wire _1982_;
wire _1983_;
wire _1984_;
wire _1985_;
wire _1986_;
wire [31:0] _1987_;
wire [31:0] _1988_;
wire [31:0] _1989_;
wire [1:0] _1990_;
wire _1991_;
wire [2:0] _1992_;
wire [2:0] _1993_;
wire [2:0] _1994_;
wire [2:0] _1995_;
wire [2:0] _1996_;
wire [2:0] _1997_;
wire [2:0] _1998_;
wire [2:0] _1999_;
wire [2:0] _2000_;
wire _2001_;
wire _2002_;
wire _2003_;
wire _2004_;
wire _2005_;
wire _2006_;
wire _2007_;
wire _2008_;
wire _2009_;
wire _2010_;
wire _2011_;
wire _2012_;
wire _2013_;
wire _2014_;
wire _2015_;
wire _2016_;
wire [1:0] _2017_;
wire [1:0] _2018_;
wire [1:0] _2019_;
wire [6:0] _2020_;
wire [6:0] _2021_;
wire [6:0] _2022_;
wire [31:0] _2023_;
wire [31:0] _2024_;
wire [31:0] _2025_;
wire _2026_;
wire [1:0] _2027_;
wire _2028_;
wire [31:0] _2029_;
wire _2030_;
wire _2031_;
wire [31:0] _2032_;
wire [31:0] _2033_;
wire [31:0] _2034_;
wire [2:0] _2035_;
wire [2:0] _2036_;
wire [2:0] _2037_;
wire [1:0] _2038_;
wire [1:0] _2039_;
wire [1:0] _2040_;
wire _2041_;
wire [1:0] _2042_;
wire _2043_;
wire [31:0] _2044_;
wire _2045_;
wire [6:0] _2046_;
wire [6:0] _2047_;
wire [6:0] _2048_;
wire _2049_;
wire [31:0] _2050_;
wire _2051_;
wire [3:0] _2052_;
wire [3:0] _2053_;
wire [3:0] _2054_;
wire [31:0] _2055_;
wire [31:0] _2056_;
wire [31:0] _2057_;
wire [31:0] _2058_;
wire [31:0] _2059_;
wire [31:0] _2060_;
wire [31:0] _2061_;
wire [31:0] _2062_;
wire [31:0] _2063_;
wire _2064_;
wire _2065_;
wire _2066_;
wire _2067_;
wire _2068_;
wire [31:0] _2069_;
wire [31:0] _2070_;
wire [31:0] _2071_;
wire _2072_;
wire [2:0] _2073_;
wire [1:0] _2074_;
wire [1:0] _2075_;
wire [1:0] _2076_;
wire _2077_;
wire [31:0] _2078_;
wire _2079_;
wire _2080_;
wire _2081_;
wire [6:0] _2082_;
wire [6:0] _2083_;
wire [6:0] _2084_;
wire [6:0] _2085_;
wire [6:0] _2086_;
wire [6:0] _2087_;
wire [6:0] _2088_;
wire [6:0] _2089_;
wire [6:0] _2090_;
wire _2091_;
wire _2092_;
wire _2093_;
wire [31:0] _2094_;
wire [31:0] _2095_;
wire [31:0] _2096_;
wire [31:0] _2097_;
wire [31:0] _2098_;
wire [31:0] _2099_;
wire [31:0] _2100_;
wire _2101_;
wire _2102_;
wire [6:0] _2103_;
wire [6:0] _2104_;
wire [6:0] _2105_;
wire [1:0] _2106_;
wire [1:0] _2107_;
wire [1:0] _2108_;
wire [1:0] _2109_;
wire [3:0] _2110_;
wire [1:0] _2111_;
wire [1:0] _2112_;
wire [1:0] _2113_;
wire [1:0] _2114_;
wire _2115_;
wire [11:0] _2116_;
wire [1:0] _2117_;
wire [1:0] _2118_;
wire [1:0] _2119_;
wire [1:0] _2120_;
wire _2121_;
wire [1:0] _2122_;
wire [1:0] _2123_;
wire [1:0] _2124_;
wire [7:0] _2125_;
wire [7:0] _2126_;
wire [7:0] _2127_;
wire [31:0] _2128_;
wire [31:0] _2129_;
wire _2130_;
wire _2131_;
wire [7:0] _2132_;
wire [7:0] _2133_;
wire [7:0] _2134_;
wire [31:0] _2135_;
wire [31:0] _2136_;
wire [31:0] _2137_;
wire _2138_;
wire [5:0] _2139_;
wire [5:0] _2140_;
wire [5:0] _2141_;
wire _2142_;
wire [31:0] _2143_;
wire [31:0] _2144_;
wire [31:0] _2145_;
wire [1:0] _2146_;
wire [1:0] _2147_;
wire [1:0] _2148_;
wire [63:0] _2149_;
wire [63:0] _2150_;
wire [63:0] _2151_;
wire _2152_;
/* cellift = 32'd1 */
wire _2153_;
wire [1:0] _2154_;
wire [1:0] _2155_;
wire _2156_;
wire _2157_;
wire _2158_;
wire _2159_;
wire _2160_;
wire _2161_;
wire _2162_;
wire _2163_;
wire _2164_;
wire _2165_;
wire _2166_;
wire _2167_;
wire _2168_;
wire _2169_;
wire _2170_;
wire _2171_;
wire [2:0] _2172_;
wire [2:0] _2173_;
wire [2:0] _2174_;
wire [2:0] _2175_;
wire [2:0] _2176_;
wire [2:0] _2177_;
wire [2:0] _2178_;
wire [2:0] _2179_;
wire [2:0] _2180_;
wire [2:0] _2181_;
wire [2:0] _2182_;
wire [2:0] _2183_;
wire [2:0] _2184_;
wire [2:0] _2185_;
wire [2:0] _2186_;
wire [2:0] _2187_;
wire [2:0] _2188_;
wire [2:0] _2189_;
wire [2:0] _2190_;
wire [2:0] _2191_;
wire [2:0] _2192_;
wire [2:0] _2193_;
wire [2:0] _2194_;
wire [2:0] _2195_;
wire [2:0] _2196_;
wire [2:0] _2197_;
wire [2:0] _2198_;
wire [2:0] _2199_;
wire [2:0] _2200_;
wire [2:0] _2201_;
wire [2:0] _2202_;
wire [2:0] _2203_;
wire [2:0] _2204_;
wire [2:0] _2205_;
wire [2:0] _2206_;
wire [2:0] _2207_;
wire [2:0] _2208_;
wire [2:0] _2209_;
wire [2:0] _2210_;
wire [2:0] _2211_;
wire [2:0] _2212_;
wire [2:0] _2213_;
wire _2214_;
wire _2215_;
wire _2216_;
wire _2217_;
wire _2218_;
wire _2219_;
wire _2220_;
wire _2221_;
wire _2222_;
wire _2223_;
wire _2224_;
wire _2225_;
wire _2226_;
wire _2227_;
wire _2228_;
wire _2229_;
wire _2230_;
wire _2231_;
wire _2232_;
wire _2233_;
wire _2234_;
wire _2235_;
wire _2236_;
wire _2237_;
wire _2238_;
wire _2239_;
wire _2240_;
wire _2241_;
wire [2:0] _2242_;
wire [2:0] _2243_;
wire [2:0] _2244_;
wire [2:0] _2245_;
wire [2:0] _2246_;
wire [2:0] _2247_;
wire [2:0] _2248_;
wire [2:0] _2249_;
wire [2:0] _2250_;
wire [2:0] _2251_;
wire [2:0] _2252_;
wire [2:0] _2253_;
wire _2254_;
wire _2255_;
wire _2256_;
wire _2257_;
wire _2258_;
wire _2259_;
wire _2260_;
wire _2261_;
wire _2262_;
wire _2263_;
wire _2264_;
wire _2265_;
wire _2266_;
wire _2267_;
wire [8:0] _2268_;
wire [8:0] _2269_;
wire [8:0] _2270_;
wire [8:0] _2271_;
wire [8:0] _2272_;
wire [8:0] _2273_;
wire [8:0] _2274_;
wire [8:0] _2275_;
wire [8:0] _2276_;
wire [8:0] _2277_;
wire [8:0] _2278_;
wire [8:0] _2279_;
wire [8:0] _2280_;
wire [8:0] _2281_;
wire [8:0] _2282_;
wire _2283_;
wire _2284_;
wire _2285_;
wire _2286_;
wire _2287_;
wire _2288_;
wire _2289_;
wire _2290_;
wire _2291_;
wire _2292_;
wire _2293_;
wire _2294_;
wire _2295_;
wire _2296_;
wire _2297_;
wire [63:0] _2298_;
wire [63:0] _2299_;
wire _2300_;
wire _2301_;
wire _2302_;
wire _2303_;
wire _2304_;
wire _2305_;
wire _2306_;
wire _2307_;
wire _2308_;
wire _2309_;
wire _2310_;
wire _2311_;
wire _2312_;
wire _2313_;
wire _2314_;
wire [31:0] _2315_;
wire [31:0] _2316_;
wire _2317_;
wire _2318_;
wire _2319_;
wire _2320_;
wire _2321_;
wire _2322_;
wire _2323_;
wire _2324_;
wire _2325_;
wire _2326_;
wire _2327_;
wire _2328_;
wire _2329_;
wire _2330_;
wire _2331_;
wire _2332_;
wire _2333_;
wire _2334_;
wire _2335_;
wire _2336_;
wire _2337_;
wire _2338_;
wire _2339_;
wire _2340_;
wire _2341_;
wire _2342_;
wire _2343_;
wire _2344_;
wire [2:0] _2345_;
wire [2:0] _2346_;
wire [2:0] _2347_;
wire [2:0] _2348_;
wire [2:0] _2349_;
wire [2:0] _2350_;
wire [2:0] _2351_;
wire [2:0] _2352_;
wire [2:0] _2353_;
wire [2:0] _2354_;
wire [2:0] _2355_;
wire [2:0] _2356_;
wire [2:0] _2357_;
wire [2:0] _2358_;
wire [31:0] _2359_;
wire _2360_;
wire [31:0] _2361_;
wire [2:0] _2362_;
wire [2:0] _2363_;
wire [2:0] _2364_;
wire _2365_;
wire _2366_;
wire _2367_;
wire _2368_;
wire _2369_;
wire _2370_;
wire _2371_;
wire [1:0] _2372_;
wire [6:0] _2373_;
wire [31:0] _2374_;
wire _2375_;
wire [1:0] _2376_;
wire _2377_;
wire [31:0] _2378_;
wire [2:0] _2379_;
wire [1:0] _2380_;
wire _2381_;
wire [1:0] _2382_;
wire _2383_;
wire [31:0] _2384_;
wire _2385_;
wire [6:0] _2386_;
wire _2387_;
wire [31:0] _2388_;
wire _2389_;
wire [3:0] _2390_;
wire [31:0] _2391_;
wire [31:0] _2392_;
wire [31:0] _2393_;
wire _2394_;
wire _2395_;
wire _2396_;
wire _2397_;
wire _2398_;
wire [31:0] _2399_;
wire _2400_;
wire [2:0] _2401_;
wire [1:0] _2402_;
wire _2403_;
wire [31:0] _2404_;
wire _2405_;
wire _2406_;
wire _2407_;
wire [6:0] _2408_;
wire [6:0] _2409_;
wire [6:0] _2410_;
wire _2411_;
wire _2412_;
wire _2413_;
wire [31:0] _2414_;
wire [31:0] _2415_;
wire [31:0] _2416_;
wire _2417_;
wire _2418_;
wire [6:0] _2419_;
wire [1:0] _2420_;
wire [1:0] _2421_;
wire [1:0] _2422_;
wire _2423_;
wire [1:0] _2424_;
wire [1:0] _2425_;
wire _2426_;
wire [1:0] _2427_;
wire [7:0] _2428_;
wire [31:0] _2429_;
wire [7:0] _2430_;
wire [31:0] _2431_;
wire _2432_;
wire [5:0] _2433_;
wire [31:0] _2434_;
wire [1:0] _2435_;
wire [63:0] _2436_;
wire _2437_;
wire _2438_;
wire _2439_;
wire _2440_;
wire _2441_;
wire _2442_;
wire _2443_;
wire _2444_;
wire _2445_;
wire _2446_;
wire _2447_;
wire _2448_;
wire _2449_;
wire _2450_;
wire _2451_;
wire _2452_;
wire _2453_;
wire _2454_;
wire _2455_;
wire _2456_;
wire _2457_;
wire _2458_;
wire _2459_;
wire _2460_;
wire _2461_;
wire _2462_;
wire _2463_;
wire _2464_;
wire _2465_;
wire _2466_;
wire _2467_;
wire _2468_;
wire _2469_;
wire _2470_;
wire _2471_;
wire _2472_;
wire _2473_;
wire _2474_;
wire _2475_;
wire _2476_;
wire _2477_;
wire _2478_;
wire _2479_;
wire _2480_;
wire _2481_;
wire _2482_;
wire _2483_;
wire _2484_;
wire _2485_;
wire _2486_;
wire _2487_;
wire _2488_;
wire _2489_;
wire _2490_;
wire _2491_;
wire _2492_;
wire _2493_;
wire _2494_;
wire _2495_;
wire _2496_;
wire _2497_;
wire _2498_;
wire _2499_;
wire _2500_;
wire _2501_;
wire _2502_;
wire _2503_;
wire _2504_;
wire _2505_;
wire _2506_;
wire _2507_;
wire _2508_;
wire _2509_;
wire _2510_;
wire _2511_;
wire _2512_;
wire _2513_;
wire _2514_;
wire _2515_;
wire _2516_;
wire _2517_;
wire _2518_;
wire _2519_;
wire _2520_;
wire _2521_;
wire _2522_;
wire _2523_;
wire _2524_;
wire _2525_;
wire _2526_;
wire _2527_;
wire _2528_;
wire _2529_;
wire _2530_;
wire _2531_;
wire _2532_;
wire _2533_;
wire _2534_;
wire _2535_;
wire _2536_;
wire _2537_;
wire _2538_;
wire _2539_;
wire _2540_;
wire _2541_;
wire _2542_;
wire _2543_;
wire _2544_;
wire _2545_;
wire _2546_;
wire _2547_;
wire _2548_;
wire _2549_;
wire _2550_;
wire _2551_;
wire _2552_;
wire _2553_;
wire _2554_;
wire _2555_;
wire _2556_;
wire _2557_;
wire _2558_;
wire _2559_;
wire _2560_;
wire _2561_;
wire _2562_;
wire _2563_;
wire _2564_;
wire _2565_;
wire _2566_;
wire _2567_;
wire _2568_;
wire _2569_;
wire _2570_;
wire _2571_;
wire _2572_;
wire _2573_;
wire _2574_;
wire _2575_;
wire _2576_;
wire _2577_;
wire _2578_;
wire _2579_;
wire _2580_;
wire _2581_;
wire _2582_;
wire _2583_;
wire _2584_;
wire _2585_;
wire _2586_;
wire _2587_;
wire _2588_;
wire _2589_;
wire _2590_;
wire _2591_;
wire _2592_;
wire _2593_;
wire _2594_;
wire _2595_;
wire _2596_;
wire _2597_;
wire _2598_;
wire _2599_;
wire _2600_;
wire _2601_;
wire _2602_;
wire _2603_;
wire _2604_;
wire _2605_;
wire _2606_;
wire _2607_;
wire _2608_;
wire _2609_;
wire _2610_;
wire _2611_;
wire _2612_;
wire _2613_;
/* cellift = 32'd1 */
wire _2614_;
wire _2615_;
/* cellift = 32'd1 */
wire _2616_;
wire _2617_;
/* cellift = 32'd1 */
wire _2618_;
wire _2619_;
/* cellift = 32'd1 */
wire _2620_;
wire _2621_;
/* cellift = 32'd1 */
wire _2622_;
wire _2623_;
/* cellift = 32'd1 */
wire _2624_;
wire _2625_;
/* cellift = 32'd1 */
wire _2626_;
wire _2627_;
/* cellift = 32'd1 */
wire _2628_;
wire _2629_;
/* cellift = 32'd1 */
wire _2630_;
wire _2631_;
/* cellift = 32'd1 */
wire _2632_;
wire _2633_;
/* cellift = 32'd1 */
wire _2634_;
wire _2635_;
/* cellift = 32'd1 */
wire _2636_;
wire _2637_;
/* cellift = 32'd1 */
wire _2638_;
wire _2639_;
/* cellift = 32'd1 */
wire _2640_;
wire _2641_;
/* cellift = 32'd1 */
wire _2642_;
wire _2643_;
/* cellift = 32'd1 */
wire _2644_;
wire [2:0] _2645_;
/* cellift = 32'd1 */
wire [2:0] _2646_;
wire [2:0] _2647_;
/* cellift = 32'd1 */
wire [2:0] _2648_;
wire [2:0] _2649_;
/* cellift = 32'd1 */
wire [2:0] _2650_;
wire [2:0] _2651_;
/* cellift = 32'd1 */
wire [2:0] _2652_;
wire [2:0] _2653_;
/* cellift = 32'd1 */
wire [2:0] _2654_;
wire [2:0] _2655_;
/* cellift = 32'd1 */
wire [2:0] _2656_;
wire [2:0] _2657_;
/* cellift = 32'd1 */
wire [2:0] _2658_;
wire [2:0] _2659_;
/* cellift = 32'd1 */
wire [2:0] _2660_;
wire [2:0] _2661_;
/* cellift = 32'd1 */
wire [2:0] _2662_;
wire [2:0] _2663_;
/* cellift = 32'd1 */
wire [2:0] _2664_;
wire [2:0] _2665_;
/* cellift = 32'd1 */
wire [2:0] _2666_;
wire [2:0] _2667_;
/* cellift = 32'd1 */
wire [2:0] _2668_;
wire [2:0] _2669_;
/* cellift = 32'd1 */
wire [2:0] _2670_;
wire [2:0] _2671_;
/* cellift = 32'd1 */
wire [2:0] _2672_;
wire [2:0] _2673_;
/* cellift = 32'd1 */
wire [2:0] _2674_;
wire [2:0] _2675_;
/* cellift = 32'd1 */
wire [2:0] _2676_;
wire [2:0] _2677_;
/* cellift = 32'd1 */
wire [2:0] _2678_;
wire [2:0] _2679_;
/* cellift = 32'd1 */
wire [2:0] _2680_;
wire [2:0] _2681_;
/* cellift = 32'd1 */
wire [2:0] _2682_;
wire [2:0] _2683_;
/* cellift = 32'd1 */
wire [2:0] _2684_;
wire [2:0] _2685_;
/* cellift = 32'd1 */
wire [2:0] _2686_;
wire [2:0] _2687_;
/* cellift = 32'd1 */
wire [2:0] _2688_;
wire [2:0] _2689_;
/* cellift = 32'd1 */
wire [2:0] _2690_;
wire [2:0] _2691_;
/* cellift = 32'd1 */
wire [2:0] _2692_;
wire [2:0] _2693_;
/* cellift = 32'd1 */
wire [2:0] _2694_;
wire [2:0] _2695_;
/* cellift = 32'd1 */
wire [2:0] _2696_;
wire [2:0] _2697_;
/* cellift = 32'd1 */
wire [2:0] _2698_;
wire [2:0] _2699_;
/* cellift = 32'd1 */
wire [2:0] _2700_;
wire [2:0] _2701_;
/* cellift = 32'd1 */
wire [2:0] _2702_;
wire [2:0] _2703_;
/* cellift = 32'd1 */
wire [2:0] _2704_;
wire [2:0] _2705_;
/* cellift = 32'd1 */
wire [2:0] _2706_;
wire [2:0] _2707_;
/* cellift = 32'd1 */
wire [2:0] _2708_;
wire [2:0] _2709_;
/* cellift = 32'd1 */
wire [2:0] _2710_;
wire [2:0] _2711_;
/* cellift = 32'd1 */
wire [2:0] _2712_;
wire [2:0] _2713_;
/* cellift = 32'd1 */
wire [2:0] _2714_;
wire [2:0] _2715_;
/* cellift = 32'd1 */
wire [2:0] _2716_;
wire [2:0] _2717_;
/* cellift = 32'd1 */
wire [2:0] _2718_;
wire [2:0] _2719_;
/* cellift = 32'd1 */
wire [2:0] _2720_;
wire [2:0] _2721_;
/* cellift = 32'd1 */
wire [2:0] _2722_;
wire [2:0] _2723_;
/* cellift = 32'd1 */
wire [2:0] _2724_;
wire [2:0] _2725_;
/* cellift = 32'd1 */
wire [2:0] _2726_;
wire [2:0] _2727_;
/* cellift = 32'd1 */
wire [2:0] _2728_;
wire [2:0] _2729_;
/* cellift = 32'd1 */
wire [2:0] _2730_;
wire [2:0] _2731_;
/* cellift = 32'd1 */
wire [2:0] _2732_;
wire _2733_;
/* cellift = 32'd1 */
wire _2734_;
wire _2735_;
/* cellift = 32'd1 */
wire _2736_;
wire _2737_;
/* cellift = 32'd1 */
wire _2738_;
wire _2739_;
/* cellift = 32'd1 */
wire _2740_;
wire _2741_;
/* cellift = 32'd1 */
wire _2742_;
wire _2743_;
/* cellift = 32'd1 */
wire _2744_;
wire _2745_;
/* cellift = 32'd1 */
wire _2746_;
wire _2747_;
/* cellift = 32'd1 */
wire _2748_;
wire _2749_;
/* cellift = 32'd1 */
wire _2750_;
wire _2751_;
/* cellift = 32'd1 */
wire _2752_;
wire _2753_;
/* cellift = 32'd1 */
wire _2754_;
wire _2755_;
/* cellift = 32'd1 */
wire _2756_;
wire _2757_;
/* cellift = 32'd1 */
wire _2758_;
wire _2759_;
/* cellift = 32'd1 */
wire _2760_;
wire _2761_;
/* cellift = 32'd1 */
wire _2762_;
wire _2763_;
/* cellift = 32'd1 */
wire _2764_;
wire _2765_;
/* cellift = 32'd1 */
wire _2766_;
wire _2767_;
/* cellift = 32'd1 */
wire _2768_;
wire _2769_;
/* cellift = 32'd1 */
wire _2770_;
wire _2771_;
/* cellift = 32'd1 */
wire _2772_;
wire _2773_;
/* cellift = 32'd1 */
wire _2774_;
wire _2775_;
/* cellift = 32'd1 */
wire _2776_;
wire _2777_;
/* cellift = 32'd1 */
wire _2778_;
wire _2779_;
/* cellift = 32'd1 */
wire _2780_;
wire _2781_;
/* cellift = 32'd1 */
wire _2782_;
wire _2783_;
/* cellift = 32'd1 */
wire _2784_;
wire _2785_;
/* cellift = 32'd1 */
wire _2786_;
wire _2787_;
/* cellift = 32'd1 */
wire _2788_;
wire _2789_;
/* cellift = 32'd1 */
wire _2790_;
wire [2:0] _2791_;
/* cellift = 32'd1 */
wire [2:0] _2792_;
wire [2:0] _2793_;
/* cellift = 32'd1 */
wire [2:0] _2794_;
wire [2:0] _2795_;
/* cellift = 32'd1 */
wire [2:0] _2796_;
wire [2:0] _2797_;
/* cellift = 32'd1 */
wire [2:0] _2798_;
wire [2:0] _2799_;
/* cellift = 32'd1 */
wire [2:0] _2800_;
wire [2:0] _2801_;
/* cellift = 32'd1 */
wire [2:0] _2802_;
wire [2:0] _2803_;
/* cellift = 32'd1 */
wire [2:0] _2804_;
wire [2:0] _2805_;
/* cellift = 32'd1 */
wire [2:0] _2806_;
wire [2:0] _2807_;
/* cellift = 32'd1 */
wire [2:0] _2808_;
wire [2:0] _2809_;
/* cellift = 32'd1 */
wire [2:0] _2810_;
wire [2:0] _2811_;
/* cellift = 32'd1 */
wire [2:0] _2812_;
wire [2:0] _2813_;
/* cellift = 32'd1 */
wire [2:0] _2814_;
wire _2815_;
/* cellift = 32'd1 */
wire _2816_;
wire _2817_;
/* cellift = 32'd1 */
wire _2818_;
wire _2819_;
/* cellift = 32'd1 */
wire _2820_;
wire _2821_;
/* cellift = 32'd1 */
wire _2822_;
wire _2823_;
/* cellift = 32'd1 */
wire _2824_;
wire _2825_;
/* cellift = 32'd1 */
wire _2826_;
wire _2827_;
/* cellift = 32'd1 */
wire _2828_;
wire _2829_;
/* cellift = 32'd1 */
wire _2830_;
wire _2831_;
/* cellift = 32'd1 */
wire _2832_;
wire _2833_;
/* cellift = 32'd1 */
wire _2834_;
wire _2835_;
/* cellift = 32'd1 */
wire _2836_;
wire _2837_;
/* cellift = 32'd1 */
wire _2838_;
wire _2839_;
/* cellift = 32'd1 */
wire _2840_;
wire _2841_;
/* cellift = 32'd1 */
wire _2842_;
wire [8:0] _2843_;
/* cellift = 32'd1 */
wire [8:0] _2844_;
wire [8:0] _2845_;
/* cellift = 32'd1 */
wire [8:0] _2846_;
wire [8:0] _2847_;
/* cellift = 32'd1 */
wire [8:0] _2848_;
wire [8:0] _2849_;
/* cellift = 32'd1 */
wire [8:0] _2850_;
wire [8:0] _2851_;
/* cellift = 32'd1 */
wire [8:0] _2852_;
wire [8:0] _2853_;
/* cellift = 32'd1 */
wire [8:0] _2854_;
wire [8:0] _2855_;
/* cellift = 32'd1 */
wire [8:0] _2856_;
wire [8:0] _2857_;
/* cellift = 32'd1 */
wire [8:0] _2858_;
wire [8:0] _2859_;
/* cellift = 32'd1 */
wire [8:0] _2860_;
wire [8:0] _2861_;
/* cellift = 32'd1 */
wire [8:0] _2862_;
wire [8:0] _2863_;
/* cellift = 32'd1 */
wire [8:0] _2864_;
wire [8:0] _2865_;
/* cellift = 32'd1 */
wire [8:0] _2866_;
wire [8:0] _2867_;
/* cellift = 32'd1 */
wire [8:0] _2868_;
wire [8:0] _2869_;
/* cellift = 32'd1 */
wire [8:0] _2870_;
wire [8:0] _2871_;
/* cellift = 32'd1 */
wire [8:0] _2872_;
wire _2873_;
/* cellift = 32'd1 */
wire _2874_;
wire _2875_;
/* cellift = 32'd1 */
wire _2876_;
wire _2877_;
/* cellift = 32'd1 */
wire _2878_;
wire _2879_;
/* cellift = 32'd1 */
wire _2880_;
wire _2881_;
/* cellift = 32'd1 */
wire _2882_;
wire _2883_;
/* cellift = 32'd1 */
wire _2884_;
wire _2885_;
/* cellift = 32'd1 */
wire _2886_;
wire _2887_;
/* cellift = 32'd1 */
wire _2888_;
wire _2889_;
/* cellift = 32'd1 */
wire _2890_;
wire _2891_;
/* cellift = 32'd1 */
wire _2892_;
wire _2893_;
/* cellift = 32'd1 */
wire _2894_;
wire _2895_;
/* cellift = 32'd1 */
wire _2896_;
wire _2897_;
/* cellift = 32'd1 */
wire _2898_;
wire _2899_;
/* cellift = 32'd1 */
wire _2900_;
wire _2901_;
/* cellift = 32'd1 */
wire _2902_;
/* cellift = 32'd1 */
wire [63:0] _2903_;
wire _2904_;
/* cellift = 32'd1 */
wire _2905_;
wire _2906_;
/* cellift = 32'd1 */
wire _2907_;
wire _2908_;
/* cellift = 32'd1 */
wire _2909_;
wire _2910_;
/* cellift = 32'd1 */
wire _2911_;
wire _2912_;
/* cellift = 32'd1 */
wire _2913_;
wire _2914_;
/* cellift = 32'd1 */
wire _2915_;
wire _2916_;
/* cellift = 32'd1 */
wire _2917_;
wire _2918_;
/* cellift = 32'd1 */
wire _2919_;
wire _2920_;
/* cellift = 32'd1 */
wire _2921_;
wire _2922_;
/* cellift = 32'd1 */
wire _2923_;
wire _2924_;
/* cellift = 32'd1 */
wire _2925_;
wire _2926_;
/* cellift = 32'd1 */
wire _2927_;
wire _2928_;
/* cellift = 32'd1 */
wire _2929_;
wire _2930_;
/* cellift = 32'd1 */
wire _2931_;
wire _2932_;
/* cellift = 32'd1 */
wire _2933_;
wire [31:0] _2934_;
/* cellift = 32'd1 */
wire [31:0] _2935_;
wire _2936_;
/* cellift = 32'd1 */
wire _2937_;
wire _2938_;
/* cellift = 32'd1 */
wire _2939_;
wire _2940_;
/* cellift = 32'd1 */
wire _2941_;
wire _2942_;
/* cellift = 32'd1 */
wire _2943_;
wire _2944_;
/* cellift = 32'd1 */
wire _2945_;
wire _2946_;
/* cellift = 32'd1 */
wire _2947_;
wire _2948_;
/* cellift = 32'd1 */
wire _2949_;
wire _2950_;
/* cellift = 32'd1 */
wire _2951_;
wire _2952_;
/* cellift = 32'd1 */
wire _2953_;
wire _2954_;
/* cellift = 32'd1 */
wire _2955_;
wire _2956_;
/* cellift = 32'd1 */
wire _2957_;
wire _2958_;
/* cellift = 32'd1 */
wire _2959_;
wire _2960_;
/* cellift = 32'd1 */
wire _2961_;
wire _2962_;
/* cellift = 32'd1 */
wire _2963_;
wire _2964_;
/* cellift = 32'd1 */
wire _2965_;
wire _2966_;
/* cellift = 32'd1 */
wire _2967_;
wire _2968_;
/* cellift = 32'd1 */
wire _2969_;
wire _2970_;
/* cellift = 32'd1 */
wire _2971_;
wire _2972_;
/* cellift = 32'd1 */
wire _2973_;
wire _2974_;
/* cellift = 32'd1 */
wire _2975_;
wire _2976_;
/* cellift = 32'd1 */
wire _2977_;
wire _2978_;
/* cellift = 32'd1 */
wire _2979_;
wire _2980_;
/* cellift = 32'd1 */
wire _2981_;
wire _2982_;
/* cellift = 32'd1 */
wire _2983_;
wire _2984_;
/* cellift = 32'd1 */
wire _2985_;
wire _2986_;
/* cellift = 32'd1 */
wire _2987_;
wire _2988_;
/* cellift = 32'd1 */
wire _2989_;
wire _2990_;
/* cellift = 32'd1 */
wire _2991_;
wire [2:0] _2992_;
/* cellift = 32'd1 */
wire [2:0] _2993_;
wire [2:0] _2994_;
/* cellift = 32'd1 */
wire [2:0] _2995_;
wire [2:0] _2996_;
/* cellift = 32'd1 */
wire [2:0] _2997_;
wire [2:0] _2998_;
/* cellift = 32'd1 */
wire [2:0] _2999_;
wire [2:0] _3000_;
/* cellift = 32'd1 */
wire [2:0] _3001_;
wire [2:0] _3002_;
/* cellift = 32'd1 */
wire [2:0] _3003_;
wire [2:0] _3004_;
/* cellift = 32'd1 */
wire [2:0] _3005_;
wire [2:0] _3006_;
/* cellift = 32'd1 */
wire [2:0] _3007_;
wire [2:0] _3008_;
/* cellift = 32'd1 */
wire [2:0] _3009_;
wire [2:0] _3010_;
/* cellift = 32'd1 */
wire [2:0] _3011_;
wire [2:0] _3012_;
/* cellift = 32'd1 */
wire [2:0] _3013_;
wire [2:0] _3014_;
wire [2:0] _3015_;
/* cellift = 32'd1 */
wire [2:0] _3016_;
wire [2:0] _3017_;
/* cellift = 32'd1 */
wire [2:0] _3018_;
wire [31:0] _3019_;
/* src = "generated/sv2v_out.v:13935.30-13935.54" */
wire _3020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13935.30-13935.54" */
wire _3021_;
/* src = "generated/sv2v_out.v:14087.409-14087.428" */
wire _3022_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.409-14087.428" */
wire _3023_;
/* src = "generated/sv2v_out.v:14087.388-14087.407" */
wire _3024_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.388-14087.407" */
wire _3025_;
/* src = "generated/sv2v_out.v:14087.367-14087.386" */
wire _3026_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.367-14087.386" */
wire _3027_;
/* src = "generated/sv2v_out.v:14087.346-14087.365" */
wire _3028_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.346-14087.365" */
wire _3029_;
/* src = "generated/sv2v_out.v:14087.325-14087.344" */
wire _3030_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.325-14087.344" */
wire _3031_;
/* src = "generated/sv2v_out.v:14087.304-14087.323" */
wire _3032_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.304-14087.323" */
wire _3033_;
/* src = "generated/sv2v_out.v:14087.283-14087.302" */
wire _3034_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.283-14087.302" */
wire _3035_;
/* src = "generated/sv2v_out.v:14087.262-14087.281" */
wire _3036_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.262-14087.281" */
wire _3037_;
/* src = "generated/sv2v_out.v:14087.241-14087.260" */
wire _3038_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.241-14087.260" */
wire _3039_;
/* src = "generated/sv2v_out.v:14087.220-14087.239" */
wire _3040_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.220-14087.239" */
wire _3041_;
/* src = "generated/sv2v_out.v:14087.199-14087.218" */
wire _3042_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.199-14087.218" */
wire _3043_;
/* src = "generated/sv2v_out.v:14087.178-14087.197" */
wire _3044_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.178-14087.197" */
wire _3045_;
/* src = "generated/sv2v_out.v:14087.157-14087.176" */
wire _3046_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.157-14087.176" */
wire _3047_;
/* src = "generated/sv2v_out.v:14087.136-14087.155" */
wire _3048_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.136-14087.155" */
wire _3049_;
/* src = "generated/sv2v_out.v:14087.115-14087.134" */
wire _3050_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.115-14087.134" */
wire _3051_;
/* src = "generated/sv2v_out.v:14087.94-14087.113" */
wire _3052_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.94-14087.113" */
wire _3053_;
/* src = "generated/sv2v_out.v:14087.73-14087.92" */
wire _3054_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.73-14087.92" */
wire _3055_;
/* src = "generated/sv2v_out.v:14087.52-14087.71" */
wire _3056_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.52-14087.71" */
wire _3057_;
/* src = "generated/sv2v_out.v:14087.31-14087.50" */
wire _3058_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.31-14087.50" */
wire _3059_;
/* src = "generated/sv2v_out.v:14087.10-14087.29" */
wire _3060_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14087.10-14087.29" */
wire _3061_;
/* src = "generated/sv2v_out.v:14104.46-14104.75" */
wire _3062_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14104.46-14104.75" */
wire _3063_;
/* src = "generated/sv2v_out.v:14104.15-14104.44" */
wire _3064_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14104.15-14104.44" */
wire _3065_;
/* src = "generated/sv2v_out.v:14249.56-14249.72" */
wire _3066_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14249.56-14249.72" */
wire _3067_;
/* src = "generated/sv2v_out.v:14249.38-14249.54" */
wire _3068_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14249.38-14249.54" */
wire _3069_;
/* src = "generated/sv2v_out.v:14249.20-14249.36" */
wire _3070_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14249.20-14249.36" */
wire _3071_;
/* src = "generated/sv2v_out.v:14801.50-14801.69" */
wire _3072_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14801.50-14801.69" */
wire _3073_;
/* src = "generated/sv2v_out.v:14131.10-14131.66" */
wire _3074_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14131.10-14131.66" */
wire _3075_;
/* src = "generated/sv2v_out.v:14143.10-14143.60" */
wire _3076_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14143.10-14143.60" */
wire _3077_;
/* src = "generated/sv2v_out.v:14198.12-14198.38" */
wire _3078_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14198.12-14198.38" */
wire _3079_;
/* src = "generated/sv2v_out.v:14131.11-14131.35" */
wire _3080_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14131.11-14131.35" */
wire _3081_;
/* src = "generated/sv2v_out.v:14131.41-14131.65" */
wire _3082_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14131.41-14131.65" */
wire _3083_;
/* src = "generated/sv2v_out.v:14143.11-14143.32" */
wire _3084_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14143.11-14143.32" */
wire _3085_;
/* src = "generated/sv2v_out.v:14143.38-14143.59" */
wire _3086_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14143.38-14143.59" */
wire _3087_;
/* src = "generated/sv2v_out.v:14213.9-14213.33" */
wire _3088_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14213.9-14213.33" */
wire _3089_;
/* src = "generated/sv2v_out.v:0.0-0.0" */
wire [31:0] _3090_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:0.0-0.0" */
wire [31:0] _3091_;
/* src = "generated/sv2v_out.v:14250.47-14250.66" */
wire _3092_;
/* src = "generated/sv2v_out.v:14634.40-14634.57" */
wire _3093_;
/* src = "generated/sv2v_out.v:14845.50-14845.89" */
wire _3094_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14845.50-14845.89" */
wire _3095_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:0.0-0.0" */
wire [31:0] _3096_;
/* src = "generated/sv2v_out.v:13936.48-13936.79" */
wire _3097_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13936.48-13936.79" */
wire _3098_;
/* src = "generated/sv2v_out.v:13936.47-13936.99" */
wire _3099_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13936.47-13936.99" */
wire _3100_;
/* src = "generated/sv2v_out.v:13936.46-13936.118" */
wire _3101_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13936.46-13936.118" */
wire _3102_;
/* src = "generated/sv2v_out.v:13991.30-13991.55" */
wire _3103_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13991.30-13991.55" */
wire _3104_;
/* src = "generated/sv2v_out.v:14244.26-14244.51" */
wire [31:0] _3105_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14244.26-14244.51" */
wire [31:0] _3106_;
/* src = "generated/sv2v_out.v:14845.52-14845.88" */
wire _3107_;
/* src = "generated/sv2v_out.v:14858.31-14858.54" */
wire _3108_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:14858.31-14858.54" */
wire _3109_;
wire _3110_;
/* cellift = 32'd1 */
wire _3111_;
wire [2:0] _3112_;
/* cellift = 32'd1 */
wire [2:0] _3113_;
wire [2:0] _3114_;
/* cellift = 32'd1 */
wire [2:0] _3115_;
wire _3116_;
/* cellift = 32'd1 */
wire _3117_;
wire _3118_;
/* cellift = 32'd1 */
wire _3119_;
wire _3120_;
/* cellift = 32'd1 */
wire _3121_;
wire _3122_;
/* cellift = 32'd1 */
wire _3123_;
wire [31:0] _3124_;
/* cellift = 32'd1 */
wire [31:0] _3125_;
wire [31:0] _3126_;
/* cellift = 32'd1 */
wire [31:0] _3127_;
wire _3128_;
/* cellift = 32'd1 */
wire _3129_;
wire _3130_;
/* cellift = 32'd1 */
wire _3131_;
wire _3132_;
/* cellift = 32'd1 */
wire _3133_;
wire _3134_;
/* cellift = 32'd1 */
wire _3135_;
wire _3136_;
/* cellift = 32'd1 */
wire _3137_;
wire _3138_;
/* cellift = 32'd1 */
wire _3139_;
wire [6:0] _3140_;
/* cellift = 32'd1 */
wire [6:0] _3141_;
wire [6:0] _3142_;
/* cellift = 32'd1 */
wire [6:0] _3143_;
wire _3144_;
/* cellift = 32'd1 */
wire _3145_;
wire _3146_;
/* cellift = 32'd1 */
wire _3147_;
wire [31:0] _3148_;
/* cellift = 32'd1 */
wire [31:0] _3149_;
wire [31:0] _3150_;
/* cellift = 32'd1 */
wire [31:0] _3151_;
wire _3152_;
/* cellift = 32'd1 */
wire _3153_;
wire _3154_;
/* cellift = 32'd1 */
wire _3155_;
wire [1:0] _3156_;
/* cellift = 32'd1 */
wire [1:0] _3157_;
wire [1:0] _3158_;
/* cellift = 32'd1 */
wire [1:0] _3159_;
wire _3160_;
wire _3161_;
wire [30:0] _3162_;
/* cellift = 32'd1 */
wire [30:0] _3163_;
wire _3164_;
/* cellift = 32'd1 */
wire _3165_;
wire [30:0] _3166_;
/* cellift = 32'd1 */
wire [30:0] _3167_;
wire _3168_;
/* cellift = 32'd1 */
wire _3169_;
wire _3170_;
wire _3171_;
wire _3172_;
wire _3173_;
wire _3174_;
wire _3175_;
/* cellift = 32'd1 */
wire _3176_;
wire _3177_;
wire _3178_;
wire _3179_;
wire _3180_;
wire _3181_;
wire _3182_;
/* cellift = 32'd1 */
wire _3183_;
wire [28:0] _3184_;
/* cellift = 32'd1 */
wire [28:0] _3185_;
wire _3186_;
/* cellift = 32'd1 */
wire _3187_;
wire _3188_;
/* cellift = 32'd1 */
wire _3189_;
wire _3190_;
/* cellift = 32'd1 */
wire _3191_;
wire _3192_;
wire _3193_;
/* cellift = 32'd1 */
wire _3194_;
wire _3195_;
/* cellift = 32'd1 */
wire _3196_;
wire _3197_;
/* cellift = 32'd1 */
wire _3198_;
wire _3199_;
/* cellift = 32'd1 */
wire _3200_;
wire _3201_;
/* cellift = 32'd1 */
wire _3202_;
wire _3203_;
/* cellift = 32'd1 */
wire _3204_;
wire _3205_;
/* cellift = 32'd1 */
wire _3206_;
wire _3207_;
/* cellift = 32'd1 */
wire _3208_;
wire _3209_;
/* cellift = 32'd1 */
wire _3210_;
wire _3211_;
/* cellift = 32'd1 */
wire _3212_;
wire _3213_;
/* cellift = 32'd1 */
wire _3214_;
wire _3215_;
/* cellift = 32'd1 */
wire _3216_;
wire _3217_;
/* cellift = 32'd1 */
wire _3218_;
wire _3219_;
/* cellift = 32'd1 */
wire _3220_;
wire _3221_;
/* cellift = 32'd1 */
wire _3222_;
wire _3223_;
/* cellift = 32'd1 */
wire _3224_;
wire _3225_;
/* cellift = 32'd1 */
wire _3226_;
wire _3227_;
/* cellift = 32'd1 */
wire _3228_;
wire _3229_;
/* cellift = 32'd1 */
wire _3230_;
wire _3231_;
/* cellift = 32'd1 */
wire _3232_;
wire _3233_;
/* cellift = 32'd1 */
wire _3234_;
wire _3235_;
/* cellift = 32'd1 */
wire _3236_;
wire _3237_;
/* cellift = 32'd1 */
wire _3238_;
wire _3239_;
/* cellift = 32'd1 */
wire _3240_;
wire _3241_;
/* cellift = 32'd1 */
wire _3242_;
wire _3243_;
/* cellift = 32'd1 */
wire _3244_;
wire _3245_;
/* cellift = 32'd1 */
wire _3246_;
wire _3247_;
/* cellift = 32'd1 */
wire _3248_;
wire _3249_;
/* cellift = 32'd1 */
wire _3250_;
wire _3251_;
/* cellift = 32'd1 */
wire _3252_;
wire _3253_;
/* cellift = 32'd1 */
wire _3254_;
wire _3255_;
wire _3256_;
/* cellift = 32'd1 */
wire _3257_;
wire _3258_;
/* cellift = 32'd1 */
wire _3259_;
wire [1:0] _3260_;
/* cellift = 32'd1 */
wire [1:0] _3261_;
wire _3262_;
/* cellift = 32'd1 */
wire _3263_;
wire _3264_;
/* cellift = 32'd1 */
wire _3265_;
wire _3266_;
/* cellift = 32'd1 */
wire _3267_;
wire _3268_;
/* cellift = 32'd1 */
wire _3269_;
/* src = "generated/sv2v_out.v:13991.58-13991.116" */
wire [25:0] _3270_;
/* src = "generated/sv2v_out.v:13755.20-13755.31" */
input [31:0] boot_addr_i;
wire [31:0] boot_addr_i;
/* cellift = 32'd1 */
input [31:0] boot_addr_i_t0;
wire [31:0] boot_addr_i_t0;
/* src = "generated/sv2v_out.v:13811.13-13811.21" */
input branch_i;
wire branch_i;
/* cellift = 32'd1 */
input branch_i_t0;
wire branch_i_t0;
/* src = "generated/sv2v_out.v:13812.13-13812.27" */
input branch_taken_i;
wire branch_taken_i;
/* cellift = 32'd1 */
input branch_taken_i_t0;
wire branch_taken_i_t0;
/* src = "generated/sv2v_out.v:13747.13-13747.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:13910.12-13910.29" */
wire [7:0] cpuctrlsts_part_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13910.12-13910.29" */
wire [7:0] cpuctrlsts_part_d_t0;
/* src = "generated/sv2v_out.v:13914.7-13914.26" */
wire cpuctrlsts_part_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13914.7-13914.26" */
wire cpuctrlsts_part_err_t0;
/* src = "generated/sv2v_out.v:13909.13-13909.30" */
wire [7:0] cpuctrlsts_part_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13909.13-13909.30" */
wire [7:0] cpuctrlsts_part_q_t0;
/* src = "generated/sv2v_out.v:13913.6-13913.24" */
wire cpuctrlsts_part_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13913.6-13913.24" */
wire cpuctrlsts_part_we_t0;
/* src = "generated/sv2v_out.v:13756.13-13756.25" */
input csr_access_i;
wire csr_access_i;
/* cellift = 32'd1 */
input csr_access_i_t0;
wire csr_access_i_t0;
/* src = "generated/sv2v_out.v:13757.20-13757.30" */
input [11:0] csr_addr_i;
wire [11:0] csr_addr_i;
/* cellift = 32'd1 */
input [11:0] csr_addr_i_t0;
wire [11:0] csr_addr_i_t0;
/* src = "generated/sv2v_out.v:13779.21-13779.31" */
output [31:0] csr_depc_o;
wire [31:0] csr_depc_o;
/* cellift = 32'd1 */
output [31:0] csr_depc_o_t0;
wire [31:0] csr_depc_o_t0;
/* src = "generated/sv2v_out.v:13801.19-13801.31" */
input [6:0] csr_mcause_i;
wire [6:0] csr_mcause_i;
/* cellift = 32'd1 */
input [6:0] csr_mcause_i_t0;
wire [6:0] csr_mcause_i_t0;
/* src = "generated/sv2v_out.v:13770.21-13770.31" */
output [31:0] csr_mepc_o;
wire [31:0] csr_mepc_o;
/* cellift = 32'd1 */
output [31:0] csr_mepc_o_t0;
wire [31:0] csr_mepc_o_t0;
/* src = "generated/sv2v_out.v:13769.14-13769.31" */
output csr_mstatus_mie_o;
wire csr_mstatus_mie_o;
/* cellift = 32'd1 */
output csr_mstatus_mie_o_t0;
wire csr_mstatus_mie_o_t0;
/* src = "generated/sv2v_out.v:13752.14-13752.30" */
output csr_mstatus_tw_o;
wire csr_mstatus_tw_o;
/* cellift = 32'd1 */
output csr_mstatus_tw_o_t0;
wire csr_mstatus_tw_o_t0;
/* src = "generated/sv2v_out.v:13802.20-13802.31" */
input [31:0] csr_mtval_i;
wire [31:0] csr_mtval_i;
/* cellift = 32'd1 */
input [31:0] csr_mtval_i_t0;
wire [31:0] csr_mtval_i_t0;
/* src = "generated/sv2v_out.v:13771.21-13771.32" */
output [31:0] csr_mtval_o;
wire [31:0] csr_mtval_o;
/* cellift = 32'd1 */
output [31:0] csr_mtval_o_t0;
wire [31:0] csr_mtval_o_t0;
/* src = "generated/sv2v_out.v:13754.13-13754.29" */
input csr_mtvec_init_i;
wire csr_mtvec_init_i;
/* cellift = 32'd1 */
input csr_mtvec_init_i_t0;
wire csr_mtvec_init_i_t0;
/* src = "generated/sv2v_out.v:13753.21-13753.32" */
output [31:0] csr_mtvec_o;
wire [31:0] csr_mtvec_o;
/* cellift = 32'd1 */
output [31:0] csr_mtvec_o_t0;
wire [31:0] csr_mtvec_o_t0;
/* src = "generated/sv2v_out.v:13760.8-13760.19" */
input csr_op_en_i;
wire csr_op_en_i;
/* cellift = 32'd1 */
input csr_op_en_i_t0;
wire csr_op_en_i_t0;
/* src = "generated/sv2v_out.v:13759.19-13759.27" */
input [1:0] csr_op_i;
wire [1:0] csr_op_i;
/* cellift = 32'd1 */
input [1:0] csr_op_i_t0;
wire [1:0] csr_op_i_t0;
/* src = "generated/sv2v_out.v:13773.43-13773.57" */
output [135:0] csr_pmp_addr_o;
wire [135:0] csr_pmp_addr_o;
/* cellift = 32'd1 */
output [135:0] csr_pmp_addr_o_t0;
wire [135:0] csr_pmp_addr_o_t0;
/* src = "generated/sv2v_out.v:13772.42-13772.55" */
output [23:0] csr_pmp_cfg_o;
wire [23:0] csr_pmp_cfg_o;
/* cellift = 32'd1 */
output [23:0] csr_pmp_cfg_o_t0;
wire [23:0] csr_pmp_cfg_o_t0;
/* src = "generated/sv2v_out.v:13774.20-13774.37" */
output [2:0] csr_pmp_mseccfg_o;
wire [2:0] csr_pmp_mseccfg_o;
/* cellift = 32'd1 */
output [2:0] csr_pmp_mseccfg_o_t0;
wire [2:0] csr_pmp_mseccfg_o_t0;
/* src = "generated/sv2v_out.v:13761.21-13761.32" */
output [31:0] csr_rdata_o;
wire [31:0] csr_rdata_o;
/* cellift = 32'd1 */
output [31:0] csr_rdata_o_t0;
wire [31:0] csr_rdata_o_t0;
/* src = "generated/sv2v_out.v:13799.13-13799.31" */
input csr_restore_dret_i;
wire csr_restore_dret_i;
/* cellift = 32'd1 */
input csr_restore_dret_i_t0;
wire csr_restore_dret_i_t0;
/* src = "generated/sv2v_out.v:13798.13-13798.31" */
input csr_restore_mret_i;
wire csr_restore_mret_i;
/* cellift = 32'd1 */
input csr_restore_mret_i_t0;
wire csr_restore_mret_i_t0;
/* src = "generated/sv2v_out.v:13800.13-13800.29" */
input csr_save_cause_i;
wire csr_save_cause_i;
/* cellift = 32'd1 */
input csr_save_cause_i_t0;
wire csr_save_cause_i_t0;
/* src = "generated/sv2v_out.v:13796.13-13796.26" */
input csr_save_id_i;
wire csr_save_id_i;
/* cellift = 32'd1 */
input csr_save_id_i_t0;
wire csr_save_id_i_t0;
/* src = "generated/sv2v_out.v:13795.13-13795.26" */
input csr_save_if_i;
wire csr_save_if_i;
/* cellift = 32'd1 */
input csr_save_if_i_t0;
wire csr_save_if_i_t0;
/* src = "generated/sv2v_out.v:13797.13-13797.26" */
input csr_save_wb_i;
wire csr_save_wb_i;
/* cellift = 32'd1 */
input csr_save_wb_i_t0;
wire csr_save_wb_i_t0;
/* src = "generated/sv2v_out.v:13793.14-13793.30" */
output csr_shadow_err_o;
wire csr_shadow_err_o;
/* cellift = 32'd1 */
output csr_shadow_err_o_t0;
wire csr_shadow_err_o_t0;
/* src = "generated/sv2v_out.v:13758.20-13758.31" */
input [31:0] csr_wdata_i;
wire [31:0] csr_wdata_i;
/* cellift = 32'd1 */
input [31:0] csr_wdata_i_t0;
wire [31:0] csr_wdata_i_t0;
/* src = "generated/sv2v_out.v:13919.7-13919.17" */
wire csr_we_int;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13919.7-13919.17" */
wire csr_we_int_t0;
/* src = "generated/sv2v_out.v:13920.7-13920.13" */
wire csr_wr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13920.7-13920.13" */
wire csr_wr_t0;
/* src = "generated/sv2v_out.v:13787.14-13787.31" */
output data_ind_timing_o;
wire data_ind_timing_o;
/* cellift = 32'd1 */
output data_ind_timing_o_t0;
wire data_ind_timing_o_t0;
/* src = "generated/sv2v_out.v:13921.6-13921.13" */
wire dbg_csr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13921.6-13921.13" */
wire dbg_csr_t0;
/* src = "generated/sv2v_out.v:13869.13-13869.19" */
wire [31:0] dcsr_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13869.13-13869.19" */
wire [31:0] dcsr_d_t0;
/* src = "generated/sv2v_out.v:13870.6-13870.13" */
wire dcsr_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13870.6-13870.13" */
wire dcsr_en_t0;
/* src = "generated/sv2v_out.v:13868.14-13868.20" */
wire [31:0] dcsr_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13868.14-13868.20" */
wire [31:0] dcsr_q_t0;
/* src = "generated/sv2v_out.v:13777.19-13777.32" */
input [2:0] debug_cause_i;
wire [2:0] debug_cause_i;
/* cellift = 32'd1 */
input [2:0] debug_cause_i_t0;
wire [2:0] debug_cause_i_t0;
/* src = "generated/sv2v_out.v:13778.13-13778.29" */
input debug_csr_save_i;
wire debug_csr_save_i;
/* cellift = 32'd1 */
input debug_csr_save_i_t0;
wire debug_csr_save_i_t0;
/* src = "generated/sv2v_out.v:13781.14-13781.29" */
output debug_ebreakm_o;
wire debug_ebreakm_o;
/* cellift = 32'd1 */
output debug_ebreakm_o_t0;
wire debug_ebreakm_o_t0;
/* src = "generated/sv2v_out.v:13782.14-13782.29" */
output debug_ebreaku_o;
wire debug_ebreaku_o;
/* cellift = 32'd1 */
output debug_ebreaku_o_t0;
wire debug_ebreaku_o_t0;
/* src = "generated/sv2v_out.v:13776.13-13776.34" */
input debug_mode_entering_i;
wire debug_mode_entering_i;
/* cellift = 32'd1 */
input debug_mode_entering_i_t0;
wire debug_mode_entering_i_t0;
/* src = "generated/sv2v_out.v:13775.13-13775.25" */
input debug_mode_i;
wire debug_mode_i;
/* cellift = 32'd1 */
input debug_mode_i_t0;
wire debug_mode_i_t0;
/* src = "generated/sv2v_out.v:13780.14-13780.33" */
output debug_single_step_o;
wire debug_single_step_o;
/* cellift = 32'd1 */
output debug_single_step_o_t0;
wire debug_single_step_o_t0;
/* src = "generated/sv2v_out.v:13872.13-13872.19" */
wire [31:0] depc_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13872.13-13872.19" */
wire [31:0] depc_d_t0;
/* src = "generated/sv2v_out.v:13873.6-13873.13" */
wire depc_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13873.6-13873.13" */
wire depc_en_t0;
/* src = "generated/sv2v_out.v:13817.13-13817.23" */
input div_wait_i;
wire div_wait_i;
/* cellift = 32'd1 */
input div_wait_i_t0;
wire div_wait_i_t0;
/* src = "generated/sv2v_out.v:13804.13-13804.32" */
output double_fault_seen_o;
wire double_fault_seen_o;
/* cellift = 32'd1 */
output double_fault_seen_o_t0;
wire double_fault_seen_o_t0;
/* src = "generated/sv2v_out.v:13876.6-13876.18" */
wire dscratch0_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13876.6-13876.18" */
wire dscratch0_en_t0;
/* src = "generated/sv2v_out.v:13874.14-13874.25" */
wire [31:0] dscratch0_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13874.14-13874.25" */
wire [31:0] dscratch0_q_t0;
/* src = "generated/sv2v_out.v:13877.6-13877.18" */
wire dscratch1_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13877.6-13877.18" */
wire dscratch1_en_t0;
/* src = "generated/sv2v_out.v:13875.14-13875.25" */
wire [31:0] dscratch1_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13875.14-13875.25" */
wire [31:0] dscratch1_q_t0;
/* src = "generated/sv2v_out.v:13815.13-13815.25" */
input dside_wait_i;
wire dside_wait_i;
/* cellift = 32'd1 */
input dside_wait_i_t0;
wire dside_wait_i_t0;
/* src = "generated/sv2v_out.v:13788.14-13788.30" */
output dummy_instr_en_o;
wire dummy_instr_en_o;
/* cellift = 32'd1 */
output dummy_instr_en_o_t0;
wire dummy_instr_en_o_t0;
/* src = "generated/sv2v_out.v:13789.20-13789.38" */
output [2:0] dummy_instr_mask_o;
wire [2:0] dummy_instr_mask_o;
/* cellift = 32'd1 */
output [2:0] dummy_instr_mask_o_t0;
wire [2:0] dummy_instr_mask_o_t0;
/* src = "generated/sv2v_out.v:13790.14-13790.35" */
output dummy_instr_seed_en_o;
wire dummy_instr_seed_en_o;
/* cellift = 32'd1 */
output dummy_instr_seed_en_o_t0;
wire dummy_instr_seed_en_o_t0;
/* src = "generated/sv2v_out.v:13791.21-13791.39" */
output [31:0] dummy_instr_seed_o;
wire [31:0] dummy_instr_seed_o;
/* cellift = 32'd1 */
output [31:0] dummy_instr_seed_o_t0;
wire [31:0] dummy_instr_seed_o_t0;
/* src = "generated/sv2v_out.v:13749.20-13749.29" */
input [31:0] hart_id_i;
wire [31:0] hart_id_i;
/* cellift = 32'd1 */
input [31:0] hart_id_i_t0;
wire [31:0] hart_id_i_t0;
/* src = "generated/sv2v_out.v:13794.13-13794.31" */
input ic_scr_key_valid_i;
wire ic_scr_key_valid_i;
/* cellift = 32'd1 */
input ic_scr_key_valid_i_t0;
wire ic_scr_key_valid_i_t0;
/* src = "generated/sv2v_out.v:13792.14-13792.29" */
output icache_enable_o;
wire icache_enable_o;
/* cellift = 32'd1 */
output icache_enable_o_t0;
wire icache_enable_o_t0;
/* src = "generated/sv2v_out.v:13922.6-13922.17" */
wire illegal_csr;
/* src = "generated/sv2v_out.v:13924.7-13924.22" */
wire illegal_csr_dbg;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13924.7-13924.22" */
wire illegal_csr_dbg_t0;
/* src = "generated/sv2v_out.v:13803.14-13803.32" */
output illegal_csr_insn_o;
wire illegal_csr_insn_o;
/* cellift = 32'd1 */
output illegal_csr_insn_o_t0;
wire illegal_csr_insn_o_t0;
/* src = "generated/sv2v_out.v:13923.7-13923.23" */
wire illegal_csr_priv;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13923.7-13923.23" */
wire illegal_csr_priv_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13922.6-13922.17" */
wire illegal_csr_t0;
/* src = "generated/sv2v_out.v:13925.7-13925.24" */
wire illegal_csr_write;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13925.7-13925.24" */
wire illegal_csr_write_t0;
/* src = "generated/sv2v_out.v:13806.13-13806.35" */
input instr_ret_compressed_i;
wire instr_ret_compressed_i;
/* cellift = 32'd1 */
input instr_ret_compressed_i_t0;
wire instr_ret_compressed_i_t0;
/* src = "generated/sv2v_out.v:13808.13-13808.40" */
input instr_ret_compressed_spec_i;
wire instr_ret_compressed_spec_i;
/* cellift = 32'd1 */
input instr_ret_compressed_spec_i_t0;
wire instr_ret_compressed_spec_i_t0;
/* src = "generated/sv2v_out.v:13805.13-13805.24" */
input instr_ret_i;
wire instr_ret_i;
/* cellift = 32'd1 */
input instr_ret_i_t0;
wire instr_ret_i_t0;
/* src = "generated/sv2v_out.v:13807.13-13807.29" */
input instr_ret_spec_i;
wire instr_ret_spec_i;
/* cellift = 32'd1 */
input instr_ret_spec_i_t0;
wire instr_ret_spec_i_t0;
/* src = "generated/sv2v_out.v:13764.13-13764.27" */
input irq_external_i;
wire irq_external_i;
/* cellift = 32'd1 */
input irq_external_i_t0;
wire irq_external_i_t0;
/* src = "generated/sv2v_out.v:13765.20-13765.30" */
input [14:0] irq_fast_i;
wire [14:0] irq_fast_i;
/* cellift = 32'd1 */
input [14:0] irq_fast_i_t0;
wire [14:0] irq_fast_i_t0;
/* src = "generated/sv2v_out.v:13767.14-13767.27" */
output irq_pending_o;
wire irq_pending_o;
/* cellift = 32'd1 */
output irq_pending_o_t0;
wire irq_pending_o_t0;
/* src = "generated/sv2v_out.v:13762.13-13762.27" */
input irq_software_i;
wire irq_software_i;
/* cellift = 32'd1 */
input irq_software_i_t0;
wire irq_software_i_t0;
/* src = "generated/sv2v_out.v:13763.13-13763.24" */
input irq_timer_i;
wire irq_timer_i;
/* cellift = 32'd1 */
input irq_timer_i_t0;
wire irq_timer_i_t0;
/* src = "generated/sv2v_out.v:13768.21-13768.27" */
output [17:0] irqs_o;
wire [17:0] irqs_o;
/* cellift = 32'd1 */
output [17:0] irqs_o_t0;
wire [17:0] irqs_o_t0;
/* src = "generated/sv2v_out.v:13809.13-13809.25" */
input iside_wait_i;
wire iside_wait_i;
/* cellift = 32'd1 */
input iside_wait_i_t0;
wire iside_wait_i_t0;
/* src = "generated/sv2v_out.v:13810.13-13810.19" */
input jump_i;
wire jump_i;
/* cellift = 32'd1 */
input jump_i_t0;
wire jump_i_t0;
/* src = "generated/sv2v_out.v:13858.12-13858.20" */
wire [6:0] mcause_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13858.12-13858.20" */
wire [6:0] mcause_d_t0;
/* src = "generated/sv2v_out.v:13859.6-13859.15" */
wire mcause_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13859.6-13859.15" */
wire mcause_en_t0;
/* src = "generated/sv2v_out.v:13857.13-13857.21" */
wire [6:0] mcause_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13857.13-13857.21" */
wire [6:0] mcause_q_t0;
/* src = "generated/sv2v_out.v:13891.14-13891.27" */
wire [31:0] mcountinhibit;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13891.14-13891.27" */
wire [31:0] mcountinhibit_t0;
/* src = "generated/sv2v_out.v:13894.6-13894.22" */
wire mcountinhibit_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13894.6-13894.22" */
wire mcountinhibit_we_t0;
/* src = "generated/sv2v_out.v:13813.13-13813.23" */
input mem_load_i;
wire mem_load_i;
/* cellift = 32'd1 */
input mem_load_i_t0;
wire mem_load_i_t0;
/* src = "generated/sv2v_out.v:13814.13-13814.24" */
input mem_store_i;
wire mem_store_i;
/* cellift = 32'd1 */
input mem_store_i_t0;
wire mem_store_i_t0;
/* src = "generated/sv2v_out.v:13855.13-13855.19" */
wire [31:0] mepc_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13855.13-13855.19" */
wire [31:0] mepc_d_t0;
/* src = "generated/sv2v_out.v:13856.6-13856.13" */
wire mepc_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13856.6-13856.13" */
wire mepc_en_t0;
/* src = "generated/sv2v_out.v:13895.14-13895.25" */
wire [63:0] \mhpmcounter[0] ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13895.14-13895.25" */
wire [63:0] \mhpmcounter[0]_t0 ;
/* src = "generated/sv2v_out.v:13895.14-13895.25" */
wire [63:0] \mhpmcounter[2] ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13895.14-13895.25" */
wire [63:0] \mhpmcounter[2]_t0 ;
/* src = "generated/sv2v_out.v:13896.13-13896.27" */
/* unused_bits = "1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] mhpmcounter_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13896.13-13896.27" */
/* unused_bits = "1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] mhpmcounter_we_t0;
/* src = "generated/sv2v_out.v:13897.13-13897.28" */
/* unused_bits = "1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] mhpmcounterh_we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13897.13-13897.28" */
/* unused_bits = "1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] mhpmcounterh_we_t0;
/* src = "generated/sv2v_out.v:13851.6-13851.12" */
wire mie_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13851.6-13851.12" */
wire mie_en_t0;
/* src = "generated/sv2v_out.v:13849.14-13849.19" */
wire [17:0] mie_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13849.14-13849.19" */
wire [17:0] mie_q_t0;
/* src = "generated/sv2v_out.v:13904.14-13904.27" */
wire [63:0] minstret_next;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13904.14-13904.27" */
wire [63:0] minstret_next_t0;
/* src = "generated/sv2v_out.v:13905.14-13905.26" */
wire [63:0] minstret_raw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13905.14-13905.26" */
wire [63:0] minstret_raw_t0;
/* src = "generated/sv2v_out.v:13853.6-13853.17" */
wire mscratch_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13853.6-13853.17" */
wire mscratch_en_t0;
/* src = "generated/sv2v_out.v:13852.14-13852.24" */
wire [31:0] mscratch_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13852.14-13852.24" */
wire [31:0] mscratch_q_t0;
/* src = "generated/sv2v_out.v:13883.13-13883.27" */
wire [6:0] mstack_cause_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13883.13-13883.27" */
wire [6:0] mstack_cause_q_t0;
/* src = "generated/sv2v_out.v:13880.6-13880.15" */
wire mstack_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13880.6-13880.15" */
wire mstack_en_t0;
/* src = "generated/sv2v_out.v:13881.14-13881.26" */
wire [31:0] mstack_epc_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13881.14-13881.26" */
wire [31:0] mstack_epc_q_t0;
/* src = "generated/sv2v_out.v:13878.13-13878.21" */
wire [2:0] mstack_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13878.13-13878.21" */
wire [2:0] mstack_q_t0;
/* src = "generated/sv2v_out.v:13846.12-13846.21" */
wire [5:0] mstatus_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13846.12-13846.21" */
wire [5:0] mstatus_d_t0;
/* src = "generated/sv2v_out.v:13848.6-13848.16" */
wire mstatus_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13848.6-13848.16" */
wire mstatus_en_t0;
/* src = "generated/sv2v_out.v:13847.7-13847.18" */
wire mstatus_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13847.7-13847.18" */
wire mstatus_err_t0;
/* src = "generated/sv2v_out.v:13845.13-13845.22" */
wire [5:0] mstatus_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13845.13-13845.22" */
wire [5:0] mstatus_q_t0;
/* src = "generated/sv2v_out.v:13861.13-13861.20" */
wire [31:0] mtval_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13861.13-13861.20" */
wire [31:0] mtval_d_t0;
/* src = "generated/sv2v_out.v:13862.6-13862.14" */
wire mtval_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13862.6-13862.14" */
wire mtval_en_t0;
/* src = "generated/sv2v_out.v:13864.13-13864.20" */
wire [31:0] mtvec_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13864.13-13864.20" */
wire [31:0] mtvec_d_t0;
/* src = "generated/sv2v_out.v:13866.6-13866.14" */
wire mtvec_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13866.6-13866.14" */
wire mtvec_en_t0;
/* src = "generated/sv2v_out.v:13865.7-13865.16" */
wire mtvec_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13865.7-13865.16" */
wire mtvec_err_t0;
/* src = "generated/sv2v_out.v:13816.13-13816.23" */
input mul_wait_i;
wire mul_wait_i;
/* cellift = 32'd1 */
input mul_wait_i_t0;
wire mul_wait_i_t0;
/* src = "generated/sv2v_out.v:13766.13-13766.23" */
input nmi_mode_i;
wire nmi_mode_i;
/* cellift = 32'd1 */
input nmi_mode_i_t0;
wire nmi_mode_i_t0;
/* src = "generated/sv2v_out.v:13785.20-13785.27" */
input [31:0] pc_id_i;
wire [31:0] pc_id_i;
/* cellift = 32'd1 */
input [31:0] pc_id_i_t0;
wire [31:0] pc_id_i_t0;
/* src = "generated/sv2v_out.v:13784.20-13784.27" */
input [31:0] pc_if_i;
wire [31:0] pc_if_i;
/* cellift = 32'd1 */
input [31:0] pc_if_i_t0;
wire [31:0] pc_if_i_t0;
/* src = "generated/sv2v_out.v:13786.20-13786.27" */
input [31:0] pc_wb_i;
wire [31:0] pc_wb_i;
/* cellift = 32'd1 */
input [31:0] pc_wb_i_t0;
wire [31:0] pc_wb_i_t0;
/* src = "generated/sv2v_out.v:13844.12-13844.22" */
wire [1:0] priv_lvl_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13844.12-13844.22" */
wire [1:0] priv_lvl_d_t0;
/* src = "generated/sv2v_out.v:13750.20-13750.34" */
output [1:0] priv_mode_id_o;
reg [1:0] priv_mode_id_o;
/* cellift = 32'd1 */
output [1:0] priv_mode_id_o_t0;
reg [1:0] priv_mode_id_o_t0;
/* src = "generated/sv2v_out.v:13751.20-13751.35" */
output [1:0] priv_mode_lsu_o;
wire [1:0] priv_mode_lsu_o;
/* cellift = 32'd1 */
output [1:0] priv_mode_lsu_o_t0;
wire [1:0] priv_mode_lsu_o_t0;
/* src = "generated/sv2v_out.v:13748.13-13748.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:13783.14-13783.29" */
output trigger_match_o;
wire trigger_match_o;
/* cellift = 32'd1 */
output trigger_match_o_t0;
wire trigger_match_o_t0;
assign illegal_csr_dbg = dbg_csr & /* src = "generated/sv2v_out.v:13933.27-13933.50" */ _0349_;
assign illegal_csr_insn_o = csr_access_i & /* src = "generated/sv2v_out.v:13936.30-13936.119" */ _3101_;
assign _0145_ = _0414_ & /* src = "generated/sv2v_out.v:14245.26-14245.52" */ csr_rdata_o;
assign _0147_ = csr_wr & /* src = "generated/sv2v_out.v:14250.23-14250.43" */ csr_op_en_i;
assign csr_we_int = _0147_ & /* src = "generated/sv2v_out.v:14250.22-14250.66" */ _3092_;
assign irqs_o = { irq_software_i, irq_timer_i, irq_external_i, irq_fast_i } & /* src = "generated/sv2v_out.v:14261.18-14261.29" */ mie_q;
assign _0150_ = instr_ret_i & /* src = "generated/sv2v_out.v:14634.18-14634.57" */ _3093_;
assign _0152_ = instr_ret_spec_i & /* src = "generated/sv2v_out.v:14641.27-14641.63" */ _3093_;
assign icache_enable_o = cpuctrlsts_part_q[0] & /* src = "generated/sv2v_out.v:14845.27-14845.89" */ _3094_;
assign _0154_ = ~ _0452_;
assign _0155_ = ~ mcountinhibit_we;
assign _2154_ = priv_lvl_d ^ priv_mode_id_o;
assign _2155_ = { dummy_instr_seed_o[2], dummy_instr_seed_o[0] } ^ { mcountinhibit[2], mcountinhibit[0] };
assign _1589_ = priv_lvl_d_t0 | priv_mode_id_o_t0;
assign _1593_ = { dummy_instr_seed_o_t0[2], dummy_instr_seed_o_t0[0] } | { mcountinhibit_t0[2], mcountinhibit_t0[0] };
assign _1590_ = _2154_ | _1589_;
assign _1594_ = _2155_ | _1593_;
assign _0487_ = { _0452_, _0452_ } & priv_lvl_d_t0;
assign _0490_ = { mcountinhibit_we, mcountinhibit_we } & { dummy_instr_seed_o_t0[2], dummy_instr_seed_o_t0[0] };
assign _0488_ = { _0154_, _0154_ } & priv_mode_id_o_t0;
assign _0491_ = { _0155_, _0155_ } & { mcountinhibit_t0[2], mcountinhibit_t0[0] };
assign _0489_ = _1590_ & { _0453_, _0453_ };
assign _0492_ = _1594_ & { mcountinhibit_we_t0, mcountinhibit_we_t0 };
assign _1591_ = _0487_ | _0488_;
assign _1595_ = _0490_ | _0491_;
assign _1592_ = _1591_ | _0489_;
assign _1596_ = _1595_ | _0492_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers  */
/* PC_TAINT_INFO STATE_NAME priv_mode_id_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) priv_mode_id_o_t0 <= 2'h0;
else priv_mode_id_o_t0 <= _1592_;
reg [1:0] _3299_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers  */
/* PC_TAINT_INFO STATE_NAME _3299_ */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) _3299_ <= 2'h0;
else _3299_ <= _1596_;
assign { mcountinhibit_t0[2], mcountinhibit_t0[0] } = _3299_;
assign _0460_ = dbg_csr_t0 & _0349_;
assign _0463_ = csr_access_i_t0 & _3101_;
assign _0466_ = csr_wdata_i_t0 & csr_rdata_o;
assign _0469_ = csr_wr_t0 & csr_op_en_i;
assign _0472_ = _0148_ & _3092_;
assign _0475_ = { irq_software_i_t0, irq_timer_i_t0, irq_external_i_t0, irq_fast_i_t0 } & mie_q;
assign _0478_ = instr_ret_i_t0 & _3093_;
assign _0481_ = instr_ret_spec_i_t0 & _3093_;
assign _0484_ = cpuctrlsts_part_q_t0[0] & _3094_;
assign _0461_ = debug_mode_i_t0 & dbg_csr;
assign _0464_ = _3102_ & csr_access_i;
assign _0467_ = csr_rdata_o_t0 & _0414_;
assign _0470_ = csr_op_en_i_t0 & csr_wr;
assign _0473_ = illegal_csr_insn_o_t0 & _0147_;
assign _0476_ = mie_q_t0 & { irq_software_i, irq_timer_i, irq_external_i, irq_fast_i };
assign _0479_ = mcountinhibit_t0[2] & instr_ret_i;
assign _0482_ = mcountinhibit_t0[2] & instr_ret_spec_i;
assign _0485_ = _3095_ & cpuctrlsts_part_q[0];
assign _0462_ = dbg_csr_t0 & debug_mode_i_t0;
assign _0465_ = csr_access_i_t0 & _3102_;
assign _0468_ = csr_wdata_i_t0 & csr_rdata_o_t0;
assign _0471_ = csr_wr_t0 & csr_op_en_i_t0;
assign _0474_ = _0148_ & illegal_csr_insn_o_t0;
assign _0477_ = { irq_software_i_t0, irq_timer_i_t0, irq_external_i_t0, irq_fast_i_t0 } & mie_q_t0;
assign _0480_ = instr_ret_i_t0 & mcountinhibit_t0[2];
assign _0483_ = instr_ret_spec_i_t0 & mcountinhibit_t0[2];
assign _0486_ = cpuctrlsts_part_q_t0[0] & _3095_;
assign _1580_ = _0460_ | _0461_;
assign _1581_ = _0463_ | _0464_;
assign _1582_ = _0466_ | _0467_;
assign _1583_ = _0469_ | _0470_;
assign _1584_ = _0472_ | _0473_;
assign _1585_ = _0475_ | _0476_;
assign _1586_ = _0478_ | _0479_;
assign _1587_ = _0481_ | _0482_;
assign _1588_ = _0484_ | _0485_;
assign illegal_csr_dbg_t0 = _1580_ | _0462_;
assign illegal_csr_insn_o_t0 = _1581_ | _0465_;
assign _0146_ = _1582_ | _0468_;
assign _0148_ = _1583_ | _0471_;
assign csr_we_int_t0 = _1584_ | _0474_;
assign irqs_o_t0 = _1585_ | _0477_;
assign _0151_ = _1586_ | _0480_;
assign _0153_ = _1587_ | _0483_;
assign icache_enable_o_t0 = _1588_ | _0486_;
assign _0156_ = | csr_addr_i_t0[11:10];
assign _0157_ = | dummy_instr_seed_o_t0[31:30];
assign _0160_ = | mstatus_q_t0[3:2];
assign _0162_ = | csr_addr_i_t0;
assign _0164_ = ~ csr_addr_i_t0[11:10];
assign _0165_ = ~ dummy_instr_seed_o_t0[31:30];
assign _0168_ = ~ mstatus_q_t0[3:2];
assign _0170_ = ~ csr_addr_i_t0;
assign _1163_ = csr_addr_i[11:10] & _0164_;
assign _1164_ = dummy_instr_seed_o[31:30] & _0165_;
assign _1186_ = mstatus_q[3:2] & _0168_;
assign _1543_ = csr_addr_i & _0170_;
assign _2437_ = _1163_ == _0164_;
assign _2438_ = _1164_ == { _0165_[1], 1'h0 };
assign _2439_ = _1164_ == _0165_;
assign _2440_ = _1184_ == _0166_;
assign _2441_ = _1185_ == _0167_;
assign _2442_ = _1186_ == _0168_;
assign _2443_ = _1210_ == _0169_;
assign _2444_ = _1210_ == { _0169_[1], 1'h0 };
assign _2445_ = _1210_ == { 1'h0, _0169_[0] };
assign _2446_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5], 5'h00 };
assign _2447_ = _1543_ == { _0170_[11:8], 3'h0, _0170_[4], 2'h0, _0170_[1], 1'h0 };
assign _2448_ = _1543_ == { 2'h0, _0170_[9:8], 7'h00, _0170_[0] };
assign _2449_ = _1545_ == _0171_;
assign _2450_ = _1545_ == { _0171_[4:1], 1'h0 };
assign _2451_ = _1545_ == { _0171_[4:2], 1'h0, _0171_[0] };
assign _2452_ = _1545_ == { _0171_[4:2], 2'h0 };
assign _2453_ = _1545_ == { _0171_[4:3], 1'h0, _0171_[1:0] };
assign _2454_ = _1545_ == { _0171_[4:3], 1'h0, _0171_[1], 1'h0 };
assign _2455_ = _1545_ == { _0171_[4:3], 2'h0, _0171_[0] };
assign _2456_ = _1545_ == { _0171_[4:3], 3'h0 };
assign _2457_ = _1545_ == { _0171_[4], 1'h0, _0171_[2:0] };
assign _2458_ = _1545_ == { _0171_[4], 1'h0, _0171_[2:1], 1'h0 };
assign _2459_ = _1545_ == { _0171_[4], 1'h0, _0171_[2], 1'h0, _0171_[0] };
assign _2460_ = _1545_ == { _0171_[4], 1'h0, _0171_[2], 2'h0 };
assign _2461_ = _1545_ == { _0171_[4], 2'h0, _0171_[1:0] };
assign _2462_ = _1545_ == { _0171_[4], 2'h0, _0171_[1], 1'h0 };
assign _2463_ = _1545_ == { _0171_[4], 3'h0, _0171_[0] };
assign _2464_ = _1545_ == { _0171_[4], 4'h0 };
assign _2465_ = _1545_ == { 1'h0, _0171_[3:0] };
assign _2466_ = _1545_ == { 1'h0, _0171_[3:1], 1'h0 };
assign _2467_ = _1545_ == { 1'h0, _0171_[3:2], 1'h0, _0171_[0] };
assign _2468_ = _1545_ == { 1'h0, _0171_[3:2], 2'h0 };
assign _2469_ = _1545_ == { 1'h0, _0171_[3], 1'h0, _0171_[1:0] };
assign _2470_ = _1545_ == { 1'h0, _0171_[3], 1'h0, _0171_[1], 1'h0 };
assign _2471_ = _1545_ == { 1'h0, _0171_[3], 2'h0, _0171_[0] };
assign _2472_ = _1545_ == { 1'h0, _0171_[3], 3'h0 };
assign _2473_ = _1545_ == { 2'h0, _0171_[2:0] };
assign _2474_ = _1545_ == { 2'h0, _0171_[2:1], 1'h0 };
assign _2475_ = _1545_ == { 2'h0, _0171_[2], 1'h0, _0171_[0] };
assign _2476_ = _1545_ == { 2'h0, _0171_[2], 2'h0 };
assign _2477_ = _1545_ == { 3'h0, _0171_[1:0] };
assign _2478_ = _1545_ == { 3'h0, _0171_[1], 1'h0 };
assign _2479_ = _1545_ == { 4'h0, _0171_[0] };
assign _2480_ = _1543_ == { 1'h0, _0170_[10:7], 1'h0, _0170_[5:4], 2'h0, _0170_[1:0] };
assign _2481_ = _1543_ == { 1'h0, _0170_[10:7], 1'h0, _0170_[5:4], 2'h0, _0170_[1], 1'h0 };
assign _2482_ = _1543_ == { 1'h0, _0170_[10:7], 1'h0, _0170_[5:4], 3'h0, _0170_[0] };
assign _2483_ = _1543_ == { 1'h0, _0170_[10:7], 1'h0, _0170_[5:4], 4'h0 };
assign _2484_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5:0] };
assign _2485_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5:1], 1'h0 };
assign _2486_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5:2], 1'h0, _0170_[0] };
assign _2487_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5:2], 2'h0 };
assign _2488_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5:3], 1'h0, _0170_[1:0] };
assign _2489_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5:3], 1'h0, _0170_[1], 1'h0 };
assign _2490_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5:3], 2'h0, _0170_[0] };
assign _2491_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5:3], 3'h0 };
assign _2492_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5:4], 1'h0, _0170_[2:0] };
assign _2493_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5:4], 1'h0, _0170_[2:1], 1'h0 };
assign _2494_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5:4], 1'h0, _0170_[2], 1'h0, _0170_[0] };
assign _2495_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5:4], 1'h0, _0170_[2], 2'h0 };
assign _2496_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5:4], 2'h0, _0170_[1:0] };
assign _2497_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5:4], 2'h0, _0170_[1], 1'h0 };
assign _2498_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5:4], 3'h0, _0170_[0] };
assign _2499_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5:4], 4'h0 };
assign _2500_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5], 3'h0, _0170_[1:0] };
assign _2501_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5], 3'h0, _0170_[1], 1'h0 };
assign _2502_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5], 4'h0, _0170_[0] };
assign _2503_ = _1543_ == { 2'h0, _0170_[9:7], 1'h0, _0170_[5], 5'h00 };
assign _2504_ = _1543_ == { 2'h0, _0170_[9:8], 1'h0, _0170_[6], 3'h0, _0170_[2], 2'h0 };
assign _2505_ = _1543_ == { 2'h0, _0170_[9:8], 1'h0, _0170_[6], 4'h0, _0170_[1:0] };
assign _2506_ = _1543_ == { 2'h0, _0170_[9:8], 1'h0, _0170_[6], 4'h0, _0170_[1], 1'h0 };
assign _2507_ = _1543_ == { 2'h0, _0170_[9:8], 1'h0, _0170_[6], 5'h00, _0170_[0] };
assign _2508_ = _1543_ == { 2'h0, _0170_[9:8], 5'h00, _0170_[2], 1'h0, _0170_[0] };
assign _2509_ = _1543_ == { 2'h0, _0170_[9:8], 1'h0, _0170_[6], 6'h00 };
assign _2510_ = _1543_ == { 2'h0, _0170_[9:8], 5'h00, _0170_[2], 2'h0 };
assign _2511_ = _1543_ == { 2'h0, _0170_[9:8], 8'h00 };
assign _2512_ = _1543_ == { _0170_[11:8], 3'h0, _0170_[4], 1'h0, _0170_[2], 2'h0 };
assign _2513_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 6'h00, _0170_[1], 1'h0 };
assign _2514_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 4'h0, _0170_[3], 1'h0, _0170_[1:0] };
assign _2515_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 4'h0, _0170_[3:2], 2'h0 };
assign _2516_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 4'h0, _0170_[3:2], 1'h0, _0170_[0] };
assign _2517_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 4'h0, _0170_[3:1], 1'h0 };
assign _2518_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 4'h0, _0170_[3:0] };
assign _2519_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 3'h0, _0170_[4], 4'h0 };
assign _2520_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 3'h0, _0170_[4], 3'h0, _0170_[0] };
assign _2521_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 3'h0, _0170_[4], 2'h0, _0170_[1], 1'h0 };
assign _2522_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 3'h0, _0170_[4], 2'h0, _0170_[1:0] };
assign _2523_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 3'h0, _0170_[4], 1'h0, _0170_[2], 2'h0 };
assign _2524_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 6'h00, _0170_[1:0] };
assign _2525_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 3'h0, _0170_[4], 1'h0, _0170_[2], 1'h0, _0170_[0] };
assign _2526_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 3'h0, _0170_[4], 1'h0, _0170_[2:1], 1'h0 };
assign _2527_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 3'h0, _0170_[4], 1'h0, _0170_[2:0] };
assign _2528_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 3'h0, _0170_[4:3], 3'h0 };
assign _2529_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 3'h0, _0170_[4:3], 2'h0, _0170_[0] };
assign _2530_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 3'h0, _0170_[4:3], 1'h0, _0170_[1], 1'h0 };
assign _2531_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 3'h0, _0170_[4:3], 1'h0, _0170_[1:0] };
assign _2532_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 3'h0, _0170_[4:2], 2'h0 };
assign _2533_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 3'h0, _0170_[4:2], 1'h0, _0170_[0] };
assign _2534_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 3'h0, _0170_[4:1], 1'h0 };
assign _2535_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 5'h00, _0170_[2], 2'h0 };
assign _2536_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 3'h0, _0170_[4:0] };
assign _2537_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 5'h00, _0170_[2], 1'h0, _0170_[0] };
assign _2538_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 5'h00, _0170_[2:1], 1'h0 };
assign _2539_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 5'h00, _0170_[2:0] };
assign _2540_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 4'h0, _0170_[3], 3'h0 };
assign _2541_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 4'h0, _0170_[3], 2'h0, _0170_[0] };
assign _2542_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 4'h0, _0170_[3], 1'h0, _0170_[1], 1'h0 };
assign _2543_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5], 3'h0, _0170_[1:0] };
assign _2544_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5], 2'h0, _0170_[2], 2'h0 };
assign _2545_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5], 1'h0, _0170_[3:2], 1'h0, _0170_[0] };
assign _2546_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5], 1'h0, _0170_[3:1], 1'h0 };
assign _2547_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5], 1'h0, _0170_[3:0] };
assign _2548_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5:4], 4'h0 };
assign _2549_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5:4], 3'h0, _0170_[0] };
assign _2550_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5:4], 2'h0, _0170_[1], 1'h0 };
assign _2551_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5:4], 2'h0, _0170_[1:0] };
assign _2552_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5:4], 1'h0, _0170_[2], 2'h0 };
assign _2553_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5:4], 1'h0, _0170_[2], 1'h0, _0170_[0] };
assign _2554_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5:4], 1'h0, _0170_[2:1], 1'h0 };
assign _2555_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5], 2'h0, _0170_[2], 1'h0, _0170_[0] };
assign _2556_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5:4], 1'h0, _0170_[2:0] };
assign _2557_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5:3], 3'h0 };
assign _2558_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5:3], 2'h0, _0170_[0] };
assign _2559_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5:3], 1'h0, _0170_[1], 1'h0 };
assign _2560_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5:3], 1'h0, _0170_[1:0] };
assign _2561_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5:2], 2'h0 };
assign _2562_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5:2], 1'h0, _0170_[0] };
assign _2563_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5:1], 1'h0 };
assign _2564_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5:0] };
assign _2565_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5], 2'h0, _0170_[2:1], 1'h0 };
assign _2566_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5], 2'h0, _0170_[2:0] };
assign _2567_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5], 1'h0, _0170_[3], 3'h0 };
assign _2568_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5], 1'h0, _0170_[3], 2'h0, _0170_[0] };
assign _2569_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5], 1'h0, _0170_[3], 1'h0, _0170_[1], 1'h0 };
assign _2570_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5], 1'h0, _0170_[3], 1'h0, _0170_[1:0] };
assign _2571_ = _1543_ == { 2'h0, _0170_[9:8], 2'h0, _0170_[5], 1'h0, _0170_[3:2], 2'h0 };
assign _2572_ = _1543_ == { 1'h0, _0170_[10:6], 5'h00, _0170_[0] };
assign _2573_ = _1543_ == { 1'h0, _0170_[10:6], 6'h00 };
assign _2574_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 7'h00 };
assign _2575_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 5'h00, _0170_[1], 1'h0 };
assign _2576_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 3'h0, _0170_[3], 1'h0, _0170_[1:0] };
assign _2577_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 3'h0, _0170_[3:2], 2'h0 };
assign _2578_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 3'h0, _0170_[3:2], 1'h0, _0170_[0] };
assign _2579_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 3'h0, _0170_[3:1], 1'h0 };
assign _2580_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 3'h0, _0170_[3:0] };
assign _2581_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 2'h0, _0170_[4], 4'h0 };
assign _2582_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 2'h0, _0170_[4], 3'h0, _0170_[0] };
assign _2583_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 2'h0, _0170_[4], 2'h0, _0170_[1], 1'h0 };
assign _2584_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 2'h0, _0170_[4], 2'h0, _0170_[1:0] };
assign _2585_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 2'h0, _0170_[4], 1'h0, _0170_[2], 2'h0 };
assign _2586_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 5'h00, _0170_[1:0] };
assign _2587_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 2'h0, _0170_[4], 1'h0, _0170_[2], 1'h0, _0170_[0] };
assign _2588_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 2'h0, _0170_[4], 1'h0, _0170_[2:1], 1'h0 };
assign _2589_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 2'h0, _0170_[4], 1'h0, _0170_[2:0] };
assign _2590_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 2'h0, _0170_[4:3], 3'h0 };
assign _2591_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 2'h0, _0170_[4:3], 2'h0, _0170_[0] };
assign _2592_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 2'h0, _0170_[4:3], 1'h0, _0170_[1], 1'h0 };
assign _2593_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 2'h0, _0170_[4:3], 1'h0, _0170_[1:0] };
assign _2594_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 2'h0, _0170_[4:2], 2'h0 };
assign _2595_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 2'h0, _0170_[4:2], 1'h0, _0170_[0] };
assign _2596_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 2'h0, _0170_[4:1], 1'h0 };
assign _2597_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 4'h0, _0170_[2], 2'h0 };
assign _2598_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 2'h0, _0170_[4:0] };
assign _2599_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 4'h0, _0170_[2], 1'h0, _0170_[0] };
assign _2600_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 4'h0, _0170_[2:1], 1'h0 };
assign _2601_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 4'h0, _0170_[2:0] };
assign _2602_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 3'h0, _0170_[3], 3'h0 };
assign _2603_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 3'h0, _0170_[3], 2'h0, _0170_[0] };
assign _2604_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:7], 3'h0, _0170_[3], 1'h0, _0170_[1], 1'h0 };
assign _2605_ = _1543_ == { _0170_[11], 1'h0, _0170_[9:8], 8'h00 };
assign _2606_ = _1543_ == { 2'h0, _0170_[9:8], 5'h00, _0170_[2:1], 1'h0 };
assign _2607_ = _1543_ == { 2'h0, _0170_[9:8], 4'h0, _0170_[3], 1'h0, _0170_[1], 1'h0 };
assign _2608_ = _1543_ == { 2'h0, _0170_[9:8], 3'h0, _0170_[4:3], 1'h0, _0170_[1], 1'h0 };
assign _2609_ = _1543_ == { 2'h0, _0170_[9:8], 3'h0, _0170_[4], 4'h0 };
assign _2610_ = _1543_ == { _0170_[11:8], 3'h0, _0170_[4], 1'h0, _0170_[2], 1'h0, _0170_[0] };
assign _2611_ = _1543_ == { _0170_[11:8], 3'h0, _0170_[4], 2'h0, _0170_[1:0] };
assign _2612_ = _1543_ == { _0170_[11:8], 3'h0, _0170_[4], 3'h0, _0170_[0] };
assign _3021_ = _2437_ & _0156_;
assign _3063_ = _2438_ & _0157_;
assign _3065_ = _2439_ & _0157_;
assign _3081_ = _2440_ & _0158_;
assign _3085_ = _2441_ & _0159_;
assign _3089_ = _2442_ & _0160_;
assign _3067_ = _2443_ & _0161_;
assign _3069_ = _2444_ & _0161_;
assign _3071_ = _2445_ & _0161_;
assign _0050_ = _2446_ & _0162_;
assign _2670_[2] = _2447_ & _0162_;
assign _3257_ = _2448_ & _0162_;
assign _3194_ = _2449_ & _0163_;
assign _3196_ = _2450_ & _0163_;
assign _3198_ = _2451_ & _0163_;
assign _3200_ = _2452_ & _0163_;
assign _3202_ = _2453_ & _0163_;
assign _3204_ = _2454_ & _0163_;
assign _3206_ = _2455_ & _0163_;
assign _3208_ = _2456_ & _0163_;
assign _3210_ = _2457_ & _0163_;
assign _3212_ = _2458_ & _0163_;
assign _3214_ = _2459_ & _0163_;
assign _3216_ = _2460_ & _0163_;
assign _3218_ = _2461_ & _0163_;
assign _3220_ = _2462_ & _0163_;
assign _3222_ = _2463_ & _0163_;
assign _3224_ = _2464_ & _0163_;
assign _3226_ = _2465_ & _0163_;
assign _3228_ = _2466_ & _0163_;
assign _3230_ = _2467_ & _0163_;
assign _3232_ = _2468_ & _0163_;
assign _3234_ = _2469_ & _0163_;
assign _3236_ = _2470_ & _0163_;
assign _3238_ = _2471_ & _0163_;
assign _3240_ = _2472_ & _0163_;
assign _3242_ = _2473_ & _0163_;
assign _3244_ = _2474_ & _0163_;
assign _3246_ = _2475_ & _0163_;
assign _3248_ = _2476_ & _0163_;
assign _3250_ = _2477_ & _0163_;
assign _3252_ = _2478_ & _0163_;
assign _3254_ = _2479_ & _0163_;
assign _0042_ = _2480_ & _0162_;
assign _0040_ = _2481_ & _0162_;
assign _0036_ = _2482_ & _0162_;
assign _0032_ = _2483_ & _0162_;
assign _3023_ = _2484_ & _0162_;
assign _3025_ = _2485_ & _0162_;
assign _3027_ = _2486_ & _0162_;
assign _3029_ = _2487_ & _0162_;
assign _3031_ = _2488_ & _0162_;
assign _3033_ = _2489_ & _0162_;
assign _3035_ = _2490_ & _0162_;
assign _3037_ = _2491_ & _0162_;
assign _3039_ = _2492_ & _0162_;
assign _3041_ = _2493_ & _0162_;
assign _3043_ = _2494_ & _0162_;
assign _3045_ = _2495_ & _0162_;
assign _3047_ = _2496_ & _0162_;
assign _3049_ = _2497_ & _0162_;
assign _3051_ = _2498_ & _0162_;
assign _3053_ = _2499_ & _0162_;
assign _3055_ = _2500_ & _0162_;
assign _3057_ = _2501_ & _0162_;
assign _3059_ = _2502_ & _0162_;
assign _3061_ = _2503_ & _0162_;
assign _3191_ = _2504_ & _0162_;
assign _0072_ = _2505_ & _0162_;
assign _0048_ = _2506_ & _0162_;
assign _0054_ = _2507_ & _0162_;
assign _3176_ = _2508_ & _0162_;
assign _0062_ = _2509_ & _0162_;
assign _0060_ = _2510_ & _0162_;
assign _0068_ = _2511_ & _0162_;
assign _3189_ = _2512_ & _0162_;
assign _3167_[1] = _2513_ & _0162_;
assign _3167_[10] = _2514_ & _0162_;
assign _3167_[11] = _2515_ & _0162_;
assign _3167_[12] = _2516_ & _0162_;
assign _3167_[13] = _2517_ & _0162_;
assign _3167_[14] = _2518_ & _0162_;
assign _3167_[15] = _2519_ & _0162_;
assign _3167_[16] = _2520_ & _0162_;
assign _3167_[17] = _2521_ & _0162_;
assign _3167_[18] = _2522_ & _0162_;
assign _3167_[19] = _2523_ & _0162_;
assign _3167_[2] = _2524_ & _0162_;
assign _3167_[20] = _2525_ & _0162_;
assign _3167_[21] = _2526_ & _0162_;
assign _3167_[22] = _2527_ & _0162_;
assign _3167_[23] = _2528_ & _0162_;
assign _3167_[24] = _2529_ & _0162_;
assign _3167_[25] = _2530_ & _0162_;
assign _3167_[26] = _2531_ & _0162_;
assign _3167_[27] = _2532_ & _0162_;
assign _3167_[28] = _2533_ & _0162_;
assign _3167_[29] = _2534_ & _0162_;
assign _3167_[3] = _2535_ & _0162_;
assign _3167_[30] = _2536_ & _0162_;
assign _3167_[4] = _2537_ & _0162_;
assign _3167_[5] = _2538_ & _0162_;
assign _3167_[6] = _2539_ & _0162_;
assign _3167_[7] = _2540_ & _0162_;
assign _3167_[8] = _2541_ & _0162_;
assign _3167_[9] = _2542_ & _0162_;
assign _3185_[0] = _2543_ & _0162_;
assign _3185_[1] = _2544_ & _0162_;
assign _3185_[10] = _2545_ & _0162_;
assign _3185_[11] = _2546_ & _0162_;
assign _3185_[12] = _2547_ & _0162_;
assign _3185_[13] = _2548_ & _0162_;
assign _3185_[14] = _2549_ & _0162_;
assign _3185_[15] = _2550_ & _0162_;
assign _3185_[16] = _2551_ & _0162_;
assign _3185_[17] = _2552_ & _0162_;
assign _3185_[18] = _2553_ & _0162_;
assign _3185_[19] = _2554_ & _0162_;
assign _3185_[2] = _2555_ & _0162_;
assign _3185_[20] = _2556_ & _0162_;
assign _3185_[21] = _2557_ & _0162_;
assign _3185_[22] = _2558_ & _0162_;
assign _3185_[23] = _2559_ & _0162_;
assign _3185_[24] = _2560_ & _0162_;
assign _3185_[25] = _2561_ & _0162_;
assign _3185_[26] = _2562_ & _0162_;
assign _3185_[27] = _2563_ & _0162_;
assign _3185_[28] = _2564_ & _0162_;
assign _3185_[3] = _2565_ & _0162_;
assign _3185_[4] = _2566_ & _0162_;
assign _3185_[5] = _2567_ & _0162_;
assign _3185_[6] = _2568_ & _0162_;
assign _3185_[7] = _2569_ & _0162_;
assign _3185_[8] = _2570_ & _0162_;
assign _3185_[9] = _2571_ & _0162_;
assign _3073_ = _2572_ & _0162_;
assign _0028_ = _2573_ & _0162_;
assign _3163_[0] = _2574_ & _0162_;
assign _3163_[1] = _2575_ & _0162_;
assign _3163_[10] = _2576_ & _0162_;
assign _3163_[11] = _2577_ & _0162_;
assign _3163_[12] = _2578_ & _0162_;
assign _3163_[13] = _2579_ & _0162_;
assign _3163_[14] = _2580_ & _0162_;
assign _3163_[15] = _2581_ & _0162_;
assign _3163_[16] = _2582_ & _0162_;
assign _3163_[17] = _2583_ & _0162_;
assign _3163_[18] = _2584_ & _0162_;
assign _3163_[19] = _2585_ & _0162_;
assign _3163_[2] = _2586_ & _0162_;
assign _3163_[20] = _2587_ & _0162_;
assign _3163_[21] = _2588_ & _0162_;
assign _3163_[22] = _2589_ & _0162_;
assign _3163_[23] = _2590_ & _0162_;
assign _3163_[24] = _2591_ & _0162_;
assign _3163_[25] = _2592_ & _0162_;
assign _3163_[26] = _2593_ & _0162_;
assign _3163_[27] = _2594_ & _0162_;
assign _3163_[28] = _2595_ & _0162_;
assign _3163_[29] = _2596_ & _0162_;
assign _3163_[3] = _2597_ & _0162_;
assign _3163_[30] = _2598_ & _0162_;
assign _3163_[4] = _2599_ & _0162_;
assign _3163_[5] = _2600_ & _0162_;
assign _3163_[6] = _2601_ & _0162_;
assign _3163_[7] = _2602_ & _0162_;
assign _3163_[8] = _2603_ & _0162_;
assign _3163_[9] = _2604_ & _0162_;
assign _3167_[0] = _2605_ & _0162_;
assign _3259_ = _2606_ & _0162_;
assign _3261_[0] = _2607_ & _0162_;
assign _3261_[1] = _2608_ & _0162_;
assign _3263_ = _2609_ & _0162_;
assign _3265_ = _2610_ & _0162_;
assign _3267_ = _2611_ & _0162_;
assign _3269_ = _2612_ & _0162_;
/* src = "generated/sv2v_out.v:14234.2-14238.29" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers  */
/* PC_TAINT_INFO STATE_NAME priv_mode_id_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) priv_mode_id_o <= 2'h3;
else if (_0452_) priv_mode_id_o <= priv_lvl_d;
reg [1:0] _3710_;
/* src = "generated/sv2v_out.v:14696.2-14700.39" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c15e0aa98717c0c04f1cca2ff0d3e7c6727de751\ibex_cs_registers  */
/* PC_TAINT_INFO STATE_NAME _3710_ */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) _3710_ <= 2'h0;
else if (mcountinhibit_we) _3710_ <= { dummy_instr_seed_o[2], dummy_instr_seed_o[0] };
assign { mcountinhibit[2], mcountinhibit[0] } = _3710_;
assign _0450_ = { _1165_, _1167_ } > { _1965_, _1967_ };
assign _0451_ = { _1964_, _1966_ } > { _1166_, _1168_ };
assign illegal_csr_priv_t0 = _0450_ ^ _0451_;
assign _0172_ = ~ csr_addr_i_t0[8];
assign _0173_ = ~ csr_addr_i_t0[9];
assign _0174_ = ~ priv_mode_id_o_t0[0];
assign _0175_ = ~ priv_mode_id_o_t0[1];
assign _1165_ = csr_addr_i[9] & _0173_;
assign _1166_ = priv_mode_id_o[1] & _0175_;
assign _1964_ = csr_addr_i[9] | csr_addr_i_t0[9];
assign _1965_ = priv_mode_id_o[1] | priv_mode_id_o_t0[1];
assign _1167_ = csr_addr_i[8] & _0172_;
assign _1168_ = priv_mode_id_o[0] & _0174_;
assign _1966_ = csr_addr_i[8] | csr_addr_i_t0[8];
assign _1967_ = priv_mode_id_o[0] | priv_mode_id_o_t0[0];
assign _1169_ = _3021_ & csr_wr;
assign _1172_ = _3081_ & _3082_;
assign _1175_ = _3085_ & _3086_;
assign _1178_ = csr_we_int_t0 & _3072_;
assign _1170_ = csr_wr_t0 & _3020_;
assign _1173_ = _3083_ & _3080_;
assign _1176_ = _3087_ & _3084_;
assign _1179_ = _3073_ & csr_we_int;
assign _1171_ = _3021_ & csr_wr_t0;
assign _1174_ = _3081_ & _3083_;
assign _1177_ = _3085_ & _3087_;
assign _1180_ = csr_we_int_t0 & _3073_;
assign _1968_ = _1169_ | _1170_;
assign _1969_ = _1172_ | _1173_;
assign _1970_ = _1175_ | _1176_;
assign _1971_ = _1178_ | _1179_;
assign illegal_csr_write_t0 = _1968_ | _1171_;
assign _3075_ = _1969_ | _1174_;
assign _3077_ = _1970_ | _1177_;
assign dummy_instr_seed_en_o_t0 = _1971_ | _1180_;
assign _0176_ = | { csr_save_cause_i_t0, csr_restore_mret_i_t0, csr_restore_dret_i_t0 };
assign _0177_ = | { _0060_, _0062_, _0054_, _0048_, _0072_, _0032_, _0036_, _0040_, _0042_, _0050_, _0028_, _0068_, _2670_[2], _3269_, _3267_, _3265_, _3263_, _3261_, _3259_, _3257_, _3191_, _3189_, _3185_, _3176_, _3167_, _3163_, _3073_, _3061_, _3059_, _3057_, _3055_, _3053_, _3051_, _3049_, _3047_, _3045_, _3043_, _3041_, _3039_, _3037_, _3035_, _3033_, _3031_, _3029_, _3027_, _3025_, _3023_ };
assign _0178_ = | { _0032_, _0036_, _0040_, _0042_ };
assign _0179_ = | { _3071_, _3111_ };
assign _0180_ = | { _3254_, _3250_, _3248_, _3246_, _3244_, _3242_, _3240_, _3238_, _3236_, _3234_, _3232_, _3230_, _3228_, _3226_, _3224_, _3222_, _3220_, _3218_, _3216_, _3214_, _3212_, _3210_, _3208_, _3206_, _3204_, _3202_, _3200_, _3198_, _3196_, _3194_ };
assign _0181_ = | { _0032_, _0036_, _1561_, _1559_, _3191_, _3185_, _3167_ };
assign _0182_ = | { _1559_, _3185_, _3167_ };
assign _0183_ = | { _0032_, _0036_, _0040_, _1567_, _1559_, _3185_, _3167_ };
assign _0184_ = | { _0062_, _1575_, _3176_ };
assign _0185_ = | { _0072_, _0032_, _0042_, _1573_, _1571_, _3185_ };
assign _0186_ = | { _0032_, _0042_, _1573_, _1571_, _3191_, _3185_ };
assign _0187_ = | { _3185_, _3167_, _3163_ };
assign _0188_ = | { _0054_, _0048_, _0072_ };
assign _0189_ = | { _0032_, _0036_, _1561_, _3185_, _3167_, _3163_ };
assign _0190_ = | { _0042_, _1571_, _3185_ };
assign _0191_ = | { _0054_, _1563_, _3176_ };
assign _0192_ = | { _0032_, _0036_, _1561_, _1559_, _3185_, _3167_ };
assign _0158_ = | dummy_instr_seed_o_t0[12:11];
assign _0159_ = | dummy_instr_seed_o_t0[1:0];
assign _0161_ = | csr_op_i_t0;
assign _0193_ = | _3167_;
assign _0194_ = | _3163_;
assign _0195_ = | _3185_;
assign _0163_ = | csr_addr_i_t0[4:0];
assign _0196_ = | { _3061_, _3059_, _3057_, _3055_, _3053_, _3051_, _3049_, _3047_, _3045_, _3043_, _3041_, _3039_, _3037_, _3035_, _3033_, _3031_, _3029_, _3027_, _3025_, _3023_ };
assign _0197_ = | { _3069_, _3067_, _3071_ };
assign _0198_ = | irqs_o_t0;
assign _0199_ = ~ { csr_save_cause_i_t0, csr_restore_dret_i_t0, csr_restore_mret_i_t0 };
assign _0200_ = ~ { _3269_, _3267_, _3265_, _3263_, _3261_, _3259_, _3257_, _2670_[2], _3191_, _3189_, _3185_, _0060_, _0062_, _0054_, _0048_, _0072_, _3176_, _0036_, _0040_, _0042_, _0050_, _0028_, _3167_, _3163_, _0068_, _0032_, _3073_, _3061_, _3059_, _3057_, _3055_, _3053_, _3051_, _3049_, _3047_, _3045_, _3043_, _3041_, _3039_, _3037_, _3035_, _3033_, _3031_, _3029_, _3027_, _3025_, _3023_ };
assign _0201_ = ~ { _0036_, _0040_, _0042_, _0032_ };
assign _0202_ = ~ { _3071_, _3111_ };
assign _0203_ = ~ { _3254_, _3250_, _3248_, _3246_, _3244_, _3242_, _3240_, _3238_, _3236_, _3234_, _3232_, _3230_, _3228_, _3226_, _3224_, _3222_, _3220_, _3218_, _3216_, _3214_, _3212_, _3210_, _3208_, _3206_, _3204_, _3202_, _3200_, _3198_, _3196_, _3194_ };
assign _0204_ = ~ { _1559_, _1561_, _3191_, _3185_, _0036_, _3167_, _0032_ };
assign _0205_ = ~ { _1559_, _3185_, _3167_ };
assign _0206_ = ~ { _1559_, _1567_, _3185_, _0036_, _0040_, _3167_, _0032_ };
assign _0207_ = ~ { _0062_, _3176_, _1575_ };
assign _0208_ = ~ { _1571_, _1573_, _3185_, _0072_, _0042_, _0032_ };
assign _0209_ = ~ { _1571_, _1573_, _3191_, _3185_, _0042_, _0032_ };
assign _0210_ = ~ { _3185_, _3167_, _3163_ };
assign _0211_ = ~ { _0054_, _0048_, _0072_ };
assign _0212_ = ~ { _1561_, _3185_, _0036_, _3167_, _3163_, _0032_ };
assign _0213_ = ~ { _1571_, _3185_, _0042_ };
assign _0214_ = ~ { _1563_, _0054_, _3176_ };
assign _0215_ = ~ { _1559_, _1561_, _3185_, _0036_, _3167_, _0032_ };
assign _0166_ = ~ dummy_instr_seed_o_t0[12:11];
assign _0167_ = ~ dummy_instr_seed_o_t0[1:0];
assign _0169_ = ~ csr_op_i_t0;
assign _0216_ = ~ _3167_;
assign _0217_ = ~ _3163_;
assign _0218_ = ~ _3185_;
assign _0171_ = ~ csr_addr_i_t0[4:0];
assign _0219_ = ~ { _3061_, _3059_, _3057_, _3055_, _3053_, _3051_, _3049_, _3047_, _3045_, _3043_, _3041_, _3039_, _3037_, _3035_, _3033_, _3031_, _3029_, _3027_, _3025_, _3023_ };
assign _0220_ = ~ { _3071_, _3069_, _3067_ };
assign _0221_ = ~ irqs_o_t0;
assign _0493_ = { csr_save_cause_i, csr_restore_dret_i, csr_restore_mret_i } & _0199_;
assign _0494_ = { _3268_, _3266_, _3264_, _3262_, _3260_, _3258_, _3256_, _3192_, _3190_, _3188_, _3184_, _3181_, _3180_, _3179_, _3178_, _3177_, _3175_, _3174_, _3173_, _3172_, _3171_, _3170_, _3166_, _3162_, _3161_, _3160_, _3072_, _3060_, _3058_, _3056_, _3054_, _3052_, _3050_, _3048_, _3046_, _3044_, _3042_, _3040_, _3038_, _3036_, _3034_, _3032_, _3030_, _3028_, _3026_, _3024_, _3022_ } & _0200_;
assign _0495_ = { _3174_, _3173_, _3172_, _3160_ } & _0201_;
assign _0496_ = { _3070_, _3110_ } & _0202_;
assign _0497_ = { _3253_, _3249_, _3247_, _3245_, _3243_, _3241_, _3239_, _3237_, _3235_, _3233_, _3231_, _3229_, _3227_, _3225_, _3223_, _3221_, _3219_, _3217_, _3215_, _3213_, _3211_, _3209_, _3207_, _3205_, _3203_, _3201_, _3199_, _3197_, _3195_, _3193_ } & _0203_;
assign _0534_ = { _1558_, _1560_, _3190_, _3184_, _3174_, _3166_, _3160_ } & _0204_;
assign _0535_ = { _1558_, _3184_, _3166_ } & _0205_;
assign _0536_ = { _1558_, _1566_, _3184_, _3174_, _3173_, _3166_, _3160_ } & _0206_;
assign _0537_ = { _3180_, _3175_, _1574_ } & _0207_;
assign _0538_ = { _1570_, _1572_, _3184_, _3177_, _3172_, _3160_ } & _0208_;
assign _0539_ = { _1570_, _1572_, _3190_, _3184_, _3172_, _3160_ } & _0209_;
assign _0540_ = { _3184_, _3166_, _3162_ } & _0210_;
assign _0541_ = { _3179_, _3178_, _3177_ } & _0211_;
assign _0542_ = { _1560_, _3184_, _3174_, _3166_, _3162_, _3160_ } & _0212_;
assign _0543_ = { _1570_, _3184_, _3172_ } & _0213_;
assign _0544_ = { _1562_, _3179_, _3175_ } & _0214_;
assign _0545_ = { _1558_, _1560_, _3184_, _3174_, _3166_, _3160_ } & _0215_;
assign _1184_ = dummy_instr_seed_o[12:11] & _0166_;
assign _1185_ = dummy_instr_seed_o[1:0] & _0167_;
assign _1210_ = csr_op_i & _0169_;
assign _1488_ = _3166_ & _0216_;
assign _1542_ = _3162_ & _0217_;
assign _1544_ = _3184_ & _0218_;
assign _1545_ = csr_addr_i[4:0] & _0171_;
assign _1546_ = { _3060_, _3058_, _3056_, _3054_, _3052_, _3050_, _3048_, _3046_, _3044_, _3042_, _3040_, _3038_, _3036_, _3034_, _3032_, _3030_, _3028_, _3026_, _3024_, _3022_ } & _0219_;
assign _1547_ = { _3070_, _3068_, _3066_ } & _0220_;
assign _1548_ = irqs_o & _0221_;
assign _0222_ = ! _0493_;
assign _0223_ = ! _0494_;
assign _0224_ = ! _0495_;
assign _0225_ = ! _0496_;
assign _0226_ = ! _0497_;
assign _0227_ = ! _0534_;
assign _0228_ = ! _0535_;
assign _0229_ = ! _0536_;
assign _0230_ = ! _0537_;
assign _0231_ = ! _0538_;
assign _0232_ = ! _0539_;
assign _0233_ = ! _0540_;
assign _0234_ = ! _0541_;
assign _0235_ = ! _0542_;
assign _0236_ = ! _0543_;
assign _0237_ = ! _0544_;
assign _0238_ = ! _0545_;
assign _0239_ = ! _1184_;
assign _0240_ = ! _1185_;
assign _0241_ = ! _1210_;
assign _0242_ = ! _1488_;
assign _0243_ = ! _1542_;
assign _0244_ = ! _1544_;
assign _0245_ = ! _1546_;
assign _0246_ = ! _1547_;
assign _0247_ = ! _1548_;
assign _0453_ = _0222_ & _0176_;
assign _0011_ = _0223_ & _0177_;
assign dbg_csr_t0 = _0224_ & _0178_;
assign _0457_ = _0225_ & _0179_;
assign _0459_ = _0226_ & _0180_;
assign _0430_ = _0227_ & _0181_;
assign _0426_ = _0228_ & _0182_;
assign _0432_ = _0229_ & _0183_;
assign _0442_ = _0230_ & _0184_;
assign _0444_ = _0231_ & _0185_;
assign _0440_ = _0232_ & _0186_;
assign _0434_ = _0233_ & _0187_;
assign _0446_ = _0234_ & _0188_;
assign _0436_ = _0235_ & _0189_;
assign _0438_ = _0236_ & _0190_;
assign _0428_ = _0237_ & _0191_;
assign _0448_ = _0238_ & _0192_;
assign _3083_ = _0239_ & _0158_;
assign _3087_ = _0240_ & _0159_;
assign _3111_ = _0241_ & _0161_;
assign _3169_ = _0242_ & _0193_;
assign _3165_ = _0243_ & _0194_;
assign _3187_ = _0244_ & _0195_;
assign _3183_ = _0245_ & _0196_;
assign csr_wr_t0 = _0246_ & _0197_;
assign irq_pending_o_t0 = _0247_ & _0198_;
assign _0248_ = ~ csr_mcause_i[5];
assign _0249_ = ~ csr_mcause_i[6];
assign _1181_ = csr_mcause_i_t0[5] & _0249_;
assign _1182_ = csr_mcause_i_t0[6] & _0248_;
assign _1183_ = csr_mcause_i_t0[5] & csr_mcause_i_t0[6];
assign _1972_ = _1181_ | _1182_;
assign _3079_ = _1972_ | _1183_;
assign _0250_ = ~ _3170_;
assign _0251_ = ~ _3168_;
assign _0252_ = ~ _1558_;
assign _0253_ = ~ _3172_;
assign _0254_ = ~ _3160_;
assign _0255_ = ~ _3174_;
assign _0256_ = ~ _1560_;
assign _0257_ = ~ _0425_;
assign _0258_ = ~ _3177_;
assign _0259_ = ~ _3179_;
assign _0260_ = ~ _1562_;
assign _0261_ = ~ _3180_;
assign _0262_ = ~ _3188_;
assign _0263_ = ~ _3161_;
assign _0264_ = ~ _1564_;
assign _0265_ = ~ _0427_;
assign _0266_ = ~ _0429_;
assign _0267_ = ~ { _3170_, _3170_, _3170_ };
assign _0268_ = ~ { _1558_, _1558_, _1558_ };
assign _0269_ = ~ { _3171_, _3171_, _3171_ };
assign _0270_ = ~ { _3174_, _3174_, _3174_ };
assign _0271_ = ~ { _3173_, _3173_, _3173_ };
assign _0272_ = ~ { _1566_, _1566_, _1566_ };
assign _0273_ = ~ { _0425_, _0425_, _0425_ };
assign _0274_ = ~ { _3177_, _3177_, _3177_ };
assign _0275_ = ~ { _3179_, _3179_, _3179_ };
assign _0276_ = ~ { _1562_, _1562_, _1562_ };
assign _0277_ = ~ { _3180_, _3180_, _3180_ };
assign _0278_ = ~ { _3188_, _3188_, _3188_ };
assign _0279_ = ~ { _1568_, _1568_, _1568_ };
assign _0280_ = ~ { _0427_, _0427_, _0427_ };
assign _0281_ = ~ { _0431_, _0431_, _0431_ };
assign _0282_ = ~ { _3164_, _3164_, _3164_ };
assign _0283_ = ~ { _3172_, _3172_, _3172_ };
assign _0284_ = ~ { _1560_, _1560_, _1560_ };
assign _0285_ = ~ { _0433_, _0433_, _0433_ };
assign _0286_ = ~ { _0435_, _0435_, _0435_ };
assign _0287_ = ~ { _3186_, _3186_, _3186_ };
assign _0288_ = ~ { _1570_, _1570_, _1570_ };
assign _0289_ = ~ { _3160_, _3160_, _3160_ };
assign _0290_ = ~ { _1572_, _1572_, _1572_ };
assign _0291_ = ~ { _0437_, _0437_, _0437_ };
assign _0292_ = ~ { _3256_, _3256_, _3256_ };
assign _0293_ = ~ { _1564_, _1564_, _1564_ };
assign _0294_ = ~ { _0439_, _0439_, _0439_ };
assign _0295_ = ~ _3164_;
assign _0296_ = ~ _3186_;
assign _0297_ = ~ _1570_;
assign _0298_ = ~ _3173_;
assign _0299_ = ~ _1572_;
assign _0300_ = ~ _0437_;
assign _0301_ = ~ _3178_;
assign _0302_ = ~ _3175_;
assign _0303_ = ~ _1574_;
assign _0304_ = ~ _3256_;
assign _0305_ = ~ _1576_;
assign _0306_ = ~ _0441_;
assign _0307_ = ~ _0443_;
assign _0308_ = ~ _0439_;
assign _0309_ = ~ { _3178_, _3178_, _3178_ };
assign _0310_ = ~ { _3175_, _3175_, _3175_ };
assign _0311_ = ~ { _1578_, _1578_, _1578_ };
assign _0312_ = ~ { _0445_, _0445_, _0445_ };
assign _0313_ = ~ { _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_ };
assign _0314_ = ~ { _3186_, _3186_, _3186_, _3186_, _3186_, _3186_, _3186_, _3186_, _3186_ };
assign _0315_ = ~ { _1570_, _1570_, _1570_, _1570_, _1570_, _1570_, _1570_, _1570_, _1570_ };
assign _0316_ = ~ { _3173_, _3173_, _3173_, _3173_, _3173_, _3173_, _3173_, _3173_, _3173_ };
assign _0317_ = ~ { _3160_, _3160_, _3160_, _3160_, _3160_, _3160_, _3160_, _3160_, _3160_ };
assign _0318_ = ~ { _1572_, _1572_, _1572_, _1572_, _1572_, _1572_, _1572_, _1572_, _1572_ };
assign _0319_ = ~ { _0437_, _0437_, _0437_, _0437_, _0437_, _0437_, _0437_, _0437_, _0437_ };
assign _0320_ = ~ { _3177_, _3177_, _3177_, _3177_, _3177_, _3177_, _3177_, _3177_, _3177_ };
assign _0321_ = ~ { _3179_, _3179_, _3179_, _3179_, _3179_, _3179_, _3179_, _3179_, _3179_ };
assign _0322_ = ~ { _1562_, _1562_, _1562_, _1562_, _1562_, _1562_, _1562_, _1562_, _1562_ };
assign _0323_ = ~ { _3180_, _3180_, _3180_, _3180_, _3180_, _3180_, _3180_, _3180_, _3180_ };
assign _0324_ = ~ { _3256_, _3256_, _3256_, _3256_, _3256_, _3256_, _3256_, _3256_, _3256_ };
assign _0325_ = ~ { _1564_, _1564_, _1564_, _1564_, _1564_, _1564_, _1564_, _1564_, _1564_ };
assign _0326_ = ~ { _0427_, _0427_, _0427_, _0427_, _0427_, _0427_, _0427_, _0427_, _0427_ };
assign _0327_ = ~ { _0439_, _0439_, _0439_, _0439_, _0439_, _0439_, _0439_, _0439_, _0439_ };
assign _0328_ = ~ { _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_ };
assign _0329_ = ~ { _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_ };
assign _0330_ = ~ { _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_ };
assign _0331_ = ~ { _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_ };
assign _0332_ = ~ _0433_;
assign _0333_ = ~ _1578_;
assign _0334_ = ~ _0445_;
assign _0335_ = ~ _0435_;
assign _0336_ = ~ { _2152_, _2152_, _2152_ };
assign _0337_ = ~ { _0447_, _0447_, _0447_ };
assign _0338_ = ~ csr_save_cause_i;
assign _0339_ = ~ nmi_mode_i;
assign _0340_ = ~ { nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i };
assign _0341_ = ~ _3088_;
assign _0342_ = ~ { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
assign _0343_ = ~ { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
assign _0344_ = ~ { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
assign _0345_ = ~ csr_restore_mret_i;
assign _0346_ = ~ csr_restore_dret_i;
assign _0347_ = ~ cpuctrlsts_part_q[6];
assign _0348_ = ~ _3078_;
assign _0349_ = ~ debug_mode_i;
assign _0350_ = ~ { debug_mode_i, debug_mode_i };
assign _0351_ = ~ { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i };
assign _0352_ = ~ { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i };
assign _0353_ = ~ debug_csr_save_i;
assign _0354_ = ~ { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
assign _0355_ = ~ { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
assign _0356_ = ~ { debug_csr_save_i, debug_csr_save_i };
assign _0357_ = ~ { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
assign _0358_ = ~ { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
assign _0359_ = ~ { csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i };
assign _0360_ = ~ { csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i };
assign _0361_ = ~ { csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i };
assign _0362_ = ~ { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
assign _0363_ = ~ { csr_save_cause_i, csr_save_cause_i };
assign _0364_ = ~ { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
assign _0365_ = ~ { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
assign _0366_ = ~ { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
assign _0367_ = ~ { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
assign _0368_ = ~ { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
assign _0369_ = ~ { nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i };
assign _0370_ = ~ { csr_restore_dret_i, csr_restore_dret_i };
assign _0371_ = ~ { _3160_, _3160_, _3160_, _3160_ };
assign _0372_ = ~ { _3161_, _3161_ };
assign _0373_ = ~ { _3160_, _3160_, _3160_, _3160_, _3160_, _3160_, _3160_, _3160_, _3160_, _3160_, _3160_, _3160_ };
assign _0374_ = ~ { _3160_, _3160_ };
assign _0375_ = ~ { _3076_, _3076_ };
assign _0376_ = ~ { _3074_, _3074_ };
assign _0377_ = ~ { _3170_, _3170_, _3170_, _3170_, _3170_, _3170_, _3170_, _3170_ };
assign _0378_ = ~ _3171_;
assign _0379_ = ~ _3181_;
assign _0380_ = ~ csr_we_int;
assign _0381_ = ~ { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int };
assign _0382_ = ~ { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int };
assign _0383_ = ~ { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int };
assign _0384_ = ~ _3182_;
assign _0385_ = ~ { csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i };
assign _0386_ = ~ { mstatus_q[1], mstatus_q[1] };
assign _0387_ = ~ { _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_ };
assign _1609_ = _0028_ | _0250_;
assign _1613_ = _1559_ | _0252_;
assign _1616_ = _0042_ | _0253_;
assign _1619_ = _0032_ | _0254_;
assign _1622_ = _0036_ | _0255_;
assign _1625_ = _1561_ | _0256_;
assign _1628_ = _0426_ | _0257_;
assign _1631_ = _0072_ | _0258_;
assign _1634_ = _0054_ | _0259_;
assign _1637_ = _1563_ | _0260_;
assign _1640_ = _0062_ | _0261_;
assign _1644_ = _0068_ | _0263_;
assign _1647_ = _1565_ | _0264_;
assign _1650_ = _0428_ | _0265_;
assign _1653_ = _0430_ | _0266_;
assign _1656_ = { _0028_, _0028_, _0028_ } | _0267_;
assign _1660_ = { _1559_, _1559_, _1559_ } | _0268_;
assign _1663_ = { _0050_, _0050_, _0050_ } | _0269_;
assign _1666_ = { _0036_, _0036_, _0036_ } | _0270_;
assign _1669_ = { _0040_, _0040_, _0040_ } | _0271_;
assign _1672_ = { _1567_, _1567_, _1567_ } | _0272_;
assign _1675_ = { _0426_, _0426_, _0426_ } | _0273_;
assign _1678_ = { _0072_, _0072_, _0072_ } | _0274_;
assign _1681_ = { _0054_, _0054_, _0054_ } | _0275_;
assign _1684_ = { _1563_, _1563_, _1563_ } | _0276_;
assign _1687_ = { _0062_, _0062_, _0062_ } | _0277_;
assign _1689_ = { _3189_, _3189_, _3189_ } | _0278_;
assign _1692_ = { _1569_, _1569_, _1569_ } | _0279_;
assign _1695_ = { _0428_, _0428_, _0428_ } | _0280_;
assign _1698_ = { _0432_, _0432_, _0432_ } | _0281_;
assign _1701_ = { _3165_, _3165_, _3165_ } | _0282_;
assign _1704_ = { _0042_, _0042_, _0042_ } | _0283_;
assign _1708_ = { _1561_, _1561_, _1561_ } | _0284_;
assign _1711_ = { _0434_, _0434_, _0434_ } | _0285_;
assign _1719_ = { _0436_, _0436_, _0436_ } | _0286_;
assign _1723_ = { _3187_, _3187_, _3187_ } | _0287_;
assign _1724_ = { _1571_, _1571_, _1571_ } | _0288_;
assign _1728_ = { _0032_, _0032_, _0032_ } | _0289_;
assign _1731_ = { _1573_, _1573_, _1573_ } | _0290_;
assign _1734_ = { _0438_, _0438_, _0438_ } | _0291_;
assign _1741_ = { _3257_, _3257_, _3257_ } | _0292_;
assign _1742_ = { _1565_, _1565_, _1565_ } | _0293_;
assign _1746_ = { _0440_, _0440_, _0440_ } | _0294_;
assign _1749_ = _3165_ | _0295_;
assign _1752_ = _3187_ | _0296_;
assign _1753_ = _1571_ | _0297_;
assign _1756_ = _0040_ | _0298_;
assign _1760_ = _1573_ | _0299_;
assign _1763_ = _0438_ | _0300_;
assign _1766_ = _0048_ | _0301_;
assign _1769_ = _3176_ | _0302_;
assign _1772_ = _1575_ | _0303_;
assign _1775_ = _3257_ | _0304_;
assign _1776_ = _1577_ | _0305_;
assign _1779_ = _0442_ | _0306_;
assign _1782_ = _0444_ | _0307_;
assign _1798_ = _0440_ | _0308_;
assign _1806_ = { _0048_, _0048_, _0048_ } | _0309_;
assign _1810_ = { _3176_, _3176_, _3176_ } | _0310_;
assign _1813_ = { _1579_, _1579_, _1579_ } | _0311_;
assign _1816_ = { _0446_, _0446_, _0446_ } | _0312_;
assign _1833_ = { _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_ } | _0313_;
assign _1836_ = { _3187_, _3187_, _3187_, _3187_, _3187_, _3187_, _3187_, _3187_, _3187_ } | _0314_;
assign _1837_ = { _1571_, _1571_, _1571_, _1571_, _1571_, _1571_, _1571_, _1571_, _1571_ } | _0315_;
assign _1840_ = { _0040_, _0040_, _0040_, _0040_, _0040_, _0040_, _0040_, _0040_, _0040_ } | _0316_;
assign _1843_ = { _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_ } | _0317_;
assign _1846_ = { _1573_, _1573_, _1573_, _1573_, _1573_, _1573_, _1573_, _1573_, _1573_ } | _0318_;
assign _1849_ = { _0438_, _0438_, _0438_, _0438_, _0438_, _0438_, _0438_, _0438_, _0438_ } | _0319_;
assign _1852_ = { _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_ } | _0320_;
assign _1855_ = { _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_ } | _0321_;
assign _1858_ = { _1563_, _1563_, _1563_, _1563_, _1563_, _1563_, _1563_, _1563_, _1563_ } | _0322_;
assign _1861_ = { _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_ } | _0323_;
assign _1865_ = { _3257_, _3257_, _3257_, _3257_, _3257_, _3257_, _3257_, _3257_, _3257_ } | _0324_;
assign _1866_ = { _1565_, _1565_, _1565_, _1565_, _1565_, _1565_, _1565_, _1565_, _1565_ } | _0325_;
assign _1869_ = { _0428_, _0428_, _0428_, _0428_, _0428_, _0428_, _0428_, _0428_, _0428_ } | _0326_;
assign _1872_ = { _0440_, _0440_, _0440_, _0440_, _0440_, _0440_, _0440_, _0440_, _0440_ } | _0327_;
assign _1889_ = { _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_ } | _0328_;
assign _1892_ = { _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_ } | _0329_;
assign _1907_ = { _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_ } | _0330_;
assign _1910_ = { _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_ } | _0331_;
assign _1917_ = _0434_ | _0332_;
assign _1923_ = _1579_ | _0333_;
assign _1926_ = _0446_ | _0334_;
assign _1929_ = _0436_ | _0335_;
assign _1957_ = { _2153_, _2153_, _2153_ } | _0336_;
assign _1961_ = { _0448_, _0448_, _0448_ } | _0337_;
assign _1982_ = csr_save_cause_i_t0 | _0338_;
assign _1985_ = nmi_mode_i_t0 | _0339_;
assign _1987_ = { nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0 } | _0340_;
assign _1991_ = _3089_ | _0341_;
assign _1992_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } | _0342_;
assign _1995_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } | _0343_;
assign _1998_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } | _0344_;
assign _2001_ = csr_restore_mret_i_t0 | _0345_;
assign _2004_ = csr_restore_dret_i_t0 | _0346_;
assign _2011_ = cpuctrlsts_part_q_t0[6] | _0347_;
assign _2012_ = _3079_ | _0348_;
assign _2014_ = debug_mode_i_t0 | _0349_;
assign _2017_ = { debug_mode_i_t0, debug_mode_i_t0 } | _0350_;
assign _2020_ = { debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0 } | _0351_;
assign _2023_ = { debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0 } | _0352_;
assign _2030_ = debug_csr_save_i_t0 | _0353_;
assign _2032_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } | _0354_;
assign _2035_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } | _0355_;
assign _2038_ = { debug_csr_save_i_t0, debug_csr_save_i_t0 } | _0356_;
assign _2046_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } | _0357_;
assign _2052_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } | _0358_;
assign _2055_ = { csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0 } | _0359_;
assign _2058_ = { csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0 } | _0360_;
assign _2061_ = { csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0 } | _0361_;
assign _2069_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } | _0362_;
assign _2074_ = { csr_save_cause_i_t0, csr_save_cause_i_t0 } | _0363_;
assign _2082_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } | _0364_;
assign _2085_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } | _0365_;
assign _2088_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } | _0366_;
assign _2094_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } | _0367_;
assign _2097_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } | _0368_;
assign _2103_ = { nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0 } | _0369_;
assign _2107_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0 } | _0370_;
assign _2110_ = { _0032_, _0032_, _0032_, _0032_ } | _0371_;
assign _2111_ = { _0068_, _0068_ } | _0372_;
assign _2116_ = { _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_ } | _0373_;
assign _2118_ = { _0032_, _0032_ } | _0374_;
assign _2123_ = { _3077_, _3077_ } | _0375_;
assign _2124_ = { _3075_, _3075_ } | _0376_;
assign _2125_ = { _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_ } | _0377_;
assign _2130_ = csr_we_int_t0 | _0380_;
assign _2132_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } | _0381_;
assign _2135_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } | _0382_;
assign _2139_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } | _0383_;
assign _2142_ = _3183_ | _0384_;
assign _2143_ = { csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0 } | _0385_;
assign _2146_ = { mstatus_q_t0[1], mstatus_q_t0[1] } | _0386_;
assign _2149_ = { _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_ } | _0387_;
assign _1610_ = _0028_ | _3170_;
assign _1612_ = _3169_ | _3168_;
assign _1614_ = _1559_ | _1558_;
assign _1617_ = _0042_ | _3172_;
assign _1620_ = _0032_ | _3160_;
assign _1623_ = _0036_ | _3174_;
assign _1626_ = _1561_ | _1560_;
assign _1629_ = _0426_ | _0425_;
assign _1632_ = _0072_ | _3177_;
assign _1635_ = _0054_ | _3179_;
assign _1638_ = _1563_ | _1562_;
assign _1641_ = _0062_ | _3180_;
assign _1643_ = _3189_ | _3188_;
assign _1645_ = _0068_ | _3161_;
assign _1648_ = _1565_ | _1564_;
assign _1651_ = _0428_ | _0427_;
assign _1654_ = _0430_ | _0429_;
assign _1657_ = { _0028_, _0028_, _0028_ } | { _3170_, _3170_, _3170_ };
assign _1659_ = { _3169_, _3169_, _3169_ } | { _3168_, _3168_, _3168_ };
assign _1661_ = { _1559_, _1559_, _1559_ } | { _1558_, _1558_, _1558_ };
assign _1664_ = { _0050_, _0050_, _0050_ } | { _3171_, _3171_, _3171_ };
assign _1667_ = { _0036_, _0036_, _0036_ } | { _3174_, _3174_, _3174_ };
assign _1670_ = { _0040_, _0040_, _0040_ } | { _3173_, _3173_, _3173_ };
assign _1673_ = { _1567_, _1567_, _1567_ } | { _1566_, _1566_, _1566_ };
assign _1676_ = { _0426_, _0426_, _0426_ } | { _0425_, _0425_, _0425_ };
assign _1679_ = { _0072_, _0072_, _0072_ } | { _3177_, _3177_, _3177_ };
assign _1682_ = { _0054_, _0054_, _0054_ } | { _3179_, _3179_, _3179_ };
assign _1685_ = { _1563_, _1563_, _1563_ } | { _1562_, _1562_, _1562_ };
assign _1688_ = { _0062_, _0062_, _0062_ } | { _3180_, _3180_, _3180_ };
assign _1690_ = { _3189_, _3189_, _3189_ } | { _3188_, _3188_, _3188_ };
assign _1693_ = { _1569_, _1569_, _1569_ } | { _1568_, _1568_, _1568_ };
assign _1696_ = { _0428_, _0428_, _0428_ } | { _0427_, _0427_, _0427_ };
assign _1699_ = { _0432_, _0432_, _0432_ } | { _0431_, _0431_, _0431_ };
assign _1702_ = { _3165_, _3165_, _3165_ } | { _3164_, _3164_, _3164_ };
assign _1705_ = { _0042_, _0042_, _0042_ } | { _3172_, _3172_, _3172_ };
assign _1709_ = { _1561_, _1561_, _1561_ } | { _1560_, _1560_, _1560_ };
assign _1712_ = { _0434_, _0434_, _0434_ } | { _0433_, _0433_, _0433_ };
assign _1720_ = { _0436_, _0436_, _0436_ } | { _0435_, _0435_, _0435_ };
assign _1725_ = { _1571_, _1571_, _1571_ } | { _1570_, _1570_, _1570_ };
assign _1729_ = { _0032_, _0032_, _0032_ } | { _3160_, _3160_, _3160_ };
assign _1732_ = { _1573_, _1573_, _1573_ } | { _1572_, _1572_, _1572_ };
assign _1735_ = { _0438_, _0438_, _0438_ } | { _0437_, _0437_, _0437_ };
assign _1743_ = { _1565_, _1565_, _1565_ } | { _1564_, _1564_, _1564_ };
assign _1747_ = { _0440_, _0440_, _0440_ } | { _0439_, _0439_, _0439_ };
assign _1750_ = _3165_ | _3164_;
assign _1754_ = _1571_ | _1570_;
assign _1757_ = _0040_ | _3173_;
assign _1761_ = _1573_ | _1572_;
assign _1764_ = _0438_ | _0437_;
assign _1767_ = _0048_ | _3178_;
assign _1770_ = _3176_ | _3175_;
assign _1773_ = _1575_ | _1574_;
assign _1777_ = _1577_ | _1576_;
assign _1780_ = _0442_ | _0441_;
assign _1783_ = _0444_ | _0443_;
assign _1799_ = _0440_ | _0439_;
assign _1807_ = { _0048_, _0048_, _0048_ } | { _3178_, _3178_, _3178_ };
assign _1811_ = { _3176_, _3176_, _3176_ } | { _3175_, _3175_, _3175_ };
assign _1814_ = { _1579_, _1579_, _1579_ } | { _1578_, _1578_, _1578_ };
assign _1817_ = { _0446_, _0446_, _0446_ } | { _0445_, _0445_, _0445_ };
assign _1834_ = { _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_ } | { _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_ };
assign _1838_ = { _1571_, _1571_, _1571_, _1571_, _1571_, _1571_, _1571_, _1571_, _1571_ } | { _1570_, _1570_, _1570_, _1570_, _1570_, _1570_, _1570_, _1570_, _1570_ };
assign _1841_ = { _0040_, _0040_, _0040_, _0040_, _0040_, _0040_, _0040_, _0040_, _0040_ } | { _3173_, _3173_, _3173_, _3173_, _3173_, _3173_, _3173_, _3173_, _3173_ };
assign _1844_ = { _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_ } | { _3160_, _3160_, _3160_, _3160_, _3160_, _3160_, _3160_, _3160_, _3160_ };
assign _1847_ = { _1573_, _1573_, _1573_, _1573_, _1573_, _1573_, _1573_, _1573_, _1573_ } | { _1572_, _1572_, _1572_, _1572_, _1572_, _1572_, _1572_, _1572_, _1572_ };
assign _1850_ = { _0438_, _0438_, _0438_, _0438_, _0438_, _0438_, _0438_, _0438_, _0438_ } | { _0437_, _0437_, _0437_, _0437_, _0437_, _0437_, _0437_, _0437_, _0437_ };
assign _1853_ = { _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_ } | { _3177_, _3177_, _3177_, _3177_, _3177_, _3177_, _3177_, _3177_, _3177_ };
assign _1856_ = { _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_ } | { _3179_, _3179_, _3179_, _3179_, _3179_, _3179_, _3179_, _3179_, _3179_ };
assign _1859_ = { _1563_, _1563_, _1563_, _1563_, _1563_, _1563_, _1563_, _1563_, _1563_ } | { _1562_, _1562_, _1562_, _1562_, _1562_, _1562_, _1562_, _1562_, _1562_ };
assign _1862_ = { _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_ } | { _3180_, _3180_, _3180_, _3180_, _3180_, _3180_, _3180_, _3180_, _3180_ };
assign _1864_ = { _3189_, _3189_, _3189_, _3189_, _3189_, _3189_, _3189_, _3189_, _3189_ } | { _3188_, _3188_, _3188_, _3188_, _3188_, _3188_, _3188_, _3188_, _3188_ };
assign _1867_ = { _1565_, _1565_, _1565_, _1565_, _1565_, _1565_, _1565_, _1565_, _1565_ } | { _1564_, _1564_, _1564_, _1564_, _1564_, _1564_, _1564_, _1564_, _1564_ };
assign _1870_ = { _0428_, _0428_, _0428_, _0428_, _0428_, _0428_, _0428_, _0428_, _0428_ } | { _0427_, _0427_, _0427_, _0427_, _0427_, _0427_, _0427_, _0427_, _0427_ };
assign _1873_ = { _0440_, _0440_, _0440_, _0440_, _0440_, _0440_, _0440_, _0440_, _0440_ } | { _0439_, _0439_, _0439_, _0439_, _0439_, _0439_, _0439_, _0439_, _0439_ };
assign _1890_ = { _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_ } | { _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_, _3251_ };
assign _1908_ = { _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_ } | { _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_, _3066_ };
assign _1911_ = { _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_ } | { _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_, _0456_ };
assign _1918_ = _0434_ | _0433_;
assign _1924_ = _1579_ | _1578_;
assign _1927_ = _0446_ | _0445_;
assign _1930_ = _0436_ | _0435_;
assign _1958_ = { _2153_, _2153_, _2153_ } | { _2152_, _2152_, _2152_ };
assign _1962_ = { _0448_, _0448_, _0448_ } | { _0447_, _0447_, _0447_ };
assign _1983_ = csr_save_cause_i_t0 | csr_save_cause_i;
assign _1986_ = nmi_mode_i_t0 | nmi_mode_i;
assign _1988_ = { nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0 } | { nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i };
assign _1990_ = { nmi_mode_i_t0, nmi_mode_i_t0 } | { nmi_mode_i, nmi_mode_i };
assign _1993_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } | { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
assign _1996_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } | { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
assign _1999_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } | { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
assign _2002_ = csr_restore_mret_i_t0 | csr_restore_mret_i;
assign _2005_ = csr_restore_dret_i_t0 | csr_restore_dret_i;
assign _2013_ = _3079_ | _3078_;
assign _2015_ = debug_mode_i_t0 | debug_mode_i;
assign _2018_ = { debug_mode_i_t0, debug_mode_i_t0 } | { debug_mode_i, debug_mode_i };
assign _2021_ = { debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0 } | { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i };
assign _2024_ = { debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0 } | { debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i, debug_mode_i };
assign _2031_ = debug_csr_save_i_t0 | debug_csr_save_i;
assign _2033_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } | { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
assign _2036_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } | { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
assign _2039_ = { debug_csr_save_i_t0, debug_csr_save_i_t0 } | { debug_csr_save_i, debug_csr_save_i };
assign _2047_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } | { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
assign _2053_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } | { debug_csr_save_i, debug_csr_save_i, debug_csr_save_i, debug_csr_save_i };
assign _2056_ = { csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0 } | { csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i, csr_save_wb_i };
assign _2059_ = { csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0 } | { csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i, csr_save_id_i };
assign _2062_ = { csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0 } | { csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i, csr_save_if_i };
assign _2070_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } | { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
assign _2075_ = { csr_save_cause_i_t0, csr_save_cause_i_t0 } | { csr_save_cause_i, csr_save_cause_i };
assign _2083_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } | { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
assign _2086_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } | { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
assign _2089_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } | { csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i, csr_save_cause_i };
assign _2095_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } | { csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i, csr_restore_mret_i };
assign _2098_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } | { csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i, csr_restore_dret_i };
assign _2104_ = { nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0 } | { nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i, nmi_mode_i };
assign _2106_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0 } | { csr_restore_mret_i, csr_restore_mret_i };
assign _2108_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0 } | { csr_restore_dret_i, csr_restore_dret_i };
assign _2112_ = { _0068_, _0068_ } | { _3161_, _3161_ };
assign _2119_ = { _0032_, _0032_ } | { _3160_, _3160_ };
assign _2126_ = { _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_ } | { _3170_, _3170_, _3170_, _3170_, _3170_, _3170_, _3170_, _3170_ };
assign _2128_ = { _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_ } | { _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_, _3164_ };
assign _2129_ = { _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_ } | { _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_, _3168_ };
assign _2131_ = csr_we_int_t0 | csr_we_int;
assign _2133_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } | { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int };
assign _2136_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } | { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int };
assign _2140_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } | { csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int, csr_we_int };
assign _2144_ = { csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0 } | { csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i, csr_mtvec_init_i };
assign _2147_ = { mstatus_q_t0[1], mstatus_q_t0[1] } | { mstatus_q[1], mstatus_q[1] };
assign _2150_ = { _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_ } | { _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_, _0152_ };
assign _0546_ = _0023_[35] & _1609_;
assign _0551_ = _2616_ & _1613_;
assign _0554_ = dscratch0_q_t0[3] & _1616_;
assign _0557_ = irq_software_i_t0 & _1619_;
assign _0560_ = _2622_ & _1622_;
assign _0563_ = _2624_ & _1625_;
assign _0566_ = _2626_ & _1628_;
assign _0569_ = mcause_q_t0[3] & _1631_;
assign _0572_ = csr_mtvec_o_t0[3] & _1634_;
assign _0575_ = _2632_ & _1637_;
assign _0578_ = mie_q_t0[17] & _1640_;
assign _0583_ = _2638_ & _1644_;
assign _0586_ = _2640_ & _1647_;
assign _0589_ = _2642_ & _1650_;
assign _0592_ = _2644_ & _1653_;
assign _0595_ = _0023_[34:32] & _1656_;
assign _0600_ = _2648_ & _1660_;
assign _0603_ = dscratch1_q_t0[2:0] & _1663_;
assign _0606_ = dcsr_q_t0[2:0] & _1666_;
assign _0609_ = _2654_ & _1669_;
assign _0612_ = _2656_ & _1672_;
assign _0615_ = _2658_ & _1675_;
assign _0618_ = mcause_q_t0[2:0] & _1678_;
assign _0621_ = csr_mtvec_o_t0[2:0] & _1681_;
assign _0624_ = _2664_ & _1684_;
assign _0629_ = { _2670_[2], _2670_[2], 1'h0 } & _1689_;
assign _0632_ = _2672_ & _1692_;
assign _0635_ = _2674_ & _1695_;
assign _0638_ = _2676_ & _1698_;
assign _0643_ = _2678_ & _1701_;
assign _0646_ = dscratch0_q_t0[10:8] & _1704_;
assign _0649_ = dcsr_q_t0[10:8] & _1666_;
assign _0652_ = _2684_ & _1708_;
assign _0655_ = _2686_ & _1711_;
assign _0658_ = { mcause_q_t0[6], mcause_q_t0[6], mcause_q_t0[6] } & _1678_;
assign _0661_ = csr_mtvec_o_t0[10:8] & _1681_;
assign _0664_ = _2692_ & _1684_;
assign _0671_ = _2698_ & _1692_;
assign _0674_ = _2700_ & _1695_;
assign _0677_ = _2702_ & _1719_;
assign _0680_ = _0023_[20:18] & _1701_;
assign _0683_ = dscratch1_q_t0[20:18] & _1723_;
assign _0685_ = _2706_ & _1724_;
assign _0688_ = csr_depc_o_t0[20:18] & _1669_;
assign _0691_ = irq_fast_i_t0[4:2] & _1728_;
assign _0694_ = _2712_ & _1731_;
assign _0697_ = _2714_ & _1734_;
assign _0702_ = csr_mtvec_o_t0[20:18] & _1681_;
assign _0705_ = _2720_ & _1684_;
assign _0708_ = mie_q_t0[4:2] & _1687_;
assign _0713_ = _2726_ & _1741_;
assign _0715_ = _2728_ & _1742_;
assign _0718_ = _2730_ & _1695_;
assign _0721_ = _2732_ & _1746_;
assign _0724_ = _0023_[12] & _1749_;
assign _0727_ = dscratch1_q_t0[12] & _1752_;
assign _0729_ = _2736_ & _1753_;
assign _0732_ = csr_depc_o_t0[12] & _1756_;
assign _0735_ = csr_mtval_o_t0[12] & _1619_;
assign _0738_ = _2742_ & _1760_;
assign _0741_ = _2744_ & _1763_;
assign _0744_ = csr_mepc_o_t0[12] & _1766_;
assign _0747_ = mscratch_q_t0[12] & _1769_;
assign _0750_ = _2750_ & _1772_;
assign _0753_ = mstatus_q_t0[3] & _1775_;
assign _0757_ = _2756_ & _1776_;
assign _0760_ = _2758_ & _1779_;
assign _0763_ = _2760_ & _1782_;
assign _0766_ = _0023_[17] & _1749_;
assign _0769_ = dscratch1_q_t0[17] & _1752_;
assign _0771_ = _2764_ & _1753_;
assign _0774_ = csr_depc_o_t0[17] & _1756_;
assign _0777_ = irq_fast_i_t0[1] & _1619_;
assign _0780_ = _2770_ & _1760_;
assign _0783_ = _2772_ & _1763_;
assign _0786_ = mcause_q_t0[6] & _1631_;
assign _0789_ = csr_mtvec_o_t0[17] & _1634_;
assign _0792_ = _2778_ & _1637_;
assign _0795_ = mie_q_t0[1] & _1640_;
assign _0800_ = _2784_ & _1644_;
assign _0803_ = _2786_ & _1647_;
assign _0806_ = _2788_ & _1650_;
assign _0809_ = _2790_ & _1798_;
assign _0814_ = _2792_ & _1701_;
assign _0817_ = dscratch0_q_t0[15:13] & _1704_;
assign _0820_ = dcsr_q_t0[15:13] & _1666_;
assign _0823_ = _2798_ & _1708_;
assign _0826_ = _2800_ & _1711_;
assign _0829_ = csr_mepc_o_t0[15:13] & _1806_;
assign _0832_ = _2804_ & _1678_;
assign _0835_ = mscratch_q_t0[15:13] & _1810_;
assign _0840_ = _2810_ & _1813_;
assign _0843_ = _2812_ & _1816_;
assign _0846_ = _2814_ & _1719_;
assign _0849_ = _0023_[16] & _1749_;
assign _0852_ = dscratch1_q_t0[16] & _1752_;
assign _0854_ = _2818_ & _1753_;
assign _0857_ = csr_depc_o_t0[16] & _1756_;
assign _0860_ = irq_fast_i_t0[0] & _1619_;
assign _0863_ = _2824_ & _1760_;
assign _0866_ = _2826_ & _1763_;
assign _0871_ = csr_mtvec_o_t0[16] & _1634_;
assign _0874_ = _2832_ & _1637_;
assign _0877_ = mie_q_t0[0] & _1640_;
assign _0882_ = _2838_ & _1647_;
assign _0885_ = _2840_ & _1650_;
assign _0888_ = _2842_ & _1798_;
assign _0891_ = _0023_[30:22] & _1833_;
assign _0894_ = dscratch1_q_t0[30:22] & _1836_;
assign _0896_ = _2846_ & _1837_;
assign _0899_ = csr_depc_o_t0[30:22] & _1840_;
assign _0902_ = irq_fast_i_t0[14:6] & _1843_;
assign _0905_ = _2852_ & _1846_;
assign _0908_ = _2854_ & _1849_;
assign _0911_ = { mcause_q_t0[6], mcause_q_t0[6], mcause_q_t0[6], mcause_q_t0[6], mcause_q_t0[6], mcause_q_t0[6], mcause_q_t0[6], mcause_q_t0[6], mcause_q_t0[6] } & _1852_;
assign _0914_ = csr_mtvec_o_t0[30:22] & _1855_;
assign _0917_ = _2860_ & _1858_;
assign _0920_ = mie_q_t0[14:6] & _1861_;
assign _0925_ = _2866_ & _1865_;
assign _0927_ = _2868_ & _1866_;
assign _0930_ = _2870_ & _1869_;
assign _0933_ = _2872_ & _1872_;
assign _0936_ = _0023_[11] & _1749_;
assign _0939_ = dscratch1_q_t0[11] & _1752_;
assign _0941_ = _2876_ & _1753_;
assign _0944_ = csr_depc_o_t0[11] & _1756_;
assign _0947_ = irq_external_i_t0 & _1619_;
assign _0950_ = _2882_ & _1760_;
assign _0953_ = _2884_ & _1763_;
assign _0958_ = csr_mtvec_o_t0[11] & _1634_;
assign _0961_ = _2890_ & _1637_;
assign _0964_ = mie_q_t0[15] & _1640_;
assign _0969_ = _2896_ & _1644_;
assign _0972_ = _2898_ & _1647_;
assign _0975_ = _2900_ & _1650_;
assign _0978_ = _2902_ & _1798_;
assign _0981_ = \mhpmcounter[0]_t0  & _1889_;
assign _0984_ = _2903_ & _1892_;
assign _0986_ = _0023_[21] & _1749_;
assign _0989_ = dscratch1_q_t0[21] & _1752_;
assign _0991_ = _2907_ & _1753_;
assign _0994_ = csr_depc_o_t0[21] & _1756_;
assign _0997_ = irq_fast_i_t0[5] & _1619_;
assign _1000_ = _2913_ & _1760_;
assign _1003_ = _2915_ & _1763_;
assign _1008_ = csr_mtvec_o_t0[21] & _1634_;
assign _1011_ = _2921_ & _1637_;
assign _1014_ = mie_q_t0[5] & _1640_;
assign _1019_ = _2927_ & _1644_;
assign _1022_ = _2929_ & _1647_;
assign _1025_ = _2931_ & _1650_;
assign _1028_ = _2933_ & _1798_;
assign _1031_ = _3106_ & _1907_;
assign _1034_ = _2935_ & _1910_;
assign _1039_ = _2937_ & _1749_;
assign _1042_ = dscratch0_q_t0[31] & _1616_;
assign _1045_ = dcsr_q_t0[31] & _1622_;
assign _1048_ = _2943_ & _1625_;
assign _1051_ = _2945_ & _1917_;
assign _1054_ = csr_mepc_o_t0[31] & _1766_;
assign _1057_ = _2949_ & _1631_;
assign _1060_ = mscratch_q_t0[31] & _1769_;
assign _1065_ = _2955_ & _1923_;
assign _1068_ = _2957_ & _1926_;
assign _1071_ = _2959_ & _1929_;
assign _1074_ = _0023_[39] & _1609_;
assign _1079_ = _2963_ & _1613_;
assign _1082_ = dscratch0_q_t0[7] & _1616_;
assign _1085_ = irq_timer_i_t0 & _1619_;
assign _1088_ = _2969_ & _1622_;
assign _1091_ = _2971_ & _1625_;
assign _1094_ = _2973_ & _1628_;
assign _1099_ = csr_mtvec_o_t0[7] & _1634_;
assign _1102_ = _2979_ & _1637_;
assign _1105_ = mie_q_t0[16] & _1640_;
assign _1110_ = _2985_ & _1644_;
assign _1113_ = _2987_ & _1647_;
assign _1116_ = _2989_ & _1650_;
assign _1119_ = _2991_ & _1653_;
assign _1122_ = _0023_[38:36] & _1656_;
assign _1127_ = _2995_ & _1660_;
assign _1130_ = dscratch0_q_t0[6:4] & _1704_;
assign _1133_ = dcsr_q_t0[6:4] & _1666_;
assign _1136_ = _3001_ & _1708_;
assign _1139_ = _3003_ & _1675_;
assign _1142_ = { mcause_q_t0[6], mcause_q_t0[6], mcause_q_t0[4] } & _1678_;
assign _1145_ = csr_mtvec_o_t0[6:4] & _1681_;
assign _1148_ = _3009_ & _1684_;
assign _1151_ = hart_id_i_t0[6:4] & _1687_;
assign _1154_ = { 2'h0, _2670_[2] } & _1957_;
assign _1157_ = _3016_ & _1695_;
assign _1160_ = _3018_ & _1961_;
assign _1211_ = _0001_[7] & _1982_;
assign _1214_ = _0013_ & _1985_;
assign _1216_ = { dummy_instr_seed_o_t0[31:1], 1'h0 } & _1987_;
assign _1219_ = _0015_ & _1985_;
assign _1225_ = _0017_[1] & _1991_;
assign _1227_ = _0017_[4:2] & _1992_;
assign _1230_ = _3113_ & _1995_;
assign _1233_ = _3115_ & _1998_;
assign _1236_ = _0017_[1] & _2001_;
assign _1239_ = _3117_ & _2004_;
assign _1242_ = _3119_ & _1982_;
assign _1245_ = _0017_[5] & _2001_;
assign _1248_ = _3121_ & _2004_;
assign _1251_ = _3123_ & _1982_;
assign _1256_ = cpuctrlsts_part_q_t0[6] & _2012_;
assign _1258_ = _0001_[7] & _2011_;
assign _1262_ = _0128_ & _2014_;
assign _1265_ = _0126_ & _2017_;
assign _1268_ = _0097_ & _2014_;
assign _1270_ = csr_mcause_i_t0 & _2020_;
assign _1275_ = _0044_ & _2023_;
assign _1280_ = _0138_ & _2012_;
assign _1283_ = priv_mode_id_o_t0 & _2017_;
assign _1286_ = mstatus_q_t0[5] & _2014_;
assign _1291_ = csr_mtval_i_t0 & _2023_;
assign _1296_ = _0009_ & _2030_;
assign _1298_ = { dummy_instr_seed_o_t0[31:1], 1'h0 } & _2032_;
assign _1301_ = _0007_ & _2030_;
assign _1303_ = _0005_[8:6] & _2035_;
assign _1306_ = _0005_[1:0] & _2038_;
assign _1309_ = _0113_ & _2030_;
assign _1312_ = _0111_ & _2038_;
assign _1315_ = debug_mode_i_t0 & _2030_;
assign _1317_ = _0124_ & _2030_;
assign _1320_ = _0087_ & _2032_;
assign _1323_ = _0116_ & _2030_;
assign _1326_ = _0080_ & _2046_;
assign _1329_ = _0118_ & _2030_;
assign _1332_ = _0082_ & _2032_;
assign _1335_ = _0122_ & _2030_;
assign _1338_ = _0136_ & _2052_;
assign _1341_ = _0078_ & _2030_;
assign _1343_ = pc_id_i_t0 & _2055_;
assign _1346_ = _3125_ & _2058_;
assign _1349_ = _3127_ & _2061_;
assign _1352_ = _0003_ & _2001_;
assign _1354_ = _3129_ & _2004_;
assign _1357_ = _3131_ & _1982_;
assign _1360_ = _0001_[6] & _2001_;
assign _1362_ = _3133_ & _2004_;
assign _1365_ = _3135_ & _1982_;
assign _1370_ = _0009_ & _1982_;
assign _1373_ = { dummy_instr_seed_o_t0[31:1], 1'h0 } & _2069_;
assign _1376_ = _0007_ & _1982_;
assign _1379_ = _0005_[8:6] & _1998_;
assign _1382_ = _0005_[1:0] & _2074_;
assign _1385_ = _0021_ & _1982_;
assign _1388_ = dummy_instr_seed_o_t0 & _2069_;
assign _1391_ = _0013_ & _2001_;
assign _1394_ = _3137_ & _2004_;
assign _1397_ = _3139_ & _1982_;
assign _1400_ = { _3065_, _3063_, dummy_instr_seed_o_t0[4:0] } & _2082_;
assign _1403_ = _3141_ & _2085_;
assign _1406_ = _3143_ & _2088_;
assign _1409_ = _0015_ & _2001_;
assign _1412_ = _3145_ & _2004_;
assign _1415_ = _3147_ & _1982_;
assign _1418_ = { dummy_instr_seed_o_t0[31:1], 1'h0 } & _2094_;
assign _1421_ = _3149_ & _2097_;
assign _1424_ = _3151_ & _2069_;
assign _1427_ = _0019_ & _2001_;
assign _1429_ = _3153_ & _2004_;
assign _1432_ = _3155_ & _1982_;
assign _1435_ = { _3065_, _3063_, dummy_instr_seed_o_t0[4:0] } & _2103_;
assign _1440_ = _3157_ & _2107_;
assign _1443_ = _3159_ & _2074_;
assign _1447_ = dcsr_q_t0[31:28] & _2110_;
assign _1449_ = mstatus_q_t0[5:4] & _2111_;
assign _1452_ = mstatus_q_t0[3:2] & _2111_;
assign _1455_ = dcsr_q_t0[15] & _1619_;
assign _1458_ = dcsr_q_t0[14] & _1619_;
assign _1460_ = dcsr_q_t0[27:16] & _2116_;
assign _1462_ = mstatus_q_t0[1:0] & _2111_;
assign _1465_ = dcsr_q_t0[1:0] & _2118_;
assign _1468_ = dcsr_q_t0[5] & _1619_;
assign _1470_ = dcsr_q_t0[4] & _1619_;
assign _1472_ = dcsr_q_t0[3] & _1619_;
assign _1474_ = dcsr_q_t0[2] & _1619_;
assign _1477_ = dcsr_q_t0[13:12] & _2118_;
assign _1480_ = dcsr_q_t0[11] & _1619_;
assign _1482_ = dummy_instr_seed_o_t0[1:0] & _2123_;
assign _1484_ = dcsr_q_t0[9] & _1619_;
assign _1486_ = dummy_instr_seed_o_t0[12:11] & _2124_;
assign _1489_ = cpuctrlsts_part_q_t0 & _2125_;
assign _1496_ = dcsr_q_t0[10] & _1619_;
assign _1498_ = csr_mtvec_init_i_t0 & _1769_;
assign _1502_ = cpuctrlsts_part_q_t0 & _2132_;
assign _1519_ = dcsr_q_t0 & _2135_;
assign _1522_ = csr_mtvec_init_i_t0 & _2130_;
assign _1537_ = mstatus_q_t0 & _2139_;
assign _1540_ = _0011_ & _2142_;
assign _1549_ = { dummy_instr_seed_o_t0[31:8], 8'h00 } & _2143_;
assign _1552_ = priv_mode_id_o_t0 & _2146_;
assign _1555_ = minstret_raw_t0 & _2149_;
assign _0547_ = cpuctrlsts_part_q_t0[3] & _1610_;
assign _0549_ = _0023_[3] & _1612_;
assign _0552_ = _2614_ & _1614_;
assign _0555_ = dscratch1_q_t0[3] & _1617_;
assign _0558_ = dcsr_q_t0[3] & _1620_;
assign _0561_ = csr_depc_o_t0[3] & _1623_;
assign _0564_ = _2620_ & _1626_;
assign _0567_ = _2618_ & _1629_;
assign _0570_ = csr_mtval_o_t0[3] & _1632_;
assign _0573_ = csr_mepc_o_t0[3] & _1635_;
assign _0576_ = _2630_ & _1638_;
assign _0579_ = mscratch_q_t0[3] & _1641_;
assign _0581_ = hart_id_i_t0[3] & _1643_;
assign _0584_ = mstatus_q_t0[5] & _1645_;
assign _0587_ = _2636_ & _1648_;
assign _0590_ = _2634_ & _1651_;
assign _0593_ = _2628_ & _1654_;
assign _0596_ = cpuctrlsts_part_q_t0[2:0] & _1657_;
assign _0598_ = _0023_[2:0] & _1659_;
assign _0601_ = _2646_ & _1661_;
assign _0604_ = { mcountinhibit_t0[2], 1'h0, mcountinhibit_t0[0] } & _1664_;
assign _0607_ = csr_depc_o_t0[2:0] & _1667_;
assign _0610_ = dscratch0_q_t0[2:0] & _1670_;
assign _0613_ = _2652_ & _1673_;
assign _0616_ = _2650_ & _1676_;
assign _0619_ = csr_mtval_o_t0[2:0] & _1679_;
assign _0622_ = csr_mepc_o_t0[2:0] & _1682_;
assign _0625_ = _2662_ & _1685_;
assign _0627_ = mscratch_q_t0[2:0] & _1688_;
assign _0630_ = hart_id_i_t0[2:0] & _1690_;
assign _0633_ = _2668_ & _1693_;
assign _0636_ = _2666_ & _1696_;
assign _0639_ = _2660_ & _1699_;
assign _0641_ = _0023_[10:8] & _1659_;
assign _0644_ = _0023_[42:40] & _1702_;
assign _0647_ = dscratch1_q_t0[10:8] & _1705_;
assign _0650_ = csr_depc_o_t0[10:8] & _1667_;
assign _0653_ = _2682_ & _1709_;
assign _0656_ = _2680_ & _1712_;
assign _0659_ = csr_mtval_o_t0[10:8] & _1679_;
assign _0662_ = csr_mepc_o_t0[10:8] & _1682_;
assign _0665_ = _2690_ & _1685_;
assign _0667_ = mscratch_q_t0[10:8] & _1688_;
assign _0669_ = hart_id_i_t0[10:8] & _1690_;
assign _0672_ = _2696_ & _1693_;
assign _0675_ = _2694_ & _1696_;
assign _0678_ = _2688_ & _1720_;
assign _0681_ = _0023_[52:50] & _1702_;
assign _0686_ = _2704_ & _1725_;
assign _0689_ = dscratch0_q_t0[20:18] & _1670_;
assign _0692_ = dcsr_q_t0[20:18] & _1729_;
assign _0695_ = _2710_ & _1732_;
assign _0698_ = _2708_ & _1735_;
assign _0700_ = csr_mtval_o_t0[20:18] & _1679_;
assign _0703_ = csr_mepc_o_t0[20:18] & _1682_;
assign _0706_ = _2718_ & _1685_;
assign _0709_ = mscratch_q_t0[20:18] & _1688_;
assign _0711_ = hart_id_i_t0[20:18] & _1690_;
assign _0716_ = _2724_ & _1743_;
assign _0719_ = _2722_ & _1696_;
assign _0722_ = _2716_ & _1747_;
assign _0725_ = _0023_[44] & _1750_;
assign _0730_ = _2734_ & _1754_;
assign _0733_ = dscratch0_q_t0[12] & _1757_;
assign _0736_ = dcsr_q_t0[12] & _1620_;
assign _0739_ = _2740_ & _1761_;
assign _0742_ = _2738_ & _1764_;
assign _0745_ = mcause_q_t0[6] & _1767_;
assign _0748_ = csr_mtvec_o_t0[12] & _1770_;
assign _0751_ = _2748_ & _1773_;
assign _0755_ = hart_id_i_t0[12] & _1643_;
assign _0758_ = _2754_ & _1777_;
assign _0761_ = _2752_ & _1780_;
assign _0764_ = _2746_ & _1783_;
assign _0767_ = _0023_[49] & _1750_;
assign _0772_ = _2762_ & _1754_;
assign _0775_ = dscratch0_q_t0[17] & _1757_;
assign _0778_ = dcsr_q_t0[17] & _1620_;
assign _0781_ = _2768_ & _1761_;
assign _0784_ = _2766_ & _1764_;
assign _0787_ = csr_mtval_o_t0[17] & _1632_;
assign _0790_ = csr_mepc_o_t0[17] & _1635_;
assign _0793_ = _2776_ & _1638_;
assign _0796_ = mscratch_q_t0[17] & _1641_;
assign _0798_ = hart_id_i_t0[17] & _1643_;
assign _0801_ = mstatus_q_t0[1] & _1645_;
assign _0804_ = _2782_ & _1648_;
assign _0807_ = _2780_ & _1651_;
assign _0810_ = _2774_ & _1799_;
assign _0812_ = _0023_[15:13] & _1659_;
assign _0815_ = _0023_[47:45] & _1702_;
assign _0818_ = dscratch1_q_t0[15:13] & _1705_;
assign _0821_ = csr_depc_o_t0[15:13] & _1667_;
assign _0824_ = _2796_ & _1709_;
assign _0827_ = _2794_ & _1712_;
assign _0830_ = { mcause_q_t0[6], mcause_q_t0[6], mcause_q_t0[6] } & _1807_;
assign _0833_ = csr_mtval_o_t0[15:13] & _1679_;
assign _0836_ = csr_mtvec_o_t0[15:13] & _1811_;
assign _0838_ = hart_id_i_t0[15:13] & _1690_;
assign _0841_ = _2808_ & _1814_;
assign _0844_ = _2806_ & _1817_;
assign _0847_ = _2802_ & _1720_;
assign _0850_ = _0023_[48] & _1750_;
assign _0855_ = _2816_ & _1754_;
assign _0858_ = dscratch0_q_t0[16] & _1757_;
assign _0861_ = dcsr_q_t0[16] & _1620_;
assign _0864_ = _2822_ & _1761_;
assign _0867_ = _2820_ & _1764_;
assign _0869_ = csr_mtval_o_t0[16] & _1632_;
assign _0872_ = csr_mepc_o_t0[16] & _1635_;
assign _0875_ = _2830_ & _1638_;
assign _0878_ = mscratch_q_t0[16] & _1641_;
assign _0880_ = hart_id_i_t0[16] & _1643_;
assign _0883_ = _2836_ & _1648_;
assign _0886_ = _2834_ & _1651_;
assign _0889_ = _2828_ & _1799_;
assign _0892_ = _0023_[62:54] & _1834_;
assign _0897_ = _2844_ & _1838_;
assign _0900_ = dscratch0_q_t0[30:22] & _1841_;
assign _0903_ = dcsr_q_t0[30:22] & _1844_;
assign _0906_ = _2850_ & _1847_;
assign _0909_ = _2848_ & _1850_;
assign _0912_ = csr_mtval_o_t0[30:22] & _1853_;
assign _0915_ = csr_mepc_o_t0[30:22] & _1856_;
assign _0918_ = _2858_ & _1859_;
assign _0921_ = mscratch_q_t0[30:22] & _1862_;
assign _0923_ = hart_id_i_t0[30:22] & _1864_;
assign _0928_ = _2864_ & _1867_;
assign _0931_ = _2862_ & _1870_;
assign _0934_ = _2856_ & _1873_;
assign _0937_ = _0023_[43] & _1750_;
assign _0942_ = _2874_ & _1754_;
assign _0945_ = dscratch0_q_t0[11] & _1757_;
assign _0948_ = dcsr_q_t0[11] & _1620_;
assign _0951_ = _2880_ & _1761_;
assign _0954_ = _2878_ & _1764_;
assign _0956_ = csr_mtval_o_t0[11] & _1632_;
assign _0959_ = csr_mepc_o_t0[11] & _1635_;
assign _0962_ = _2888_ & _1638_;
assign _0965_ = mscratch_q_t0[11] & _1641_;
assign _0967_ = hart_id_i_t0[11] & _1643_;
assign _0970_ = mstatus_q_t0[2] & _1645_;
assign _0973_ = _2894_ & _1648_;
assign _0976_ = _2892_ & _1651_;
assign _0979_ = _2886_ & _1799_;
assign _0982_ = \mhpmcounter[2]_t0  & _1890_;
assign _0987_ = _0023_[53] & _1750_;
assign _0992_ = _2905_ & _1754_;
assign _0995_ = dscratch0_q_t0[21] & _1757_;
assign _0998_ = dcsr_q_t0[21] & _1620_;
assign _1001_ = _2911_ & _1761_;
assign _1004_ = _2909_ & _1764_;
assign _1006_ = csr_mtval_o_t0[21] & _1632_;
assign _1009_ = csr_mepc_o_t0[21] & _1635_;
assign _1012_ = _2919_ & _1638_;
assign _1015_ = mscratch_q_t0[21] & _1641_;
assign _1017_ = hart_id_i_t0[21] & _1643_;
assign _1020_ = mstatus_q_t0[0] & _1645_;
assign _1023_ = _2925_ & _1648_;
assign _1026_ = _2923_ & _1651_;
assign _1029_ = _2917_ & _1799_;
assign _1032_ = _0146_ & _1908_;
assign _1035_ = csr_wdata_i_t0 & _1911_;
assign _1037_ = _0023_[31] & _1612_;
assign _1040_ = _0023_[63] & _1750_;
assign _1043_ = dscratch1_q_t0[31] & _1617_;
assign _1046_ = csr_depc_o_t0[31] & _1623_;
assign _1049_ = _2941_ & _1626_;
assign _1052_ = _2939_ & _1918_;
assign _1055_ = _3104_ & _1767_;
assign _1058_ = csr_mtval_o_t0[31] & _1632_;
assign _1061_ = csr_mtvec_o_t0[31] & _1770_;
assign _1063_ = hart_id_i_t0[31] & _1643_;
assign _1066_ = _2953_ & _1924_;
assign _1069_ = _2951_ & _1927_;
assign _1072_ = _2947_ & _1930_;
assign _1075_ = cpuctrlsts_part_q_t0[7] & _1610_;
assign _1077_ = _0023_[7] & _1612_;
assign _1080_ = _2961_ & _1614_;
assign _1083_ = dscratch1_q_t0[7] & _1617_;
assign _1086_ = dcsr_q_t0[7] & _1620_;
assign _1089_ = csr_depc_o_t0[7] & _1623_;
assign _1092_ = _2967_ & _1626_;
assign _1095_ = _2965_ & _1629_;
assign _1097_ = csr_mtval_o_t0[7] & _1632_;
assign _1100_ = csr_mepc_o_t0[7] & _1635_;
assign _1103_ = _2977_ & _1638_;
assign _1106_ = mscratch_q_t0[7] & _1641_;
assign _1108_ = hart_id_i_t0[7] & _1643_;
assign _1111_ = mstatus_q_t0[4] & _1645_;
assign _1114_ = _2983_ & _1648_;
assign _1117_ = _2981_ & _1651_;
assign _1120_ = _2975_ & _1654_;
assign _1123_ = cpuctrlsts_part_q_t0[6:4] & _1657_;
assign _1125_ = _0023_[6:4] & _1659_;
assign _1128_ = _2993_ & _1661_;
assign _1131_ = dscratch1_q_t0[6:4] & _1705_;
assign _1134_ = csr_depc_o_t0[6:4] & _1667_;
assign _1137_ = _2999_ & _1709_;
assign _1140_ = _2997_ & _1676_;
assign _1143_ = csr_mtval_o_t0[6:4] & _1679_;
assign _1146_ = csr_mepc_o_t0[6:4] & _1682_;
assign _1149_ = _3007_ & _1685_;
assign _1152_ = mscratch_q_t0[6:4] & _1688_;
assign _1155_ = _3013_ & _1958_;
assign _1158_ = _3011_ & _1696_;
assign _1161_ = _3005_ & _1962_;
assign _1212_ = _0089_[1] & _1983_;
assign _1217_ = mstack_epc_q_t0 & _1988_;
assign _1221_ = mstack_q_t0[1:0] & _1990_;
assign _1223_ = mstack_q_t0[2] & _1986_;
assign _1228_ = _0144_ & _1993_;
assign _1231_ = _0017_[4:2] & _1996_;
assign _1234_ = _0120_[2:0] & _1999_;
assign _1237_ = _0142_ & _2002_;
assign _1240_ = _0017_[1] & _2005_;
assign _1243_ = _0017_[1] & _1983_;
assign _1246_ = mstatus_q_t0[4] & _2002_;
assign _1249_ = _0017_[5] & _2005_;
assign _1252_ = _0120_[3] & _1983_;
assign _1254_ = _0001_[6] & _2013_;
assign _1260_ = _0003_ & _2013_;
assign _1263_ = _0003_ & _2015_;
assign _1266_ = _0001_[7:6] & _2018_;
assign _1271_ = { _3065_, _3063_, dummy_instr_seed_o_t0[4:0] } & _2021_;
assign _1273_ = _0013_ & _2015_;
assign _1276_ = { dummy_instr_seed_o_t0[31:1], 1'h0 } & _2024_;
assign _1278_ = _0015_ & _2015_;
assign _1281_ = _0001_[7] & _2013_;
assign _1284_ = _0017_[3:2] & _2018_;
assign _1287_ = _0017_[4] & _2015_;
assign _1289_ = _0019_ & _2015_;
assign _1292_ = dummy_instr_seed_o_t0 & _2024_;
assign _1294_ = _0021_ & _2015_;
assign _1299_ = _0044_ & _2033_;
assign _1304_ = debug_cause_i_t0 & _2036_;
assign _1307_ = priv_mode_id_o_t0 & _2039_;
assign _1310_ = _0003_ & _2031_;
assign _1313_ = _0001_[7:6] & _2039_;
assign _1318_ = _0021_ & _2031_;
assign _1321_ = dummy_instr_seed_o_t0 & _2033_;
assign _1324_ = _0013_ & _2031_;
assign _1327_ = { _3065_, _3063_, dummy_instr_seed_o_t0[4:0] } & _2047_;
assign _1330_ = _0015_ & _2031_;
assign _1333_ = { dummy_instr_seed_o_t0[31:1], 1'h0 } & _2033_;
assign _1336_ = _0019_ & _2031_;
assign _1339_ = _0017_[5:2] & _2053_;
assign _1344_ = pc_wb_i_t0 & _2056_;
assign _1347_ = pc_id_i_t0 & _2059_;
assign _1350_ = pc_if_i_t0 & _2062_;
assign _1355_ = _0003_ & _2005_;
assign _1358_ = _0091_ & _1983_;
assign _1363_ = _0001_[6] & _2005_;
assign _1366_ = _0089_[0] & _1983_;
assign _1368_ = _0064_ & _1983_;
assign _1371_ = _0095_ & _1983_;
assign _1374_ = _0034_ & _2070_;
assign _1377_ = _0093_ & _1983_;
assign _1380_ = _0140_ & _1999_;
assign _1383_ = _0130_ & _2075_;
assign _1386_ = _0109_ & _1983_;
assign _1389_ = _0070_ & _2070_;
assign _1392_ = _0132_ & _2002_;
assign _1395_ = _0013_ & _2005_;
assign _1398_ = _0101_ & _1983_;
assign _1401_ = _0099_ & _2083_;
assign _1404_ = { _3065_, _3063_, dummy_instr_seed_o_t0[4:0] } & _2086_;
assign _1407_ = _0046_ & _2089_;
assign _1410_ = _0134_ & _2002_;
assign _1413_ = _0015_ & _2005_;
assign _1416_ = _0105_ & _1983_;
assign _1419_ = _0103_ & _2095_;
assign _1422_ = { dummy_instr_seed_o_t0[31:1], 1'h0 } & _2098_;
assign _1425_ = _0052_ & _2070_;
assign _1430_ = _0019_ & _2005_;
assign _1433_ = _0107_ & _1983_;
assign _1436_ = mstack_cause_q_t0 & _2104_;
assign _1438_ = _0038_ & _1983_;
assign _3157_ = mstatus_q_t0[3:2] & _2106_;
assign _1441_ = dcsr_q_t0[1:0] & _2108_;
assign _1445_ = _0017_[5] & _2015_;
assign _1450_ = { dummy_instr_seed_o_t0[3], dummy_instr_seed_o_t0[7] } & _2112_;
assign _1453_ = _0085_ & _2112_;
assign _1456_ = dummy_instr_seed_o_t0[15] & _1620_;
assign _1463_ = { dummy_instr_seed_o_t0[17], dummy_instr_seed_o_t0[21] } & _2112_;
assign _1466_ = _0076_ & _2119_;
assign _1475_ = dummy_instr_seed_o_t0[2] & _1620_;
assign _1478_ = dummy_instr_seed_o_t0[13:12] & _2119_;
assign _1490_ = { dummy_instr_seed_o_t0[7:1], 1'h0 } & _2126_;
assign _1492_ = _3096_ & _2128_;
assign _1494_ = _3096_ & _2129_;
assign _1500_ = _0028_ & _2131_;
assign _1503_ = _0026_ & _2133_;
assign _1505_ = _0058_ & _2136_;
assign _1507_ = _0056_ & _2136_;
assign _1509_ = _0050_ & _2131_;
assign _1511_ = _0042_ & _2131_;
assign _1513_ = _0040_ & _2131_;
assign _1515_ = _0036_ & _2131_;
assign _1517_ = _0032_ & _2131_;
assign _1520_ = { _0030_[31:9], dcsr_q_t0[8:6], _0030_[5:0] } & _2136_;
assign _1523_ = _0074_ & _2131_;
assign _1525_ = _0072_ & _2131_;
assign _1527_ = _0048_ & _2131_;
assign _1529_ = _0054_ & _2131_;
assign _1531_ = _0062_ & _2131_;
assign _1533_ = _0060_ & _2131_;
assign _1535_ = _0068_ & _2131_;
assign _1538_ = _0066_ & _2140_;
assign _1550_ = { boot_addr_i_t0[31:8], 8'h00 } & _2144_;
assign _1553_ = mstatus_q_t0[3:2] & _2147_;
assign _1556_ = minstret_next_t0 & _2150_;
assign _1611_ = _0546_ | _0547_;
assign _1615_ = _0551_ | _0552_;
assign _1618_ = _0554_ | _0555_;
assign _1621_ = _0557_ | _0558_;
assign _1624_ = _0560_ | _0561_;
assign _1627_ = _0563_ | _0564_;
assign _1630_ = _0566_ | _0567_;
assign _1633_ = _0569_ | _0570_;
assign _1636_ = _0572_ | _0573_;
assign _1639_ = _0575_ | _0576_;
assign _1642_ = _0578_ | _0579_;
assign _1646_ = _0583_ | _0584_;
assign _1649_ = _0586_ | _0587_;
assign _1652_ = _0589_ | _0590_;
assign _1655_ = _0592_ | _0593_;
assign _1658_ = _0595_ | _0596_;
assign _1662_ = _0600_ | _0601_;
assign _1665_ = _0603_ | _0604_;
assign _1668_ = _0606_ | _0607_;
assign _1671_ = _0609_ | _0610_;
assign _1674_ = _0612_ | _0613_;
assign _1677_ = _0615_ | _0616_;
assign _1680_ = _0618_ | _0619_;
assign _1683_ = _0621_ | _0622_;
assign _1686_ = _0624_ | _0625_;
assign _1691_ = _0629_ | _0630_;
assign _1694_ = _0632_ | _0633_;
assign _1697_ = _0635_ | _0636_;
assign _1700_ = _0638_ | _0639_;
assign _1703_ = _0643_ | _0644_;
assign _1706_ = _0646_ | _0647_;
assign _1707_ = _0649_ | _0650_;
assign _1710_ = _0652_ | _0653_;
assign _1713_ = _0655_ | _0656_;
assign _1714_ = _0658_ | _0659_;
assign _1715_ = _0661_ | _0662_;
assign _1716_ = _0664_ | _0665_;
assign _1717_ = _0671_ | _0672_;
assign _1718_ = _0674_ | _0675_;
assign _1721_ = _0677_ | _0678_;
assign _1722_ = _0680_ | _0681_;
assign _1726_ = _0685_ | _0686_;
assign _1727_ = _0688_ | _0689_;
assign _1730_ = _0691_ | _0692_;
assign _1733_ = _0694_ | _0695_;
assign _1736_ = _0697_ | _0698_;
assign _1737_ = _0658_ | _0700_;
assign _1738_ = _0702_ | _0703_;
assign _1739_ = _0705_ | _0706_;
assign _1740_ = _0708_ | _0709_;
assign _1744_ = _0715_ | _0716_;
assign _1745_ = _0718_ | _0719_;
assign _1748_ = _0721_ | _0722_;
assign _1751_ = _0724_ | _0725_;
assign _1755_ = _0729_ | _0730_;
assign _1758_ = _0732_ | _0733_;
assign _1759_ = _0735_ | _0736_;
assign _1762_ = _0738_ | _0739_;
assign _1765_ = _0741_ | _0742_;
assign _1768_ = _0744_ | _0745_;
assign _1771_ = _0747_ | _0748_;
assign _1774_ = _0750_ | _0751_;
assign _1778_ = _0757_ | _0758_;
assign _1781_ = _0760_ | _0761_;
assign _1784_ = _0763_ | _0764_;
assign _1785_ = _0766_ | _0767_;
assign _1786_ = _0771_ | _0772_;
assign _1787_ = _0774_ | _0775_;
assign _1788_ = _0777_ | _0778_;
assign _1789_ = _0780_ | _0781_;
assign _1790_ = _0783_ | _0784_;
assign _1791_ = _0786_ | _0787_;
assign _1792_ = _0789_ | _0790_;
assign _1793_ = _0792_ | _0793_;
assign _1794_ = _0795_ | _0796_;
assign _1795_ = _0800_ | _0801_;
assign _1796_ = _0803_ | _0804_;
assign _1797_ = _0806_ | _0807_;
assign _1800_ = _0809_ | _0810_;
assign _1801_ = _0814_ | _0815_;
assign _1802_ = _0817_ | _0818_;
assign _1803_ = _0820_ | _0821_;
assign _1804_ = _0823_ | _0824_;
assign _1805_ = _0826_ | _0827_;
assign _1808_ = _0829_ | _0830_;
assign _1809_ = _0832_ | _0833_;
assign _1812_ = _0835_ | _0836_;
assign _1815_ = _0840_ | _0841_;
assign _1818_ = _0843_ | _0844_;
assign _1819_ = _0846_ | _0847_;
assign _1820_ = _0849_ | _0850_;
assign _1821_ = _0854_ | _0855_;
assign _1822_ = _0857_ | _0858_;
assign _1823_ = _0860_ | _0861_;
assign _1824_ = _0863_ | _0864_;
assign _1825_ = _0866_ | _0867_;
assign _1826_ = _0786_ | _0869_;
assign _1827_ = _0871_ | _0872_;
assign _1828_ = _0874_ | _0875_;
assign _1829_ = _0877_ | _0878_;
assign _1830_ = _0882_ | _0883_;
assign _1831_ = _0885_ | _0886_;
assign _1832_ = _0888_ | _0889_;
assign _1835_ = _0891_ | _0892_;
assign _1839_ = _0896_ | _0897_;
assign _1842_ = _0899_ | _0900_;
assign _1845_ = _0902_ | _0903_;
assign _1848_ = _0905_ | _0906_;
assign _1851_ = _0908_ | _0909_;
assign _1854_ = _0911_ | _0912_;
assign _1857_ = _0914_ | _0915_;
assign _1860_ = _0917_ | _0918_;
assign _1863_ = _0920_ | _0921_;
assign _1868_ = _0927_ | _0928_;
assign _1871_ = _0930_ | _0931_;
assign _1874_ = _0933_ | _0934_;
assign _1875_ = _0936_ | _0937_;
assign _1876_ = _0941_ | _0942_;
assign _1877_ = _0944_ | _0945_;
assign _1878_ = _0947_ | _0948_;
assign _1879_ = _0950_ | _0951_;
assign _1880_ = _0953_ | _0954_;
assign _1881_ = _0786_ | _0956_;
assign _1882_ = _0958_ | _0959_;
assign _1883_ = _0961_ | _0962_;
assign _1884_ = _0964_ | _0965_;
assign _1885_ = _0969_ | _0970_;
assign _1886_ = _0972_ | _0973_;
assign _1887_ = _0975_ | _0976_;
assign _1888_ = _0978_ | _0979_;
assign _1891_ = _0981_ | _0982_;
assign _1893_ = _0986_ | _0987_;
assign _1894_ = _0991_ | _0992_;
assign _1895_ = _0994_ | _0995_;
assign _1896_ = _0997_ | _0998_;
assign _1897_ = _1000_ | _1001_;
assign _1898_ = _1003_ | _1004_;
assign _1899_ = _0786_ | _1006_;
assign _1900_ = _1008_ | _1009_;
assign _1901_ = _1011_ | _1012_;
assign _1902_ = _1014_ | _1015_;
assign _1903_ = _1019_ | _1020_;
assign _1904_ = _1022_ | _1023_;
assign _1905_ = _1025_ | _1026_;
assign _1906_ = _1028_ | _1029_;
assign _1909_ = _1031_ | _1032_;
assign _1912_ = _1034_ | _1035_;
assign _1913_ = _1039_ | _1040_;
assign _1914_ = _1042_ | _1043_;
assign _1915_ = _1045_ | _1046_;
assign _1916_ = _1048_ | _1049_;
assign _1919_ = _1051_ | _1052_;
assign _1920_ = _1054_ | _1055_;
assign _1921_ = _1057_ | _1058_;
assign _1922_ = _1060_ | _1061_;
assign _1925_ = _1065_ | _1066_;
assign _1928_ = _1068_ | _1069_;
assign _1931_ = _1071_ | _1072_;
assign _1932_ = _1074_ | _1075_;
assign _1933_ = _1079_ | _1080_;
assign _1934_ = _1082_ | _1083_;
assign _1935_ = _1085_ | _1086_;
assign _1936_ = _1088_ | _1089_;
assign _1937_ = _1091_ | _1092_;
assign _1938_ = _1094_ | _1095_;
assign _1939_ = _0786_ | _1097_;
assign _1940_ = _1099_ | _1100_;
assign _1941_ = _1102_ | _1103_;
assign _1942_ = _1105_ | _1106_;
assign _1943_ = _1110_ | _1111_;
assign _1944_ = _1113_ | _1114_;
assign _1945_ = _1116_ | _1117_;
assign _1946_ = _1119_ | _1120_;
assign _1947_ = _1122_ | _1123_;
assign _1948_ = _1127_ | _1128_;
assign _1949_ = _1130_ | _1131_;
assign _1950_ = _1133_ | _1134_;
assign _1951_ = _1136_ | _1137_;
assign _1952_ = _1139_ | _1140_;
assign _1953_ = _1142_ | _1143_;
assign _1954_ = _1145_ | _1146_;
assign _1955_ = _1148_ | _1149_;
assign _1956_ = _1151_ | _1152_;
assign _1959_ = _1154_ | _1155_;
assign _1960_ = _1157_ | _1158_;
assign _1963_ = _1160_ | _1161_;
assign _1984_ = _1211_ | _1212_;
assign _1989_ = _1216_ | _1217_;
assign _1994_ = _1227_ | _1228_;
assign _1997_ = _1230_ | _1231_;
assign _2000_ = _1233_ | _1234_;
assign _2003_ = _1236_ | _1237_;
assign _2006_ = _1239_ | _1240_;
assign _2007_ = _1242_ | _1243_;
assign _2008_ = _1245_ | _1246_;
assign _2009_ = _1248_ | _1249_;
assign _2010_ = _1251_ | _1252_;
assign _2016_ = _1262_ | _1263_;
assign _2019_ = _1265_ | _1266_;
assign _2022_ = _1270_ | _1271_;
assign _2025_ = _1275_ | _1276_;
assign _2026_ = _1280_ | _1281_;
assign _2027_ = _1283_ | _1284_;
assign _2028_ = _1286_ | _1287_;
assign _2029_ = _1291_ | _1292_;
assign _2034_ = _1298_ | _1299_;
assign _2037_ = _1303_ | _1304_;
assign _2040_ = _1306_ | _1307_;
assign _2041_ = _1309_ | _1310_;
assign _2042_ = _1312_ | _1313_;
assign _2043_ = _1317_ | _1318_;
assign _2044_ = _1320_ | _1321_;
assign _2045_ = _1323_ | _1324_;
assign _2048_ = _1326_ | _1327_;
assign _2049_ = _1329_ | _1330_;
assign _2050_ = _1332_ | _1333_;
assign _2051_ = _1335_ | _1336_;
assign _2054_ = _1338_ | _1339_;
assign _2057_ = _1343_ | _1344_;
assign _2060_ = _1346_ | _1347_;
assign _2063_ = _1349_ | _1350_;
assign _2064_ = _1354_ | _1355_;
assign _2065_ = _1357_ | _1358_;
assign _2066_ = _1362_ | _1363_;
assign _2067_ = _1365_ | _1366_;
assign _2068_ = _1370_ | _1371_;
assign _2071_ = _1373_ | _1374_;
assign _2072_ = _1376_ | _1377_;
assign _2073_ = _1379_ | _1380_;
assign _2076_ = _1382_ | _1383_;
assign _2077_ = _1385_ | _1386_;
assign _2078_ = _1388_ | _1389_;
assign _2079_ = _1391_ | _1392_;
assign _2080_ = _1394_ | _1395_;
assign _2081_ = _1397_ | _1398_;
assign _2084_ = _1400_ | _1401_;
assign _2087_ = _1403_ | _1404_;
assign _2090_ = _1406_ | _1407_;
assign _2091_ = _1409_ | _1410_;
assign _2092_ = _1412_ | _1413_;
assign _2093_ = _1415_ | _1416_;
assign _2096_ = _1418_ | _1419_;
assign _2099_ = _1421_ | _1422_;
assign _2100_ = _1424_ | _1425_;
assign _2101_ = _1429_ | _1430_;
assign _2102_ = _1432_ | _1433_;
assign _2105_ = _1435_ | _1436_;
assign _2109_ = _1440_ | _1441_;
assign _2113_ = _1449_ | _1450_;
assign _2114_ = _1452_ | _1453_;
assign _2115_ = _1455_ | _1456_;
assign _2117_ = _1462_ | _1463_;
assign _2120_ = _1465_ | _1466_;
assign _2121_ = _1474_ | _1475_;
assign _2122_ = _1477_ | _1478_;
assign _2127_ = _1489_ | _1490_;
assign _2134_ = _1502_ | _1503_;
assign _2137_ = _1519_ | _1520_;
assign _2138_ = _1522_ | _1523_;
assign _2141_ = _1537_ | _1538_;
assign _2145_ = _1549_ | _1550_;
assign _2148_ = _1552_ | _1553_;
assign _2151_ = _1555_ | _1556_;
assign _2156_ = _0022_[35] ^ cpuctrlsts_part_q[3];
assign _2157_ = _0024_[3] ^ _0022_[3];
assign _2158_ = _2615_ ^ _2613_;
assign _2159_ = dscratch0_q[3] ^ dscratch1_q[3];
assign _2160_ = irq_software_i ^ dcsr_q[3];
assign _2161_ = _2621_ ^ csr_depc_o[3];
assign _2162_ = _2623_ ^ _2619_;
assign _2163_ = _2625_ ^ _2617_;
assign _2164_ = mcause_q[3] ^ csr_mtval_o[3];
assign _2165_ = csr_mtvec_o[3] ^ csr_mepc_o[3];
assign _2166_ = _2631_ ^ _2629_;
assign _2167_ = mie_q[17] ^ mscratch_q[3];
assign _2168_ = _2637_ ^ mstatus_q[5];
assign _2169_ = _2639_ ^ _2635_;
assign _2170_ = _2641_ ^ _2633_;
assign _2171_ = _2643_ ^ _2627_;
assign _2172_ = _0022_[34:32] ^ cpuctrlsts_part_q[2:0];
assign _2173_ = _0024_[2:0] ^ _0022_[2:0];
assign _2174_ = _2647_ ^ _2645_;
assign _2175_ = dscratch1_q[2:0] ^ { mcountinhibit[2], 1'h0, mcountinhibit[0] };
assign _2176_ = dcsr_q[2:0] ^ csr_depc_o[2:0];
assign _2177_ = _2653_ ^ dscratch0_q[2:0];
assign _2178_ = _2655_ ^ _2651_;
assign _2179_ = _2657_ ^ _2649_;
assign _2180_ = mcause_q[2:0] ^ csr_mtval_o[2:0];
assign _2181_ = csr_mtvec_o[2:0] ^ csr_mepc_o[2:0];
assign _2182_ = _2663_ ^ _2661_;
assign _2183_ = _2669_ ^ hart_id_i[2:0];
assign _2184_ = _2671_ ^ _2667_;
assign _2185_ = _2673_ ^ _2665_;
assign _2186_ = _2675_ ^ _2659_;
assign _2187_ = _0024_[10:8] ^ _0022_[10:8];
assign _2188_ = _2677_ ^ _0022_[42:40];
assign _2189_ = dscratch0_q[10:8] ^ dscratch1_q[10:8];
assign _2190_ = dcsr_q[10:8] ^ csr_depc_o[10:8];
assign _2191_ = _2683_ ^ _2681_;
assign _2192_ = _2685_ ^ _2679_;
assign _2193_ = _3270_[5:3] ^ csr_mtval_o[10:8];
assign _2194_ = csr_mtvec_o[10:8] ^ csr_mepc_o[10:8];
assign _2195_ = _2691_ ^ _2689_;
assign _2196_ = _2697_ ^ _2695_;
assign _2197_ = _2699_ ^ _2693_;
assign _2198_ = _2701_ ^ _2687_;
assign _2199_ = _0022_[20:18] ^ _0022_[52:50];
assign _2200_ = dscratch1_q[20:18] ^ _0024_[20:18];
assign _2201_ = _2705_ ^ _2703_;
assign _2202_ = csr_depc_o[20:18] ^ dscratch0_q[20:18];
assign _2203_ = irq_fast_i[4:2] ^ dcsr_q[20:18];
assign _2204_ = _2711_ ^ _2709_;
assign _2205_ = _2713_ ^ _2707_;
assign _2206_ = _3270_[15:13] ^ csr_mtval_o[20:18];
assign _2207_ = csr_mtvec_o[20:18] ^ csr_mepc_o[20:18];
assign _2208_ = _2719_ ^ _2717_;
assign _2209_ = mie_q[4:2] ^ mscratch_q[20:18];
assign _2211_ = _2727_ ^ _2723_;
assign _2212_ = _2729_ ^ _2721_;
assign _2213_ = _2731_ ^ _2715_;
assign _2214_ = _0022_[12] ^ _0022_[44];
assign _2215_ = dscratch1_q[12] ^ _0024_[12];
assign _2216_ = _2735_ ^ _2733_;
assign _2217_ = csr_depc_o[12] ^ dscratch0_q[12];
assign _2218_ = csr_mtval_o[12] ^ dcsr_q[12];
assign _2219_ = _2741_ ^ _2739_;
assign _2220_ = _2743_ ^ _2737_;
assign _2221_ = csr_mepc_o[12] ^ _3270_[7];
assign _2222_ = mscratch_q[12] ^ csr_mtvec_o[12];
assign _2223_ = _2749_ ^ _2747_;
assign _2224_ = _2755_ ^ _2753_;
assign _2225_ = _2757_ ^ _2751_;
assign _2226_ = _2759_ ^ _2745_;
assign _2227_ = _0022_[17] ^ _0022_[49];
assign _2228_ = dscratch1_q[17] ^ _0024_[17];
assign _2229_ = _2763_ ^ _2761_;
assign _2230_ = csr_depc_o[17] ^ dscratch0_q[17];
assign _2231_ = irq_fast_i[1] ^ dcsr_q[17];
assign _2232_ = _2769_ ^ _2767_;
assign _2233_ = _2771_ ^ _2765_;
assign _2234_ = _3270_[12] ^ csr_mtval_o[17];
assign _2235_ = csr_mtvec_o[17] ^ csr_mepc_o[17];
assign _2236_ = _2777_ ^ _2775_;
assign _2237_ = mie_q[1] ^ mscratch_q[17];
assign _2238_ = _2783_ ^ mstatus_q[1];
assign _2239_ = _2785_ ^ _2781_;
assign _2240_ = _2787_ ^ _2779_;
assign _2241_ = _2789_ ^ _2773_;
assign _2242_ = _0024_[15:13] ^ _0022_[15:13];
assign _2243_ = _2791_ ^ _0022_[47:45];
assign _2244_ = dscratch0_q[15:13] ^ dscratch1_q[15:13];
assign _2245_ = dcsr_q[15:13] ^ csr_depc_o[15:13];
assign _2246_ = _2797_ ^ _2795_;
assign _2247_ = _2799_ ^ _2793_;
assign _2248_ = csr_mepc_o[15:13] ^ _3270_[10:8];
assign _2249_ = _2803_ ^ csr_mtval_o[15:13];
assign _2250_ = mscratch_q[15:13] ^ csr_mtvec_o[15:13];
assign _2251_ = _2809_ ^ _2807_;
assign _2252_ = _2811_ ^ _2805_;
assign _2253_ = _2813_ ^ _2801_;
assign _2254_ = _0022_[16] ^ _0022_[48];
assign _2255_ = dscratch1_q[16] ^ _0024_[16];
assign _2256_ = _2817_ ^ _2815_;
assign _2257_ = csr_depc_o[16] ^ dscratch0_q[16];
assign _2258_ = irq_fast_i[0] ^ dcsr_q[16];
assign _2259_ = _2823_ ^ _2821_;
assign _2260_ = _2825_ ^ _2819_;
assign _2261_ = _3270_[11] ^ csr_mtval_o[16];
assign _2262_ = csr_mtvec_o[16] ^ csr_mepc_o[16];
assign _2263_ = _2831_ ^ _2829_;
assign _2264_ = mie_q[0] ^ mscratch_q[16];
assign _2265_ = _2837_ ^ _2835_;
assign _2266_ = _2839_ ^ _2833_;
assign _2267_ = _2841_ ^ _2827_;
assign _2268_ = _0022_[30:22] ^ _0022_[62:54];
assign _2269_ = dscratch1_q[30:22] ^ _0024_[30:22];
assign _2270_ = _2845_ ^ _2843_;
assign _2271_ = csr_depc_o[30:22] ^ dscratch0_q[30:22];
assign _2272_ = irq_fast_i[14:6] ^ dcsr_q[30:22];
assign _2273_ = _2851_ ^ _2849_;
assign _2274_ = _2853_ ^ _2847_;
assign _2275_ = _3270_[25:17] ^ csr_mtval_o[30:22];
assign _2276_ = csr_mtvec_o[30:22] ^ csr_mepc_o[30:22];
assign _2277_ = _2859_ ^ _2857_;
assign _2278_ = mie_q[14:6] ^ mscratch_q[30:22];
assign _2280_ = _2867_ ^ _2863_;
assign _2281_ = _2869_ ^ _2861_;
assign _2282_ = _2871_ ^ _2855_;
assign _2283_ = _0022_[11] ^ _0022_[43];
assign _2284_ = dscratch1_q[11] ^ _0024_[11];
assign _2285_ = _2875_ ^ _2873_;
assign _2286_ = csr_depc_o[11] ^ dscratch0_q[11];
assign _2287_ = irq_external_i ^ dcsr_q[11];
assign _2288_ = _2881_ ^ _2879_;
assign _2289_ = _2883_ ^ _2877_;
assign _2290_ = _3270_[6] ^ csr_mtval_o[11];
assign _2291_ = csr_mtvec_o[11] ^ csr_mepc_o[11];
assign _2292_ = _2889_ ^ _2887_;
assign _2293_ = mie_q[15] ^ mscratch_q[11];
assign _2294_ = _2895_ ^ mstatus_q[2];
assign _2295_ = _2897_ ^ _2893_;
assign _2296_ = _2899_ ^ _2891_;
assign _2297_ = _2901_ ^ _2885_;
assign _2298_ = \mhpmcounter[0]  ^ \mhpmcounter[2] ;
assign _2300_ = _0022_[21] ^ _0022_[53];
assign _2301_ = dscratch1_q[21] ^ _0024_[21];
assign _2302_ = _2906_ ^ _2904_;
assign _2303_ = csr_depc_o[21] ^ dscratch0_q[21];
assign _2304_ = irq_fast_i[5] ^ dcsr_q[21];
assign _2305_ = _2912_ ^ _2910_;
assign _2306_ = _2914_ ^ _2908_;
assign _2307_ = _3270_[16] ^ csr_mtval_o[21];
assign _2308_ = csr_mtvec_o[21] ^ csr_mepc_o[21];
assign _2309_ = _2920_ ^ _2918_;
assign _2310_ = mie_q[5] ^ mscratch_q[21];
assign _2311_ = _2926_ ^ mstatus_q[0];
assign _2312_ = _2928_ ^ _2924_;
assign _2313_ = _2930_ ^ _2922_;
assign _2314_ = _2932_ ^ _2916_;
assign _2315_ = _3105_ ^ _0145_;
assign _2316_ = _2934_ ^ csr_wdata_i;
assign _2317_ = _0024_[31] ^ _0022_[31];
assign _2318_ = _2936_ ^ _0022_[63];
assign _2319_ = dscratch0_q[31] ^ dscratch1_q[31];
assign _2320_ = dcsr_q[31] ^ csr_depc_o[31];
assign _2321_ = _2942_ ^ _2940_;
assign _2322_ = _2944_ ^ _2938_;
assign _2323_ = csr_mepc_o[31] ^ _3103_;
assign _2324_ = _2948_ ^ csr_mtval_o[31];
assign _2325_ = mscratch_q[31] ^ csr_mtvec_o[31];
assign _2326_ = _2954_ ^ _2952_;
assign _2327_ = _2956_ ^ _2950_;
assign _2328_ = _2958_ ^ _2946_;
assign _2329_ = _0022_[39] ^ cpuctrlsts_part_q[7];
assign _2330_ = _0024_[7] ^ _0022_[7];
assign _2331_ = _2962_ ^ _2960_;
assign _2332_ = dscratch0_q[7] ^ dscratch1_q[7];
assign _2333_ = irq_timer_i ^ dcsr_q[7];
assign _2334_ = _2968_ ^ csr_depc_o[7];
assign _2335_ = _2970_ ^ _2966_;
assign _2336_ = _2972_ ^ _2964_;
assign _2337_ = _3270_[2] ^ csr_mtval_o[7];
assign _2338_ = csr_mtvec_o[7] ^ csr_mepc_o[7];
assign _2339_ = _2978_ ^ _2976_;
assign _2340_ = mie_q[16] ^ mscratch_q[7];
assign _2341_ = _2984_ ^ mstatus_q[4];
assign _2342_ = _2986_ ^ _2982_;
assign _2343_ = _2988_ ^ _2980_;
assign _2344_ = _2990_ ^ _2974_;
assign _2345_ = _0022_[38:36] ^ cpuctrlsts_part_q[6:4];
assign _2346_ = _0024_[6:4] ^ _0022_[6:4];
assign _2347_ = _2994_ ^ _2992_;
assign _2348_ = dscratch0_q[6:4] ^ dscratch1_q[6:4];
assign _2349_ = dcsr_q[6:4] ^ csr_depc_o[6:4];
assign _2350_ = _3000_ ^ _2998_;
assign _2351_ = _3002_ ^ _2996_;
assign _2352_ = { _3270_[1:0], mcause_q[4] } ^ csr_mtval_o[6:4];
assign _2353_ = csr_mtvec_o[6:4] ^ csr_mepc_o[6:4];
assign _2354_ = _3008_ ^ _3006_;
assign _2355_ = hart_id_i[6:4] ^ mscratch_q[6:4];
assign _2356_ = _3014_ ^ _3012_;
assign _2357_ = _3015_ ^ _3010_;
assign _2358_ = _3017_ ^ _3004_;
assign _2360_ = _0000_[7] ^ _0088_[1];
assign _2361_ = { dummy_instr_seed_o[31:1], 1'h0 } ^ mstack_epc_q;
assign _2362_ = _0016_[4:2] ^ _0143_;
assign _2363_ = _3112_ ^ _0016_[4:2];
assign _2364_ = _3114_ ^ _0119_[2:0];
assign _2365_ = _0016_[1] ^ _0141_;
assign _2366_ = _3116_ ^ _0016_[1];
assign _2367_ = _3118_ ^ _0016_[1];
assign _2368_ = _0016_[5] ^ mstatus_q[4];
assign _2369_ = _3120_ ^ _0016_[5];
assign _2370_ = _3122_ ^ _0119_[3];
assign _2371_ = _0127_ ^ _0002_;
assign _2372_ = _0125_ ^ _0000_[7:6];
assign _2373_ = csr_mcause_i ^ { _3064_, _3062_, dummy_instr_seed_o[4:0] };
assign _2374_ = _0043_ ^ { dummy_instr_seed_o[31:1], 1'h0 };
assign _2375_ = _0137_ ^ _0000_[7];
assign _2376_ = priv_mode_id_o ^ _0016_[3:2];
assign _2377_ = mstatus_q[5] ^ _0016_[4];
assign _2378_ = csr_mtval_i ^ dummy_instr_seed_o;
assign _2379_ = _0004_[8:6] ^ debug_cause_i;
assign _2380_ = _0004_[1:0] ^ priv_mode_id_o;
assign _2381_ = _0112_ ^ _0002_;
assign _2382_ = _0110_ ^ _0000_[7:6];
assign _2383_ = _0123_ ^ _0020_;
assign _2384_ = _0086_ ^ dummy_instr_seed_o;
assign _2385_ = _0115_ ^ _0012_;
assign _2386_ = _0079_ ^ { _3064_, _3062_, dummy_instr_seed_o[4:0] };
assign _2387_ = _0117_ ^ _0014_;
assign _2388_ = _0081_ ^ { dummy_instr_seed_o[31:1], 1'h0 };
assign _2389_ = _0121_ ^ _0018_;
assign _2390_ = _0135_ ^ _0016_[5:2];
assign _2391_ = pc_id_i ^ pc_wb_i;
assign _2392_ = _3124_ ^ pc_id_i;
assign _2393_ = _3126_ ^ pc_if_i;
assign _2394_ = _3128_ ^ _0002_;
assign _2395_ = _3130_ ^ _0090_;
assign _2396_ = _3132_ ^ _0000_[6];
assign _2397_ = _3134_ ^ _0088_[0];
assign _2398_ = _0008_ ^ _0094_;
assign _2399_ = { dummy_instr_seed_o[31:1], 1'h0 } ^ _0033_;
assign _2400_ = _0006_ ^ _0092_;
assign _2401_ = _0004_[8:6] ^ _0139_;
assign _2402_ = _0004_[1:0] ^ _0129_;
assign _2403_ = _0020_ ^ _0108_;
assign _2404_ = dummy_instr_seed_o ^ _0069_;
assign _2405_ = _0012_ ^ _0131_;
assign _2406_ = _3136_ ^ _0012_;
assign _2407_ = _3138_ ^ _0100_;
assign _2408_ = { _3064_, _3062_, dummy_instr_seed_o[4:0] } ^ _0098_;
assign _2409_ = _3140_ ^ { _3064_, _3062_, dummy_instr_seed_o[4:0] };
assign _2410_ = _3142_ ^ _0045_;
assign _2411_ = _0014_ ^ _0133_;
assign _2412_ = _3144_ ^ _0014_;
assign _2413_ = _3146_ ^ _0104_;
assign _2414_ = { dummy_instr_seed_o[31:1], 1'h0 } ^ _0102_;
assign _2415_ = _3148_ ^ { dummy_instr_seed_o[31:1], 1'h0 };
assign _2416_ = _3150_ ^ _0051_;
assign _2417_ = _3152_ ^ _0018_;
assign _2418_ = _3154_ ^ _0106_;
assign _2419_ = { _3064_, _3062_, dummy_instr_seed_o[4:0] } ^ mstack_cause_q;
assign _2420_ = _3156_ ^ dcsr_q[1:0];
assign _2421_ = mstatus_q[5:4] ^ { dummy_instr_seed_o[3], dummy_instr_seed_o[7] };
assign _2422_ = mstatus_q[3:2] ^ _0084_;
assign _2423_ = dcsr_q[15] ^ dummy_instr_seed_o[15];
assign _2424_ = mstatus_q[1:0] ^ { dummy_instr_seed_o[17], dummy_instr_seed_o[21] };
assign _2425_ = dcsr_q[1:0] ^ _0075_;
assign _2426_ = dcsr_q[2] ^ dummy_instr_seed_o[2];
assign _2427_ = dcsr_q[13:12] ^ dummy_instr_seed_o[13:12];
assign _2428_ = cpuctrlsts_part_q ^ { dummy_instr_seed_o[7:1], 1'h0 };
assign _2430_ = cpuctrlsts_part_q ^ _0025_;
assign _2431_ = dcsr_q ^ { _0029_[31:9], dcsr_q[8:6], _0029_[5:0] };
assign _2432_ = csr_mtvec_init_i ^ _0073_;
assign _2433_ = mstatus_q ^ _0065_;
assign _2434_ = { dummy_instr_seed_o[31:8], 8'h01 } ^ { boot_addr_i[31:8], 8'h01 };
assign _2435_ = priv_mode_id_o ^ mstatus_q[3:2];
assign _2436_ = minstret_raw ^ minstret_next;
assign _0548_ = _0028_ & _2156_;
assign _0550_ = _3169_ & _2157_;
assign _0553_ = _1559_ & _2158_;
assign _0556_ = _0042_ & _2159_;
assign _0559_ = _0032_ & _2160_;
assign _0562_ = _0036_ & _2161_;
assign _0565_ = _1561_ & _2162_;
assign _0568_ = _0426_ & _2163_;
assign _0571_ = _0072_ & _2164_;
assign _0574_ = _0054_ & _2165_;
assign _0577_ = _1563_ & _2166_;
assign _0580_ = _0062_ & _2167_;
assign _0582_ = _3189_ & hart_id_i[3];
assign _0585_ = _0068_ & _2168_;
assign _0588_ = _1565_ & _2169_;
assign _0591_ = _0428_ & _2170_;
assign _0594_ = _0430_ & _2171_;
assign _0597_ = { _0028_, _0028_, _0028_ } & _2172_;
assign _0599_ = { _3169_, _3169_, _3169_ } & _2173_;
assign _0602_ = { _1559_, _1559_, _1559_ } & _2174_;
assign _0605_ = { _0050_, _0050_, _0050_ } & _2175_;
assign _0608_ = { _0036_, _0036_, _0036_ } & _2176_;
assign _0611_ = { _0040_, _0040_, _0040_ } & _2177_;
assign _0614_ = { _1567_, _1567_, _1567_ } & _2178_;
assign _0617_ = { _0426_, _0426_, _0426_ } & _2179_;
assign _0620_ = { _0072_, _0072_, _0072_ } & _2180_;
assign _0623_ = { _0054_, _0054_, _0054_ } & _2181_;
assign _0626_ = { _1563_, _1563_, _1563_ } & _2182_;
assign _0628_ = { _0062_, _0062_, _0062_ } & { _0404_, mscratch_q[1:0] };
assign _0631_ = { _3189_, _3189_, _3189_ } & _2183_;
assign _0634_ = { _1569_, _1569_, _1569_ } & _2184_;
assign _0637_ = { _0428_, _0428_, _0428_ } & _2185_;
assign _0640_ = { _0432_, _0432_, _0432_ } & _2186_;
assign _0642_ = { _3169_, _3169_, _3169_ } & _2187_;
assign _0645_ = { _3165_, _3165_, _3165_ } & _2188_;
assign _0648_ = { _0042_, _0042_, _0042_ } & _2189_;
assign _0651_ = { _0036_, _0036_, _0036_ } & _2190_;
assign _0654_ = { _1561_, _1561_, _1561_ } & _2191_;
assign _0657_ = { _0434_, _0434_, _0434_ } & _2192_;
assign _0660_ = { _0072_, _0072_, _0072_ } & _2193_;
assign _0663_ = { _0054_, _0054_, _0054_ } & _2194_;
assign _0666_ = { _1563_, _1563_, _1563_ } & _2195_;
assign _0668_ = { _0062_, _0062_, _0062_ } & { mscratch_q[10:9], _0405_ };
assign _0670_ = { _3189_, _3189_, _3189_ } & hart_id_i[10:8];
assign _0673_ = { _1569_, _1569_, _1569_ } & _2196_;
assign _0676_ = { _0428_, _0428_, _0428_ } & _2197_;
assign _0679_ = { _0436_, _0436_, _0436_ } & _2198_;
assign _0682_ = { _3165_, _3165_, _3165_ } & _2199_;
assign _0684_ = { _3187_, _3187_, _3187_ } & _2200_;
assign _0687_ = { _1571_, _1571_, _1571_ } & _2201_;
assign _0690_ = { _0040_, _0040_, _0040_ } & _2202_;
assign _0693_ = { _0032_, _0032_, _0032_ } & _2203_;
assign _0696_ = { _1573_, _1573_, _1573_ } & _2204_;
assign _0699_ = { _0438_, _0438_, _0438_ } & _2205_;
assign _0701_ = { _0072_, _0072_, _0072_ } & _2206_;
assign _0704_ = { _0054_, _0054_, _0054_ } & _2207_;
assign _0707_ = { _1563_, _1563_, _1563_ } & _2208_;
assign _0710_ = { _0062_, _0062_, _0062_ } & _2209_;
assign _0712_ = { _3189_, _3189_, _3189_ } & hart_id_i[20:18];
assign _0714_ = { _3257_, _3257_, _3257_ } & { _0406_, _2210_[1:0] };
assign _0717_ = { _1565_, _1565_, _1565_ } & _2211_;
assign _0720_ = { _0428_, _0428_, _0428_ } & _2212_;
assign _0723_ = { _0440_, _0440_, _0440_ } & _2213_;
assign _0726_ = _3165_ & _2214_;
assign _0728_ = _3187_ & _2215_;
assign _0731_ = _1571_ & _2216_;
assign _0734_ = _0040_ & _2217_;
assign _0737_ = _0032_ & _2218_;
assign _0740_ = _1573_ & _2219_;
assign _0743_ = _0438_ & _2220_;
assign _0746_ = _0048_ & _2221_;
assign _0749_ = _3176_ & _2222_;
assign _0752_ = _1575_ & _2223_;
assign _0754_ = _3257_ & _0392_;
assign _0756_ = _3189_ & hart_id_i[12];
assign _0759_ = _1577_ & _2224_;
assign _0762_ = _0442_ & _2225_;
assign _0765_ = _0444_ & _2226_;
assign _0768_ = _3165_ & _2227_;
assign _0770_ = _3187_ & _2228_;
assign _0773_ = _1571_ & _2229_;
assign _0776_ = _0040_ & _2230_;
assign _0779_ = _0032_ & _2231_;
assign _0782_ = _1573_ & _2232_;
assign _0785_ = _0438_ & _2233_;
assign _0788_ = _0072_ & _2234_;
assign _0791_ = _0054_ & _2235_;
assign _0794_ = _1563_ & _2236_;
assign _0797_ = _0062_ & _2237_;
assign _0799_ = _3189_ & hart_id_i[17];
assign _0802_ = _0068_ & _2238_;
assign _0805_ = _1565_ & _2239_;
assign _0808_ = _0428_ & _2240_;
assign _0811_ = _0440_ & _2241_;
assign _0813_ = { _3169_, _3169_, _3169_ } & _2242_;
assign _0816_ = { _3165_, _3165_, _3165_ } & _2243_;
assign _0819_ = { _0042_, _0042_, _0042_ } & _2244_;
assign _0822_ = { _0036_, _0036_, _0036_ } & _2245_;
assign _0825_ = { _1561_, _1561_, _1561_ } & _2246_;
assign _0828_ = { _0434_, _0434_, _0434_ } & _2247_;
assign _0831_ = { _0048_, _0048_, _0048_ } & _2248_;
assign _0834_ = { _0072_, _0072_, _0072_ } & _2249_;
assign _0837_ = { _3176_, _3176_, _3176_ } & _2250_;
assign _0839_ = { _3189_, _3189_, _3189_ } & hart_id_i[15:13];
assign _0842_ = { _1579_, _1579_, _1579_ } & _2251_;
assign _0845_ = { _0446_, _0446_, _0446_ } & _2252_;
assign _0848_ = { _0436_, _0436_, _0436_ } & _2253_;
assign _0851_ = _3165_ & _2254_;
assign _0853_ = _3187_ & _2255_;
assign _0856_ = _1571_ & _2256_;
assign _0859_ = _0040_ & _2257_;
assign _0862_ = _0032_ & _2258_;
assign _0865_ = _1573_ & _2259_;
assign _0868_ = _0438_ & _2260_;
assign _0870_ = _0072_ & _2261_;
assign _0873_ = _0054_ & _2262_;
assign _0876_ = _1563_ & _2263_;
assign _0879_ = _0062_ & _2264_;
assign _0881_ = _3189_ & hart_id_i[16];
assign _0884_ = _1565_ & _2265_;
assign _0887_ = _0428_ & _2266_;
assign _0890_ = _0440_ & _2267_;
assign _0893_ = { _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_ } & _2268_;
assign _0895_ = { _3187_, _3187_, _3187_, _3187_, _3187_, _3187_, _3187_, _3187_, _3187_ } & _2269_;
assign _0898_ = { _1571_, _1571_, _1571_, _1571_, _1571_, _1571_, _1571_, _1571_, _1571_ } & _2270_;
assign _0901_ = { _0040_, _0040_, _0040_, _0040_, _0040_, _0040_, _0040_, _0040_, _0040_ } & _2271_;
assign _0904_ = { _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_ } & _2272_;
assign _0907_ = { _1573_, _1573_, _1573_, _1573_, _1573_, _1573_, _1573_, _1573_, _1573_ } & _2273_;
assign _0910_ = { _0438_, _0438_, _0438_, _0438_, _0438_, _0438_, _0438_, _0438_, _0438_ } & _2274_;
assign _0913_ = { _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_, _0072_ } & _2275_;
assign _0916_ = { _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_ } & _2276_;
assign _0919_ = { _1563_, _1563_, _1563_, _1563_, _1563_, _1563_, _1563_, _1563_, _1563_ } & _2277_;
assign _0922_ = { _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_, _0062_ } & _2278_;
assign _0924_ = { _3189_, _3189_, _3189_, _3189_, _3189_, _3189_, _3189_, _3189_, _3189_ } & hart_id_i[30:22];
assign _0926_ = { _3257_, _3257_, _3257_, _3257_, _3257_, _3257_, _3257_, _3257_, _3257_ } & { _0407_, _2279_[7:0] };
assign _0929_ = { _1565_, _1565_, _1565_, _1565_, _1565_, _1565_, _1565_, _1565_, _1565_ } & _2280_;
assign _0932_ = { _0428_, _0428_, _0428_, _0428_, _0428_, _0428_, _0428_, _0428_, _0428_ } & _2281_;
assign _0935_ = { _0440_, _0440_, _0440_, _0440_, _0440_, _0440_, _0440_, _0440_, _0440_ } & _2282_;
assign _0938_ = _3165_ & _2283_;
assign _0940_ = _3187_ & _2284_;
assign _0943_ = _1571_ & _2285_;
assign _0946_ = _0040_ & _2286_;
assign _0949_ = _0032_ & _2287_;
assign _0952_ = _1573_ & _2288_;
assign _0955_ = _0438_ & _2289_;
assign _0957_ = _0072_ & _2290_;
assign _0960_ = _0054_ & _2291_;
assign _0963_ = _1563_ & _2292_;
assign _0966_ = _0062_ & _2293_;
assign _0968_ = _3189_ & hart_id_i[11];
assign _0971_ = _0068_ & _2294_;
assign _0974_ = _1565_ & _2295_;
assign _0977_ = _0428_ & _2296_;
assign _0980_ = _0440_ & _2297_;
assign _0983_ = { _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_, _3252_ } & _2298_;
assign _0985_ = { _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_ } & _2299_;
assign _0988_ = _3165_ & _2300_;
assign _0990_ = _3187_ & _2301_;
assign _0993_ = _1571_ & _2302_;
assign _0996_ = _0040_ & _2303_;
assign _0999_ = _0032_ & _2304_;
assign _1002_ = _1573_ & _2305_;
assign _1005_ = _0438_ & _2306_;
assign _1007_ = _0072_ & _2307_;
assign _1010_ = _0054_ & _2308_;
assign _1013_ = _1563_ & _2309_;
assign _1016_ = _0062_ & _2310_;
assign _1018_ = _3189_ & hart_id_i[21];
assign _1021_ = _0068_ & _2311_;
assign _1024_ = _1565_ & _2312_;
assign _1027_ = _0428_ & _2313_;
assign _1030_ = _0440_ & _2314_;
assign _1033_ = { _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_, _3067_ } & _2315_;
assign _1036_ = { _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_, _0457_ } & _2316_;
assign _1038_ = _3169_ & _2317_;
assign _1041_ = _3165_ & _2318_;
assign _1044_ = _0042_ & _2319_;
assign _1047_ = _0036_ & _2320_;
assign _1050_ = _1561_ & _2321_;
assign _1053_ = _0434_ & _2322_;
assign _1056_ = _0048_ & _2323_;
assign _1059_ = _0072_ & _2324_;
assign _1062_ = _3176_ & _2325_;
assign _1064_ = _3189_ & hart_id_i[31];
assign _1067_ = _1579_ & _2326_;
assign _1070_ = _0446_ & _2327_;
assign _1073_ = _0436_ & _2328_;
assign _1076_ = _0028_ & _2329_;
assign _1078_ = _3169_ & _2330_;
assign _1081_ = _1559_ & _2331_;
assign _1084_ = _0042_ & _2332_;
assign _1087_ = _0032_ & _2333_;
assign _1090_ = _0036_ & _2334_;
assign _1093_ = _1561_ & _2335_;
assign _1096_ = _0426_ & _2336_;
assign _1098_ = _0072_ & _2337_;
assign _1101_ = _0054_ & _2338_;
assign _1104_ = _1563_ & _2339_;
assign _1107_ = _0062_ & _2340_;
assign _1109_ = _3189_ & hart_id_i[7];
assign _1112_ = _0068_ & _2341_;
assign _1115_ = _1565_ & _2342_;
assign _1118_ = _0428_ & _2343_;
assign _1121_ = _0430_ & _2344_;
assign _1124_ = { _0028_, _0028_, _0028_ } & _2345_;
assign _1126_ = { _3169_, _3169_, _3169_ } & _2346_;
assign _1129_ = { _1559_, _1559_, _1559_ } & _2347_;
assign _1132_ = { _0042_, _0042_, _0042_ } & _2348_;
assign _1135_ = { _0036_, _0036_, _0036_ } & _2349_;
assign _1138_ = { _1561_, _1561_, _1561_ } & _2350_;
assign _1141_ = { _0426_, _0426_, _0426_ } & _2351_;
assign _1144_ = { _0072_, _0072_, _0072_ } & _2352_;
assign _1147_ = { _0054_, _0054_, _0054_ } & _2353_;
assign _1150_ = { _1563_, _1563_, _1563_ } & _2354_;
assign _1153_ = { _0062_, _0062_, _0062_ } & _2355_;
assign _1156_ = { _2153_, _2153_, _2153_ } & _2356_;
assign _1159_ = { _0428_, _0428_, _0428_ } & _2357_;
assign _1162_ = { _0448_, _0448_, _0448_ } & _2358_;
assign _1213_ = csr_save_cause_i_t0 & _2360_;
assign _1215_ = nmi_mode_i_t0 & _0395_;
assign _1218_ = { nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0 } & _2361_;
assign _1220_ = nmi_mode_i_t0 & _0396_;
assign _1222_ = { nmi_mode_i_t0, nmi_mode_i_t0 } & mstack_q[1:0];
assign _1224_ = nmi_mode_i_t0 & _0397_;
assign _1226_ = _3089_ & _0016_[1];
assign _1229_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } & _2362_;
assign _1232_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } & _2363_;
assign _1235_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } & _2364_;
assign _1238_ = csr_restore_mret_i_t0 & _2365_;
assign _1241_ = csr_restore_dret_i_t0 & _2366_;
assign _1244_ = csr_save_cause_i_t0 & _2367_;
assign _1247_ = csr_restore_mret_i_t0 & _2368_;
assign _1250_ = csr_restore_dret_i_t0 & _2369_;
assign _1253_ = csr_save_cause_i_t0 & _2370_;
assign _1255_ = _3079_ & _0393_;
assign _1257_ = _3079_ & _0114_;
assign _1259_ = cpuctrlsts_part_q_t0[6] & _0394_;
assign _1261_ = _3079_ & _0398_;
assign _1264_ = debug_mode_i_t0 & _2371_;
assign _1267_ = { debug_mode_i_t0, debug_mode_i_t0 } & _2372_;
assign _1269_ = debug_mode_i_t0 & _0096_;
assign _1272_ = { debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0 } & _2373_;
assign _1274_ = debug_mode_i_t0 & _0395_;
assign _1277_ = { debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0 } & _2374_;
assign _1279_ = debug_mode_i_t0 & _0396_;
assign _1282_ = _3079_ & _2375_;
assign _1285_ = { debug_mode_i_t0, debug_mode_i_t0 } & _2376_;
assign _1288_ = debug_mode_i_t0 & _2377_;
assign _1290_ = debug_mode_i_t0 & _0399_;
assign _1293_ = { debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0, debug_mode_i_t0 } & _2378_;
assign _1295_ = debug_mode_i_t0 & _0400_;
assign _1297_ = debug_csr_save_i_t0 & _0401_;
assign _1300_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } & _2374_;
assign _1302_ = debug_csr_save_i_t0 & _0402_;
assign _1305_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } & _2379_;
assign _1308_ = { debug_csr_save_i_t0, debug_csr_save_i_t0 } & _2380_;
assign _1311_ = debug_csr_save_i_t0 & _2381_;
assign _1314_ = { debug_csr_save_i_t0, debug_csr_save_i_t0 } & _2382_;
assign _1316_ = debug_csr_save_i_t0 & _0083_;
assign _1319_ = debug_csr_save_i_t0 & _2383_;
assign _1322_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } & _2384_;
assign _1325_ = debug_csr_save_i_t0 & _2385_;
assign _1328_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } & _2386_;
assign _1331_ = debug_csr_save_i_t0 & _2387_;
assign _1334_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } & _2388_;
assign _1337_ = debug_csr_save_i_t0 & _2389_;
assign _1340_ = { debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0, debug_csr_save_i_t0 } & _2390_;
assign _1342_ = debug_csr_save_i_t0 & _0077_;
assign _1345_ = { csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0, csr_save_wb_i_t0 } & _2391_;
assign _1348_ = { csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0, csr_save_id_i_t0 } & _2392_;
assign _1351_ = { csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0, csr_save_if_i_t0 } & _2393_;
assign _1353_ = csr_restore_mret_i_t0 & _0398_;
assign _1356_ = csr_restore_dret_i_t0 & _2394_;
assign _1359_ = csr_save_cause_i_t0 & _2395_;
assign _1361_ = csr_restore_mret_i_t0 & _0000_[6];
assign _1364_ = csr_restore_dret_i_t0 & _2396_;
assign _1367_ = csr_save_cause_i_t0 & _2397_;
assign _1369_ = csr_save_cause_i_t0 & _0063_;
assign _1372_ = csr_save_cause_i_t0 & _2398_;
assign _1375_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } & _2399_;
assign _1378_ = csr_save_cause_i_t0 & _2400_;
assign _1381_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } & _2401_;
assign _1384_ = { csr_save_cause_i_t0, csr_save_cause_i_t0 } & _2402_;
assign _1387_ = csr_save_cause_i_t0 & _2403_;
assign _1390_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } & _2404_;
assign _1393_ = csr_restore_mret_i_t0 & _2405_;
assign _1396_ = csr_restore_dret_i_t0 & _2406_;
assign _1399_ = csr_save_cause_i_t0 & _2407_;
assign _1402_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } & _2408_;
assign _1405_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } & _2409_;
assign _1408_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } & _2410_;
assign _1411_ = csr_restore_mret_i_t0 & _2411_;
assign _1414_ = csr_restore_dret_i_t0 & _2412_;
assign _1417_ = csr_save_cause_i_t0 & _2413_;
assign _1420_ = { csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0, csr_restore_mret_i_t0 } & _2414_;
assign _1423_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0, csr_restore_dret_i_t0 } & _2415_;
assign _1426_ = { csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0, csr_save_cause_i_t0 } & _2416_;
assign _1428_ = csr_restore_mret_i_t0 & _0399_;
assign _1431_ = csr_restore_dret_i_t0 & _2417_;
assign _1434_ = csr_save_cause_i_t0 & _2418_;
assign _1437_ = { nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0, nmi_mode_i_t0 } & _2419_;
assign _1439_ = csr_save_cause_i_t0 & _0037_;
assign _1442_ = { csr_restore_dret_i_t0, csr_restore_dret_i_t0 } & _2420_;
assign _1444_ = { csr_save_cause_i_t0, csr_save_cause_i_t0 } & _0408_;
assign _1446_ = debug_mode_i_t0 & _0016_[5];
assign _1448_ = { _0032_, _0032_, _0032_, _0032_ } & { dcsr_q[31], _0409_, dcsr_q[29:28] };
assign _1451_ = { _0068_, _0068_ } & _2421_;
assign _1454_ = { _0068_, _0068_ } & _2422_;
assign _1457_ = _0032_ & _2423_;
assign _1459_ = _0032_ & dcsr_q[14];
assign _1461_ = { _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_, _0032_ } & dcsr_q[27:16];
assign _1464_ = { _0068_, _0068_ } & _2424_;
assign _1467_ = { _0032_, _0032_ } & _2425_;
assign _1469_ = _0032_ & dcsr_q[5];
assign _1471_ = _0032_ & dcsr_q[4];
assign _1473_ = _0032_ & dcsr_q[3];
assign _1476_ = _0032_ & _2426_;
assign _1479_ = { _0032_, _0032_ } & _2427_;
assign _1481_ = _0032_ & dcsr_q[11];
assign _1483_ = { _3077_, _3077_ } & dummy_instr_seed_o[1:0];
assign _1485_ = _0032_ & dcsr_q[9];
assign _1487_ = { _3075_, _3075_ } & dummy_instr_seed_o[12:11];
assign _1491_ = { _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_, _0028_ } & _2428_;
assign _1493_ = { _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_, _3165_ } & _2429_;
assign _1495_ = { _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_, _3169_ } & _2429_;
assign _1497_ = _0032_ & dcsr_q[10];
assign _1499_ = _3176_ & _0403_;
assign _1501_ = csr_we_int_t0 & _0027_;
assign _1504_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } & _2430_;
assign _1506_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } & _0057_;
assign _1508_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } & _0055_;
assign _1510_ = csr_we_int_t0 & _0049_;
assign _1512_ = csr_we_int_t0 & _0041_;
assign _1514_ = csr_we_int_t0 & _0039_;
assign _1516_ = csr_we_int_t0 & _0035_;
assign _1518_ = csr_we_int_t0 & _0031_;
assign _1521_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } & _2431_;
assign _1524_ = csr_we_int_t0 & _2432_;
assign _1526_ = csr_we_int_t0 & _0071_;
assign _1528_ = csr_we_int_t0 & _0047_;
assign _1530_ = csr_we_int_t0 & _0053_;
assign _1532_ = csr_we_int_t0 & _0061_;
assign _1534_ = csr_we_int_t0 & _0059_;
assign _1536_ = csr_we_int_t0 & _0067_;
assign _1539_ = { csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0, csr_we_int_t0 } & _2433_;
assign _1541_ = _3183_ & _0391_;
assign _1551_ = { csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0, csr_mtvec_init_i_t0 } & _2434_;
assign _1554_ = { mstatus_q_t0[1], mstatus_q_t0[1] } & _2435_;
assign _1557_ = { _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_, _0153_ } & _2436_;
assign _2614_ = _0548_ | _1611_;
assign _2616_ = _0550_ | _0549_;
assign _2618_ = _0553_ | _1615_;
assign _2620_ = _0556_ | _1618_;
assign _2622_ = _0559_ | _1621_;
assign _2624_ = _0562_ | _1624_;
assign _2626_ = _0565_ | _1627_;
assign _2628_ = _0568_ | _1630_;
assign _2630_ = _0571_ | _1633_;
assign _2632_ = _0574_ | _1636_;
assign _2634_ = _0577_ | _1639_;
assign _2636_ = _0580_ | _1642_;
assign _2638_ = _0582_ | _0581_;
assign _2640_ = _0585_ | _1646_;
assign _2642_ = _0588_ | _1649_;
assign _2644_ = _0591_ | _1652_;
assign csr_rdata_o_t0[3] = _0594_ | _1655_;
assign _2646_ = _0597_ | _1658_;
assign _2648_ = _0599_ | _0598_;
assign _2650_ = _0602_ | _1662_;
assign _2652_ = _0605_ | _1665_;
assign _2654_ = _0608_ | _1668_;
assign _2656_ = _0611_ | _1671_;
assign _2658_ = _0614_ | _1674_;
assign _2660_ = _0617_ | _1677_;
assign _2662_ = _0620_ | _1680_;
assign _2664_ = _0623_ | _1683_;
assign _2666_ = _0626_ | _1686_;
assign _2668_ = _0628_ | _0627_;
assign _2672_ = _0631_ | _1691_;
assign _2674_ = _0634_ | _1694_;
assign _2676_ = _0637_ | _1697_;
assign csr_rdata_o_t0[2:0] = _0640_ | _1700_;
assign _2678_ = _0642_ | _0641_;
assign _2680_ = _0645_ | _1703_;
assign _2682_ = _0648_ | _1706_;
assign _2684_ = _0651_ | _1707_;
assign _2686_ = _0654_ | _1710_;
assign _2688_ = _0657_ | _1713_;
assign _2690_ = _0660_ | _1714_;
assign _2692_ = _0663_ | _1715_;
assign _2694_ = _0666_ | _1716_;
assign _2696_ = _0668_ | _0667_;
assign _2698_ = _0670_ | _0669_;
assign _2700_ = _0673_ | _1717_;
assign _2702_ = _0676_ | _1718_;
assign csr_rdata_o_t0[10:8] = _0679_ | _1721_;
assign _2704_ = _0682_ | _1722_;
assign _2706_ = _0684_ | _0683_;
assign _2708_ = _0687_ | _1726_;
assign _2710_ = _0690_ | _1727_;
assign _2712_ = _0693_ | _1730_;
assign _2714_ = _0696_ | _1733_;
assign _2716_ = _0699_ | _1736_;
assign _2718_ = _0701_ | _1737_;
assign _2720_ = _0704_ | _1738_;
assign _2722_ = _0707_ | _1739_;
assign _2724_ = _0710_ | _1740_;
assign _2726_ = _0712_ | _0711_;
assign _2728_ = _0714_ | _0713_;
assign _2730_ = _0717_ | _1744_;
assign _2732_ = _0720_ | _1745_;
assign csr_rdata_o_t0[20:18] = _0723_ | _1748_;
assign _2734_ = _0726_ | _1751_;
assign _2736_ = _0728_ | _0727_;
assign _2738_ = _0731_ | _1755_;
assign _2740_ = _0734_ | _1758_;
assign _2742_ = _0737_ | _1759_;
assign _2744_ = _0740_ | _1762_;
assign _2746_ = _0743_ | _1765_;
assign _2748_ = _0746_ | _1768_;
assign _2750_ = _0749_ | _1771_;
assign _2752_ = _0752_ | _1774_;
assign _2754_ = _0754_ | _0753_;
assign _2756_ = _0756_ | _0755_;
assign _2758_ = _0759_ | _1778_;
assign _2760_ = _0762_ | _1781_;
assign csr_rdata_o_t0[12] = _0765_ | _1784_;
assign _2762_ = _0768_ | _1785_;
assign _2764_ = _0770_ | _0769_;
assign _2766_ = _0773_ | _1786_;
assign _2768_ = _0776_ | _1787_;
assign _2770_ = _0779_ | _1788_;
assign _2772_ = _0782_ | _1789_;
assign _2774_ = _0785_ | _1790_;
assign _2776_ = _0788_ | _1791_;
assign _2778_ = _0791_ | _1792_;
assign _2780_ = _0794_ | _1793_;
assign _2782_ = _0797_ | _1794_;
assign _2784_ = _0799_ | _0798_;
assign _2786_ = _0802_ | _1795_;
assign _2788_ = _0805_ | _1796_;
assign _2790_ = _0808_ | _1797_;
assign csr_rdata_o_t0[17] = _0811_ | _1800_;
assign _2792_ = _0813_ | _0812_;
assign _2794_ = _0816_ | _1801_;
assign _2796_ = _0819_ | _1802_;
assign _2798_ = _0822_ | _1803_;
assign _2800_ = _0825_ | _1804_;
assign _2802_ = _0828_ | _1805_;
assign _2804_ = _0831_ | _1808_;
assign _2806_ = _0834_ | _1809_;
assign _2808_ = _0837_ | _1812_;
assign _2810_ = _0839_ | _0838_;
assign _2812_ = _0842_ | _1815_;
assign _2814_ = _0845_ | _1818_;
assign csr_rdata_o_t0[15:13] = _0848_ | _1819_;
assign _2816_ = _0851_ | _1820_;
assign _2818_ = _0853_ | _0852_;
assign _2820_ = _0856_ | _1821_;
assign _2822_ = _0859_ | _1822_;
assign _2824_ = _0862_ | _1823_;
assign _2826_ = _0865_ | _1824_;
assign _2828_ = _0868_ | _1825_;
assign _2830_ = _0870_ | _1826_;
assign _2832_ = _0873_ | _1827_;
assign _2834_ = _0876_ | _1828_;
assign _2836_ = _0879_ | _1829_;
assign _2838_ = _0881_ | _0880_;
assign _2840_ = _0884_ | _1830_;
assign _2842_ = _0887_ | _1831_;
assign csr_rdata_o_t0[16] = _0890_ | _1832_;
assign _2844_ = _0893_ | _1835_;
assign _2846_ = _0895_ | _0894_;
assign _2848_ = _0898_ | _1839_;
assign _2850_ = _0901_ | _1842_;
assign _2852_ = _0904_ | _1845_;
assign _2854_ = _0907_ | _1848_;
assign _2856_ = _0910_ | _1851_;
assign _2858_ = _0913_ | _1854_;
assign _2860_ = _0916_ | _1857_;
assign _2862_ = _0919_ | _1860_;
assign _2864_ = _0922_ | _1863_;
assign _2866_ = _0924_ | _0923_;
assign _2868_ = _0926_ | _0925_;
assign _2870_ = _0929_ | _1868_;
assign _2872_ = _0932_ | _1871_;
assign csr_rdata_o_t0[30:22] = _0935_ | _1874_;
assign _2874_ = _0938_ | _1875_;
assign _2876_ = _0940_ | _0939_;
assign _2878_ = _0943_ | _1876_;
assign _2880_ = _0946_ | _1877_;
assign _2882_ = _0949_ | _1878_;
assign _2884_ = _0952_ | _1879_;
assign _2886_ = _0955_ | _1880_;
assign _2888_ = _0957_ | _1881_;
assign _2890_ = _0960_ | _1882_;
assign _2892_ = _0963_ | _1883_;
assign _2894_ = _0966_ | _1884_;
assign _2896_ = _0968_ | _0967_;
assign _2898_ = _0971_ | _1885_;
assign _2900_ = _0974_ | _1886_;
assign _2902_ = _0977_ | _1887_;
assign csr_rdata_o_t0[11] = _0980_ | _1888_;
assign _2903_ = _0983_ | _1891_;
assign _0023_ = _0985_ | _0984_;
assign _2905_ = _0988_ | _1893_;
assign _2907_ = _0990_ | _0989_;
assign _2909_ = _0993_ | _1894_;
assign _2911_ = _0996_ | _1895_;
assign _2913_ = _0999_ | _1896_;
assign _2915_ = _1002_ | _1897_;
assign _2917_ = _1005_ | _1898_;
assign _2919_ = _1007_ | _1899_;
assign _2921_ = _1010_ | _1900_;
assign _2923_ = _1013_ | _1901_;
assign _2925_ = _1016_ | _1902_;
assign _2927_ = _1018_ | _1017_;
assign _2929_ = _1021_ | _1903_;
assign _2931_ = _1024_ | _1904_;
assign _2933_ = _1027_ | _1905_;
assign csr_rdata_o_t0[21] = _1030_ | _1906_;
assign _2935_ = _1033_ | _1909_;
assign dummy_instr_seed_o_t0 = _1036_ | _1912_;
assign _2937_ = _1038_ | _1037_;
assign _2939_ = _1041_ | _1913_;
assign _2941_ = _1044_ | _1914_;
assign _2943_ = _1047_ | _1915_;
assign _2945_ = _1050_ | _1916_;
assign _2947_ = _1053_ | _1919_;
assign _2949_ = _1056_ | _1920_;
assign _2951_ = _1059_ | _1921_;
assign _2953_ = _1062_ | _1922_;
assign _2955_ = _1064_ | _1063_;
assign _2957_ = _1067_ | _1925_;
assign _2959_ = _1070_ | _1928_;
assign csr_rdata_o_t0[31] = _1073_ | _1931_;
assign _2961_ = _1076_ | _1932_;
assign _2963_ = _1078_ | _1077_;
assign _2965_ = _1081_ | _1933_;
assign _2967_ = _1084_ | _1934_;
assign _2969_ = _1087_ | _1935_;
assign _2971_ = _1090_ | _1936_;
assign _2973_ = _1093_ | _1937_;
assign _2975_ = _1096_ | _1938_;
assign _2977_ = _1098_ | _1939_;
assign _2979_ = _1101_ | _1940_;
assign _2981_ = _1104_ | _1941_;
assign _2983_ = _1107_ | _1942_;
assign _2985_ = _1109_ | _1108_;
assign _2987_ = _1112_ | _1943_;
assign _2989_ = _1115_ | _1944_;
assign _2991_ = _1118_ | _1945_;
assign csr_rdata_o_t0[7] = _1121_ | _1946_;
assign _2993_ = _1124_ | _1947_;
assign _2995_ = _1126_ | _1125_;
assign _2997_ = _1129_ | _1948_;
assign _2999_ = _1132_ | _1949_;
assign _3001_ = _1135_ | _1950_;
assign _3003_ = _1138_ | _1951_;
assign _3005_ = _1141_ | _1952_;
assign _3007_ = _1144_ | _1953_;
assign _3009_ = _1147_ | _1954_;
assign _3011_ = _1150_ | _1955_;
assign _3013_ = _1153_ | _1956_;
assign _3016_ = _1156_ | _1959_;
assign _3018_ = _1159_ | _1960_;
assign csr_rdata_o_t0[6:4] = _1162_ | _1963_;
assign cpuctrlsts_part_d_t0[7] = _1213_ | _1984_;
assign _0132_ = _1215_ | _1214_;
assign _0103_ = _1218_ | _1989_;
assign _0134_ = _1220_ | _1219_;
assign _0144_[1:0] = _1222_ | _1221_;
assign _0144_[2] = _1224_ | _1223_;
assign _0142_ = _1226_ | _1225_;
assign _3113_ = _1229_ | _1994_;
assign _3115_ = _1232_ | _1997_;
assign mstatus_d_t0[4:2] = _1235_ | _2000_;
assign _3117_ = _1238_ | _2003_;
assign _3119_ = _1241_ | _2006_;
assign mstatus_d_t0[1] = _1244_ | _2007_;
assign _3121_ = _1247_ | _2008_;
assign _3123_ = _1250_ | _2009_;
assign mstatus_d_t0[5] = _1253_ | _2010_;
assign _0126_[0] = _1255_ | _1254_;
assign _0097_ = _1257_ | _1256_;
assign _0138_ = _1259_ | _1258_;
assign _0128_ = _1261_ | _1260_;
assign _0113_ = _1264_ | _2016_;
assign _0111_ = _1267_ | _2019_;
assign _0078_ = _1269_ | _1268_;
assign _0080_ = _1272_ | _2022_;
assign _0116_ = _1274_ | _1273_;
assign _0082_ = _1277_ | _2025_;
assign _0118_ = _1279_ | _1278_;
assign _0126_[1] = _1282_ | _2026_;
assign _0136_[1:0] = _1285_ | _2027_;
assign _0136_[2] = _1288_ | _2028_;
assign _0122_ = _1290_ | _1289_;
assign _0087_ = _1293_ | _2029_;
assign _0124_ = _1295_ | _1294_;
assign _0095_ = _1297_ | _1296_;
assign _0034_ = _1300_ | _2034_;
assign _0093_ = _1302_ | _1301_;
assign _0140_ = _1305_ | _2037_;
assign _0130_ = _1308_ | _2040_;
assign _0091_ = _1311_ | _2041_;
assign _0089_ = _1314_ | _2042_;
assign _0064_ = _1316_ | _1315_;
assign _0109_ = _1319_ | _2043_;
assign _0070_ = _1322_ | _2044_;
assign _0101_ = _1325_ | _2045_;
assign _0046_ = _1328_ | _2048_;
assign _0105_ = _1331_ | _2049_;
assign _0052_ = _1334_ | _2050_;
assign _0107_ = _1337_ | _2051_;
assign _0120_ = _1340_ | _2054_;
assign _0038_ = _1342_ | _1341_;
assign _3125_ = _1345_ | _2057_;
assign _3127_ = _1348_ | _2060_;
assign _0044_ = _1351_ | _2063_;
assign _3129_ = _1353_ | _1352_;
assign _3131_ = _1356_ | _2064_;
assign cpuctrlsts_part_we_t0 = _1359_ | _2065_;
assign _3133_ = _1361_ | _1360_;
assign _3135_ = _1364_ | _2066_;
assign cpuctrlsts_part_d_t0[6] = _1367_ | _2067_;
assign mstack_en_t0 = _1369_ | _1368_;
assign depc_en_t0 = _1372_ | _2068_;
assign depc_d_t0 = _1375_ | _2071_;
assign dcsr_en_t0 = _1378_ | _2072_;
assign dcsr_d_t0[8:6] = _1381_ | _2073_;
assign dcsr_d_t0[1:0] = _1384_ | _2076_;
assign mtval_en_t0 = _1387_ | _2077_;
assign mtval_d_t0 = _1390_ | _2078_;
assign _3137_ = _1393_ | _2079_;
assign _3139_ = _1396_ | _2080_;
assign mcause_en_t0 = _1399_ | _2081_;
assign _3141_ = _1402_ | _2084_;
assign _3143_ = _1405_ | _2087_;
assign mcause_d_t0 = _1408_ | _2090_;
assign _3145_ = _1411_ | _2091_;
assign _3147_ = _1414_ | _2092_;
assign mepc_en_t0 = _1417_ | _2093_;
assign _3149_ = _1420_ | _2096_;
assign _3151_ = _1423_ | _2099_;
assign mepc_d_t0 = _1426_ | _2100_;
assign _3153_ = _1428_ | _1427_;
assign _3155_ = _1431_ | _2101_;
assign mstatus_en_t0 = _1434_ | _2102_;
assign _0099_ = _1437_ | _2105_;
assign double_fault_seen_o_t0 = _1439_ | _1438_;
assign _3159_ = _1442_ | _2109_;
assign priv_lvl_d_t0 = _1444_ | _1443_;
assign _0136_[3] = _1446_ | _1445_;
assign _0030_[31:28] = _1448_ | _1447_;
assign _0066_[5:4] = _1451_ | _2113_;
assign _0066_[3:2] = _1454_ | _2114_;
assign _0030_[15] = _1457_ | _2115_;
assign _0030_[14] = _1459_ | _1458_;
assign _0030_[27:16] = _1461_ | _1460_;
assign _0066_[1:0] = _1464_ | _2117_;
assign _0030_[1:0] = _1467_ | _2120_;
assign _0030_[5] = _1469_ | _1468_;
assign _0030_[4] = _1471_ | _1470_;
assign _0030_[3] = _1473_ | _1472_;
assign _0030_[2] = _1476_ | _2121_;
assign _0030_[13:12] = _1479_ | _2122_;
assign _0030_[11] = _1481_ | _1480_;
assign _0076_ = _1483_ | _1482_;
assign _0030_[9] = _1485_ | _1484_;
assign _0085_ = _1487_ | _1486_;
assign _0026_ = _1491_ | _2127_;
assign _0058_ = _1493_ | _1492_;
assign _0056_ = _1495_ | _1494_;
assign _0030_[10] = _1497_ | _1496_;
assign _0074_ = _1499_ | _1498_;
assign _0003_ = _1501_ | _1500_;
assign { _0001_[7:6], cpuctrlsts_part_d_t0[5:0] } = _1504_ | _2134_;
assign mhpmcounterh_we_t0 = _1506_ | _1505_;
assign mhpmcounter_we_t0 = _1508_ | _1507_;
assign mcountinhibit_we_t0 = _1510_ | _1509_;
assign dscratch1_en_t0 = _1512_ | _1511_;
assign dscratch0_en_t0 = _1514_ | _1513_;
assign _0009_ = _1516_ | _1515_;
assign _0007_ = _1518_ | _1517_;
assign { dcsr_d_t0[31:9], _0005_[8:6], dcsr_d_t0[5:2], _0005_[1:0] } = _1521_ | _2137_;
assign mtvec_en_t0 = _1524_ | _2138_;
assign _0021_ = _1526_ | _1525_;
assign _0013_ = _1528_ | _1527_;
assign _0015_ = _1530_ | _1529_;
assign mscratch_en_t0 = _1532_ | _1531_;
assign mie_en_t0 = _1534_ | _1533_;
assign _0019_ = _1536_ | _1535_;
assign { _0017_[5:1], mstatus_d_t0[0] } = _1539_ | _2141_;
assign illegal_csr_t0 = _1541_ | _1540_;
assign mtvec_d_t0 = _1551_ | _2145_;
assign priv_mode_lsu_o_t0 = _1554_ | _2148_;
assign \mhpmcounter[2]_t0  = _1557_ | _2151_;
assign _0388_ = ~ { 27'h0000000, csr_addr_i_t0[4:0] };
assign _1187_ = { 27'h0000000, csr_addr_i[4:0] } & _0388_;
assign _1973_ = { 27'h0000000, csr_addr_i[4:0] } | { 27'h0000000, csr_addr_i_t0[4:0] };
assign _0389_ = - _1187_;
assign _0390_ = - _1973_;
assign _2359_ = _0389_ ^ _0390_;
assign _3091_ = _2359_ | { 27'h0000000, csr_addr_i_t0[4:0] };
assign _0452_ = | { csr_save_cause_i, csr_restore_dret_i, csr_restore_mret_i };
assign _0392_ = ~ mstatus_q[3];
assign _0393_ = ~ _0000_[6];
assign _0394_ = ~ _0000_[7];
assign _0395_ = ~ _0012_;
assign _0396_ = ~ _0014_;
assign _0397_ = ~ mstack_q[2];
assign _0398_ = ~ _0002_;
assign _0399_ = ~ _0018_;
assign _0400_ = ~ _0020_;
assign _0401_ = ~ _0008_;
assign _0402_ = ~ _0006_;
assign _0403_ = ~ csr_mtvec_init_i;
assign _0404_ = ~ mscratch_q[2];
assign _0405_ = ~ mscratch_q[8];
assign _0406_ = ~ _2725_[2];
assign _0407_ = ~ _2865_[8];
assign _0408_ = ~ _3158_;
assign _0409_ = ~ dcsr_q[30];
assign _0391_ = | { _3268_, _3266_, _3264_, _3262_, _3260_, _3258_, _3256_, _3192_, _3190_, _3188_, _3184_, _3181_, _3180_, _3179_, _3178_, _3177_, _3175_, _3174_, _3173_, _3172_, _3171_, _3170_, _3166_, _3162_, _3161_, _3160_, _3072_, _3060_, _3058_, _3056_, _3054_, _3052_, _3050_, _3048_, _3046_, _3044_, _3042_, _3040_, _3038_, _3036_, _3034_, _3032_, _3030_, _3028_, _3026_, _3024_, _3022_ };
assign _0454_ = | { _3255_, _3253_, _3251_, _3249_, _3247_, _3245_, _3243_, _3241_, _3239_, _3237_, _3235_, _3233_, _3231_, _3229_, _3227_, _3225_, _3223_, _3221_, _3219_, _3217_, _3215_, _3213_, _3211_, _3209_, _3207_, _3205_, _3203_, _3201_, _3199_, _3197_, _3195_, _3193_ };
assign _0455_ = | { _3174_, _3173_, _3172_, _3160_ };
assign _0456_ = | { _3070_, _3110_ };
assign _0458_ = | { _3253_, _3249_, _3247_, _3245_, _3243_, _3241_, _3239_, _3237_, _3235_, _3233_, _3231_, _3229_, _3227_, _3225_, _3223_, _3221_, _3219_, _3217_, _3215_, _3213_, _3211_, _3209_, _3207_, _3205_, _3203_, _3201_, _3199_, _3197_, _3195_, _3193_ };
assign _0410_ = ~ illegal_csr;
assign _0411_ = ~ _3097_;
assign _0412_ = ~ _3099_;
assign _0413_ = ~ mcause_q[5];
assign _0414_ = ~ csr_wdata_i;
assign _0415_ = ~ mstatus_err;
assign _0416_ = ~ _3108_;
assign _0417_ = ~ illegal_csr_write;
assign _0418_ = ~ illegal_csr_priv;
assign _0419_ = ~ illegal_csr_dbg;
assign _0420_ = ~ mcause_q[6];
assign _0421_ = ~ csr_rdata_o;
assign _0422_ = ~ debug_mode_entering_i;
assign _0423_ = ~ mtvec_err;
assign _0424_ = ~ cpuctrlsts_part_err;
assign _0498_ = _3165_ & _0250_;
assign _0501_ = _0042_ & _0378_;
assign _0504_ = _3257_ & _0261_;
assign _0507_ = _0054_ & _0301_;
assign _0510_ = _0068_ & _0304_;
assign _0513_ = _0040_ & _0253_;
assign _0516_ = _0062_ & _0302_;
assign _0519_ = _3169_ & _0295_;
assign _0522_ = _0036_ & _0298_;
assign _0525_ = _0048_ & _0258_;
assign _0528_ = _0060_ & _0261_;
assign _0531_ = _3189_ & _0261_;
assign _1188_ = illegal_csr_t0 & _0417_;
assign _1191_ = _3098_ & _0418_;
assign _1194_ = _3100_ & _0419_;
assign _1197_ = mcause_q_t0[5] & _0420_;
assign _1200_ = csr_wdata_i_t0 & _0421_;
assign _1201_ = debug_mode_i_t0 & _0422_;
assign _1204_ = mstatus_err_t0 & _0423_;
assign _1207_ = _3109_ & _0424_;
assign _0499_ = _0028_ & _0295_;
assign _0502_ = _0050_ & _0253_;
assign _0505_ = _0062_ & _0304_;
assign _0508_ = _0048_ & _0259_;
assign _0511_ = _3257_ & _0263_;
assign _0514_ = _0042_ & _0298_;
assign _0517_ = _3176_ & _0261_;
assign _0520_ = _3165_ & _0251_;
assign _0523_ = _0040_ & _0255_;
assign _0526_ = _0072_ & _0301_;
assign _0529_ = _0062_ & _0379_;
assign _0532_ = _0062_ & _0262_;
assign _1189_ = illegal_csr_write_t0 & _0410_;
assign _1192_ = illegal_csr_priv_t0 & _0411_;
assign _1195_ = illegal_csr_dbg_t0 & _0412_;
assign _1198_ = mcause_q_t0[6] & _0413_;
assign _1202_ = debug_mode_entering_i_t0 & _0349_;
assign _1205_ = mtvec_err_t0 & _0415_;
assign _1208_ = cpuctrlsts_part_err_t0 & _0416_;
assign _0500_ = _3165_ & _0028_;
assign _0503_ = _0042_ & _0050_;
assign _0506_ = _3257_ & _0062_;
assign _0509_ = _0054_ & _0048_;
assign _0512_ = _0068_ & _3257_;
assign _0515_ = _0040_ & _0042_;
assign _0518_ = _0062_ & _3176_;
assign _0521_ = _3169_ & _3165_;
assign _0524_ = _0036_ & _0040_;
assign _0527_ = _0048_ & _0072_;
assign _0530_ = _0060_ & _0062_;
assign _0533_ = _3189_ & _0062_;
assign _1190_ = illegal_csr_t0 & illegal_csr_write_t0;
assign _1193_ = _3098_ & illegal_csr_priv_t0;
assign _1196_ = _3100_ & illegal_csr_dbg_t0;
assign _1199_ = mcause_q_t0[5] & mcause_q_t0[6];
assign _1203_ = debug_mode_i_t0 & debug_mode_entering_i_t0;
assign _1206_ = mstatus_err_t0 & mtvec_err_t0;
assign _1209_ = _3109_ & cpuctrlsts_part_err_t0;
assign _1597_ = _0498_ | _0499_;
assign _1598_ = _0501_ | _0502_;
assign _1599_ = _0504_ | _0505_;
assign _1600_ = _0507_ | _0508_;
assign _1601_ = _0510_ | _0511_;
assign _1602_ = _0513_ | _0514_;
assign _1603_ = _0516_ | _0517_;
assign _1604_ = _0519_ | _0520_;
assign _1605_ = _0522_ | _0523_;
assign _1606_ = _0525_ | _0526_;
assign _1607_ = _0528_ | _0529_;
assign _1608_ = _0531_ | _0532_;
assign _1974_ = _1188_ | _1189_;
assign _1975_ = _1191_ | _1192_;
assign _1976_ = _1194_ | _1195_;
assign _1977_ = _1197_ | _1198_;
assign _1978_ = _1200_ | _0467_;
assign _1979_ = _1201_ | _1202_;
assign _1980_ = _1204_ | _1205_;
assign _1981_ = _1207_ | _1208_;
assign _1559_ = _1597_ | _0500_;
assign _1567_ = _1598_ | _0503_;
assign _1569_ = _1599_ | _0506_;
assign _1575_ = _1600_ | _0509_;
assign _1577_ = _1601_ | _0512_;
assign _1561_ = _1602_ | _0515_;
assign _1579_ = _1603_ | _0518_;
assign _1571_ = _1604_ | _0521_;
assign _1573_ = _1605_ | _0524_;
assign _1563_ = _1606_ | _0527_;
assign _1565_ = _1607_ | _0530_;
assign _2153_ = _1608_ | _0533_;
assign _3098_ = _1974_ | _1190_;
assign _3100_ = _1975_ | _1193_;
assign _3102_ = _1976_ | _1196_;
assign _3104_ = _1977_ | _1199_;
assign _3106_ = _1978_ | _0468_;
assign _3095_ = _1979_ | _1203_;
assign _3109_ = _1980_ | _1206_;
assign csr_shadow_err_o_t0 = _1981_ | _1209_;
assign _1558_ = _3164_ | _3170_;
assign _1566_ = _3172_ | _3171_;
assign _1568_ = _3256_ | _3180_;
assign _1574_ = _3179_ | _3178_;
assign _1576_ = _3161_ | _3256_;
assign _1560_ = _3173_ | _3172_;
assign _1578_ = _3180_ | _3175_;
assign _1570_ = _3168_ | _3164_;
assign _1572_ = _3174_ | _3173_;
assign _1562_ = _3178_ | _3177_;
assign _1564_ = _3181_ | _3180_;
assign _2152_ = _3188_ | _3180_;
assign _0429_ = | { _1558_, _1560_, _3190_, _3184_, _3174_, _3166_, _3160_ };
assign _0425_ = | { _1558_, _3184_, _3166_ };
assign _0431_ = | { _1558_, _1566_, _3184_, _3174_, _3173_, _3166_, _3160_ };
assign _0441_ = | { _3180_, _3175_, _1574_ };
assign _0443_ = | { _1570_, _1572_, _3184_, _3177_, _3172_, _3160_ };
assign _0439_ = | { _1570_, _1572_, _3190_, _3184_, _3172_, _3160_ };
assign _0433_ = | { _3184_, _3166_, _3162_ };
assign _0445_ = | { _3179_, _3178_, _3177_ };
assign _0435_ = | { _1560_, _3184_, _3174_, _3166_, _3162_, _3160_ };
assign _0437_ = | { _1570_, _3184_, _3172_ };
assign _0427_ = | { _1562_, _3179_, _3175_ };
assign _0447_ = | { _1558_, _1560_, _3184_, _3174_, _3166_, _3160_ };
assign _2613_ = _3170_ ? cpuctrlsts_part_q[3] : _0022_[35];
assign _2615_ = _3168_ ? _0022_[3] : _0024_[3];
assign _2617_ = _1558_ ? _2613_ : _2615_;
assign _2619_ = _3172_ ? dscratch1_q[3] : dscratch0_q[3];
assign _2621_ = _3160_ ? dcsr_q[3] : irq_software_i;
assign _2623_ = _3174_ ? csr_depc_o[3] : _2621_;
assign _2625_ = _1560_ ? _2619_ : _2623_;
assign _2627_ = _0425_ ? _2617_ : _2625_;
assign _2629_ = _3177_ ? csr_mtval_o[3] : mcause_q[3];
assign _2631_ = _3179_ ? csr_mepc_o[3] : csr_mtvec_o[3];
assign _2633_ = _1562_ ? _2629_ : _2631_;
assign _2635_ = _3180_ ? mscratch_q[3] : mie_q[17];
assign _2637_ = _3188_ ? hart_id_i[3] : 1'h0;
assign _2639_ = _3161_ ? mstatus_q[5] : _2637_;
assign _2641_ = _1564_ ? _2635_ : _2639_;
assign _2643_ = _0427_ ? _2633_ : _2641_;
assign csr_rdata_o[3] = _0429_ ? _2627_ : _2643_;
assign _2645_ = _3170_ ? cpuctrlsts_part_q[2:0] : _0022_[34:32];
assign _2647_ = _3168_ ? _0022_[2:0] : _0024_[2:0];
assign _2649_ = _1558_ ? _2645_ : _2647_;
assign _2651_ = _3171_ ? { mcountinhibit[2], 1'h0, mcountinhibit[0] } : dscratch1_q[2:0];
assign _2653_ = _3174_ ? csr_depc_o[2:0] : dcsr_q[2:0];
assign _2655_ = _3173_ ? dscratch0_q[2:0] : _2653_;
assign _2657_ = _1566_ ? _2651_ : _2655_;
assign _2659_ = _0425_ ? _2649_ : _2657_;
assign _2661_ = _3177_ ? csr_mtval_o[2:0] : mcause_q[2:0];
assign _2663_ = _3179_ ? csr_mepc_o[2:0] : csr_mtvec_o[2:0];
assign _2665_ = _1562_ ? _2661_ : _2663_;
assign _2667_ = _3180_ ? mscratch_q[2:0] : 3'h4;
assign _2669_ = _3192_ ? 3'h6 : 3'h0;
assign _2671_ = _3188_ ? hart_id_i[2:0] : _2669_;
assign _2673_ = _1568_ ? _2667_ : _2671_;
assign _2675_ = _0427_ ? _2665_ : _2673_;
assign csr_rdata_o[2:0] = _0431_ ? _2659_ : _2675_;
assign _2677_ = _3168_ ? _0022_[10:8] : _0024_[10:8];
assign _2679_ = _3164_ ? _0022_[42:40] : _2677_;
assign _2681_ = _3172_ ? dscratch1_q[10:8] : dscratch0_q[10:8];
assign _2683_ = _3174_ ? csr_depc_o[10:8] : dcsr_q[10:8];
assign _2685_ = _1560_ ? _2681_ : _2683_;
assign _2687_ = _0433_ ? _2679_ : _2685_;
assign _2689_ = _3177_ ? csr_mtval_o[10:8] : _3270_[5:3];
assign _2691_ = _3179_ ? csr_mepc_o[10:8] : csr_mtvec_o[10:8];
assign _2693_ = _1562_ ? _2689_ : _2691_;
assign _2695_ = _3180_ ? mscratch_q[10:8] : 3'h1;
assign _2697_ = _3188_ ? hart_id_i[10:8] : 3'h0;
assign _2699_ = _1568_ ? _2695_ : _2697_;
assign _2701_ = _0427_ ? _2693_ : _2699_;
assign csr_rdata_o[10:8] = _0435_ ? _2687_ : _2701_;
assign _2703_ = _3164_ ? _0022_[52:50] : _0022_[20:18];
assign _2705_ = _3186_ ? _0024_[20:18] : dscratch1_q[20:18];
assign _2707_ = _1570_ ? _2703_ : _2705_;
assign _2709_ = _3173_ ? dscratch0_q[20:18] : csr_depc_o[20:18];
assign _2711_ = _3160_ ? dcsr_q[20:18] : irq_fast_i[4:2];
assign _2713_ = _1572_ ? _2709_ : _2711_;
assign _2715_ = _0437_ ? _2707_ : _2713_;
assign _2717_ = _3177_ ? csr_mtval_o[20:18] : _3270_[15:13];
assign _2719_ = _3179_ ? csr_mepc_o[20:18] : csr_mtvec_o[20:18];
assign _2721_ = _1562_ ? _2717_ : _2719_;
assign _2723_ = _3180_ ? mscratch_q[20:18] : mie_q[4:2];
assign { _2725_[2], _2210_[1:0] } = _3188_ ? hart_id_i[20:18] : 3'h0;
assign _2727_ = _3256_ ? 3'h4 : { _2725_[2], _2210_[1:0] };
assign _2729_ = _1564_ ? _2723_ : _2727_;
assign _2731_ = _0427_ ? _2721_ : _2729_;
assign csr_rdata_o[20:18] = _0439_ ? _2715_ : _2731_;
assign _2733_ = _3164_ ? _0022_[44] : _0022_[12];
assign _2735_ = _3186_ ? _0024_[12] : dscratch1_q[12];
assign _2737_ = _1570_ ? _2733_ : _2735_;
assign _2739_ = _3173_ ? dscratch0_q[12] : csr_depc_o[12];
assign _2741_ = _3160_ ? dcsr_q[12] : csr_mtval_o[12];
assign _2743_ = _1572_ ? _2739_ : _2741_;
assign _2745_ = _0437_ ? _2737_ : _2743_;
assign _2747_ = _3178_ ? _3270_[7] : csr_mepc_o[12];
assign _2749_ = _3175_ ? csr_mtvec_o[12] : mscratch_q[12];
assign _2751_ = _1574_ ? _2747_ : _2749_;
assign _2753_ = _3256_ ? 1'h1 : mstatus_q[3];
assign _2755_ = _3188_ ? hart_id_i[12] : 1'h0;
assign _2757_ = _1576_ ? _2753_ : _2755_;
assign _2759_ = _0441_ ? _2751_ : _2757_;
assign csr_rdata_o[12] = _0443_ ? _2745_ : _2759_;
assign _2761_ = _3164_ ? _0022_[49] : _0022_[17];
assign _2763_ = _3186_ ? _0024_[17] : dscratch1_q[17];
assign _2765_ = _1570_ ? _2761_ : _2763_;
assign _2767_ = _3173_ ? dscratch0_q[17] : csr_depc_o[17];
assign _2769_ = _3160_ ? dcsr_q[17] : irq_fast_i[1];
assign _2771_ = _1572_ ? _2767_ : _2769_;
assign _2773_ = _0437_ ? _2765_ : _2771_;
assign _2775_ = _3177_ ? csr_mtval_o[17] : _3270_[12];
assign _2777_ = _3179_ ? csr_mepc_o[17] : csr_mtvec_o[17];
assign _2779_ = _1562_ ? _2775_ : _2777_;
assign _2781_ = _3180_ ? mscratch_q[17] : mie_q[1];
assign _2783_ = _3188_ ? hart_id_i[17] : 1'h0;
assign _2785_ = _3161_ ? mstatus_q[1] : _2783_;
assign _2787_ = _1564_ ? _2781_ : _2785_;
assign _2789_ = _0427_ ? _2779_ : _2787_;
assign csr_rdata_o[17] = _0439_ ? _2773_ : _2789_;
assign _2791_ = _3168_ ? _0022_[15:13] : _0024_[15:13];
assign _2793_ = _3164_ ? _0022_[47:45] : _2791_;
assign _2795_ = _3172_ ? dscratch1_q[15:13] : dscratch0_q[15:13];
assign _2797_ = _3174_ ? csr_depc_o[15:13] : dcsr_q[15:13];
assign _2799_ = _1560_ ? _2795_ : _2797_;
assign _2801_ = _0433_ ? _2793_ : _2799_;
assign _2803_ = _3178_ ? _3270_[10:8] : csr_mepc_o[15:13];
assign _2805_ = _3177_ ? csr_mtval_o[15:13] : _2803_;
assign _2807_ = _3175_ ? csr_mtvec_o[15:13] : mscratch_q[15:13];
assign _2809_ = _3188_ ? hart_id_i[15:13] : 3'h0;
assign _2811_ = _1578_ ? _2807_ : _2809_;
assign _2813_ = _0445_ ? _2805_ : _2811_;
assign csr_rdata_o[15:13] = _0435_ ? _2801_ : _2813_;
assign _2815_ = _3164_ ? _0022_[48] : _0022_[16];
assign _2817_ = _3186_ ? _0024_[16] : dscratch1_q[16];
assign _2819_ = _1570_ ? _2815_ : _2817_;
assign _2821_ = _3173_ ? dscratch0_q[16] : csr_depc_o[16];
assign _2823_ = _3160_ ? dcsr_q[16] : irq_fast_i[0];
assign _2825_ = _1572_ ? _2821_ : _2823_;
assign _2827_ = _0437_ ? _2819_ : _2825_;
assign _2829_ = _3177_ ? csr_mtval_o[16] : _3270_[11];
assign _2831_ = _3179_ ? csr_mepc_o[16] : csr_mtvec_o[16];
assign _2833_ = _1562_ ? _2829_ : _2831_;
assign _2835_ = _3180_ ? mscratch_q[16] : mie_q[0];
assign _2837_ = _3188_ ? hart_id_i[16] : 1'h0;
assign _2839_ = _1564_ ? _2835_ : _2837_;
assign _2841_ = _0427_ ? _2833_ : _2839_;
assign csr_rdata_o[16] = _0439_ ? _2827_ : _2841_;
assign _2843_ = _3164_ ? _0022_[62:54] : _0022_[30:22];
assign _2845_ = _3186_ ? _0024_[30:22] : dscratch1_q[30:22];
assign _2847_ = _1570_ ? _2843_ : _2845_;
assign _2849_ = _3173_ ? dscratch0_q[30:22] : csr_depc_o[30:22];
assign _2851_ = _3160_ ? dcsr_q[30:22] : irq_fast_i[14:6];
assign _2853_ = _1572_ ? _2849_ : _2851_;
assign _2855_ = _0437_ ? _2847_ : _2853_;
assign _2857_ = _3177_ ? csr_mtval_o[30:22] : _3270_[25:17];
assign _2859_ = _3179_ ? csr_mepc_o[30:22] : csr_mtvec_o[30:22];
assign _2861_ = _1562_ ? _2857_ : _2859_;
assign _2863_ = _3180_ ? mscratch_q[30:22] : mie_q[14:6];
assign { _2865_[8], _2279_[7:0] } = _3188_ ? hart_id_i[30:22] : 9'h000;
assign _2867_ = _3256_ ? 9'h100 : { _2865_[8], _2279_[7:0] };
assign _2869_ = _1564_ ? _2863_ : _2867_;
assign _2871_ = _0427_ ? _2861_ : _2869_;
assign csr_rdata_o[30:22] = _0439_ ? _2855_ : _2871_;
assign _2873_ = _3164_ ? _0022_[43] : _0022_[11];
assign _2875_ = _3186_ ? _0024_[11] : dscratch1_q[11];
assign _2877_ = _1570_ ? _2873_ : _2875_;
assign _2879_ = _3173_ ? dscratch0_q[11] : csr_depc_o[11];
assign _2881_ = _3160_ ? dcsr_q[11] : irq_external_i;
assign _2883_ = _1572_ ? _2879_ : _2881_;
assign _2885_ = _0437_ ? _2877_ : _2883_;
assign _2887_ = _3177_ ? csr_mtval_o[11] : _3270_[6];
assign _2889_ = _3179_ ? csr_mepc_o[11] : csr_mtvec_o[11];
assign _2891_ = _1562_ ? _2887_ : _2889_;
assign _2893_ = _3180_ ? mscratch_q[11] : mie_q[15];
assign _2895_ = _3188_ ? hart_id_i[11] : 1'h0;
assign _2897_ = _3161_ ? mstatus_q[2] : _2895_;
assign _2899_ = _1564_ ? _2893_ : _2897_;
assign _2901_ = _0427_ ? _2891_ : _2899_;
assign csr_rdata_o[11] = _0439_ ? _2885_ : _2901_;
assign _2299_ = _3251_ ? \mhpmcounter[2]  : \mhpmcounter[0] ;
assign _0022_ = _0458_ ? 64'h0000000000000000 : _2299_;
assign _2904_ = _3164_ ? _0022_[53] : _0022_[21];
assign _2906_ = _3186_ ? _0024_[21] : dscratch1_q[21];
assign _2908_ = _1570_ ? _2904_ : _2906_;
assign _2910_ = _3173_ ? dscratch0_q[21] : csr_depc_o[21];
assign _2912_ = _3160_ ? dcsr_q[21] : irq_fast_i[5];
assign _2914_ = _1572_ ? _2910_ : _2912_;
assign _2916_ = _0437_ ? _2908_ : _2914_;
assign _2918_ = _3177_ ? csr_mtval_o[21] : _3270_[16];
assign _2920_ = _3179_ ? csr_mepc_o[21] : csr_mtvec_o[21];
assign _2922_ = _1562_ ? _2918_ : _2920_;
assign _2924_ = _3180_ ? mscratch_q[21] : mie_q[5];
assign _2926_ = _3188_ ? hart_id_i[21] : 1'h0;
assign _2928_ = _3161_ ? mstatus_q[0] : _2926_;
assign _2930_ = _1564_ ? _2924_ : _2928_;
assign _2932_ = _0427_ ? _2922_ : _2930_;
assign csr_rdata_o[21] = _0439_ ? _2916_ : _2932_;
assign _2934_ = _3066_ ? _0145_ : _3105_;
assign dummy_instr_seed_o = _0456_ ? csr_wdata_i : _2934_;
assign _2936_ = _3168_ ? _0022_[31] : _0024_[31];
assign _2938_ = _3164_ ? _0022_[63] : _2936_;
assign _2940_ = _3172_ ? dscratch1_q[31] : dscratch0_q[31];
assign _2942_ = _3174_ ? csr_depc_o[31] : dcsr_q[31];
assign _2944_ = _1560_ ? _2940_ : _2942_;
assign _2946_ = _0433_ ? _2938_ : _2944_;
assign _2948_ = _3178_ ? _3103_ : csr_mepc_o[31];
assign _2950_ = _3177_ ? csr_mtval_o[31] : _2948_;
assign _2952_ = _3175_ ? csr_mtvec_o[31] : mscratch_q[31];
assign _2954_ = _3188_ ? hart_id_i[31] : 1'h0;
assign _2956_ = _1578_ ? _2952_ : _2954_;
assign _2958_ = _0445_ ? _2950_ : _2956_;
assign csr_rdata_o[31] = _0435_ ? _2946_ : _2958_;
assign _2960_ = _3170_ ? cpuctrlsts_part_q[7] : _0022_[39];
assign _2962_ = _3168_ ? _0022_[7] : _0024_[7];
assign _2964_ = _1558_ ? _2960_ : _2962_;
assign _2966_ = _3172_ ? dscratch1_q[7] : dscratch0_q[7];
assign _2968_ = _3160_ ? dcsr_q[7] : irq_timer_i;
assign _2970_ = _3174_ ? csr_depc_o[7] : _2968_;
assign _2972_ = _1560_ ? _2966_ : _2970_;
assign _2974_ = _0425_ ? _2964_ : _2972_;
assign _2976_ = _3177_ ? csr_mtval_o[7] : _3270_[2];
assign _2978_ = _3179_ ? csr_mepc_o[7] : csr_mtvec_o[7];
assign _2980_ = _1562_ ? _2976_ : _2978_;
assign _2982_ = _3180_ ? mscratch_q[7] : mie_q[16];
assign _2984_ = _3188_ ? hart_id_i[7] : 1'h0;
assign _2986_ = _3161_ ? mstatus_q[4] : _2984_;
assign _2988_ = _1564_ ? _2982_ : _2986_;
assign _2990_ = _0427_ ? _2980_ : _2988_;
assign csr_rdata_o[7] = _0429_ ? _2974_ : _2990_;
assign _2992_ = _3170_ ? cpuctrlsts_part_q[6:4] : _0022_[38:36];
assign _2994_ = _3168_ ? _0022_[6:4] : _0024_[6:4];
assign _2996_ = _1558_ ? _2992_ : _2994_;
assign _2998_ = _3172_ ? dscratch1_q[6:4] : dscratch0_q[6:4];
assign _3000_ = _3174_ ? csr_depc_o[6:4] : dcsr_q[6:4];
assign _3002_ = _1560_ ? _2998_ : _3000_;
assign _3004_ = _0425_ ? _2996_ : _3002_;
assign _3006_ = _3177_ ? csr_mtval_o[6:4] : { _3270_[1:0], mcause_q[4] };
assign _3008_ = _3179_ ? csr_mepc_o[6:4] : csr_mtvec_o[6:4];
assign _3010_ = _1562_ ? _3006_ : _3008_;
assign _3012_ = _3180_ ? mscratch_q[6:4] : hart_id_i[6:4];
assign _3014_ = _3192_ ? 3'h1 : 3'h0;
assign _3015_ = _2152_ ? _3012_ : _3014_;
assign _3017_ = _0427_ ? _3010_ : _3015_;
assign csr_rdata_o[6:4] = _0447_ ? _3004_ : _3017_;
assign _0449_ = | _3091_;
assign _3019_ = $signed(_3090_) < 0 ? 1'h0 << - _3090_ : 1'h0 >> _3090_;
assign _3096_ = { _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_, _0449_ } | _3019_;
assign _3020_ = csr_addr_i[11:10] == /* src = "generated/sv2v_out.v:13935.30-13935.54" */ 2'h3;
assign _3062_ = dummy_instr_seed_o[31:30] == /* src = "generated/sv2v_out.v:14104.46-14104.75" */ 2'h2;
assign _3064_ = dummy_instr_seed_o[31:30] == /* src = "generated/sv2v_out.v:14104.15-14104.44" */ 2'h3;
assign illegal_csr_priv = csr_addr_i[9:8] > /* src = "generated/sv2v_out.v:13934.28-13934.56" */ priv_mode_id_o;
assign illegal_csr_write = _3020_ && /* src = "generated/sv2v_out.v:13935.29-13935.65" */ csr_wr;
assign _3074_ = _3080_ && /* src = "generated/sv2v_out.v:14131.10-14131.66" */ _3082_;
assign _3076_ = _3084_ && /* src = "generated/sv2v_out.v:14143.10-14143.60" */ _3086_;
assign dummy_instr_seed_en_o = csr_we_int && /* src = "generated/sv2v_out.v:14801.35-14801.70" */ _3072_;
assign _3078_ = csr_mcause_i[5] || /* src = "generated/sv2v_out.v:14198.12-14198.38" */ csr_mcause_i[6];
assign _3080_ = dummy_instr_seed_o[12:11] != /* src = "generated/sv2v_out.v:14131.11-14131.35" */ 2'h3;
assign _3082_ = | /* src = "generated/sv2v_out.v:14131.41-14131.65" */ dummy_instr_seed_o[12:11];
assign _3084_ = dummy_instr_seed_o[1:0] != /* src = "generated/sv2v_out.v:14143.11-14143.32" */ 2'h3;
assign _3086_ = | /* src = "generated/sv2v_out.v:14143.38-14143.59" */ dummy_instr_seed_o[1:0];
assign _3088_ = mstatus_q[3:2] != /* src = "generated/sv2v_out.v:14213.9-14213.33" */ 2'h3;
assign _3090_ = - /* src = "generated/sv2v_out.v:0.0-0.0" */ $signed({ 27'h0000000, csr_addr_i[4:0] });
assign _3092_ = ~ /* src = "generated/sv2v_out.v:14250.47-14250.66" */ illegal_csr_insn_o;
assign _0149_ = ~ /* src = "generated/sv2v_out.v:14622.40-14622.57" */ mcountinhibit[0];
assign _3093_ = ~ /* src = "generated/sv2v_out.v:14641.46-14641.63" */ mcountinhibit[2];
assign _3094_ = ~ /* src = "generated/sv2v_out.v:14845.50-14845.89" */ _3107_;
assign _3097_ = illegal_csr | /* src = "generated/sv2v_out.v:13936.48-13936.79" */ illegal_csr_write;
assign _3099_ = _3097_ | /* src = "generated/sv2v_out.v:13936.47-13936.99" */ illegal_csr_priv;
assign _3101_ = _3099_ | /* src = "generated/sv2v_out.v:13936.46-13936.118" */ illegal_csr_dbg;
assign _3103_ = mcause_q[5] | /* src = "generated/sv2v_out.v:13991.30-13991.55" */ mcause_q[6];
assign _3105_ = csr_wdata_i | /* src = "generated/sv2v_out.v:14244.26-14244.51" */ csr_rdata_o;
assign _3107_ = debug_mode_i | /* src = "generated/sv2v_out.v:14845.52-14845.88" */ debug_mode_entering_i;
assign _3108_ = mstatus_err | /* src = "generated/sv2v_out.v:14858.31-14858.54" */ mtvec_err;
assign csr_shadow_err_o = _3108_ | /* src = "generated/sv2v_out.v:14858.29-14858.92" */ cpuctrlsts_part_err;
assign _3110_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14242.3-14248.10" */ csr_op_i;
assign _3066_ = csr_op_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14242.3-14248.10" */ 2'h3;
assign _3068_ = csr_op_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14242.3-14248.10" */ 2'h2;
assign _3070_ = csr_op_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14242.3-14248.10" */ 2'h1;
assign cpuctrlsts_part_d[7] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0088_[1] : _0000_[7];
assign _0131_ = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14217.9-14217.19|generated/sv2v_out.v:14217.5-14228.8" */ 1'h1 : _0012_;
assign _0102_ = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14217.9-14217.19|generated/sv2v_out.v:14217.5-14228.8" */ mstack_epc_q : { dummy_instr_seed_o[31:1], 1'h0 };
assign _0133_ = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14217.9-14217.19|generated/sv2v_out.v:14217.5-14228.8" */ 1'h1 : _0014_;
assign _0143_[1:0] = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14217.9-14217.19|generated/sv2v_out.v:14217.5-14228.8" */ mstack_q[1:0] : 2'h0;
assign _0143_[2] = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14217.9-14217.19|generated/sv2v_out.v:14217.5-14228.8" */ mstack_q[2] : 1'h1;
assign _0141_ = _3088_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14213.9-14213.33|generated/sv2v_out.v:14213.5-14214.26" */ 1'h0 : _0016_[1];
assign _3112_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0143_ : _0016_[4:2];
assign _3114_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0016_[4:2] : _3112_;
assign mstatus_d[4:2] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0119_[2:0] : _3114_;
assign _3116_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0141_ : _0016_[1];
assign _3118_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0016_[1] : _3116_;
assign mstatus_d[1] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0016_[1] : _3118_;
assign _3120_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ mstatus_q[4] : _0016_[5];
assign _3122_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0016_[5] : _3120_;
assign mstatus_d[5] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0119_[3] : _3122_;
assign _0114_ = cpuctrlsts_part_q[6] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14201.11-14201.31|generated/sv2v_out.v:14201.7-14204.10" */ 1'h1 : 1'h0;
assign _0125_[0] = _3078_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14198.10-14198.39|generated/sv2v_out.v:14198.6-14205.9" */ _0000_[6] : 1'h1;
assign _0096_ = _3078_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14198.10-14198.39|generated/sv2v_out.v:14198.6-14205.9" */ 1'h0 : _0114_;
assign _0137_ = cpuctrlsts_part_q[6] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14201.11-14201.31|generated/sv2v_out.v:14201.7-14204.10" */ 1'h1 : _0000_[7];
assign _0127_ = _3078_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14198.10-14198.39|generated/sv2v_out.v:14198.6-14205.9" */ _0002_ : 1'h1;
assign _0112_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14186.14-14186.27|generated/sv2v_out.v:14186.10-14206.8" */ _0002_ : _0127_;
assign _0110_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14186.14-14186.27|generated/sv2v_out.v:14186.10-14206.8" */ _0000_[7:6] : _0125_;
assign _0077_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14186.14-14186.27|generated/sv2v_out.v:14186.10-14206.8" */ 1'h0 : _0096_;
assign _0083_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14186.14-14186.27|generated/sv2v_out.v:14186.10-14206.8" */ 1'h0 : 1'h1;
assign _0079_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14186.14-14186.27|generated/sv2v_out.v:14186.10-14206.8" */ { _3064_, _3062_, dummy_instr_seed_o[4:0] } : csr_mcause_i;
assign _0115_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14186.14-14186.27|generated/sv2v_out.v:14186.10-14206.8" */ _0012_ : 1'h1;
assign _0081_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14186.14-14186.27|generated/sv2v_out.v:14186.10-14206.8" */ { dummy_instr_seed_o[31:1], 1'h0 } : _0043_;
assign _0117_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14186.14-14186.27|generated/sv2v_out.v:14186.10-14206.8" */ _0014_ : 1'h1;
assign _0125_[1] = _3078_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14198.10-14198.39|generated/sv2v_out.v:14198.6-14205.9" */ _0000_[7] : _0137_;
assign _0135_[1:0] = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14186.14-14186.27|generated/sv2v_out.v:14186.10-14206.8" */ _0016_[3:2] : priv_mode_id_o;
assign _0135_[2] = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14186.14-14186.27|generated/sv2v_out.v:14186.10-14206.8" */ _0016_[4] : mstatus_q[5];
assign _0121_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14186.14-14186.27|generated/sv2v_out.v:14186.10-14206.8" */ _0018_ : 1'h1;
assign _0086_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14186.14-14186.27|generated/sv2v_out.v:14186.10-14206.8" */ dummy_instr_seed_o : csr_mtval_i;
assign _0123_ = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14186.14-14186.27|generated/sv2v_out.v:14186.10-14206.8" */ _0020_ : 1'h1;
assign _0094_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ 1'h1 : _0008_;
assign _0033_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ _0043_ : { dummy_instr_seed_o[31:1], 1'h0 };
assign _0092_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ 1'h1 : _0006_;
assign _0139_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ debug_cause_i : _0004_[8:6];
assign _0129_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ priv_mode_id_o : _0004_[1:0];
assign _0090_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ _0002_ : _0112_;
assign _0088_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ _0000_[7:6] : _0110_;
assign _0063_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ 1'h0 : _0083_;
assign _0108_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ _0020_ : _0123_;
assign _0069_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ dummy_instr_seed_o : _0086_;
assign _0100_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ _0012_ : _0115_;
assign _0045_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ { _3064_, _3062_, dummy_instr_seed_o[4:0] } : _0079_;
assign _0104_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ _0014_ : _0117_;
assign _0051_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ { dummy_instr_seed_o[31:1], 1'h0 } : _0081_;
assign _0106_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ _0018_ : _0121_;
assign _0119_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ _0016_[5:2] : _0135_;
assign _0037_ = debug_csr_save_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14179.9-14179.25|generated/sv2v_out.v:14179.5-14206.8" */ 1'h0 : _0077_;
assign _3124_ = csr_save_wb_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14171.5-14177.12" */ pc_wb_i : pc_id_i;
assign _3126_ = csr_save_id_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14171.5-14177.12" */ pc_id_i : _3124_;
assign _0043_ = csr_save_if_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14171.5-14177.12" */ pc_if_i : _3126_;
assign _3128_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ 1'h1 : _0002_;
assign _3130_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0002_ : _3128_;
assign cpuctrlsts_part_we = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0090_ : _3130_;
assign _3132_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ 1'h0 : _0000_[6];
assign _3134_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0000_[6] : _3132_;
assign cpuctrlsts_part_d[6] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0088_[0] : _3134_;
assign mstack_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0063_ : 1'h0;
assign depc_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0094_ : _0008_;
assign depc_d = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0033_ : { dummy_instr_seed_o[31:1], 1'h0 };
assign dcsr_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0092_ : _0006_;
assign dcsr_d[8:6] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0139_ : _0004_[8:6];
assign dcsr_d[1:0] = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0129_ : _0004_[1:0];
assign mtval_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0108_ : _0020_;
assign mtval_d = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0069_ : dummy_instr_seed_o;
assign _3136_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0131_ : _0012_;
assign _3138_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0012_ : _3136_;
assign mcause_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0100_ : _3138_;
assign _3140_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0098_ : { _3064_, _3062_, dummy_instr_seed_o[4:0] };
assign _3142_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ { _3064_, _3062_, dummy_instr_seed_o[4:0] } : _3140_;
assign mcause_d = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0045_ : _3142_;
assign _3144_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0133_ : _0014_;
assign _3146_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0014_ : _3144_;
assign mepc_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0104_ : _3146_;
assign _3148_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0102_ : { dummy_instr_seed_o[31:1], 1'h0 };
assign _3150_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ { dummy_instr_seed_o[31:1], 1'h0 } : _3148_;
assign mepc_d = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0051_ : _3150_;
assign _3152_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ 1'h1 : _0018_;
assign _3154_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0018_ : _3152_;
assign mstatus_en = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0106_ : _3154_;
assign _0098_ = nmi_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14217.9-14217.19|generated/sv2v_out.v:14217.5-14228.8" */ mstack_cause_q : { _3064_, _3062_, dummy_instr_seed_o[4:0] };
assign double_fault_seen_o = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ _0037_ : 1'h0;
assign _3156_ = csr_restore_mret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ mstatus_q[3:2] : 2'hx;
assign _3158_ = csr_restore_dret_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ dcsr_q[1:0] : _3156_;
assign priv_lvl_d = csr_save_cause_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14169.3-14232.10" */ 2'h3 : _3158_;
assign _0135_[3] = debug_mode_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14186.14-14186.27|generated/sv2v_out.v:14186.10-14206.8" */ _0016_[5] : 1'h0;
assign _0029_[31:28] = _3160_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 4'h4 : dcsr_q[31:28];
assign _0065_[5:4] = _3161_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ { dummy_instr_seed_o[3], dummy_instr_seed_o[7] } : mstatus_q[5:4];
assign _0065_[3:2] = _3161_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ _0084_ : mstatus_q[3:2];
assign _0029_[15] = _3160_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ dummy_instr_seed_o[15] : dcsr_q[15];
assign _0029_[14] = _3160_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h0 : dcsr_q[14];
assign _0029_[27:16] = _3160_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 12'h000 : dcsr_q[27:16];
assign _0065_[1:0] = _3161_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ { dummy_instr_seed_o[17], dummy_instr_seed_o[21] } : mstatus_q[1:0];
assign _0029_[1:0] = _3160_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ _0075_ : dcsr_q[1:0];
assign _0029_[5] = _3160_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h0 : dcsr_q[5];
assign _0029_[4] = _3160_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h0 : dcsr_q[4];
assign _0029_[3] = _3160_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h0 : dcsr_q[3];
assign _0029_[2] = _3160_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ dummy_instr_seed_o[2] : dcsr_q[2];
assign _0029_[13:12] = _3160_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ dummy_instr_seed_o[13:12] : dcsr_q[13:12];
assign _0029_[11] = _3160_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h0 : dcsr_q[11];
assign _0075_ = _3076_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14143.10-14143.60|generated/sv2v_out.v:14143.6-14144.28" */ 2'h0 : dummy_instr_seed_o[1:0];
assign _0029_[9] = _3160_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h0 : dcsr_q[9];
assign _0084_ = _3074_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14131.10-14131.66|generated/sv2v_out.v:14131.6-14132.31" */ 2'h0 : dummy_instr_seed_o[12:11];
assign _0067_ = _3161_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h1 : 1'h0;
assign _3168_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ _3166_;
assign _0027_ = _3170_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h1 : 1'h0;
assign _0025_ = _3170_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ { dummy_instr_seed_o[7:1], 1'h0 } : cpuctrlsts_part_q;
assign _0057_ = _3164_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ _2429_ : 32'd0;
assign _0055_ = _3168_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ _2429_ : 32'd0;
assign _0049_ = _3171_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h1 : 1'h0;
assign _0041_ = _3172_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h1 : 1'h0;
assign _0039_ = _3173_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h1 : 1'h0;
assign _0035_ = _3174_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h1 : 1'h0;
assign _0031_ = _3160_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h1 : 1'h0;
assign _0029_[10] = _3160_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h0 : dcsr_q[10];
assign _0073_ = _3175_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h1 : csr_mtvec_init_i;
assign _0071_ = _3177_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h1 : 1'h0;
assign _0047_ = _3178_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h1 : 1'h0;
assign _0053_ = _3179_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h1 : 1'h0;
assign _0061_ = _3180_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h1 : 1'h0;
assign _0059_ = _3181_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:14127.4-14168.11" */ 1'h1 : 1'h0;
assign _0002_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0027_ : 1'h0;
assign { _0000_[7:6], cpuctrlsts_part_d[5:0] } = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0025_ : cpuctrlsts_part_q;
assign mhpmcounterh_we = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0057_ : 32'd0;
assign mhpmcounter_we = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0055_ : 32'd0;
assign mcountinhibit_we = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0049_ : 1'h0;
assign dscratch1_en = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0041_ : 1'h0;
assign dscratch0_en = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0039_ : 1'h0;
assign _0008_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0035_ : 1'h0;
assign _0006_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0031_ : 1'h0;
assign { dcsr_d[31:9], _0004_[8:6], dcsr_d[5:2], _0004_[1:0] } = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ { _0029_[31:9], dcsr_q[8:6], _0029_[5:0] } : dcsr_q;
assign mtvec_en = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0073_ : csr_mtvec_init_i;
assign _0020_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0071_ : 1'h0;
assign _0012_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0047_ : 1'h0;
assign _0014_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0053_ : 1'h0;
assign mscratch_en = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0061_ : 1'h0;
assign mie_en = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0059_ : 1'h0;
assign _0018_ = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0067_ : 1'h0;
assign { _0016_[5:1], mstatus_d[0] } = csr_we_int ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14126.7-14126.17|generated/sv2v_out.v:14126.3-14168.11" */ _0065_ : mstatus_q;
assign illegal_csr = _3182_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:14087.8-14087.429|generated/sv2v_out.v:14087.4-14088.24" */ 1'h1 : _0010_;
assign _0024_ = _0454_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 32'd0 : 32'hxxxxxxxx;
assign _3164_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ _3162_;
assign _3171_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h320;
assign _3192_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hf12;
assign _3186_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ _3184_;
assign _3256_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h301;
assign _3193_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1f;
assign _3195_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1e;
assign _3197_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1d;
assign _3199_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1c;
assign _3201_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1b;
assign _3203_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h1a;
assign _3205_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h19;
assign _3207_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h18;
assign _3209_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h17;
assign _3211_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h16;
assign _3213_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h15;
assign _3215_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h14;
assign _3217_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h13;
assign _3219_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h12;
assign _3221_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h11;
assign _3223_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h10;
assign _3225_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0f;
assign _3227_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0e;
assign _3229_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0d;
assign _3231_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0c;
assign _3233_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0b;
assign _3235_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h0a;
assign _3237_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h09;
assign _3239_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h08;
assign _3241_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h07;
assign _3243_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h06;
assign _3245_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h05;
assign _3247_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h04;
assign _3249_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h03;
assign _3251_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h02;
assign _3253_ = csr_addr_i[4:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ 5'h01;
assign _3255_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0" */ csr_addr_i[4:0];
assign _3172_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h7b3;
assign _3173_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h7b2;
assign _3174_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h7b1;
assign _3160_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h7b0;
assign _3022_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3bf;
assign _3024_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3be;
assign _3026_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3bd;
assign _3028_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3bc;
assign _3030_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3bb;
assign _3032_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3ba;
assign _3034_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3b9;
assign _3036_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3b8;
assign _3038_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3b7;
assign _3040_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3b6;
assign _3042_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3b5;
assign _3044_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3b4;
assign _3046_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3b3;
assign _3048_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3b2;
assign _3050_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3b1;
assign _3052_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3b0;
assign _3054_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3a3;
assign _3056_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3a2;
assign _3058_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3a1;
assign _3060_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h3a0;
assign _3190_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h344;
assign _3177_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h343;
assign _3178_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h342;
assign _3179_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h341;
assign _3175_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h305;
assign _3180_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h340;
assign _3181_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h304;
assign _3161_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h300;
assign _3188_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hf14;
assign _3166_[1] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb02;
assign _3166_[10] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb0b;
assign _3166_[11] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb0c;
assign _3166_[12] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb0d;
assign _3166_[13] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb0e;
assign _3166_[14] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb0f;
assign _3166_[15] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb10;
assign _3166_[16] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb11;
assign _3166_[17] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb12;
assign _3166_[18] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb13;
assign _3166_[19] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb14;
assign _3166_[2] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb03;
assign _3166_[20] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb15;
assign _3166_[21] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb16;
assign _3166_[22] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb17;
assign _3166_[23] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb18;
assign _3166_[24] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb19;
assign _3166_[25] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb1a;
assign _3166_[26] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb1b;
assign _3166_[27] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb1c;
assign _3166_[28] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb1d;
assign _3166_[29] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb1e;
assign _3166_[3] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb04;
assign _3166_[30] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb1f;
assign _3166_[4] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb05;
assign _3166_[5] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb06;
assign _3166_[6] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb07;
assign _3166_[7] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb08;
assign _3166_[8] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb09;
assign _3166_[9] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb0a;
assign _3184_[0] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h323;
assign _3184_[1] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h324;
assign _3184_[10] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h32d;
assign _3184_[11] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h32e;
assign _3184_[12] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h32f;
assign _3184_[13] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h330;
assign _3184_[14] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h331;
assign _3184_[15] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h332;
assign _3184_[16] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h333;
assign _3184_[17] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h334;
assign _3184_[18] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h335;
assign _3184_[19] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h336;
assign _3184_[2] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h325;
assign _3184_[20] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h337;
assign _3184_[21] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h338;
assign _3184_[22] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h339;
assign _3184_[23] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h33a;
assign _3184_[24] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h33b;
assign _3184_[25] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h33c;
assign _3184_[26] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h33d;
assign _3184_[27] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h33e;
assign _3184_[28] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h33f;
assign _3184_[3] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h326;
assign _3184_[4] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h327;
assign _3184_[5] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h328;
assign _3184_[6] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h329;
assign _3184_[7] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h32a;
assign _3184_[8] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h32b;
assign _3184_[9] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h32c;
assign _0010_ = _0391_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 1'h0 : 1'h1;
assign _3072_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h7c1;
assign _3170_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h7c0;
assign _3162_[0] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb80;
assign _3162_[1] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb82;
assign _3162_[10] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb8b;
assign _3162_[11] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb8c;
assign _3162_[12] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb8d;
assign _3162_[13] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb8e;
assign _3162_[14] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb8f;
assign _3162_[15] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb90;
assign _3162_[16] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb91;
assign _3162_[17] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb92;
assign _3162_[18] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb93;
assign _3162_[19] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb94;
assign _3162_[2] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb83;
assign _3162_[20] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb95;
assign _3162_[21] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb96;
assign _3162_[22] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb97;
assign _3162_[23] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb98;
assign _3162_[24] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb99;
assign _3162_[25] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb9a;
assign _3162_[26] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb9b;
assign _3162_[27] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb9c;
assign _3162_[28] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb9d;
assign _3162_[29] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb9e;
assign _3162_[3] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb84;
assign _3162_[30] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb9f;
assign _3162_[4] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb85;
assign _3162_[5] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb86;
assign _3162_[6] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb87;
assign _3162_[7] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb88;
assign _3162_[8] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb89;
assign _3162_[9] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb8a;
assign _3166_[0] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hb00;
assign _3258_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h306;
assign _3260_[0] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h30a;
assign _3260_[1] = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h31a;
assign _3262_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'h310;
assign _3264_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hf15;
assign _3266_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hf13;
assign _3268_ = csr_addr_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 12'hf11;
assign dbg_csr = _0455_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:13963.3-14085.10" */ 1'h1 : 1'h0;
assign _3182_ = | /* src = "generated/sv2v_out.v:14087.8-14087.429" */ { _3060_, _3058_, _3056_, _3054_, _3052_, _3050_, _3048_, _3046_, _3044_, _3042_, _3040_, _3038_, _3036_, _3034_, _3032_, _3030_, _3028_, _3026_, _3024_, _3022_ };
assign csr_wr = | /* src = "generated/sv2v_out.v:14249.18-14249.73" */ { _3070_, _3068_, _3066_ };
assign irq_pending_o = | /* src = "generated/sv2v_out.v:14262.25-14262.32" */ irqs_o;
assign _2429_ = $signed(_3090_) < 0 ? 1'h1 << - _3090_ : 1'h1 >> _3090_;
assign _3270_ = mcause_q[6] ? /* src = "generated/sv2v_out.v:13991.58-13991.116" */ 26'h3ffffff : 26'h0000000;
assign mtvec_d = csr_mtvec_init_i ? /* src = "generated/sv2v_out.v:14108.14-14108.112" */ { boot_addr_i[31:8], 8'h01 } : { dummy_instr_seed_o[31:8], 8'h01 };
assign priv_mode_lsu_o = mstatus_q[1] ? /* src = "generated/sv2v_out.v:14240.28-14240.71" */ mstatus_q[3:2] : priv_mode_id_o;
assign \mhpmcounter[2]  = _0152_ ? /* src = "generated/sv2v_out.v:14641.27-14641.94" */ minstret_next : minstret_raw;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14619.36-14627.3" */
\$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000  mcycle_counter_i (
.clk_i(clk_i),
.counter_inc_i(_0149_),
.counter_inc_i_t0(mcountinhibit_t0[0]),
.counter_val_i(dummy_instr_seed_o),
.counter_val_i_t0(dummy_instr_seed_o_t0),
.counter_val_o(\mhpmcounter[0] ),
.counter_val_o_t0(\mhpmcounter[0]_t0 ),
.counter_we_i(mhpmcounter_we[0]),
.counter_we_i_t0(mhpmcounter_we_t0[0]),
.counterh_we_i(mhpmcounterh_we[0]),
.counterh_we_i_t0(mhpmcounterh_we_t0[0]),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14631.4-14640.3" */
\$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter  minstret_counter_i (
.clk_i(clk_i),
.counter_inc_i(_0150_),
.counter_inc_i_t0(_0151_),
.counter_val_i(dummy_instr_seed_o),
.counter_val_i_t0(dummy_instr_seed_o_t0),
.counter_val_o(minstret_raw),
.counter_val_o_t0(minstret_raw_t0),
.counter_val_upd_o(minstret_next),
.counter_val_upd_o_t0(minstret_next_t0),
.counter_we_i(mhpmcounter_we[2]),
.counter_we_i_t0(mhpmcounter_we_t0[2]),
.counterh_we_i(mhpmcounterh_we[2]),
.counterh_we_i_t0(mhpmcounterh_we_t0[2]),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14850.4-14857.3" */
\$paramod$a088b13b9337f1e1fba58a671f47d7c7701ffa49\ibex_csr  u_cpuctrlsts_part_csr (
.clk_i(clk_i),
.rd_data_o(cpuctrlsts_part_q),
.rd_data_o_t0(cpuctrlsts_part_q_t0),
.rd_error_o(cpuctrlsts_part_err),
.rd_error_o_t0(cpuctrlsts_part_err_t0),
.rst_ni(rst_ni),
.wr_data_i(cpuctrlsts_part_d),
.wr_data_i_t0(cpuctrlsts_part_d_t0),
.wr_en_i(cpuctrlsts_part_we),
.wr_en_i_t0(cpuctrlsts_part_we_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14352.4-14358.3" */
\$paramod$9a435d8f6db004a67362aa9a56f32ea481a74dbe\ibex_csr  u_dcsr_csr (
.clk_i(clk_i),
.rd_data_o(dcsr_q),
.rd_data_o_t0(dcsr_q_t0),
.rst_ni(rst_ni),
.wr_data_i(dcsr_d),
.wr_data_i_t0(dcsr_d_t0),
.wr_en_i(dcsr_en),
.wr_en_i_t0(dcsr_en_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14363.4-14369.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_depc_csr (
.clk_i(clk_i),
.rd_data_o(csr_depc_o),
.rd_data_o_t0(csr_depc_o_t0),
.rst_ni(rst_ni),
.wr_data_i(depc_d),
.wr_data_i_t0(depc_d_t0),
.wr_en_i(depc_en),
.wr_en_i_t0(depc_en_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14374.4-14380.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_dscratch0_csr (
.clk_i(clk_i),
.rd_data_o(dscratch0_q),
.rd_data_o_t0(dscratch0_q_t0),
.rst_ni(rst_ni),
.wr_data_i(dummy_instr_seed_o),
.wr_data_i_t0(dummy_instr_seed_o_t0),
.wr_en_i(dscratch0_en),
.wr_en_i_t0(dscratch0_en_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14385.4-14391.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_dscratch1_csr (
.clk_i(clk_i),
.rd_data_o(dscratch1_q),
.rd_data_o_t0(dscratch1_q_t0),
.rst_ni(rst_ni),
.wr_data_i(dummy_instr_seed_o),
.wr_data_i_t0(dummy_instr_seed_o_t0),
.wr_en_i(dscratch1_en),
.wr_en_i_t0(dscratch1_en_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14317.4-14323.3" */
\$paramod$34601000fe8707ce2501f5ed778e152043201712\ibex_csr  u_mcause_csr (
.clk_i(clk_i),
.rd_data_o(mcause_q),
.rd_data_o_t0(mcause_q_t0),
.rst_ni(rst_ni),
.wr_data_i(mcause_d),
.wr_data_i_t0(mcause_d_t0),
.wr_en_i(mcause_en),
.wr_en_i_t0(mcause_en_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14280.4-14286.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_mepc_csr (
.clk_i(clk_i),
.rd_data_o(csr_mepc_o),
.rd_data_o_t0(csr_mepc_o_t0),
.rst_ni(rst_ni),
.wr_data_i(mepc_d),
.wr_data_i_t0(mepc_d_t0),
.wr_en_i(mepc_en),
.wr_en_i_t0(mepc_en_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14295.4-14301.3" */
\$paramod$e55993a14b1fbc43320d549f521b710ed37596c6\ibex_csr  u_mie_csr (
.clk_i(clk_i),
.rd_data_o(mie_q),
.rd_data_o_t0(mie_q_t0),
.rst_ni(rst_ni),
.wr_data_i({ dummy_instr_seed_o[3], dummy_instr_seed_o[7], dummy_instr_seed_o[11], dummy_instr_seed_o[30:16] }),
.wr_data_i_t0({ dummy_instr_seed_o_t0[3], dummy_instr_seed_o_t0[7], dummy_instr_seed_o_t0[11], dummy_instr_seed_o_t0[30:16] }),
.wr_en_i(mie_en),
.wr_en_i_t0(mie_en_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14306.4-14312.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_mscratch_csr (
.clk_i(clk_i),
.rd_data_o(mscratch_q),
.rd_data_o_t0(mscratch_q_t0),
.rst_ni(rst_ni),
.wr_data_i(dummy_instr_seed_o),
.wr_data_i_t0(dummy_instr_seed_o_t0),
.wr_en_i(mscratch_en),
.wr_en_i_t0(mscratch_en_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14419.4-14425.3" */
\$paramod$34601000fe8707ce2501f5ed778e152043201712\ibex_csr  u_mstack_cause_csr (
.clk_i(clk_i),
.rd_data_o(mstack_cause_q),
.rd_data_o_t0(mstack_cause_q_t0),
.rst_ni(rst_ni),
.wr_data_i(mcause_q),
.wr_data_i_t0(mcause_q_t0),
.wr_en_i(mstack_en),
.wr_en_i_t0(mstack_en_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14397.4-14403.3" */
\$paramod$410b37fbfbfa994790f1902c150d2be939cadb3b\ibex_csr  u_mstack_csr (
.clk_i(clk_i),
.rd_data_o(mstack_q),
.rd_data_o_t0(mstack_q_t0),
.rst_ni(rst_ni),
.wr_data_i(mstatus_q[4:2]),
.wr_data_i_t0(mstatus_q_t0[4:2]),
.wr_en_i(mstack_en),
.wr_en_i_t0(mstack_en_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14408.4-14414.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_mstack_epc_csr (
.clk_i(clk_i),
.rd_data_o(mstack_epc_q),
.rd_data_o_t0(mstack_epc_q_t0),
.rst_ni(rst_ni),
.wr_data_i(csr_mepc_o),
.wr_data_i_t0(csr_mepc_o_t0),
.wr_en_i(mstack_en),
.wr_en_i_t0(mstack_en_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14268.4-14275.3" */
\$paramod$5714e31d82f2b8816750797f158ebea69a089104\ibex_csr  u_mstatus_csr (
.clk_i(clk_i),
.rd_data_o(mstatus_q),
.rd_data_o_t0(mstatus_q_t0),
.rd_error_o(mstatus_err),
.rd_error_o_t0(mstatus_err_t0),
.rst_ni(rst_ni),
.wr_data_i(mstatus_d),
.wr_data_i_t0(mstatus_d_t0),
.wr_en_i(mstatus_en),
.wr_en_i_t0(mstatus_en_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14328.4-14334.3" */
\$paramod$85ba01ab5a28334786aba5877c1fe04472f39fba\ibex_csr  u_mtval_csr (
.clk_i(clk_i),
.rd_data_o(csr_mtval_o),
.rd_data_o_t0(csr_mtval_o_t0),
.rst_ni(rst_ni),
.wr_data_i(mtval_d),
.wr_data_i_t0(mtval_d_t0),
.wr_en_i(mtval_en),
.wr_en_i_t0(mtval_en_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:14339.4-14346.3" */
\$paramod$4f46e25470a27719ee9ca03cee1a0827eff766f7\ibex_csr  u_mtvec_csr (
.clk_i(clk_i),
.rd_data_o(csr_mtvec_o),
.rd_data_o_t0(csr_mtvec_o_t0),
.rd_error_o(mtvec_err),
.rd_error_o_t0(mtvec_err_t0),
.rst_ni(rst_ni),
.wr_data_i(mtvec_d),
.wr_data_i_t0(mtvec_d_t0),
.wr_en_i(mtvec_en),
.wr_en_i_t0(mtvec_en_t0)
);
assign _0000_[5:0] = cpuctrlsts_part_d[5:0];
assign _0001_[5:0] = cpuctrlsts_part_d_t0[5:0];
assign { _0004_[31:9], _0004_[5:2] } = { dcsr_d[31:9], dcsr_d[5:2] };
assign { _0005_[31:9], _0005_[5:2] } = { dcsr_d_t0[31:9], dcsr_d_t0[5:2] };
assign _0016_[0] = mstatus_d[0];
assign _0017_[0] = mstatus_d_t0[0];
assign _0029_[8:6] = dcsr_q[8:6];
assign _0030_[8:6] = dcsr_q_t0[8:6];
assign _2210_[2] = _0406_;
assign _2279_[8] = _0407_;
assign _2670_[1:0] = { _2670_[2], 1'h0 };
assign _2725_[1:0] = _2210_[1:0];
assign _2865_[7:0] = _2279_[7:0];
assign csr_mstatus_mie_o = mstatus_q[5];
assign csr_mstatus_mie_o_t0 = mstatus_q_t0[5];
assign csr_mstatus_tw_o = mstatus_q[0];
assign csr_mstatus_tw_o_t0 = mstatus_q_t0[0];
assign csr_pmp_addr_o = 136'h0000000000000000000000000000000000;
assign csr_pmp_addr_o_t0 = 136'h0000000000000000000000000000000000;
assign csr_pmp_cfg_o = 24'h000000;
assign csr_pmp_cfg_o_t0 = 24'h000000;
assign csr_pmp_mseccfg_o = 3'h0;
assign csr_pmp_mseccfg_o_t0 = 3'h0;
assign data_ind_timing_o = cpuctrlsts_part_q[1];
assign data_ind_timing_o_t0 = cpuctrlsts_part_q_t0[1];
assign debug_ebreakm_o = dcsr_q[15];
assign debug_ebreakm_o_t0 = dcsr_q_t0[15];
assign debug_ebreaku_o = dcsr_q[12];
assign debug_ebreaku_o_t0 = dcsr_q_t0[12];
assign debug_single_step_o = dcsr_q[2];
assign debug_single_step_o_t0 = dcsr_q_t0[2];
assign dummy_instr_en_o = cpuctrlsts_part_q[2];
assign dummy_instr_en_o_t0 = cpuctrlsts_part_q_t0[2];
assign dummy_instr_mask_o = cpuctrlsts_part_q[5:3];
assign dummy_instr_mask_o_t0 = cpuctrlsts_part_q_t0[5:3];
assign { mcountinhibit[31:3], mcountinhibit[1] } = 30'h00000000;
assign { mcountinhibit_t0[31:3], mcountinhibit_t0[1] } = 30'h00000000;
assign trigger_match_o = 1'h0;
assign trigger_match_o_t0 = 1'h0;
endmodule

module \$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter (clk_i, rst_ni, counter_inc_i, counterh_we_i, counter_we_i, counter_val_i, counter_val_o, counter_val_upd_o, counter_inc_i_t0, counter_val_i_t0, counter_val_o_t0, counter_val_upd_o_t0, counter_we_i_t0, counterh_we_i_t0);
/* src = "generated/sv2v_out.v:13613.2-13627.5" */
wire [63:0] _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13613.2-13627.5" */
wire [63:0] _001_;
wire [63:0] _002_;
wire _003_;
wire _004_;
wire _005_;
wire [1:0] _006_;
wire _007_;
wire [1:0] _008_;
wire _009_;
wire [63:0] _010_;
wire [31:0] _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
/* cellift = 32'd1 */
wire _019_;
wire _020_;
/* cellift = 32'd1 */
wire _021_;
wire _022_;
/* cellift = 32'd1 */
wire _023_;
wire _024_;
/* cellift = 32'd1 */
wire _025_;
wire _026_;
/* cellift = 32'd1 */
wire _027_;
wire [63:0] _028_;
wire [31:0] _029_;
wire [31:0] _030_;
wire [31:0] _031_;
wire [31:0] _032_;
wire [31:0] _033_;
wire [31:0] _034_;
wire [1:0] _035_;
wire [1:0] _036_;
wire _037_;
wire _038_;
wire _039_;
wire [63:0] _040_;
wire [63:0] _041_;
wire [63:0] _042_;
wire [63:0] _043_;
wire [31:0] _044_;
wire [31:0] _045_;
wire [31:0] _046_;
wire [31:0] _047_;
wire [31:0] _048_;
wire [31:0] _049_;
wire [31:0] _050_;
wire [31:0] _051_;
wire [1:0] _052_;
wire [1:0] _053_;
wire _054_;
wire [63:0] _055_;
wire [63:0] _056_;
wire [63:0] _057_;
wire [63:0] _058_;
wire [31:0] _059_;
wire [31:0] _060_;
wire [63:0] _061_;
wire [31:0] _062_;
wire [31:0] _063_;
wire [63:0] _064_;
wire _065_;
wire _066_;
wire [63:0] _067_;
wire [63:0] _068_;
/* src = "generated/sv2v_out.v:13599.13-13599.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:13611.27-13611.36" */
wire [63:0] counter_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13611.27-13611.36" */
wire [63:0] counter_d_t0;
/* src = "generated/sv2v_out.v:13601.13-13601.26" */
input counter_inc_i;
wire counter_inc_i;
/* cellift = 32'd1 */
input counter_inc_i_t0;
wire counter_inc_i_t0;
/* src = "generated/sv2v_out.v:13609.13-13609.25" */
wire [63:0] counter_load;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13609.13-13609.25" */
wire [63:0] counter_load_t0;
/* src = "generated/sv2v_out.v:13604.20-13604.33" */
input [31:0] counter_val_i;
wire [31:0] counter_val_i;
/* cellift = 32'd1 */
input [31:0] counter_val_i_t0;
wire [31:0] counter_val_i_t0;
/* src = "generated/sv2v_out.v:13605.21-13605.34" */
output [63:0] counter_val_o;
reg [63:0] counter_val_o;
/* cellift = 32'd1 */
output [63:0] counter_val_o_t0;
reg [63:0] counter_val_o_t0;
/* src = "generated/sv2v_out.v:13606.21-13606.38" */
output [63:0] counter_val_upd_o;
wire [63:0] counter_val_upd_o;
/* cellift = 32'd1 */
output [63:0] counter_val_upd_o_t0;
wire [63:0] counter_val_upd_o_t0;
/* src = "generated/sv2v_out.v:13603.13-13603.25" */
input counter_we_i;
wire counter_we_i;
/* cellift = 32'd1 */
input counter_we_i_t0;
wire counter_we_i_t0;
/* src = "generated/sv2v_out.v:13602.13-13602.26" */
input counterh_we_i;
wire counterh_we_i;
/* cellift = 32'd1 */
input counterh_we_i_t0;
wire counterh_we_i_t0;
/* src = "generated/sv2v_out.v:13600.13-13600.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:13610.6-13610.8" */
wire we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13610.6-13610.8" */
wire we_t0;
assign counter_val_upd_o = counter_val_o + /* src = "generated/sv2v_out.v:13612.23-13612.86" */ 64'h0000000000000001;
assign _002_ = ~ counter_val_o_t0;
assign _028_ = counter_val_o & _002_;
assign _067_ = _028_ + 64'h0000000000000001;
assign _043_ = counter_val_o | counter_val_o_t0;
assign _068_ = _043_ + 64'h0000000000000001;
assign _061_ = _067_ ^ _068_;
assign counter_val_upd_o_t0 = _061_ | counter_val_o_t0;
assign _003_ = ~ _024_;
assign _004_ = ~ _026_;
assign _062_ = counter_d[63:32] ^ counter_val_o[63:32];
assign _063_ = counter_d[31:0] ^ counter_val_o[31:0];
assign _044_ = counter_d_t0[63:32] | counter_val_o_t0[63:32];
assign _048_ = counter_d_t0[31:0] | counter_val_o_t0[31:0];
assign _045_ = _062_ | _044_;
assign _049_ = _063_ | _048_;
assign _029_ = { _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_ } & counter_d_t0[63:32];
assign _032_ = { _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_ } & counter_d_t0[31:0];
assign _030_ = { _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_ } & counter_val_o_t0[63:32];
assign _033_ = { _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_ } & counter_val_o_t0[31:0];
assign _031_ = _045_ & { _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_ };
assign _034_ = _049_ & { _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_ };
assign _046_ = _029_ | _030_;
assign _050_ = _032_ | _033_;
assign _047_ = _046_ | _031_;
assign _051_ = _050_ | _034_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter  */
/* PC_TAINT_INFO STATE_NAME counter_val_o_t0[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o_t0[63:32] <= 32'd0;
else counter_val_o_t0[63:32] <= _047_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter  */
/* PC_TAINT_INFO STATE_NAME counter_val_o_t0[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o_t0[31:0] <= 32'd0;
else counter_val_o_t0[31:0] <= _051_;
assign _005_ = | { we_t0, counterh_we_i_t0 };
assign _006_ = ~ { we_t0, counterh_we_i_t0 };
assign _036_ = { we, counterh_we_i } & _006_;
assign _065_ = _036_ == { _006_[1], 1'h0 };
assign _066_ = _036_ == _006_;
assign _021_ = _065_ & _005_;
assign _023_ = _066_ & _005_;
/* src = "generated/sv2v_out.v:13629.2-13633.27" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter  */
/* PC_TAINT_INFO STATE_NAME counter_val_o[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o[63:32] <= 32'd0;
else if (_024_) counter_val_o[63:32] <= counter_d[63:32];
/* src = "generated/sv2v_out.v:13629.2-13633.27" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$c16eccae153ba9fb8fce8498c4f7e85e78010c3f\ibex_counter  */
/* PC_TAINT_INFO STATE_NAME counter_val_o[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o[31:0] <= 32'd0;
else if (_026_) counter_val_o[31:0] <= counter_d[31:0];
assign _007_ = | { we_t0, counter_inc_i_t0 };
assign _008_ = ~ { we_t0, counter_inc_i_t0 };
assign _035_ = { we, counter_inc_i } & _008_;
assign _009_ = ! _035_;
assign _019_ = _009_ & _007_;
assign _010_ = ~ { we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we };
assign _011_ = ~ { counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i };
assign _056_ = { we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0 } | _010_;
assign _059_ = { counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0 } | _011_;
assign _055_ = { counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0 } | { counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i };
assign _057_ = { we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0 } | { we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we };
assign _060_ = { counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0 } | { counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i };
assign _040_ = _001_ & _056_;
assign counter_load_t0[31:0] = counter_val_i_t0 & _059_;
assign _001_ = counter_val_upd_o_t0 & _055_;
assign _041_ = counter_load_t0 & _057_;
assign counter_load_t0[63:32] = counter_val_i_t0 & _060_;
assign _058_ = _040_ | _041_;
assign _064_ = _000_ ^ counter_load;
assign _042_ = { we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0 } & _064_;
assign counter_d_t0 = _042_ | _058_;
assign _018_ = | { we, counter_inc_i };
assign _020_ = { we, counterh_we_i } != 2'h2;
assign _022_ = { we, counterh_we_i } != 2'h3;
assign _024_ = & { _020_, _018_ };
assign _026_ = & { _018_, _022_ };
assign _012_ = ~ counter_we_i;
assign _013_ = ~ counterh_we_i;
assign _037_ = counter_we_i_t0 & _013_;
assign _038_ = counterh_we_i_t0 & _012_;
assign _039_ = counter_we_i_t0 & counterh_we_i_t0;
assign _054_ = _037_ | _038_;
assign we_t0 = _054_ | _039_;
assign _014_ = | { _021_, _019_ };
assign _015_ = | { _023_, _019_ };
assign _052_ = { _020_, _018_ } | { _021_, _019_ };
assign _053_ = { _018_, _022_ } | { _019_, _023_ };
assign _016_ = & _052_;
assign _017_ = & _053_;
assign _025_ = _014_ & _016_;
assign _027_ = _015_ & _017_;
assign we = counter_we_i | /* src = "generated/sv2v_out.v:13614.8-13614.36" */ counterh_we_i;
assign _000_ = counter_inc_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13623.12-13623.25|generated/sv2v_out.v:13623.8-13626.44" */ counter_val_upd_o : 64'hxxxxxxxxxxxxxxxx;
assign counter_d = we ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13621.7-13621.9|generated/sv2v_out.v:13621.3-13626.44" */ counter_load : _000_;
assign counter_load[63:32] = counterh_we_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13617.7-13617.20|generated/sv2v_out.v:13617.3-13620.6" */ counter_val_i : 32'hxxxxxxxx;
assign counter_load[31:0] = counterh_we_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13617.7-13617.20|generated/sv2v_out.v:13617.3-13620.6" */ 32'hxxxxxxxx : counter_val_i;
endmodule

module \$paramod$e55993a14b1fbc43320d549f521b710ed37596c6\ibex_csr (clk_i, rst_ni, wr_data_i, wr_en_i, rd_data_o, rd_error_o, rd_data_o_t0, rd_error_o_t0, wr_data_i_t0, wr_en_i_t0);
wire _00_;
wire [17:0] _01_;
wire [17:0] _02_;
wire [17:0] _03_;
wire [17:0] _04_;
wire [17:0] _05_;
wire [17:0] _06_;
wire [17:0] _07_;
wire [17:0] _08_;
/* src = "generated/sv2v_out.v:14871.13-14871.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:14875.28-14875.37" */
output [17:0] rd_data_o;
reg [17:0] rd_data_o;
/* cellift = 32'd1 */
output [17:0] rd_data_o_t0;
reg [17:0] rd_data_o_t0;
/* src = "generated/sv2v_out.v:14876.14-14876.24" */
output rd_error_o;
wire rd_error_o;
/* cellift = 32'd1 */
output rd_error_o_t0;
wire rd_error_o_t0;
/* src = "generated/sv2v_out.v:14872.13-14872.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:14873.27-14873.36" */
input [17:0] wr_data_i;
wire [17:0] wr_data_i;
/* cellift = 32'd1 */
input [17:0] wr_data_i_t0;
wire [17:0] wr_data_i_t0;
/* src = "generated/sv2v_out.v:14874.13-14874.20" */
input wr_en_i;
wire wr_en_i;
/* cellift = 32'd1 */
input wr_en_i_t0;
wire wr_en_i_t0;
assign _00_ = ~ wr_en_i;
assign _08_ = wr_data_i ^ rd_data_o;
assign _04_ = wr_data_i_t0 | rd_data_o_t0;
assign _05_ = _08_ | _04_;
assign _01_ = { wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i, wr_en_i } & wr_data_i_t0;
assign _02_ = { _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_, _00_ } & rd_data_o_t0;
assign _03_ = _05_ & { wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0, wr_en_i_t0 };
assign _06_ = _01_ | _02_;
assign _07_ = _06_ | _03_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$e55993a14b1fbc43320d549f521b710ed37596c6\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o_t0 <= 18'h00000;
else rd_data_o_t0 <= _07_;
/* src = "generated/sv2v_out.v:14878.2-14882.25" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$e55993a14b1fbc43320d549f521b710ed37596c6\ibex_csr  */
/* PC_TAINT_INFO STATE_NAME rd_data_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rd_data_o <= 18'h00000;
else if (wr_en_i) rd_data_o <= wr_data_i;
assign rd_error_o = 1'h0;
assign rd_error_o_t0 = 1'h0;
endmodule

module \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage (clk_i, rst_ni, ctrl_busy_o, illegal_insn_o, instr_valid_i, instr_rdata_i, instr_rdata_alu_i, instr_rdata_c_i, instr_is_compressed_i, instr_bp_taken_i, instr_req_o, instr_first_cycle_id_o, instr_valid_clear_o, id_in_ready_o, instr_exec_i, icache_inval_o, branch_decision_i, pc_set_o, pc_mux_o, nt_branch_mispredict_o, nt_branch_addr_o
, exc_pc_mux_o, exc_cause_o, illegal_c_insn_i, instr_fetch_err_i, instr_fetch_err_plus2_i, pc_id_i, ex_valid_i, lsu_resp_valid_i, alu_operator_ex_o, alu_operand_a_ex_o, alu_operand_b_ex_o, imd_val_we_ex_i, imd_val_d_ex_i, imd_val_q_ex_o, bt_a_operand_o, bt_b_operand_o, mult_en_ex_o, div_en_ex_o, mult_sel_ex_o, div_sel_ex_o, multdiv_operator_ex_o
, multdiv_signed_mode_ex_o, multdiv_operand_a_ex_o, multdiv_operand_b_ex_o, multdiv_ready_id_o, csr_access_o, csr_op_o, csr_op_en_o, csr_save_if_o, csr_save_id_o, csr_save_wb_o, csr_restore_mret_id_o, csr_restore_dret_id_o, csr_save_cause_o, csr_mtval_o, priv_mode_i, csr_mstatus_tw_i, illegal_csr_insn_i, data_ind_timing_i, lsu_req_o, lsu_we_o, lsu_type_o
, lsu_sign_ext_o, lsu_wdata_o, lsu_req_done_i, lsu_addr_incr_req_i, lsu_addr_last_i, csr_mstatus_mie_i, irq_pending_i, irqs_i, irq_nm_i, nmi_mode_o, lsu_load_err_i, lsu_load_resp_intg_err_i, lsu_store_err_i, lsu_store_resp_intg_err_i, debug_mode_o, debug_mode_entering_o, debug_cause_o, debug_csr_save_o, debug_req_i, debug_single_step_i, debug_ebreakm_i
, debug_ebreaku_i, trigger_match_i, result_ex_i, csr_rdata_i, rf_raddr_a_o, rf_rdata_a_i, rf_raddr_b_o, rf_rdata_b_i, rf_ren_a_o, rf_ren_b_o, rf_waddr_id_o, rf_wdata_id_o, rf_we_id_o, rf_rd_a_wb_match_o, rf_rd_b_wb_match_o, rf_waddr_wb_i, rf_wdata_fwd_wb_i, rf_write_wb_i, en_wb_o, instr_type_wb_o, instr_perf_count_id_o
, ready_wb_i, outstanding_load_wb_i, outstanding_store_wb_i, perf_jump_o, perf_branch_o, perf_tbranch_o, perf_dside_wait_o, perf_mul_wait_o, perf_div_wait_o, instr_id_done_o, rf_ren_b_o_t0, rf_raddr_b_o_t0, rf_ren_a_o_t0, rf_raddr_a_o_t0, csr_op_o_t0, csr_access_o_t0, instr_rdata_alu_i_t0, illegal_insn_o_t0, illegal_c_insn_i_t0, icache_inval_o_t0, csr_mstatus_mie_i_t0
, csr_mtval_o_t0, csr_restore_dret_id_o_t0, csr_restore_mret_id_o_t0, csr_save_cause_o_t0, csr_save_id_o_t0, csr_save_if_o_t0, csr_save_wb_o_t0, ctrl_busy_o_t0, debug_cause_o_t0, debug_csr_save_o_t0, debug_ebreakm_i_t0, debug_ebreaku_i_t0, debug_mode_entering_o_t0, debug_mode_o_t0, debug_req_i_t0, debug_single_step_i_t0, exc_cause_o_t0, exc_pc_mux_o_t0, id_in_ready_o_t0, instr_bp_taken_i_t0, instr_exec_i_t0
, instr_fetch_err_i_t0, instr_fetch_err_plus2_i_t0, instr_is_compressed_i_t0, instr_valid_clear_o_t0, instr_valid_i_t0, irq_pending_i_t0, irqs_i_t0, lsu_addr_last_i_t0, nmi_mode_o_t0, nt_branch_mispredict_o_t0, pc_id_i_t0, pc_mux_o_t0, pc_set_o_t0, perf_jump_o_t0, perf_tbranch_o_t0, priv_mode_i_t0, ready_wb_i_t0, trigger_match_i_t0, instr_req_o_t0, instr_rdata_i_t0, alu_operand_a_ex_o_t0
, alu_operand_b_ex_o_t0, alu_operator_ex_o_t0, branch_decision_i_t0, bt_a_operand_o_t0, bt_b_operand_o_t0, csr_mstatus_tw_i_t0, csr_op_en_o_t0, csr_rdata_i_t0, data_ind_timing_i_t0, div_en_ex_o_t0, div_sel_ex_o_t0, en_wb_o_t0, ex_valid_i_t0, illegal_csr_insn_i_t0, imd_val_d_ex_i_t0, imd_val_q_ex_o_t0, imd_val_we_ex_i_t0, instr_first_cycle_id_o_t0, instr_id_done_o_t0, instr_perf_count_id_o_t0, instr_rdata_c_i_t0
, instr_type_wb_o_t0, irq_nm_i_t0, lsu_addr_incr_req_i_t0, lsu_load_err_i_t0, lsu_load_resp_intg_err_i_t0, lsu_req_done_i_t0, lsu_req_o_t0, lsu_resp_valid_i_t0, lsu_sign_ext_o_t0, lsu_store_err_i_t0, lsu_store_resp_intg_err_i_t0, lsu_type_o_t0, lsu_wdata_o_t0, lsu_we_o_t0, mult_en_ex_o_t0, mult_sel_ex_o_t0, multdiv_operand_a_ex_o_t0, multdiv_operand_b_ex_o_t0, multdiv_operator_ex_o_t0, multdiv_ready_id_o_t0, multdiv_signed_mode_ex_o_t0
, nt_branch_addr_o_t0, outstanding_load_wb_i_t0, outstanding_store_wb_i_t0, perf_branch_o_t0, perf_div_wait_o_t0, perf_dside_wait_o_t0, perf_mul_wait_o_t0, result_ex_i_t0, rf_rd_a_wb_match_o_t0, rf_rd_b_wb_match_o_t0, rf_rdata_a_i_t0, rf_rdata_b_i_t0, rf_waddr_id_o_t0, rf_waddr_wb_i_t0, rf_wdata_fwd_wb_i_t0, rf_wdata_id_o_t0, rf_we_id_o_t0, rf_write_wb_i_t0);
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0001_;
/* src = "generated/sv2v_out.v:17474.2-17483.5" */
wire _0002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17474.2-17483.5" */
wire _0003_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0005_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0007_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0009_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0011_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0013_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0015_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0016_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0017_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0018_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0019_;
/* src = "generated/sv2v_out.v:17474.2-17483.5" */
wire _0020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17474.2-17483.5" */
wire _0021_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0022_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0023_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0024_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0025_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0026_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0027_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0028_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0029_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0030_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0031_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0032_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0033_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0034_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0035_;
/* src = "generated/sv2v_out.v:17474.2-17483.5" */
wire _0036_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17474.2-17483.5" */
wire _0037_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0038_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0039_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0040_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0041_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0042_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0043_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0044_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0045_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0046_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0047_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0048_;
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0049_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17628.2-17687.5" */
wire _0050_;
/* src = "generated/sv2v_out.v:17294.22-17294.56" */
wire _0051_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17294.22-17294.56" */
wire _0052_;
/* src = "generated/sv2v_out.v:17294.21-17294.75" */
wire _0053_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17294.21-17294.75" */
wire _0054_;
/* src = "generated/sv2v_out.v:17409.23-17409.50" */
wire _0055_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17409.23-17409.50" */
wire _0056_;
/* src = "generated/sv2v_out.v:17485.73-17485.104" */
wire _0057_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17485.73-17485.104" */
wire _0058_;
/* src = "generated/sv2v_out.v:17560.38-17560.68" */
wire _0059_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17560.38-17560.68" */
wire _0060_;
/* src = "generated/sv2v_out.v:17568.24-17568.54" */
wire _0061_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17568.24-17568.54" */
wire _0062_;
/* src = "generated/sv2v_out.v:17676.19-17676.41" */
wire _0063_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17676.19-17676.41" */
wire _0064_;
/* src = "generated/sv2v_out.v:17677.10-17677.38" */
wire _0065_;
/* src = "generated/sv2v_out.v:17690.23-17690.44" */
wire _0066_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17690.23-17690.44" */
wire _0067_;
/* src = "generated/sv2v_out.v:17725.40-17725.93" */
wire _0068_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17725.40-17725.93" */
wire _0069_;
/* src = "generated/sv2v_out.v:17751.32-17751.61" */
wire _0070_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17751.32-17751.61" */
wire _0071_;
/* src = "generated/sv2v_out.v:17755.36-17755.64" */
wire _0072_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17755.36-17755.64" */
wire _0073_;
/* src = "generated/sv2v_out.v:17755.35-17755.85" */
wire _0074_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17755.35-17755.85" */
wire _0075_;
/* src = "generated/sv2v_out.v:17755.34-17755.108" */
wire _0076_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17755.34-17755.108" */
wire _0077_;
wire _0078_;
wire _0079_;
wire _0080_;
wire _0081_;
wire _0082_;
wire _0083_;
wire _0084_;
wire _0085_;
wire _0086_;
wire [1:0] _0087_;
wire [11:0] _0088_;
wire [6:0] _0089_;
wire [1:0] _0090_;
wire [2:0] _0091_;
wire [1:0] _0092_;
wire _0093_;
wire [2:0] _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire _0109_;
wire _0110_;
wire _0111_;
wire _0112_;
wire _0113_;
wire [31:0] _0114_;
wire [31:0] _0115_;
wire [31:0] _0116_;
wire [31:0] _0117_;
wire [31:0] _0118_;
wire _0119_;
wire [31:0] _0120_;
wire [31:0] _0121_;
wire [31:0] _0122_;
wire [31:0] _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire [1:0] _0131_;
wire _0132_;
wire [2:0] _0133_;
wire [31:0] _0134_;
wire [31:0] _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire [1:0] _0139_;
wire _0140_;
wire _0141_;
wire _0142_;
wire _0143_;
wire _0144_;
wire _0145_;
wire _0146_;
wire _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
wire _0152_;
wire _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
wire _0166_;
wire _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
/* cellift = 32'd1 */
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire _0186_;
wire _0187_;
wire _0188_;
wire _0189_;
wire _0190_;
wire _0191_;
wire _0192_;
wire _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire _0199_;
wire _0200_;
wire _0201_;
wire _0202_;
wire _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
wire _0221_;
wire _0222_;
wire _0223_;
wire _0224_;
wire _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire _0241_;
wire _0242_;
wire _0243_;
wire _0244_;
wire _0245_;
wire _0246_;
wire _0247_;
wire _0248_;
wire _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire [33:0] _0270_;
wire [33:0] _0271_;
wire [33:0] _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire [33:0] _0276_;
wire [33:0] _0277_;
wire [33:0] _0278_;
wire _0279_;
wire _0280_;
wire _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire [2:0] _0285_;
wire [31:0] _0286_;
wire [31:0] _0287_;
wire [31:0] _0288_;
wire [31:0] _0289_;
wire [31:0] _0290_;
wire [31:0] _0291_;
wire [31:0] _0292_;
wire [31:0] _0293_;
wire [31:0] _0294_;
wire [31:0] _0295_;
wire [31:0] _0296_;
wire [31:0] _0297_;
wire [31:0] _0298_;
wire [31:0] _0299_;
wire [31:0] _0300_;
wire [31:0] _0301_;
wire [31:0] _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire _0324_;
wire [31:0] _0325_;
wire [31:0] _0326_;
wire [31:0] _0327_;
wire [31:0] _0328_;
wire [31:0] _0329_;
wire [31:0] _0330_;
wire [31:0] _0331_;
wire [31:0] _0332_;
wire [31:0] _0333_;
wire [31:0] _0334_;
wire [31:0] _0335_;
wire [31:0] _0336_;
wire [1:0] _0337_;
wire [11:0] _0338_;
wire [6:0] _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire _0344_;
wire _0345_;
wire _0346_;
wire _0347_;
wire _0348_;
wire _0349_;
wire _0350_;
wire _0351_;
wire _0352_;
wire _0353_;
wire _0354_;
wire _0355_;
wire _0356_;
wire _0357_;
wire _0358_;
wire _0359_;
wire _0360_;
wire _0361_;
wire _0362_;
wire _0363_;
wire _0364_;
wire _0365_;
wire _0366_;
wire _0367_;
wire _0368_;
wire _0369_;
wire [1:0] _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire _0376_;
wire _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire _0382_;
wire _0383_;
wire _0384_;
wire _0385_;
wire _0386_;
wire _0387_;
wire _0388_;
wire _0389_;
wire _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire _0398_;
wire _0399_;
wire _0400_;
wire _0401_;
wire _0402_;
wire _0403_;
wire _0404_;
wire _0405_;
wire _0406_;
wire _0407_;
wire _0408_;
wire _0409_;
wire _0410_;
wire _0411_;
wire _0412_;
wire [2:0] _0413_;
wire _0414_;
wire _0415_;
wire _0416_;
wire _0417_;
wire _0418_;
wire _0419_;
wire _0420_;
wire _0421_;
wire _0422_;
wire _0423_;
wire _0424_;
wire _0425_;
wire _0426_;
wire _0427_;
wire _0428_;
wire _0429_;
wire _0430_;
wire _0431_;
wire _0432_;
wire _0433_;
wire _0434_;
wire _0435_;
wire _0436_;
wire _0437_;
wire _0438_;
wire _0439_;
wire _0440_;
wire _0441_;
wire _0442_;
wire _0443_;
wire _0444_;
wire _0445_;
wire _0446_;
wire _0447_;
wire _0448_;
wire _0449_;
wire _0450_;
wire _0451_;
wire _0452_;
wire _0453_;
wire _0454_;
wire _0455_;
wire _0456_;
wire _0457_;
wire _0458_;
wire _0459_;
wire _0460_;
wire _0461_;
wire _0462_;
wire _0463_;
wire _0464_;
wire _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire _0469_;
wire _0470_;
wire _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire _0477_;
wire _0478_;
wire _0479_;
wire _0480_;
wire _0481_;
wire _0482_;
wire _0483_;
wire _0484_;
wire _0485_;
wire _0486_;
wire _0487_;
wire _0488_;
wire _0489_;
wire _0490_;
wire _0491_;
wire _0492_;
wire _0493_;
wire _0494_;
wire _0495_;
wire _0496_;
wire _0497_;
wire _0498_;
wire _0499_;
wire _0500_;
wire _0501_;
wire _0502_;
wire [1:0] _0503_;
wire [1:0] _0504_;
wire [1:0] _0505_;
wire _0506_;
wire _0507_;
wire [2:0] _0508_;
wire [2:0] _0509_;
wire [31:0] _0510_;
wire [31:0] _0511_;
wire [31:0] _0512_;
wire [31:0] _0513_;
wire [31:0] _0514_;
wire _0515_;
wire _0516_;
wire _0517_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
/* cellift = 32'd1 */
wire _0525_;
wire _0526_;
/* cellift = 32'd1 */
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire _0534_;
wire _0535_;
wire _0536_;
wire _0537_;
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0542_;
wire _0543_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire [33:0] _0560_;
wire [33:0] _0561_;
wire [33:0] _0562_;
wire [33:0] _0563_;
wire _0564_;
wire _0565_;
wire _0566_;
wire _0567_;
wire [33:0] _0568_;
wire [33:0] _0569_;
wire [33:0] _0570_;
wire [33:0] _0571_;
wire _0572_;
wire _0573_;
wire [31:0] _0574_;
wire [31:0] _0575_;
wire [31:0] _0576_;
wire [31:0] _0577_;
wire [31:0] _0578_;
wire [31:0] _0579_;
wire [31:0] _0580_;
wire [31:0] _0581_;
wire [31:0] _0582_;
wire [31:0] _0583_;
wire [31:0] _0584_;
wire [31:0] _0585_;
wire [31:0] _0586_;
wire [31:0] _0587_;
wire [31:0] _0588_;
wire [31:0] _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire _0596_;
wire [31:0] _0597_;
wire [31:0] _0598_;
wire [31:0] _0599_;
wire [31:0] _0600_;
wire [31:0] _0601_;
wire [31:0] _0602_;
wire [31:0] _0603_;
wire [31:0] _0604_;
wire [31:0] _0605_;
wire [31:0] _0606_;
wire [31:0] _0607_;
wire [31:0] _0608_;
wire _0609_;
wire _0610_;
wire _0611_;
wire _0612_;
wire _0613_;
wire _0614_;
wire _0615_;
wire _0616_;
wire _0617_;
wire _0618_;
wire _0619_;
wire _0620_;
wire _0621_;
wire _0622_;
wire _0623_;
wire _0624_;
wire _0625_;
wire _0626_;
wire _0627_;
wire _0628_;
wire _0629_;
wire _0630_;
wire _0631_;
wire _0632_;
wire _0633_;
wire _0634_;
wire _0635_;
wire _0636_;
wire _0637_;
wire _0638_;
wire _0639_;
wire _0640_;
wire _0641_;
wire _0642_;
wire _0643_;
wire _0644_;
wire _0645_;
wire _0646_;
wire _0647_;
wire _0648_;
wire _0649_;
wire _0650_;
wire _0651_;
wire _0652_;
wire _0653_;
wire _0654_;
wire _0655_;
wire _0656_;
wire _0657_;
wire [1:0] _0658_;
wire _0659_;
wire [2:0] _0660_;
wire [31:0] _0661_;
wire [31:0] _0662_;
wire [31:0] _0663_;
wire [31:0] _0664_;
wire _0665_;
wire [33:0] _0666_;
wire _0667_;
wire [33:0] _0668_;
wire [31:0] _0669_;
wire [31:0] _0670_;
wire [31:0] _0671_;
wire [31:0] _0672_;
wire [31:0] _0673_;
wire _0674_;
wire _0675_;
wire _0676_;
wire _0677_;
wire _0678_;
wire [31:0] _0679_;
wire [31:0] _0680_;
wire [31:0] _0681_;
wire [31:0] _0682_;
wire _0683_;
wire _0684_;
wire _0685_;
wire _0686_;
wire _0687_;
wire _0688_;
wire _0689_;
wire _0690_;
wire _0691_;
wire _0692_;
wire _0693_;
wire _0694_;
wire _0695_;
wire _0696_;
wire _0697_;
wire _0698_;
wire _0699_;
wire _0700_;
wire _0701_;
wire _0702_;
wire _0703_;
wire _0704_;
wire _0705_;
wire _0706_;
wire _0707_;
wire [31:0] _0708_;
wire _0709_;
wire _0710_;
wire _0711_;
wire _0712_;
wire _0713_;
wire _0714_;
wire _0715_;
wire _0716_;
wire _0717_;
wire _0718_;
wire _0719_;
wire _0720_;
wire _0721_;
wire _0722_;
wire _0723_;
wire _0724_;
wire _0725_;
wire _0726_;
wire _0727_;
wire _0728_;
wire [31:0] _0729_;
/* cellift = 32'd1 */
wire [31:0] _0730_;
wire [31:0] _0731_;
/* cellift = 32'd1 */
wire [31:0] _0732_;
wire [31:0] _0733_;
/* cellift = 32'd1 */
wire [31:0] _0734_;
wire [31:0] _0735_;
/* cellift = 32'd1 */
wire [31:0] _0736_;
wire [31:0] _0737_;
/* cellift = 32'd1 */
wire [31:0] _0738_;
wire [31:0] _0739_;
/* cellift = 32'd1 */
wire [31:0] _0740_;
wire [31:0] _0741_;
/* cellift = 32'd1 */
wire [31:0] _0742_;
/* src = "generated/sv2v_out.v:17476.34-17476.50" */
wire _0743_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17476.34-17476.50" */
wire _0744_;
/* src = "generated/sv2v_out.v:17476.56-17476.72" */
wire _0745_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17476.56-17476.72" */
wire _0746_;
/* src = "generated/sv2v_out.v:17477.11-17477.42" */
wire _0747_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17477.11-17477.42" */
wire _0748_;
/* src = "generated/sv2v_out.v:17477.48-17477.79" */
wire _0749_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17477.48-17477.79" */
wire _0750_;
/* src = "generated/sv2v_out.v:17477.86-17477.117" */
wire _0751_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17477.86-17477.117" */
wire _0752_;
/* src = "generated/sv2v_out.v:17477.124-17477.153" */
wire _0753_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17477.124-17477.153" */
wire _0754_;
/* src = "generated/sv2v_out.v:17481.11-17481.42" */
wire _0755_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17481.11-17481.42" */
wire _0756_;
/* src = "generated/sv2v_out.v:17481.48-17481.79" */
wire _0757_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17481.48-17481.79" */
wire _0758_;
/* src = "generated/sv2v_out.v:17481.86-17481.117" */
wire _0759_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17481.86-17481.117" */
wire _0760_;
/* src = "generated/sv2v_out.v:17481.124-17481.155" */
wire _0761_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17481.124-17481.155" */
wire _0762_;
/* src = "generated/sv2v_out.v:17476.7-17476.74" */
wire _0763_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17476.7-17476.74" */
wire _0764_;
/* src = "generated/sv2v_out.v:17480.12-17480.55" */
wire _0765_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17480.12-17480.55" */
wire _0766_;
/* src = "generated/sv2v_out.v:17476.33-17476.73" */
wire _0767_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17476.33-17476.73" */
wire _0768_;
/* src = "generated/sv2v_out.v:17477.10-17477.80" */
wire _0769_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17477.10-17477.80" */
wire _0770_;
/* src = "generated/sv2v_out.v:17477.9-17477.118" */
wire _0771_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17477.9-17477.118" */
wire _0772_;
/* src = "generated/sv2v_out.v:17477.8-17477.154" */
wire _0773_;
/* src = "generated/sv2v_out.v:17481.10-17481.80" */
wire _0774_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17481.10-17481.80" */
wire _0775_;
/* src = "generated/sv2v_out.v:17481.9-17481.118" */
wire _0776_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17481.9-17481.118" */
wire _0777_;
/* src = "generated/sv2v_out.v:17481.8-17481.156" */
wire _0778_;
/* src = "generated/sv2v_out.v:17655.20-17655.80" */
wire _0779_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17655.20-17655.80" */
wire _0780_;
/* src = "generated/sv2v_out.v:17480.38-17480.54" */
wire _0781_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17480.38-17480.54" */
wire _0782_;
/* src = "generated/sv2v_out.v:17485.31-17485.51" */
wire _0783_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17485.31-17485.51" */
wire _0784_;
/* src = "generated/sv2v_out.v:17294.38-17294.56" */
wire _0785_;
/* src = "generated/sv2v_out.v:17294.60-17294.75" */
wire _0786_;
/* src = "generated/sv2v_out.v:17484.45-17484.58" */
wire _0787_;
/* src = "generated/sv2v_out.v:17592.95-17592.115" */
wire _0788_;
/* src = "generated/sv2v_out.v:17690.23-17690.32" */
wire _0789_;
/* src = "generated/sv2v_out.v:17690.35-17690.44" */
wire _0790_;
/* src = "generated/sv2v_out.v:17725.55-17725.72" */
wire _0791_;
/* src = "generated/sv2v_out.v:17755.36-17755.46" */
wire _0792_;
/* src = "generated/sv2v_out.v:17755.49-17755.64" */
wire _0793_;
/* src = "generated/sv2v_out.v:17485.56-17485.105" */
wire _0794_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17485.56-17485.105" */
wire _0795_;
/* src = "generated/sv2v_out.v:17486.45-17486.82" */
wire _0796_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17486.45-17486.82" */
wire _0797_;
/* src = "generated/sv2v_out.v:17486.44-17486.103" */
wire _0798_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17486.44-17486.103" */
wire _0799_;
/* src = "generated/sv2v_out.v:17486.43-17486.125" */
wire _0800_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17486.43-17486.125" */
wire _0801_;
/* src = "generated/sv2v_out.v:17592.36-17592.65" */
wire _0802_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17592.36-17592.65" */
wire _0803_;
/* src = "generated/sv2v_out.v:17592.35-17592.91" */
wire _0804_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17592.35-17592.91" */
wire _0805_;
/* src = "generated/sv2v_out.v:17689.23-17689.64" */
wire _0806_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17689.23-17689.64" */
wire _0807_;
/* src = "generated/sv2v_out.v:17689.22-17689.78" */
wire _0808_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17689.22-17689.78" */
wire _0809_;
/* src = "generated/sv2v_out.v:17689.21-17689.94" */
wire _0810_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17689.21-17689.94" */
wire _0811_;
/* src = "generated/sv2v_out.v:17725.55-17725.92" */
wire _0812_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17725.55-17725.92" */
wire _0813_;
wire _0814_;
/* cellift = 32'd1 */
wire _0815_;
wire _0816_;
/* cellift = 32'd1 */
wire _0817_;
wire _0818_;
/* cellift = 32'd1 */
wire _0819_;
wire _0820_;
/* cellift = 32'd1 */
wire _0821_;
wire _0822_;
/* cellift = 32'd1 */
wire _0823_;
wire _0824_;
/* cellift = 32'd1 */
wire _0825_;
wire _0826_;
/* cellift = 32'd1 */
wire _0827_;
wire _0828_;
/* cellift = 32'd1 */
wire _0829_;
wire _0830_;
/* cellift = 32'd1 */
wire _0831_;
/* cellift = 32'd1 */
wire _0832_;
/* cellift = 32'd1 */
wire _0833_;
/* cellift = 32'd1 */
wire _0834_;
wire _0835_;
/* cellift = 32'd1 */
wire _0836_;
wire _0837_;
/* cellift = 32'd1 */
wire _0838_;
wire _0839_;
/* cellift = 32'd1 */
wire _0840_;
wire _0841_;
/* cellift = 32'd1 */
wire _0842_;
/* cellift = 32'd1 */
wire _0843_;
/* cellift = 32'd1 */
wire _0844_;
/* cellift = 32'd1 */
wire _0845_;
/* cellift = 32'd1 */
wire _0846_;
/* cellift = 32'd1 */
wire _0847_;
/* cellift = 32'd1 */
wire _0848_;
/* cellift = 32'd1 */
wire _0849_;
/* cellift = 32'd1 */
wire _0850_;
/* cellift = 32'd1 */
wire _0851_;
wire _0852_;
/* cellift = 32'd1 */
wire _0853_;
wire _0854_;
/* cellift = 32'd1 */
wire _0855_;
wire _0856_;
/* cellift = 32'd1 */
wire _0857_;
/* src = "generated/sv2v_out.v:17389.21-17389.72" */
wire [31:0] _0858_;
/* src = "generated/sv2v_out.v:17655.20-17655.94" */
wire _0859_;
/* src = "generated/sv2v_out.v:17305.7-17305.25" */
wire alu_multicycle_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17305.7-17305.25" */
wire alu_multicycle_dec_t0;
/* src = "generated/sv2v_out.v:17301.13-17301.29" */
wire [1:0] alu_op_a_mux_sel;
/* src = "generated/sv2v_out.v:17302.13-17302.33" */
wire [1:0] alu_op_a_mux_sel_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17302.13-17302.33" */
wire [1:0] alu_op_a_mux_sel_dec_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17301.13-17301.29" */
wire [1:0] alu_op_a_mux_sel_t0;
/* src = "generated/sv2v_out.v:17303.7-17303.23" */
wire alu_op_b_mux_sel;
/* src = "generated/sv2v_out.v:17304.7-17304.27" */
wire alu_op_b_mux_sel_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17304.7-17304.27" */
wire alu_op_b_mux_sel_dec_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17303.7-17303.23" */
wire alu_op_b_mux_sel_t0;
/* src = "generated/sv2v_out.v:17157.21-17157.39" */
output [31:0] alu_operand_a_ex_o;
wire [31:0] alu_operand_a_ex_o;
/* cellift = 32'd1 */
output [31:0] alu_operand_a_ex_o_t0;
wire [31:0] alu_operand_a_ex_o_t0;
/* src = "generated/sv2v_out.v:17158.21-17158.39" */
output [31:0] alu_operand_b_ex_o;
wire [31:0] alu_operand_b_ex_o;
/* cellift = 32'd1 */
output [31:0] alu_operand_b_ex_o_t0;
wire [31:0] alu_operand_b_ex_o_t0;
/* src = "generated/sv2v_out.v:17156.20-17156.37" */
output [6:0] alu_operator_ex_o;
wire [6:0] alu_operator_ex_o;
/* cellift = 32'd1 */
output [6:0] alu_operator_ex_o_t0;
wire [6:0] alu_operator_ex_o_t0;
/* src = "generated/sv2v_out.v:17143.13-17143.30" */
input branch_decision_i;
wire branch_decision_i;
/* cellift = 32'd1 */
input branch_decision_i_t0;
wire branch_decision_i_t0;
/* src = "generated/sv2v_out.v:17252.7-17252.20" */
wire branch_in_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17252.7-17252.20" */
wire branch_in_dec_t0;
/* src = "generated/sv2v_out.v:17257.7-17257.29" */
wire branch_jump_set_done_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17257.7-17257.29" */
wire branch_jump_set_done_d_t0;
/* src = "generated/sv2v_out.v:17256.6-17256.28" */
reg branch_jump_set_done_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17256.6-17256.28" */
reg branch_jump_set_done_q_t0;
/* src = "generated/sv2v_out.v:17253.7-17253.17" */
wire branch_set;
/* src = "generated/sv2v_out.v:17254.7-17254.21" */
reg branch_set_raw;
/* src = "generated/sv2v_out.v:17255.6-17255.22" */
wire branch_set_raw_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17255.6-17255.22" */
wire branch_set_raw_d_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17254.7-17254.21" */
reg branch_set_raw_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17253.7-17253.17" */
wire branch_set_t0;
/* src = "generated/sv2v_out.v:17259.7-17259.19" */
wire branch_taken;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17259.7-17259.19" */
wire branch_taken_t0;
/* src = "generated/sv2v_out.v:17308.13-17308.25" */
/* unused_bits = "0 1" */
wire [1:0] bt_a_mux_sel;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17308.13-17308.25" */
/* unused_bits = "0 1" */
wire [1:0] bt_a_mux_sel_t0;
/* src = "generated/sv2v_out.v:17162.20-17162.34" */
output [31:0] bt_a_operand_o;
wire [31:0] bt_a_operand_o;
/* cellift = 32'd1 */
output [31:0] bt_a_operand_o_t0;
wire [31:0] bt_a_operand_o_t0;
/* src = "generated/sv2v_out.v:17309.13-17309.25" */
/* unused_bits = "0 1 2" */
wire [2:0] bt_b_mux_sel;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17309.13-17309.25" */
/* unused_bits = "0 1 2" */
wire [2:0] bt_b_mux_sel_t0;
/* src = "generated/sv2v_out.v:17163.20-17163.34" */
output [31:0] bt_b_operand_o;
wire [31:0] bt_b_operand_o;
/* cellift = 32'd1 */
output [31:0] bt_b_operand_o_t0;
wire [31:0] bt_b_operand_o_t0;
/* src = "generated/sv2v_out.v:17127.13-17127.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:17268.7-17268.21" */
wire controller_run;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17268.7-17268.21" */
wire controller_run_t0;
/* src = "generated/sv2v_out.v:17173.14-17173.26" */
output csr_access_o;
wire csr_access_o;
/* cellift = 32'd1 */
output csr_access_o_t0;
wire csr_access_o_t0;
/* src = "generated/sv2v_out.v:17195.13-17195.30" */
input csr_mstatus_mie_i;
wire csr_mstatus_mie_i;
/* cellift = 32'd1 */
input csr_mstatus_mie_i_t0;
wire csr_mstatus_mie_i_t0;
/* src = "generated/sv2v_out.v:17184.13-17184.29" */
input csr_mstatus_tw_i;
wire csr_mstatus_tw_i;
/* cellift = 32'd1 */
input csr_mstatus_tw_i_t0;
wire csr_mstatus_tw_i_t0;
/* src = "generated/sv2v_out.v:17182.21-17182.32" */
output [31:0] csr_mtval_o;
wire [31:0] csr_mtval_o;
/* cellift = 32'd1 */
output [31:0] csr_mtval_o_t0;
wire [31:0] csr_mtval_o_t0;
/* src = "generated/sv2v_out.v:17175.14-17175.25" */
output csr_op_en_o;
wire csr_op_en_o;
/* cellift = 32'd1 */
output csr_op_en_o_t0;
wire csr_op_en_o_t0;
/* src = "generated/sv2v_out.v:17174.20-17174.28" */
output [1:0] csr_op_o;
wire [1:0] csr_op_o;
/* cellift = 32'd1 */
output [1:0] csr_op_o_t0;
wire [1:0] csr_op_o_t0;
/* src = "generated/sv2v_out.v:17326.6-17326.20" */
wire csr_pipe_flush;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17326.6-17326.20" */
wire csr_pipe_flush_t0;
/* src = "generated/sv2v_out.v:17214.20-17214.31" */
input [31:0] csr_rdata_i;
wire [31:0] csr_rdata_i;
/* cellift = 32'd1 */
input [31:0] csr_rdata_i_t0;
wire [31:0] csr_rdata_i_t0;
/* src = "generated/sv2v_out.v:17180.14-17180.35" */
output csr_restore_dret_id_o;
wire csr_restore_dret_id_o;
/* cellift = 32'd1 */
output csr_restore_dret_id_o_t0;
wire csr_restore_dret_id_o_t0;
/* src = "generated/sv2v_out.v:17179.14-17179.35" */
output csr_restore_mret_id_o;
wire csr_restore_mret_id_o;
/* cellift = 32'd1 */
output csr_restore_mret_id_o_t0;
wire csr_restore_mret_id_o_t0;
/* src = "generated/sv2v_out.v:17181.14-17181.30" */
output csr_save_cause_o;
wire csr_save_cause_o;
/* cellift = 32'd1 */
output csr_save_cause_o_t0;
wire csr_save_cause_o_t0;
/* src = "generated/sv2v_out.v:17177.14-17177.27" */
output csr_save_id_o;
wire csr_save_id_o;
/* cellift = 32'd1 */
output csr_save_id_o_t0;
wire csr_save_id_o_t0;
/* src = "generated/sv2v_out.v:17176.14-17176.27" */
output csr_save_if_o;
wire csr_save_if_o;
/* cellift = 32'd1 */
output csr_save_if_o_t0;
wire csr_save_if_o_t0;
/* src = "generated/sv2v_out.v:17178.14-17178.27" */
output csr_save_wb_o;
wire csr_save_wb_o;
/* cellift = 32'd1 */
output csr_save_wb_o_t0;
wire csr_save_wb_o_t0;
/* src = "generated/sv2v_out.v:17129.14-17129.25" */
output ctrl_busy_o;
wire ctrl_busy_o;
/* cellift = 32'd1 */
output ctrl_busy_o_t0;
wire ctrl_busy_o_t0;
/* src = "generated/sv2v_out.v:17186.13-17186.30" */
input data_ind_timing_i;
wire data_ind_timing_i;
/* cellift = 32'd1 */
input data_ind_timing_i_t0;
wire data_ind_timing_i_t0;
/* src = "generated/sv2v_out.v:17206.20-17206.33" */
output [2:0] debug_cause_o;
wire [2:0] debug_cause_o;
/* cellift = 32'd1 */
output [2:0] debug_cause_o_t0;
wire [2:0] debug_cause_o_t0;
/* src = "generated/sv2v_out.v:17207.14-17207.30" */
output debug_csr_save_o;
wire debug_csr_save_o;
/* cellift = 32'd1 */
output debug_csr_save_o_t0;
wire debug_csr_save_o_t0;
/* src = "generated/sv2v_out.v:17210.13-17210.28" */
input debug_ebreakm_i;
wire debug_ebreakm_i;
/* cellift = 32'd1 */
input debug_ebreakm_i_t0;
wire debug_ebreakm_i_t0;
/* src = "generated/sv2v_out.v:17211.13-17211.28" */
input debug_ebreaku_i;
wire debug_ebreaku_i;
/* cellift = 32'd1 */
input debug_ebreaku_i_t0;
wire debug_ebreaku_i_t0;
/* src = "generated/sv2v_out.v:17205.14-17205.35" */
output debug_mode_entering_o;
wire debug_mode_entering_o;
/* cellift = 32'd1 */
output debug_mode_entering_o_t0;
wire debug_mode_entering_o_t0;
/* src = "generated/sv2v_out.v:17204.14-17204.26" */
output debug_mode_o;
wire debug_mode_o;
/* cellift = 32'd1 */
output debug_mode_o_t0;
wire debug_mode_o_t0;
/* src = "generated/sv2v_out.v:17208.13-17208.24" */
input debug_req_i;
wire debug_req_i;
/* cellift = 32'd1 */
input debug_req_i_t0;
wire debug_req_i_t0;
/* src = "generated/sv2v_out.v:17209.13-17209.32" */
input debug_single_step_i;
wire debug_single_step_i;
/* cellift = 32'd1 */
input debug_single_step_i_t0;
wire debug_single_step_i_t0;
/* src = "generated/sv2v_out.v:17316.7-17316.17" */
wire div_en_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17316.7-17316.17" */
wire div_en_dec_t0;
/* src = "generated/sv2v_out.v:17165.14-17165.25" */
output div_en_ex_o;
wire div_en_ex_o;
/* cellift = 32'd1 */
output div_en_ex_o_t0;
wire div_en_ex_o_t0;
/* src = "generated/sv2v_out.v:17167.14-17167.26" */
output div_sel_ex_o;
wire div_sel_ex_o;
/* cellift = 32'd1 */
output div_sel_ex_o_t0;
wire div_sel_ex_o_t0;
/* src = "generated/sv2v_out.v:17247.7-17247.20" */
wire dret_insn_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17247.7-17247.20" */
wire dret_insn_dec_t0;
/* src = "generated/sv2v_out.v:17245.7-17245.16" */
wire ebrk_insn;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17245.7-17245.16" */
wire ebrk_insn_t0;
/* src = "generated/sv2v_out.v:17248.7-17248.21" */
wire ecall_insn_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17248.7-17248.21" */
wire ecall_insn_dec_t0;
/* src = "generated/sv2v_out.v:17229.14-17229.21" */
output en_wb_o;
wire en_wb_o;
/* cellift = 32'd1 */
output en_wb_o_t0;
wire en_wb_o_t0;
/* src = "generated/sv2v_out.v:17154.13-17154.23" */
input ex_valid_i;
wire ex_valid_i;
/* cellift = 32'd1 */
input ex_valid_i_t0;
wire ex_valid_i_t0;
/* src = "generated/sv2v_out.v:17149.20-17149.31" */
output [6:0] exc_cause_o;
wire [6:0] exc_cause_o;
/* cellift = 32'd1 */
output [6:0] exc_cause_o_t0;
wire [6:0] exc_cause_o_t0;
/* src = "generated/sv2v_out.v:17148.20-17148.32" */
output [1:0] exc_pc_mux_o;
wire [1:0] exc_pc_mux_o;
/* cellift = 32'd1 */
output [1:0] exc_pc_mux_o_t0;
wire [1:0] exc_pc_mux_o_t0;
/* src = "generated/sv2v_out.v:17276.7-17276.15" */
wire flush_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17276.7-17276.15" */
wire flush_id_t0;
/* src = "generated/sv2v_out.v:17602.8-17602.22" */
reg \g_sec_branch_taken.branch_taken_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17602.8-17602.22" */
reg \g_sec_branch_taken.branch_taken_q_t0 ;
/* src = "generated/sv2v_out.v:17740.9-17740.28" */
/* unused_bits = "0" */
wire \gen_no_stall_mem.unused_id_exception ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17740.9-17740.28" */
/* unused_bits = "0" */
wire \gen_no_stall_mem.unused_id_exception_t0 ;
/* src = "generated/sv2v_out.v:17738.9-17738.28" */
/* unused_bits = "0" */
wire \gen_no_stall_mem.unused_wb_exception ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17738.9-17738.28" */
/* unused_bits = "0" */
wire \gen_no_stall_mem.unused_wb_exception_t0 ;
/* src = "generated/sv2v_out.v:17142.14-17142.28" */
output icache_inval_o;
wire icache_inval_o;
/* cellift = 32'd1 */
output icache_inval_o_t0;
wire icache_inval_o_t0;
/* src = "generated/sv2v_out.v:17621.6-17621.14" */
wire id_fsm_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17621.6-17621.14" */
wire id_fsm_d_t0;
/* src = "generated/sv2v_out.v:17620.6-17620.14" */
reg id_fsm_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17620.6-17620.14" */
reg id_fsm_q_t0;
/* src = "generated/sv2v_out.v:17140.14-17140.27" */
output id_in_ready_o;
wire id_in_ready_o;
/* cellift = 32'd1 */
output id_in_ready_o_t0;
wire id_in_ready_o_t0;
/* src = "generated/sv2v_out.v:17150.13-17150.29" */
input illegal_c_insn_i;
wire illegal_c_insn_i;
/* cellift = 32'd1 */
input illegal_c_insn_i_t0;
wire illegal_c_insn_i_t0;
/* src = "generated/sv2v_out.v:17185.13-17185.31" */
input illegal_csr_insn_i;
wire illegal_csr_insn_i;
/* cellift = 32'd1 */
input illegal_csr_insn_i_t0;
wire illegal_csr_insn_i_t0;
/* src = "generated/sv2v_out.v:17243.7-17243.24" */
wire illegal_dret_insn;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17243.7-17243.24" */
wire illegal_dret_insn_t0;
/* src = "generated/sv2v_out.v:17242.7-17242.23" */
wire illegal_insn_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17242.7-17242.23" */
wire illegal_insn_dec_t0;
/* src = "generated/sv2v_out.v:17130.14-17130.28" */
output illegal_insn_o;
wire illegal_insn_o;
/* cellift = 32'd1 */
output illegal_insn_o_t0;
wire illegal_insn_o_t0;
/* src = "generated/sv2v_out.v:17244.7-17244.25" */
wire illegal_umode_insn;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17244.7-17244.25" */
wire illegal_umode_insn_t0;
/* src = "generated/sv2v_out.v:17160.20-17160.34" */
input [67:0] imd_val_d_ex_i;
wire [67:0] imd_val_d_ex_i;
/* cellift = 32'd1 */
input [67:0] imd_val_d_ex_i_t0;
wire [67:0] imd_val_d_ex_i_t0;
/* src = "generated/sv2v_out.v:17161.21-17161.35" */
output [67:0] imd_val_q_ex_o;
reg [67:0] imd_val_q_ex_o;
/* cellift = 32'd1 */
output [67:0] imd_val_q_ex_o_t0;
reg [67:0] imd_val_q_ex_o_t0;
/* src = "generated/sv2v_out.v:17159.19-17159.34" */
input [1:0] imd_val_we_ex_i;
wire [1:0] imd_val_we_ex_i;
/* cellift = 32'd1 */
input [1:0] imd_val_we_ex_i_t0;
wire [1:0] imd_val_we_ex_i_t0;
/* src = "generated/sv2v_out.v:17285.14-17285.19" */
wire [31:0] imm_a;
/* src = "generated/sv2v_out.v:17310.7-17310.20" */
wire imm_a_mux_sel;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17310.7-17310.20" */
wire imm_a_mux_sel_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17285.14-17285.19" */
wire [31:0] imm_a_t0;
/* src = "generated/sv2v_out.v:17286.13-17286.18" */
wire [31:0] imm_b;
/* src = "generated/sv2v_out.v:17311.13-17311.26" */
wire [2:0] imm_b_mux_sel;
/* src = "generated/sv2v_out.v:17312.13-17312.30" */
wire [2:0] imm_b_mux_sel_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17312.13-17312.30" */
wire [2:0] imm_b_mux_sel_dec_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17311.13-17311.26" */
wire [2:0] imm_b_mux_sel_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17286.13-17286.18" */
wire [31:0] imm_b_t0;
/* src = "generated/sv2v_out.v:17281.14-17281.24" */
wire [31:0] imm_b_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17281.14-17281.24" */
wire [31:0] imm_b_type_t0;
/* src = "generated/sv2v_out.v:17279.14-17279.24" */
wire [31:0] imm_i_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17279.14-17279.24" */
wire [31:0] imm_i_type_t0;
/* src = "generated/sv2v_out.v:17283.14-17283.24" */
wire [31:0] imm_j_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17283.14-17283.24" */
wire [31:0] imm_j_type_t0;
/* src = "generated/sv2v_out.v:17280.14-17280.24" */
wire [31:0] imm_s_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17280.14-17280.24" */
wire [31:0] imm_s_type_t0;
/* src = "generated/sv2v_out.v:17282.14-17282.24" */
wire [31:0] imm_u_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17282.14-17282.24" */
wire [31:0] imm_u_type_t0;
/* src = "generated/sv2v_out.v:17136.13-17136.29" */
input instr_bp_taken_i;
wire instr_bp_taken_i;
/* cellift = 32'd1 */
input instr_bp_taken_i_t0;
wire instr_bp_taken_i_t0;
/* src = "generated/sv2v_out.v:17141.13-17141.25" */
input instr_exec_i;
wire instr_exec_i;
/* cellift = 32'd1 */
input instr_exec_i_t0;
wire instr_exec_i_t0;
/* src = "generated/sv2v_out.v:17266.7-17266.22" */
wire instr_executing;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17266.7-17266.22" */
wire instr_executing_t0;
/* src = "generated/sv2v_out.v:17151.13-17151.30" */
input instr_fetch_err_i;
wire instr_fetch_err_i;
/* cellift = 32'd1 */
input instr_fetch_err_i_t0;
wire instr_fetch_err_i_t0;
/* src = "generated/sv2v_out.v:17152.13-17152.36" */
input instr_fetch_err_plus2_i;
wire instr_fetch_err_plus2_i;
/* cellift = 32'd1 */
input instr_fetch_err_plus2_i_t0;
wire instr_fetch_err_plus2_i_t0;
/* src = "generated/sv2v_out.v:17138.14-17138.36" */
output instr_first_cycle_id_o;
wire instr_first_cycle_id_o;
/* cellift = 32'd1 */
output instr_first_cycle_id_o_t0;
wire instr_first_cycle_id_o_t0;
/* src = "generated/sv2v_out.v:17241.14-17241.29" */
output instr_id_done_o;
wire instr_id_done_o;
/* cellift = 32'd1 */
output instr_id_done_o_t0;
wire instr_id_done_o_t0;
/* src = "generated/sv2v_out.v:17135.13-17135.34" */
input instr_is_compressed_i;
wire instr_is_compressed_i;
/* cellift = 32'd1 */
input instr_is_compressed_i_t0;
wire instr_is_compressed_i_t0;
/* src = "generated/sv2v_out.v:17231.14-17231.35" */
output instr_perf_count_id_o;
wire instr_perf_count_id_o;
/* cellift = 32'd1 */
output instr_perf_count_id_o_t0;
wire instr_perf_count_id_o_t0;
/* src = "generated/sv2v_out.v:17133.20-17133.37" */
input [31:0] instr_rdata_alu_i;
wire [31:0] instr_rdata_alu_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_alu_i_t0;
wire [31:0] instr_rdata_alu_i_t0;
/* src = "generated/sv2v_out.v:17134.20-17134.35" */
input [15:0] instr_rdata_c_i;
wire [15:0] instr_rdata_c_i;
/* cellift = 32'd1 */
input [15:0] instr_rdata_c_i_t0;
wire [15:0] instr_rdata_c_i_t0;
/* src = "generated/sv2v_out.v:17132.20-17132.33" */
input [31:0] instr_rdata_i;
wire [31:0] instr_rdata_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_i_t0;
wire [31:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:17137.14-17137.25" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:17230.20-17230.35" */
output [1:0] instr_type_wb_o;
wire [1:0] instr_type_wb_o;
/* cellift = 32'd1 */
output [1:0] instr_type_wb_o_t0;
wire [1:0] instr_type_wb_o_t0;
/* src = "generated/sv2v_out.v:17139.14-17139.33" */
output instr_valid_clear_o;
wire instr_valid_clear_o;
/* cellift = 32'd1 */
output instr_valid_clear_o_t0;
wire instr_valid_clear_o_t0;
/* src = "generated/sv2v_out.v:17131.13-17131.26" */
input instr_valid_i;
wire instr_valid_i;
/* cellift = 32'd1 */
input instr_valid_i_t0;
wire instr_valid_i_t0;
/* src = "generated/sv2v_out.v:17198.13-17198.21" */
input irq_nm_i;
wire irq_nm_i;
/* cellift = 32'd1 */
input irq_nm_i_t0;
wire irq_nm_i_t0;
/* src = "generated/sv2v_out.v:17196.13-17196.26" */
input irq_pending_i;
wire irq_pending_i;
/* cellift = 32'd1 */
input irq_pending_i_t0;
wire irq_pending_i_t0;
/* src = "generated/sv2v_out.v:17197.20-17197.26" */
input [17:0] irqs_i;
wire [17:0] irqs_i;
/* cellift = 32'd1 */
input [17:0] irqs_i_t0;
wire [17:0] irqs_i_t0;
/* src = "generated/sv2v_out.v:17260.7-17260.18" */
wire jump_in_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17260.7-17260.18" */
wire jump_in_dec_t0;
/* src = "generated/sv2v_out.v:17262.7-17262.15" */
wire jump_set;
/* src = "generated/sv2v_out.v:17261.7-17261.19" */
wire jump_set_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17261.7-17261.19" */
wire jump_set_dec_t0;
/* src = "generated/sv2v_out.v:17263.6-17263.18" */
wire jump_set_raw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17263.6-17263.18" */
wire jump_set_raw_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17262.7-17262.15" */
wire jump_set_t0;
/* src = "generated/sv2v_out.v:17193.13-17193.32" */
input lsu_addr_incr_req_i;
wire lsu_addr_incr_req_i;
/* cellift = 32'd1 */
input lsu_addr_incr_req_i_t0;
wire lsu_addr_incr_req_i_t0;
/* src = "generated/sv2v_out.v:17194.20-17194.35" */
input [31:0] lsu_addr_last_i;
wire [31:0] lsu_addr_last_i;
/* cellift = 32'd1 */
input [31:0] lsu_addr_last_i_t0;
wire [31:0] lsu_addr_last_i_t0;
/* src = "generated/sv2v_out.v:17200.13-17200.27" */
input lsu_load_err_i;
wire lsu_load_err_i;
/* cellift = 32'd1 */
input lsu_load_err_i_t0;
wire lsu_load_err_i_t0;
/* src = "generated/sv2v_out.v:17201.13-17201.37" */
input lsu_load_resp_intg_err_i;
wire lsu_load_resp_intg_err_i;
/* cellift = 32'd1 */
input lsu_load_resp_intg_err_i_t0;
wire lsu_load_resp_intg_err_i_t0;
/* src = "generated/sv2v_out.v:17324.7-17324.18" */
wire lsu_req_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17324.7-17324.18" */
wire lsu_req_dec_t0;
/* src = "generated/sv2v_out.v:17192.13-17192.27" */
input lsu_req_done_i;
wire lsu_req_done_i;
/* cellift = 32'd1 */
input lsu_req_done_i_t0;
wire lsu_req_done_i_t0;
/* src = "generated/sv2v_out.v:17187.14-17187.23" */
output lsu_req_o;
wire lsu_req_o;
/* cellift = 32'd1 */
output lsu_req_o_t0;
wire lsu_req_o_t0;
/* src = "generated/sv2v_out.v:17155.13-17155.29" */
input lsu_resp_valid_i;
wire lsu_resp_valid_i;
/* cellift = 32'd1 */
input lsu_resp_valid_i_t0;
wire lsu_resp_valid_i_t0;
/* src = "generated/sv2v_out.v:17190.14-17190.28" */
output lsu_sign_ext_o;
wire lsu_sign_ext_o;
/* cellift = 32'd1 */
output lsu_sign_ext_o_t0;
wire lsu_sign_ext_o_t0;
/* src = "generated/sv2v_out.v:17202.13-17202.28" */
input lsu_store_err_i;
wire lsu_store_err_i;
/* cellift = 32'd1 */
input lsu_store_err_i_t0;
wire lsu_store_err_i_t0;
/* src = "generated/sv2v_out.v:17203.13-17203.38" */
input lsu_store_resp_intg_err_i;
wire lsu_store_resp_intg_err_i;
/* cellift = 32'd1 */
input lsu_store_resp_intg_err_i_t0;
wire lsu_store_resp_intg_err_i_t0;
/* src = "generated/sv2v_out.v:17189.20-17189.30" */
output [1:0] lsu_type_o;
wire [1:0] lsu_type_o;
/* cellift = 32'd1 */
output [1:0] lsu_type_o_t0;
wire [1:0] lsu_type_o_t0;
/* src = "generated/sv2v_out.v:17191.21-17191.32" */
output [31:0] lsu_wdata_o;
wire [31:0] lsu_wdata_o;
/* cellift = 32'd1 */
output [31:0] lsu_wdata_o_t0;
wire [31:0] lsu_wdata_o_t0;
/* src = "generated/sv2v_out.v:17188.14-17188.22" */
output lsu_we_o;
wire lsu_we_o;
/* cellift = 32'd1 */
output lsu_we_o_t0;
wire lsu_we_o_t0;
/* src = "generated/sv2v_out.v:17278.7-17278.24" */
wire mem_resp_intg_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17278.7-17278.24" */
wire mem_resp_intg_err_t0;
/* src = "generated/sv2v_out.v:17246.7-17246.20" */
wire mret_insn_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17246.7-17246.20" */
wire mret_insn_dec_t0;
/* src = "generated/sv2v_out.v:17314.7-17314.18" */
wire mult_en_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17314.7-17314.18" */
wire mult_en_dec_t0;
/* src = "generated/sv2v_out.v:17164.14-17164.26" */
output mult_en_ex_o;
wire mult_en_ex_o;
/* cellift = 32'd1 */
output mult_en_ex_o_t0;
wire mult_en_ex_o_t0;
/* src = "generated/sv2v_out.v:17166.14-17166.27" */
output mult_sel_ex_o;
wire mult_sel_ex_o;
/* cellift = 32'd1 */
output mult_sel_ex_o_t0;
wire mult_sel_ex_o_t0;
/* src = "generated/sv2v_out.v:17317.7-17317.21" */
wire multdiv_en_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17317.7-17317.21" */
wire multdiv_en_dec_t0;
/* src = "generated/sv2v_out.v:17170.21-17170.43" */
output [31:0] multdiv_operand_a_ex_o;
wire [31:0] multdiv_operand_a_ex_o;
/* cellift = 32'd1 */
output [31:0] multdiv_operand_a_ex_o_t0;
wire [31:0] multdiv_operand_a_ex_o_t0;
/* src = "generated/sv2v_out.v:17171.21-17171.43" */
output [31:0] multdiv_operand_b_ex_o;
wire [31:0] multdiv_operand_b_ex_o;
/* cellift = 32'd1 */
output [31:0] multdiv_operand_b_ex_o_t0;
wire [31:0] multdiv_operand_b_ex_o_t0;
/* src = "generated/sv2v_out.v:17168.20-17168.41" */
output [1:0] multdiv_operator_ex_o;
wire [1:0] multdiv_operator_ex_o;
/* cellift = 32'd1 */
output [1:0] multdiv_operator_ex_o_t0;
wire [1:0] multdiv_operator_ex_o_t0;
/* src = "generated/sv2v_out.v:17172.14-17172.32" */
output multdiv_ready_id_o;
wire multdiv_ready_id_o;
/* cellift = 32'd1 */
output multdiv_ready_id_o_t0;
wire multdiv_ready_id_o_t0;
/* src = "generated/sv2v_out.v:17169.20-17169.44" */
output [1:0] multdiv_signed_mode_ex_o;
wire [1:0] multdiv_signed_mode_ex_o;
/* cellift = 32'd1 */
output [1:0] multdiv_signed_mode_ex_o_t0;
wire [1:0] multdiv_signed_mode_ex_o_t0;
/* src = "generated/sv2v_out.v:17277.7-17277.22" */
wire multicycle_done;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17277.7-17277.22" */
wire multicycle_done_t0;
/* src = "generated/sv2v_out.v:17199.14-17199.24" */
output nmi_mode_o;
wire nmi_mode_o;
/* cellift = 32'd1 */
output nmi_mode_o_t0;
wire nmi_mode_o_t0;
/* src = "generated/sv2v_out.v:17147.21-17147.37" */
output [31:0] nt_branch_addr_o;
wire [31:0] nt_branch_addr_o;
/* cellift = 32'd1 */
output [31:0] nt_branch_addr_o_t0;
wire [31:0] nt_branch_addr_o_t0;
/* src = "generated/sv2v_out.v:17146.14-17146.36" */
output nt_branch_mispredict_o;
wire nt_branch_mispredict_o;
/* cellift = 32'd1 */
output nt_branch_mispredict_o_t0;
wire nt_branch_mispredict_o_t0;
/* src = "generated/sv2v_out.v:17233.13-17233.34" */
input outstanding_load_wb_i;
wire outstanding_load_wb_i;
/* cellift = 32'd1 */
input outstanding_load_wb_i_t0;
wire outstanding_load_wb_i_t0;
/* src = "generated/sv2v_out.v:17234.13-17234.35" */
input outstanding_store_wb_i;
wire outstanding_store_wb_i;
/* cellift = 32'd1 */
input outstanding_store_wb_i_t0;
wire outstanding_store_wb_i_t0;
/* src = "generated/sv2v_out.v:17153.20-17153.27" */
input [31:0] pc_id_i;
wire [31:0] pc_id_i;
/* cellift = 32'd1 */
input [31:0] pc_id_i_t0;
wire [31:0] pc_id_i_t0;
/* src = "generated/sv2v_out.v:17145.20-17145.28" */
output [2:0] pc_mux_o;
wire [2:0] pc_mux_o;
/* cellift = 32'd1 */
output [2:0] pc_mux_o_t0;
wire [2:0] pc_mux_o_t0;
/* src = "generated/sv2v_out.v:17144.14-17144.22" */
output pc_set_o;
wire pc_set_o;
/* cellift = 32'd1 */
output pc_set_o_t0;
wire pc_set_o_t0;
/* src = "generated/sv2v_out.v:17236.13-17236.26" */
output perf_branch_o;
wire perf_branch_o;
/* cellift = 32'd1 */
output perf_branch_o_t0;
wire perf_branch_o_t0;
/* src = "generated/sv2v_out.v:17240.14-17240.29" */
output perf_div_wait_o;
wire perf_div_wait_o;
/* cellift = 32'd1 */
output perf_div_wait_o_t0;
wire perf_div_wait_o_t0;
/* src = "generated/sv2v_out.v:17238.14-17238.31" */
output perf_dside_wait_o;
wire perf_dside_wait_o;
/* cellift = 32'd1 */
output perf_dside_wait_o_t0;
wire perf_dside_wait_o_t0;
/* src = "generated/sv2v_out.v:17235.14-17235.25" */
output perf_jump_o;
wire perf_jump_o;
/* cellift = 32'd1 */
output perf_jump_o_t0;
wire perf_jump_o_t0;
/* src = "generated/sv2v_out.v:17239.14-17239.29" */
output perf_mul_wait_o;
wire perf_mul_wait_o;
/* cellift = 32'd1 */
output perf_mul_wait_o_t0;
wire perf_mul_wait_o_t0;
/* src = "generated/sv2v_out.v:17237.14-17237.28" */
output perf_tbranch_o;
wire perf_tbranch_o;
/* cellift = 32'd1 */
output perf_tbranch_o_t0;
wire perf_tbranch_o_t0;
/* src = "generated/sv2v_out.v:17183.19-17183.30" */
input [1:0] priv_mode_i;
wire [1:0] priv_mode_i;
/* cellift = 32'd1 */
input [1:0] priv_mode_i_t0;
wire [1:0] priv_mode_i_t0;
/* src = "generated/sv2v_out.v:17232.13-17232.23" */
input ready_wb_i;
wire ready_wb_i;
/* cellift = 32'd1 */
input ready_wb_i_t0;
wire ready_wb_i_t0;
/* src = "generated/sv2v_out.v:17213.20-17213.31" */
input [31:0] result_ex_i;
wire [31:0] result_ex_i;
/* cellift = 32'd1 */
input [31:0] result_ex_i_t0;
wire [31:0] result_ex_i_t0;
/* src = "generated/sv2v_out.v:17215.20-17215.32" */
output [4:0] rf_raddr_a_o;
wire [4:0] rf_raddr_a_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_a_o_t0;
wire [4:0] rf_raddr_a_o_t0;
/* src = "generated/sv2v_out.v:17217.20-17217.32" */
output [4:0] rf_raddr_b_o;
wire [4:0] rf_raddr_b_o;
/* cellift = 32'd1 */
output [4:0] rf_raddr_b_o_t0;
wire [4:0] rf_raddr_b_o_t0;
/* src = "generated/sv2v_out.v:17224.14-17224.32" */
output rf_rd_a_wb_match_o;
wire rf_rd_a_wb_match_o;
/* cellift = 32'd1 */
output rf_rd_a_wb_match_o_t0;
wire rf_rd_a_wb_match_o_t0;
/* src = "generated/sv2v_out.v:17225.14-17225.32" */
output rf_rd_b_wb_match_o;
wire rf_rd_b_wb_match_o;
/* cellift = 32'd1 */
output rf_rd_b_wb_match_o_t0;
wire rf_rd_b_wb_match_o_t0;
/* src = "generated/sv2v_out.v:17216.20-17216.32" */
input [31:0] rf_rdata_a_i;
wire [31:0] rf_rdata_a_i;
/* cellift = 32'd1 */
input [31:0] rf_rdata_a_i_t0;
wire [31:0] rf_rdata_a_i_t0;
/* src = "generated/sv2v_out.v:17218.20-17218.32" */
input [31:0] rf_rdata_b_i;
wire [31:0] rf_rdata_b_i;
/* cellift = 32'd1 */
input [31:0] rf_rdata_b_i_t0;
wire [31:0] rf_rdata_b_i_t0;
/* src = "generated/sv2v_out.v:17292.7-17292.19" */
wire rf_ren_a_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17292.7-17292.19" */
wire rf_ren_a_dec_t0;
/* src = "generated/sv2v_out.v:17219.14-17219.24" */
output rf_ren_a_o;
wire rf_ren_a_o;
/* cellift = 32'd1 */
output rf_ren_a_o_t0;
wire rf_ren_a_o_t0;
/* src = "generated/sv2v_out.v:17293.7-17293.19" */
wire rf_ren_b_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17293.7-17293.19" */
wire rf_ren_b_dec_t0;
/* src = "generated/sv2v_out.v:17220.14-17220.24" */
output rf_ren_b_o;
wire rf_ren_b_o;
/* cellift = 32'd1 */
output rf_ren_b_o_t0;
wire rf_ren_b_o_t0;
/* src = "generated/sv2v_out.v:17221.20-17221.33" */
output [4:0] rf_waddr_id_o;
wire [4:0] rf_waddr_id_o;
/* cellift = 32'd1 */
output [4:0] rf_waddr_id_o_t0;
wire [4:0] rf_waddr_id_o_t0;
/* src = "generated/sv2v_out.v:17226.19-17226.32" */
input [4:0] rf_waddr_wb_i;
wire [4:0] rf_waddr_wb_i;
/* cellift = 32'd1 */
input [4:0] rf_waddr_wb_i_t0;
wire [4:0] rf_waddr_wb_i_t0;
/* src = "generated/sv2v_out.v:17227.20-17227.37" */
input [31:0] rf_wdata_fwd_wb_i;
wire [31:0] rf_wdata_fwd_wb_i;
/* cellift = 32'd1 */
input [31:0] rf_wdata_fwd_wb_i_t0;
wire [31:0] rf_wdata_fwd_wb_i_t0;
/* src = "generated/sv2v_out.v:17222.20-17222.33" */
output [31:0] rf_wdata_id_o;
wire [31:0] rf_wdata_id_o;
/* cellift = 32'd1 */
output [31:0] rf_wdata_id_o_t0;
wire [31:0] rf_wdata_id_o_t0;
/* src = "generated/sv2v_out.v:17287.7-17287.19" */
wire rf_wdata_sel;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17287.7-17287.19" */
wire rf_wdata_sel_t0;
/* src = "generated/sv2v_out.v:17288.7-17288.16" */
wire rf_we_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17288.7-17288.16" */
wire rf_we_dec_t0;
/* src = "generated/sv2v_out.v:17223.14-17223.24" */
output rf_we_id_o;
wire rf_we_id_o;
/* cellift = 32'd1 */
output rf_we_id_o_t0;
wire rf_we_id_o_t0;
/* src = "generated/sv2v_out.v:17289.6-17289.15" */
wire rf_we_raw;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17289.6-17289.15" */
wire rf_we_raw_t0;
/* src = "generated/sv2v_out.v:17228.13-17228.26" */
input rf_write_wb_i;
wire rf_write_wb_i;
/* cellift = 32'd1 */
input rf_write_wb_i_t0;
wire rf_write_wb_i_t0;
/* src = "generated/sv2v_out.v:17128.13-17128.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:17306.6-17306.15" */
wire stall_alu;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17306.6-17306.15" */
wire stall_alu_t0;
/* src = "generated/sv2v_out.v:17272.6-17272.18" */
wire stall_branch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17272.6-17272.18" */
wire stall_branch_t0;
/* src = "generated/sv2v_out.v:17274.7-17274.15" */
wire stall_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17274.7-17274.15" */
wire stall_id_t0;
/* src = "generated/sv2v_out.v:17273.6-17273.16" */
wire stall_jump;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17273.6-17273.16" */
wire stall_jump_t0;
/* src = "generated/sv2v_out.v:17270.7-17270.16" */
wire stall_mem;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17270.7-17270.16" */
wire stall_mem_t0;
/* src = "generated/sv2v_out.v:17271.6-17271.19" */
wire stall_multdiv;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17271.6-17271.19" */
wire stall_multdiv_t0;
/* src = "generated/sv2v_out.v:17212.13-17212.28" */
input trigger_match_i;
wire trigger_match_i;
/* cellift = 32'd1 */
input trigger_match_i_t0;
wire trigger_match_i_t0;
/* src = "generated/sv2v_out.v:17249.7-17249.19" */
wire wfi_insn_dec;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17249.7-17249.19" */
wire wfi_insn_dec_t0;
/* src = "generated/sv2v_out.v:17284.14-17284.27" */
wire [31:0] zimm_rs1_type;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:17284.14-17284.27" */
wire [31:0] zimm_rs1_type_t0;
assign rf_ren_a_o = _0053_ & /* src = "generated/sv2v_out.v:17294.20-17294.91" */ rf_ren_a_dec;
assign _0053_ = _0051_ & /* src = "generated/sv2v_out.v:17295.21-17295.75" */ _0786_;
assign rf_ren_b_o = _0053_ & /* src = "generated/sv2v_out.v:17295.20-17295.91" */ rf_ren_b_dec;
assign _0055_ = rf_we_raw & /* src = "generated/sv2v_out.v:17409.23-17409.50" */ instr_executing;
assign rf_we_id_o = _0055_ & /* src = "generated/sv2v_out.v:17409.22-17409.73" */ _0159_;
assign illegal_dret_insn = dret_insn_dec & /* src = "generated/sv2v_out.v:17484.29-17484.58" */ _0787_;
assign _0057_ = csr_mstatus_tw_i & /* src = "generated/sv2v_out.v:17485.73-17485.104" */ wfi_insn_dec;
assign illegal_umode_insn = _0783_ & /* src = "generated/sv2v_out.v:17485.30-17485.106" */ _0794_;
assign illegal_insn_o = instr_valid_i & /* src = "generated/sv2v_out.v:17486.26-17486.126" */ _0800_;
assign _0059_ = instr_first_cycle_id_o & /* src = "generated/sv2v_out.v:17560.38-17560.68" */ lsu_req_dec;
assign _0061_ = csr_access_o & /* src = "generated/sv2v_out.v:17568.24-17568.54" */ instr_executing;
assign csr_op_en_o = _0061_ & /* src = "generated/sv2v_out.v:17568.23-17568.73" */ en_wb_o;
assign branch_jump_set_done_d = _0804_ & /* src = "generated/sv2v_out.v:17592.34-17592.115" */ _0788_;
assign jump_set = jump_set_raw & /* src = "generated/sv2v_out.v:17598.20-17598.58" */ _0165_;
assign branch_set = branch_set_raw & /* src = "generated/sv2v_out.v:17599.22-17599.62" */ _0165_;
assign _0063_ = rf_we_dec & /* src = "generated/sv2v_out.v:17676.19-17676.41" */ ex_valid_i;
assign _0065_ = multicycle_done & /* src = "generated/sv2v_out.v:17677.10-17677.38" */ ready_wb_i;
assign _0066_ = _0789_ & /* src = "generated/sv2v_out.v:17690.23-17690.44" */ _0790_;
assign en_wb_o = _0066_ & /* src = "generated/sv2v_out.v:17690.22-17690.63" */ instr_executing;
assign instr_first_cycle_id_o = instr_valid_i & /* src = "generated/sv2v_out.v:17691.29-17691.63" */ _0119_;
assign _0068_ = lsu_req_dec & /* src = "generated/sv2v_out.v:17725.40-17725.93" */ _0812_;
assign stall_mem = instr_valid_i & /* src = "generated/sv2v_out.v:17725.23-17725.94" */ _0068_;
assign _0051_ = instr_valid_i & /* src = "generated/sv2v_out.v:17727.35-17727.69" */ _0785_;
assign instr_executing = _0051_ & /* src = "generated/sv2v_out.v:17727.34-17727.87" */ controller_run;
assign _0070_ = instr_executing & /* src = "generated/sv2v_out.v:17751.32-17751.61" */ lsu_req_dec;
assign perf_dside_wait_o = _0070_ & /* src = "generated/sv2v_out.v:17751.31-17751.82" */ _0791_;
assign _0072_ = _0792_ & /* src = "generated/sv2v_out.v:17755.36-17755.64" */ _0793_;
assign _0074_ = _0072_ & /* src = "generated/sv2v_out.v:17755.35-17755.85" */ _0145_;
assign _0076_ = _0074_ & /* src = "generated/sv2v_out.v:17755.34-17755.108" */ _0159_;
assign instr_perf_count_id_o = _0076_ & /* src = "generated/sv2v_out.v:17755.33-17755.130" */ _0785_;
assign perf_mul_wait_o = stall_multdiv & /* src = "generated/sv2v_out.v:17757.27-17757.54" */ mult_en_dec;
assign perf_div_wait_o = stall_multdiv & /* src = "generated/sv2v_out.v:17758.27-17758.53" */ div_en_dec;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME \g_sec_branch_taken.branch_taken_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_sec_branch_taken.branch_taken_q_t0  <= 1'h0;
else \g_sec_branch_taken.branch_taken_q_t0  <= branch_decision_i_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME branch_set_raw_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_set_raw_t0 <= 1'h0;
else branch_set_raw_t0 <= branch_set_raw_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME branch_jump_set_done_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_jump_set_done_q_t0 <= 1'h0;
else branch_jump_set_done_q_t0 <= branch_jump_set_done_d_t0;
assign _0078_ = ~ imd_val_we_ex_i[1];
assign _0080_ = ~ imd_val_we_ex_i[0];
assign _0666_ = imd_val_d_ex_i[33:0] ^ imd_val_q_ex_o[33:0];
assign _0667_ = id_fsm_d ^ id_fsm_q;
assign _0668_ = imd_val_d_ex_i[67:34] ^ imd_val_q_ex_o[67:34];
assign _0560_ = imd_val_d_ex_i_t0[33:0] | imd_val_q_ex_o_t0[33:0];
assign _0564_ = id_fsm_d_t0 | id_fsm_q_t0;
assign _0568_ = imd_val_d_ex_i_t0[67:34] | imd_val_q_ex_o_t0[67:34];
assign _0561_ = _0666_ | _0560_;
assign _0565_ = _0667_ | _0564_;
assign _0569_ = _0668_ | _0568_;
assign _0270_ = { imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1], imd_val_we_ex_i[1] } & imd_val_d_ex_i_t0[33:0];
assign _0273_ = instr_executing & id_fsm_d_t0;
assign _0276_ = { imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0], imd_val_we_ex_i[0] } & imd_val_d_ex_i_t0[67:34];
assign _0271_ = { _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_, _0078_ } & imd_val_q_ex_o_t0[33:0];
assign _0274_ = _0079_ & id_fsm_q_t0;
assign _0277_ = { _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_, _0080_ } & imd_val_q_ex_o_t0[67:34];
assign _0272_ = _0561_ & { imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1], imd_val_we_ex_i_t0[1] };
assign _0275_ = _0565_ & instr_executing_t0;
assign _0278_ = _0569_ & { imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0], imd_val_we_ex_i_t0[0] };
assign _0562_ = _0270_ | _0271_;
assign _0566_ = _0273_ | _0274_;
assign _0570_ = _0276_ | _0277_;
assign _0563_ = _0562_ | _0272_;
assign _0567_ = _0566_ | _0275_;
assign _0571_ = _0570_ | _0278_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME imd_val_q_ex_o_t0[33:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) imd_val_q_ex_o_t0[33:0] <= 34'h000000000;
else imd_val_q_ex_o_t0[33:0] <= _0563_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME id_fsm_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) id_fsm_q_t0 <= 1'h0;
else id_fsm_q_t0 <= _0567_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME imd_val_q_ex_o_t0[67:34] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) imd_val_q_ex_o_t0[67:34] <= 34'h000000000;
else imd_val_q_ex_o_t0[67:34] <= _0571_;
assign _0174_ = _0054_ & rf_ren_a_dec;
assign _0177_ = _0052_ & _0786_;
assign _0180_ = _0054_ & rf_ren_b_dec;
assign _0183_ = rf_we_raw_t0 & instr_executing;
assign _0186_ = _0056_ & _0159_;
assign _0189_ = dret_insn_dec_t0 & _0787_;
assign _0192_ = csr_mstatus_tw_i_t0 & wfi_insn_dec;
assign _0195_ = _0784_ & _0794_;
assign _0198_ = instr_valid_i_t0 & _0800_;
assign _0201_ = instr_first_cycle_id_o_t0 & lsu_req_dec;
assign _0204_ = csr_access_o_t0 & instr_executing;
assign _0207_ = _0062_ & en_wb_o;
assign _0210_ = _0805_ & _0788_;
assign _0213_ = jump_set_raw_t0 & _0165_;
assign _0216_ = branch_set_raw_t0 & _0165_;
assign _0219_ = rf_we_dec_t0 & ex_valid_i;
assign _0222_ = multicycle_done_t0 & ready_wb_i;
assign _0225_ = stall_id_t0 & _0790_;
assign _0228_ = _0067_ & instr_executing;
assign _0231_ = instr_valid_i_t0 & _0119_;
assign _0234_ = lsu_req_dec_t0 & _0812_;
assign _0237_ = instr_valid_i_t0 & _0068_;
assign _0240_ = instr_valid_i_t0 & _0785_;
assign _0243_ = _0052_ & controller_run;
assign _0246_ = instr_executing_t0 & lsu_req_dec;
assign _0249_ = _0071_ & _0791_;
assign _0252_ = ebrk_insn_t0 & _0793_;
assign _0255_ = _0073_ & _0145_;
assign _0258_ = _0075_ & _0159_;
assign _0261_ = _0077_ & _0785_;
assign _0264_ = stall_multdiv_t0 & mult_en_dec;
assign _0267_ = stall_multdiv_t0 & div_en_dec;
assign _0175_ = rf_ren_a_dec_t0 & _0053_;
assign _0178_ = illegal_insn_o_t0 & _0051_;
assign _0181_ = rf_ren_b_dec_t0 & _0053_;
assign _0184_ = instr_executing_t0 & rf_we_raw;
assign _0187_ = illegal_csr_insn_i_t0 & _0055_;
assign _0190_ = debug_mode_o_t0 & dret_insn_dec;
assign _0193_ = wfi_insn_dec_t0 & csr_mstatus_tw_i;
assign _0196_ = _0795_ & _0783_;
assign _0199_ = _0801_ & instr_valid_i;
assign _0202_ = lsu_req_dec_t0 & instr_first_cycle_id_o;
assign _0205_ = instr_executing_t0 & csr_access_o;
assign _0208_ = en_wb_o_t0 & _0061_;
assign _0211_ = instr_valid_clear_o_t0 & _0804_;
assign _0214_ = branch_jump_set_done_q_t0 & jump_set_raw;
assign _0217_ = branch_jump_set_done_q_t0 & branch_set_raw;
assign _0220_ = ex_valid_i_t0 & rf_we_dec;
assign _0223_ = ready_wb_i_t0 & multicycle_done;
assign _0226_ = flush_id_t0 & _0789_;
assign _0229_ = instr_executing_t0 & _0066_;
assign _0232_ = id_fsm_q_t0 & instr_valid_i;
assign _0235_ = _0813_ & lsu_req_dec;
assign _0238_ = _0069_ & instr_valid_i;
assign _0241_ = instr_fetch_err_i_t0 & instr_valid_i;
assign _0244_ = controller_run_t0 & _0051_;
assign _0247_ = lsu_req_dec_t0 & instr_executing;
assign _0250_ = lsu_resp_valid_i_t0 & _0070_;
assign _0253_ = ecall_insn_dec_t0 & _0792_;
assign _0256_ = illegal_insn_dec_t0 & _0072_;
assign _0259_ = illegal_csr_insn_i_t0 & _0074_;
assign _0262_ = instr_fetch_err_i_t0 & _0076_;
assign _0265_ = mult_en_dec_t0 & stall_multdiv;
assign _0268_ = div_en_dec_t0 & stall_multdiv;
assign _0176_ = _0054_ & rf_ren_a_dec_t0;
assign _0179_ = _0052_ & illegal_insn_o_t0;
assign _0182_ = _0054_ & rf_ren_b_dec_t0;
assign _0185_ = rf_we_raw_t0 & instr_executing_t0;
assign _0188_ = _0056_ & illegal_csr_insn_i_t0;
assign _0191_ = dret_insn_dec_t0 & debug_mode_o_t0;
assign _0194_ = csr_mstatus_tw_i_t0 & wfi_insn_dec_t0;
assign _0197_ = _0784_ & _0795_;
assign _0200_ = instr_valid_i_t0 & _0801_;
assign _0203_ = instr_first_cycle_id_o_t0 & lsu_req_dec_t0;
assign _0206_ = csr_access_o_t0 & instr_executing_t0;
assign _0209_ = _0062_ & en_wb_o_t0;
assign _0212_ = _0805_ & instr_valid_clear_o_t0;
assign _0215_ = jump_set_raw_t0 & branch_jump_set_done_q_t0;
assign _0218_ = branch_set_raw_t0 & branch_jump_set_done_q_t0;
assign _0221_ = rf_we_dec_t0 & ex_valid_i_t0;
assign _0224_ = multicycle_done_t0 & ready_wb_i_t0;
assign _0227_ = stall_id_t0 & flush_id_t0;
assign _0230_ = _0067_ & instr_executing_t0;
assign _0233_ = instr_valid_i_t0 & id_fsm_q_t0;
assign _0236_ = lsu_req_dec_t0 & _0813_;
assign _0239_ = instr_valid_i_t0 & _0069_;
assign _0242_ = instr_valid_i_t0 & instr_fetch_err_i_t0;
assign _0245_ = _0052_ & controller_run_t0;
assign _0248_ = instr_executing_t0 & lsu_req_dec_t0;
assign _0251_ = _0071_ & lsu_resp_valid_i_t0;
assign _0254_ = ebrk_insn_t0 & ecall_insn_dec_t0;
assign _0257_ = _0073_ & illegal_insn_dec_t0;
assign _0260_ = _0075_ & illegal_csr_insn_i_t0;
assign _0263_ = _0077_ & instr_fetch_err_i_t0;
assign _0266_ = stall_multdiv_t0 & mult_en_dec_t0;
assign _0269_ = stall_multdiv_t0 & div_en_dec_t0;
assign _0528_ = _0174_ | _0175_;
assign _0529_ = _0177_ | _0178_;
assign _0530_ = _0180_ | _0181_;
assign _0531_ = _0183_ | _0184_;
assign _0532_ = _0186_ | _0187_;
assign _0533_ = _0189_ | _0190_;
assign _0534_ = _0192_ | _0193_;
assign _0535_ = _0195_ | _0196_;
assign _0536_ = _0198_ | _0199_;
assign _0537_ = _0201_ | _0202_;
assign _0538_ = _0204_ | _0205_;
assign _0539_ = _0207_ | _0208_;
assign _0540_ = _0210_ | _0211_;
assign _0541_ = _0213_ | _0214_;
assign _0542_ = _0216_ | _0217_;
assign _0543_ = _0219_ | _0220_;
assign _0544_ = _0222_ | _0223_;
assign _0545_ = _0225_ | _0226_;
assign _0546_ = _0228_ | _0229_;
assign _0547_ = _0231_ | _0232_;
assign _0548_ = _0234_ | _0235_;
assign _0549_ = _0237_ | _0238_;
assign _0550_ = _0240_ | _0241_;
assign _0551_ = _0243_ | _0244_;
assign _0552_ = _0246_ | _0247_;
assign _0553_ = _0249_ | _0250_;
assign _0554_ = _0252_ | _0253_;
assign _0555_ = _0255_ | _0256_;
assign _0556_ = _0258_ | _0259_;
assign _0557_ = _0261_ | _0262_;
assign _0558_ = _0264_ | _0265_;
assign _0559_ = _0267_ | _0268_;
assign rf_ren_a_o_t0 = _0528_ | _0176_;
assign _0054_ = _0529_ | _0179_;
assign rf_ren_b_o_t0 = _0530_ | _0182_;
assign _0056_ = _0531_ | _0185_;
assign rf_we_id_o_t0 = _0532_ | _0188_;
assign illegal_dret_insn_t0 = _0533_ | _0191_;
assign _0058_ = _0534_ | _0194_;
assign illegal_umode_insn_t0 = _0535_ | _0197_;
assign illegal_insn_o_t0 = _0536_ | _0200_;
assign _0060_ = _0537_ | _0203_;
assign _0062_ = _0538_ | _0206_;
assign csr_op_en_o_t0 = _0539_ | _0209_;
assign branch_jump_set_done_d_t0 = _0540_ | _0212_;
assign jump_set_t0 = _0541_ | _0215_;
assign branch_set_t0 = _0542_ | _0218_;
assign _0064_ = _0543_ | _0221_;
assign _0050_ = _0544_ | _0224_;
assign _0067_ = _0545_ | _0227_;
assign en_wb_o_t0 = _0546_ | _0230_;
assign instr_first_cycle_id_o_t0 = _0547_ | _0233_;
assign _0069_ = _0548_ | _0236_;
assign stall_mem_t0 = _0549_ | _0239_;
assign _0052_ = _0550_ | _0242_;
assign instr_executing_t0 = _0551_ | _0245_;
assign _0071_ = _0552_ | _0248_;
assign perf_dside_wait_o_t0 = _0553_ | _0251_;
assign _0073_ = _0554_ | _0254_;
assign _0075_ = _0555_ | _0257_;
assign _0077_ = _0556_ | _0260_;
assign instr_perf_count_id_o_t0 = _0557_ | _0263_;
assign perf_mul_wait_o_t0 = _0558_ | _0266_;
assign perf_div_wait_o_t0 = _0559_ | _0269_;
assign _0081_ = | csr_op_o_t0;
assign _0082_ = | instr_rdata_i_t0[31:20];
assign _0083_ = | instr_rdata_i_t0[31:25];
assign _0084_ = | priv_mode_i_t0;
assign _0086_ = | alu_op_a_mux_sel_t0;
assign _0087_ = ~ csr_op_o_t0;
assign _0088_ = ~ instr_rdata_i_t0[31:20];
assign _0089_ = ~ instr_rdata_i_t0[31:25];
assign _0090_ = ~ priv_mode_i_t0;
assign _0091_ = ~ imm_b_mux_sel_t0;
assign _0092_ = ~ alu_op_a_mux_sel_t0;
assign _0337_ = csr_op_o & _0087_;
assign _0338_ = instr_rdata_i[31:20] & _0088_;
assign _0339_ = instr_rdata_i[31:25] & _0089_;
assign _0370_ = priv_mode_i & _0090_;
assign _0413_ = imm_b_mux_sel & _0091_;
assign _0503_ = alu_op_a_mux_sel & _0092_;
assign _0710_ = _0337_ == { 1'h0, _0087_[0] };
assign _0711_ = _0337_ == { _0087_[1], 1'h0 };
assign _0712_ = _0338_ == { 2'h0, _0088_[9:8], 8'h00 };
assign _0713_ = _0338_ == { 2'h0, _0088_[9:8], 5'h00, _0088_[2], 2'h0 };
assign _0714_ = _0338_ == { 1'h0, _0088_[10:8], 1'h0, _0088_[6], 3'h0, _0088_[2:0] };
assign _0715_ = _0339_ == { 2'h0, _0089_[4:2], 1'h0, _0089_[0] };
assign _0716_ = _0338_ == { 1'h0, _0088_[10:7], 1'h0, _0088_[5:4], 4'h0 };
assign _0717_ = _0338_ == { 1'h0, _0088_[10:7], 1'h0, _0088_[5:4], 3'h0, _0088_[0] };
assign _0718_ = _0338_ == { 1'h0, _0088_[10:7], 1'h0, _0088_[5:4], 2'h0, _0088_[1], 1'h0 };
assign _0719_ = _0338_ == { 1'h0, _0088_[10:7], 1'h0, _0088_[5:4], 2'h0, _0088_[1:0] };
assign _0720_ = _0370_ == _0090_;
assign _0721_ = _0413_ == { _0091_[2], 1'h0, _0091_[0] };
assign _0722_ = _0413_ == { _0091_[2], 2'h0 };
assign _0723_ = _0413_ == { 1'h0, _0091_[1:0] };
assign _0724_ = _0413_ == { 1'h0, _0091_[1], 1'h0 };
assign _0725_ = _0413_ == { 2'h0, _0091_[0] };
assign _0726_ = _0503_ == _0092_;
assign _0727_ = _0503_ == { _0092_[1], 1'h0 };
assign _0728_ = _0503_ == { 1'h0, _0092_[0] };
assign _0744_ = _0710_ & _0081_;
assign _0746_ = _0711_ & _0081_;
assign _0748_ = _0712_ & _0082_;
assign _0750_ = _0713_ & _0082_;
assign _0752_ = _0714_ & _0082_;
assign _0754_ = _0715_ & _0083_;
assign _0756_ = _0716_ & _0082_;
assign _0758_ = _0717_ & _0082_;
assign _0760_ = _0718_ & _0082_;
assign _0762_ = _0719_ & _0082_;
assign _0784_ = _0720_ & _0084_;
assign _0815_ = _0721_ & _0085_;
assign _0817_ = _0722_ & _0085_;
assign _0819_ = _0723_ & _0085_;
assign _0821_ = _0724_ & _0085_;
assign _0823_ = _0725_ & _0085_;
assign _0853_ = _0726_ & _0086_;
assign _0855_ = _0727_ & _0086_;
assign _0857_ = _0728_ & _0086_;
/* src = "generated/sv2v_out.v:17400.4-17405.7" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME imd_val_q_ex_o[33:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) imd_val_q_ex_o[33:0] <= 34'h000000000;
else if (imd_val_we_ex_i[1]) imd_val_q_ex_o[33:0] <= imd_val_d_ex_i[33:0];
/* src = "generated/sv2v_out.v:17622.2-17627.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME id_fsm_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) id_fsm_q <= 1'h0;
else if (instr_executing) id_fsm_q <= id_fsm_d;
/* src = "generated/sv2v_out.v:17400.4-17405.7" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME imd_val_q_ex_o[67:34] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) imd_val_q_ex_o[67:34] <= 34'h000000000;
else if (imd_val_we_ex_i[0]) imd_val_q_ex_o[67:34] <= imd_val_d_ex_i[67:34];
assign _0340_ = csr_op_en_o_t0 & _0767_;
assign _0343_ = csr_op_en_o_t0 & _0781_;
assign _0341_ = _0768_ & csr_op_en_o;
assign _0344_ = _0782_ & csr_op_en_o;
assign _0342_ = csr_op_en_o_t0 & _0768_;
assign _0345_ = csr_op_en_o_t0 & _0782_;
assign _0609_ = _0340_ | _0341_;
assign _0610_ = _0343_ | _0344_;
assign _0764_ = _0609_ | _0342_;
assign _0766_ = _0610_ | _0345_;
assign _0093_ = | { _0819_, _0817_, _0815_ };
assign _0085_ = | imm_b_mux_sel_t0;
assign _0094_ = ~ { _0819_, _0817_, _0815_ };
assign _0285_ = { _0818_, _0816_, _0814_ } & _0094_;
assign _0095_ = ! _0285_;
assign _0096_ = ! _0337_;
assign _0097_ = ! _0413_;
assign _0173_ = _0095_ & _0093_;
assign _0782_ = _0096_ & _0081_;
assign _0825_ = _0097_ & _0085_;
assign _0098_ = ~ _0743_;
assign _0099_ = ~ _0747_;
assign _0100_ = ~ _0769_;
assign _0101_ = ~ _0771_;
assign _0102_ = ~ _0755_;
assign _0103_ = ~ _0774_;
assign _0104_ = ~ _0776_;
assign _0105_ = ~ data_ind_timing_i;
assign _0106_ = ~ _0745_;
assign _0107_ = ~ _0749_;
assign _0108_ = ~ _0751_;
assign _0109_ = ~ _0753_;
assign _0110_ = ~ _0757_;
assign _0111_ = ~ _0759_;
assign _0112_ = ~ _0761_;
assign _0113_ = ~ branch_decision_i;
assign _0346_ = _0744_ & _0106_;
assign _0349_ = _0748_ & _0107_;
assign _0352_ = _0770_ & _0108_;
assign _0355_ = _0772_ & _0109_;
assign _0358_ = _0756_ & _0110_;
assign _0361_ = _0775_ & _0111_;
assign _0364_ = _0777_ & _0112_;
assign _0367_ = data_ind_timing_i_t0 & _0113_;
assign _0347_ = _0746_ & _0098_;
assign _0350_ = _0750_ & _0099_;
assign _0353_ = _0752_ & _0100_;
assign _0356_ = _0754_ & _0101_;
assign _0359_ = _0758_ & _0102_;
assign _0362_ = _0760_ & _0103_;
assign _0365_ = _0762_ & _0104_;
assign _0368_ = branch_decision_i_t0 & _0105_;
assign _0348_ = _0744_ & _0746_;
assign _0351_ = _0748_ & _0750_;
assign _0354_ = _0770_ & _0752_;
assign _0357_ = _0772_ & _0754_;
assign _0360_ = _0756_ & _0758_;
assign _0363_ = _0775_ & _0760_;
assign _0366_ = _0777_ & _0762_;
assign _0369_ = data_ind_timing_i_t0 & branch_decision_i_t0;
assign _0611_ = _0346_ | _0347_;
assign _0612_ = _0349_ | _0350_;
assign _0613_ = _0352_ | _0353_;
assign _0614_ = _0355_ | _0356_;
assign _0615_ = _0358_ | _0359_;
assign _0616_ = _0361_ | _0362_;
assign _0617_ = _0364_ | _0365_;
assign _0618_ = _0367_ | _0368_;
assign _0768_ = _0611_ | _0348_;
assign _0770_ = _0612_ | _0351_;
assign _0772_ = _0613_ | _0354_;
assign _0003_ = _0614_ | _0357_;
assign _0775_ = _0615_ | _0360_;
assign _0777_ = _0616_ | _0363_;
assign _0037_ = _0617_ | _0366_;
assign _0780_ = _0618_ | _0369_;
assign _0114_ = ~ { _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_ };
assign _0115_ = ~ { _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_ };
assign _0116_ = ~ { _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_ };
assign _0117_ = ~ { _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_ };
assign _0118_ = ~ { _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_ };
assign _0119_ = ~ id_fsm_q;
assign _0120_ = ~ { rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel };
assign _0121_ = ~ { _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_ };
assign _0122_ = ~ { _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_ };
assign _0123_ = ~ { _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_ };
assign _0124_ = ~ _0065_;
assign _0125_ = ~ multdiv_en_dec;
assign _0126_ = ~ alu_multicycle_dec;
assign _0127_ = ~ jump_in_dec;
assign _0128_ = ~ branch_in_dec;
assign _0129_ = ~ lsu_req_dec;
assign _0079_ = ~ instr_executing;
assign _0130_ = ~ _0763_;
assign _0131_ = ~ { lsu_addr_incr_req_i, lsu_addr_incr_req_i };
assign _0132_ = ~ lsu_addr_incr_req_i;
assign _0133_ = ~ { lsu_addr_incr_req_i, lsu_addr_incr_req_i, lsu_addr_incr_req_i };
assign _0134_ = ~ { imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel, imm_a_mux_sel };
assign _0135_ = ~ { alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel };
assign _0574_ = { _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_ } | _0114_;
assign _0577_ = { _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_ } | _0115_;
assign _0580_ = { _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_ } | _0116_;
assign _0584_ = { _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_ } | _0117_;
assign _0587_ = { _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_ } | _0118_;
assign _0590_ = id_fsm_q_t0 | _0119_;
assign _0597_ = { rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0 } | _0120_;
assign _0600_ = { _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_ } | _0121_;
assign _0603_ = { _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_ } | _0122_;
assign _0606_ = { _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_ } | _0123_;
assign _0633_ = _0050_ | _0124_;
assign _0634_ = multdiv_en_dec_t0 | _0125_;
assign _0638_ = alu_multicycle_dec_t0 | _0126_;
assign _0639_ = jump_in_dec_t0 | _0127_;
assign _0641_ = branch_in_dec_t0 | _0128_;
assign _0645_ = lsu_req_dec_t0 | _0129_;
assign _0651_ = instr_executing_t0 | _0079_;
assign _0655_ = _0764_ | _0130_;
assign _0658_ = { lsu_addr_incr_req_i_t0, lsu_addr_incr_req_i_t0 } | _0131_;
assign _0659_ = lsu_addr_incr_req_i_t0 | _0132_;
assign _0660_ = { lsu_addr_incr_req_i_t0, lsu_addr_incr_req_i_t0, lsu_addr_incr_req_i_t0 } | _0133_;
assign _0661_ = { imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0 } | _0134_;
assign _0662_ = { alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0 } | _0135_;
assign _0575_ = { _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_ } | { _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_, _0816_ };
assign _0578_ = { _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_ } | { _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_, _0814_ };
assign _0581_ = { _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_ } | { _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_, _0820_ };
assign _0583_ = { _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_ } | { _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_, _0824_ };
assign _0585_ = { _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_ } | { _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_, _0524_ };
assign _0588_ = { _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_ } | { _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_, _0172_ };
assign _0591_ = id_fsm_q_t0 | id_fsm_q;
assign _0598_ = { rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0 } | { rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel, rf_wdata_sel };
assign _0601_ = { _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_ } | { _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_, _0852_ };
assign _0604_ = { _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_ } | { _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_, _0856_ };
assign _0607_ = { _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_ } | { _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_, _0526_ };
assign _0635_ = multdiv_en_dec_t0 | multdiv_en_dec;
assign _0637_ = ex_valid_i_t0 | ex_valid_i;
assign _0640_ = jump_in_dec_t0 | jump_in_dec;
assign _0642_ = branch_in_dec_t0 | branch_in_dec;
assign _0646_ = lsu_req_dec_t0 | lsu_req_dec;
assign _0652_ = instr_executing_t0 | instr_executing;
assign _0654_ = _0766_ | _0765_;
assign _0656_ = _0764_ | _0763_;
assign _0663_ = { alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0 } | { alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel, alu_op_b_mux_sel };
assign _0286_ = imm_u_type_t0 & _0574_;
assign _0289_ = _0730_ & _0577_;
assign _0292_ = imm_s_type_t0 & _0580_;
assign _0297_ = _0736_ & _0584_;
assign _0300_ = _0738_ & _0587_;
assign _0303_ = _0023_ & _0590_;
assign _0306_ = _0031_ & _0590_;
assign _0308_ = _0029_ & _0590_;
assign _0311_ = _0033_ & _0590_;
assign _0314_ = _0019_ & _0590_;
assign _0317_ = _0035_ & _0590_;
assign _0320_ = _0025_ & _0590_;
assign _0323_ = _0027_ & _0590_;
assign _0325_ = result_ex_i_t0 & _0597_;
assign _0328_ = pc_id_i_t0 & _0600_;
assign _0331_ = rf_rdata_a_i_t0 & _0603_;
assign _0334_ = _0742_ & _0606_;
assign _0414_ = jump_in_dec_t0 & _0633_;
assign _0416_ = branch_in_dec_t0 & _0633_;
assign _0418_ = multdiv_en_dec_t0 & _0633_;
assign _0420_ = rf_we_dec_t0 & _0634_;
assign _0424_ = alu_multicycle_dec_t0 & _0639_;
assign _0426_ = _0827_ & _0641_;
assign _0429_ = _0829_ & _0634_;
assign _0432_ = _0831_ & _0645_;
assign _0435_ = _0832_ & _0641_;
assign _0437_ = _0833_ & _0634_;
assign _0439_ = _0834_ & _0645_;
assign _0441_ = rf_we_dec_t0 & _0638_;
assign _0443_ = _0836_ & _0639_;
assign _0446_ = _0838_ & _0641_;
assign _0449_ = _0840_ & _0634_;
assign _0452_ = _0842_ & _0645_;
assign _0455_ = jump_in_dec_t0 & _0641_;
assign _0457_ = _0843_ & _0634_;
assign _0459_ = _0844_ & _0645_;
assign _0462_ = _0845_ & _0634_;
assign _0464_ = _0846_ & _0645_;
assign _0467_ = _0847_ & _0645_;
assign _0471_ = _0848_ & _0641_;
assign _0473_ = _0849_ & _0634_;
assign _0475_ = _0850_ & _0645_;
assign _0477_ = branch_in_dec_t0 & _0634_;
assign _0479_ = _0851_ & _0645_;
assign _0483_ = rf_we_dec_t0 & _0651_;
assign _0500_ = _0021_ & _0655_;
assign _0504_ = alu_op_a_mux_sel_dec_t0 & _0658_;
assign _0506_ = alu_op_b_mux_sel_dec_t0 & _0659_;
assign _0508_ = imm_b_mux_sel_dec_t0 & _0660_;
assign _0510_ = zimm_rs1_type_t0 & _0661_;
assign _0512_ = rf_rdata_b_i_t0 & _0662_;
assign _0521_ = ex_valid_i_t0 & _0645_;
assign _0287_ = imm_j_type_t0 & _0575_;
assign _0290_ = { 29'h00000000, instr_is_compressed_i_t0, instr_is_compressed_i_t0, 1'h0 } & _0578_;
assign _0293_ = imm_b_type_t0 & _0581_;
assign _0295_ = imm_i_type_t0 & _0583_;
assign _0298_ = _0734_ & _0585_;
assign _0301_ = _0732_ & _0588_;
assign _0304_ = _0050_ & _0591_;
assign _0309_ = _0046_ & _0591_;
assign _0312_ = _0043_ & _0591_;
assign _0315_ = _0041_ & _0591_;
assign _0318_ = _0048_ & _0591_;
assign _0326_ = csr_rdata_i_t0 & _0598_;
assign _0329_ = imm_a_t0 & _0601_;
assign _0332_ = lsu_addr_last_i_t0 & _0604_;
assign _0335_ = _0740_ & _0607_;
assign _0421_ = _0064_ & _0635_;
assign _0423_ = rf_we_dec_t0 & _0637_;
assign _0427_ = _0780_ & _0642_;
assign _0430_ = ex_valid_i_t0 & _0635_;
assign _0444_ = rf_we_dec_t0 & _0640_;
assign _0447_ = rf_we_dec_t0 & _0642_;
assign _0450_ = _0039_ & _0635_;
assign _0453_ = rf_we_dec_t0 & _0646_;
assign _0469_ = jump_set_dec_t0 & _0640_;
assign _0481_ = _0011_ & _0652_;
assign _0484_ = _0009_ & _0652_;
assign _0486_ = _0015_ & _0652_;
assign _0488_ = _0013_ & _0652_;
assign _0490_ = _0017_ & _0652_;
assign _0492_ = _0005_ & _0652_;
assign _0494_ = _0001_ & _0652_;
assign _0496_ = _0007_ & _0652_;
assign _0498_ = _0037_ & _0654_;
assign _0501_ = _0003_ & _0656_;
assign _0513_ = imm_b_t0 & _0663_;
assign _0515_ = _0060_ & _0652_;
assign _0517_ = mult_en_dec_t0 & _0652_;
assign _0519_ = div_en_dec_t0 & _0652_;
assign _0522_ = lsu_resp_valid_i_t0 & _0646_;
assign _0576_ = _0286_ | _0287_;
assign _0579_ = _0289_ | _0290_;
assign _0582_ = _0292_ | _0293_;
assign _0586_ = _0297_ | _0298_;
assign _0589_ = _0300_ | _0301_;
assign _0592_ = _0303_ | _0304_;
assign _0593_ = _0308_ | _0309_;
assign _0594_ = _0311_ | _0312_;
assign _0595_ = _0314_ | _0315_;
assign _0596_ = _0317_ | _0318_;
assign _0599_ = _0325_ | _0326_;
assign _0602_ = _0328_ | _0329_;
assign _0605_ = _0331_ | _0332_;
assign _0608_ = _0334_ | _0335_;
assign _0636_ = _0420_ | _0421_;
assign _0643_ = _0426_ | _0427_;
assign _0644_ = _0429_ | _0430_;
assign _0647_ = _0443_ | _0444_;
assign _0648_ = _0446_ | _0447_;
assign _0649_ = _0449_ | _0450_;
assign _0650_ = _0452_ | _0453_;
assign _0653_ = _0483_ | _0484_;
assign _0657_ = _0500_ | _0501_;
assign _0664_ = _0512_ | _0513_;
assign _0665_ = _0521_ | _0522_;
assign _0669_ = imm_u_type ^ imm_j_type;
assign _0670_ = _0729_ ^ _0858_;
assign _0671_ = imm_s_type ^ imm_b_type;
assign _0672_ = _0735_ ^ _0733_;
assign _0673_ = _0737_ ^ _0731_;
assign _0674_ = _0022_ ^ _0049_;
assign _0675_ = _0028_ ^ _0045_;
assign _0676_ = _0032_ ^ _0042_;
assign _0677_ = _0018_ ^ _0040_;
assign _0678_ = _0034_ ^ _0047_;
assign _0679_ = result_ex_i ^ csr_rdata_i;
assign _0680_ = pc_id_i ^ imm_a;
assign _0681_ = rf_rdata_a_i ^ lsu_addr_last_i;
assign _0682_ = _0741_ ^ _0739_;
assign _0683_ = rf_we_dec ^ _0063_;
assign _0684_ = _0826_ ^ _0859_;
assign _0685_ = _0828_ ^ _0044_;
assign _0690_ = _0835_ ^ rf_we_dec;
assign _0691_ = _0837_ ^ rf_we_dec;
assign _0692_ = _0839_ ^ _0038_;
assign _0693_ = _0841_ ^ rf_we_dec;
assign _0706_ = rf_we_dec ^ _0008_;
assign _0707_ = _0020_ ^ _0002_;
assign _0708_ = rf_rdata_b_i ^ imm_b;
assign _0709_ = ex_valid_i ^ lsu_resp_valid_i;
assign _0288_ = { _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_, _0817_ } & _0669_;
assign _0291_ = { _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_, _0815_ } & _0670_;
assign _0294_ = { _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_, _0821_ } & _0671_;
assign _0296_ = { _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_, _0825_ } & { imm_i_type[31:3], _0141_, imm_i_type[1:0] };
assign _0299_ = { _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_, _0525_ } & _0672_;
assign _0302_ = { _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_, _0173_ } & _0673_;
assign _0305_ = id_fsm_q_t0 & _0674_;
assign _0307_ = id_fsm_q_t0 & _0030_;
assign _0310_ = id_fsm_q_t0 & _0675_;
assign _0313_ = id_fsm_q_t0 & _0676_;
assign _0316_ = id_fsm_q_t0 & _0677_;
assign _0319_ = id_fsm_q_t0 & _0678_;
assign _0321_ = id_fsm_q_t0 & _0024_;
assign _0322_ = id_fsm_q_t0 & _0018_;
assign _0324_ = id_fsm_q_t0 & _0026_;
assign _0327_ = { rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0, rf_wdata_sel_t0 } & _0679_;
assign _0330_ = { _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_, _0853_ } & _0680_;
assign _0333_ = { _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_, _0857_ } & _0681_;
assign _0336_ = { _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_, _0527_ } & _0682_;
assign _0415_ = _0050_ & jump_in_dec;
assign _0417_ = _0050_ & branch_in_dec;
assign _0419_ = _0050_ & multdiv_en_dec;
assign _0422_ = multdiv_en_dec_t0 & _0683_;
assign _0425_ = jump_in_dec_t0 & _0136_;
assign _0428_ = branch_in_dec_t0 & _0684_;
assign _0431_ = multdiv_en_dec_t0 & _0685_;
assign _0433_ = lsu_req_dec_t0 & _0137_;
assign _0434_ = jump_in_dec_t0 & _0686_;
assign _0436_ = branch_in_dec_t0 & _0687_;
assign _0438_ = multdiv_en_dec_t0 & _0688_;
assign _0440_ = lsu_req_dec_t0 & _0689_;
assign _0442_ = alu_multicycle_dec_t0 & rf_we_dec;
assign _0445_ = jump_in_dec_t0 & _0690_;
assign _0448_ = branch_in_dec_t0 & _0691_;
assign _0451_ = multdiv_en_dec_t0 & _0692_;
assign _0454_ = lsu_req_dec_t0 & _0693_;
assign _0456_ = branch_in_dec_t0 & _0694_;
assign _0458_ = multdiv_en_dec_t0 & _0695_;
assign _0460_ = lsu_req_dec_t0 & _0696_;
assign _0461_ = branch_in_dec_t0 & _0697_;
assign _0463_ = multdiv_en_dec_t0 & _0698_;
assign _0465_ = lsu_req_dec_t0 & _0699_;
assign _0466_ = multdiv_en_dec_t0 & _0044_;
assign _0468_ = lsu_req_dec_t0 & _0700_;
assign _0470_ = jump_in_dec_t0 & jump_set_dec;
assign _0472_ = branch_in_dec_t0 & _0701_;
assign _0474_ = multdiv_en_dec_t0 & _0702_;
assign _0476_ = lsu_req_dec_t0 & _0703_;
assign _0478_ = multdiv_en_dec_t0 & _0704_;
assign _0480_ = lsu_req_dec_t0 & _0705_;
assign _0482_ = instr_executing_t0 & _0010_;
assign _0485_ = instr_executing_t0 & _0706_;
assign _0487_ = instr_executing_t0 & _0014_;
assign _0489_ = instr_executing_t0 & _0012_;
assign _0491_ = instr_executing_t0 & _0016_;
assign _0493_ = instr_executing_t0 & _0004_;
assign _0495_ = instr_executing_t0 & _0000_;
assign _0497_ = instr_executing_t0 & _0006_;
assign _0499_ = _0766_ & _0036_;
assign _0502_ = _0764_ & _0707_;
assign _0505_ = { lsu_addr_incr_req_i_t0, lsu_addr_incr_req_i_t0 } & { alu_op_a_mux_sel_dec[1], _0140_ };
assign _0507_ = lsu_addr_incr_req_i_t0 & _0138_;
assign _0509_ = { lsu_addr_incr_req_i_t0, lsu_addr_incr_req_i_t0, lsu_addr_incr_req_i_t0 } & { _0139_, imm_b_mux_sel_dec[0] };
assign _0511_ = { imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0, imm_a_mux_sel_t0 } & zimm_rs1_type;
assign _0514_ = { alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0, alu_op_b_mux_sel_t0 } & _0708_;
assign _0516_ = instr_executing_t0 & _0059_;
assign _0518_ = instr_executing_t0 & mult_en_dec;
assign _0520_ = instr_executing_t0 & div_en_dec;
assign _0523_ = lsu_req_dec_t0 & _0709_;
assign _0730_ = _0288_ | _0576_;
assign _0732_ = _0291_ | _0579_;
assign _0734_ = _0294_ | _0582_;
assign _0736_ = _0296_ | _0295_;
assign _0738_ = _0299_ | _0586_;
assign imm_b_t0 = _0302_ | _0589_;
assign id_fsm_d_t0 = _0305_ | _0592_;
assign _0011_ = _0307_ | _0306_;
assign _0009_ = _0310_ | _0593_;
assign _0015_ = _0313_ | _0594_;
assign _0013_ = _0316_ | _0595_;
assign _0017_ = _0319_ | _0596_;
assign _0005_ = _0321_ | _0320_;
assign _0001_ = _0322_ | _0314_;
assign _0007_ = _0324_ | _0323_;
assign rf_wdata_id_o_t0 = _0327_ | _0599_;
assign _0740_ = _0330_ | _0602_;
assign _0742_ = _0333_ | _0605_;
assign alu_operand_a_ex_o_t0 = _0336_ | _0608_;
assign _0043_ = _0415_ | _0414_;
assign _0041_ = _0417_ | _0416_;
assign _0048_ = _0419_ | _0418_;
assign _0046_ = _0422_ | _0636_;
assign _0039_ = _0220_ | _0423_;
assign _0827_ = _0425_ | _0424_;
assign _0829_ = _0428_ | _0643_;
assign _0831_ = _0431_ | _0644_;
assign _0023_ = _0433_ | _0432_;
assign _0832_ = _0434_ | _0424_;
assign _0833_ = _0436_ | _0435_;
assign _0834_ = _0438_ | _0437_;
assign _0031_ = _0440_ | _0439_;
assign _0836_ = _0442_ | _0441_;
assign _0838_ = _0445_ | _0647_;
assign _0840_ = _0448_ | _0648_;
assign _0842_ = _0451_ | _0649_;
assign _0029_ = _0454_ | _0650_;
assign _0843_ = _0456_ | _0455_;
assign _0844_ = _0458_ | _0457_;
assign _0033_ = _0460_ | _0459_;
assign _0845_ = _0461_ | _0427_;
assign _0846_ = _0463_ | _0462_;
assign _0019_ = _0465_ | _0464_;
assign _0847_ = _0466_ | _0430_;
assign _0035_ = _0468_ | _0467_;
assign _0848_ = _0470_ | _0469_;
assign _0849_ = _0472_ | _0471_;
assign _0850_ = _0474_ | _0473_;
assign _0025_ = _0476_ | _0475_;
assign _0851_ = _0478_ | _0477_;
assign _0027_ = _0480_ | _0479_;
assign stall_alu_t0 = _0482_ | _0481_;
assign rf_we_raw_t0 = _0485_ | _0653_;
assign stall_jump_t0 = _0487_ | _0486_;
assign stall_branch_t0 = _0489_ | _0488_;
assign stall_multdiv_t0 = _0491_ | _0490_;
assign jump_set_raw_t0 = _0493_ | _0492_;
assign branch_set_raw_d_t0 = _0495_ | _0494_;
assign perf_branch_o_t0 = _0497_ | _0496_;
assign _0021_ = _0499_ | _0498_;
assign csr_pipe_flush_t0 = _0502_ | _0657_;
assign alu_op_a_mux_sel_t0 = _0505_ | _0504_;
assign alu_op_b_mux_sel_t0 = _0507_ | _0506_;
assign imm_b_mux_sel_t0 = _0509_ | _0508_;
assign imm_a_t0 = _0511_ | _0510_;
assign alu_operand_b_ex_o_t0 = _0514_ | _0664_;
assign lsu_req_o_t0 = _0516_ | _0515_;
assign mult_en_ex_o_t0 = _0518_ | _0517_;
assign div_en_ex_o_t0 = _0520_ | _0519_;
assign multicycle_done_t0 = _0523_ | _0665_;
assign _0136_ = ~ _0686_;
assign _0137_ = ~ _0830_;
assign _0138_ = ~ alu_op_b_mux_sel_dec;
assign _0139_ = ~ imm_b_mux_sel_dec[2:1];
assign _0140_ = ~ alu_op_a_mux_sel_dec[0];
assign _0141_ = ~ imm_i_type[2];
assign _0142_ = ~ _0822_;
assign _0143_ = ~ _0854_;
assign _0144_ = ~ mret_insn_dec;
assign _0145_ = ~ illegal_insn_dec;
assign _0146_ = ~ _0796_;
assign _0147_ = ~ _0798_;
assign _0148_ = ~ lsu_load_resp_intg_err_i;
assign _0149_ = ~ mult_en_dec;
assign _0150_ = ~ branch_set_raw;
assign _0151_ = ~ _0802_;
assign _0152_ = ~ stall_mem;
assign _0153_ = ~ _0806_;
assign _0154_ = ~ _0808_;
assign _0155_ = ~ _0810_;
assign _0156_ = ~ _0820_;
assign _0157_ = ~ _0852_;
assign _0158_ = ~ _0057_;
assign _0159_ = ~ illegal_csr_insn_i;
assign _0160_ = ~ illegal_dret_insn;
assign _0161_ = ~ illegal_umode_insn;
assign _0162_ = ~ lsu_store_resp_intg_err_i;
assign _0163_ = ~ div_en_dec;
assign _0164_ = ~ jump_set_raw;
assign _0165_ = ~ branch_jump_set_done_q;
assign _0166_ = ~ \g_sec_branch_taken.branch_taken_q ;
assign _0167_ = ~ stall_multdiv;
assign _0168_ = ~ stall_jump;
assign _0169_ = ~ stall_branch;
assign _0170_ = ~ stall_alu;
assign _0171_ = ~ instr_first_cycle_id_o;
assign _0279_ = _0823_ & _0156_;
assign _0282_ = _0855_ & _0157_;
assign _0371_ = mret_insn_dec_t0 & _0158_;
assign _0374_ = illegal_insn_dec_t0 & _0159_;
assign _0377_ = _0797_ & _0160_;
assign _0380_ = _0799_ & _0161_;
assign _0383_ = lsu_load_resp_intg_err_i_t0 & _0162_;
assign _0386_ = mult_en_dec_t0 & _0163_;
assign _0389_ = branch_set_raw_t0 & _0164_;
assign _0392_ = _0803_ & _0165_;
assign _0395_ = data_ind_timing_i_t0 & _0166_;
assign _0398_ = stall_mem_t0 & _0167_;
assign _0401_ = _0807_ & _0168_;
assign _0404_ = _0809_ & _0169_;
assign _0407_ = _0811_ & _0170_;
assign _0410_ = lsu_resp_valid_i_t0 & _0171_;
assign _0280_ = _0821_ & _0142_;
assign _0283_ = _0853_ & _0143_;
assign _0372_ = _0058_ & _0144_;
assign _0375_ = illegal_csr_insn_i_t0 & _0145_;
assign _0378_ = illegal_dret_insn_t0 & _0146_;
assign _0381_ = illegal_umode_insn_t0 & _0147_;
assign _0384_ = lsu_store_resp_intg_err_i_t0 & _0148_;
assign _0387_ = div_en_dec_t0 & _0149_;
assign _0390_ = jump_set_raw_t0 & _0150_;
assign _0393_ = branch_jump_set_done_q_t0 & _0151_;
assign _0396_ = \g_sec_branch_taken.branch_taken_q_t0  & data_ind_timing_i;
assign _0399_ = stall_multdiv_t0 & _0152_;
assign _0402_ = stall_jump_t0 & _0153_;
assign _0405_ = stall_branch_t0 & _0154_;
assign _0408_ = stall_alu_t0 & _0155_;
assign _0411_ = instr_first_cycle_id_o_t0 & lsu_resp_valid_i;
assign _0281_ = _0823_ & _0821_;
assign _0284_ = _0855_ & _0853_;
assign _0373_ = mret_insn_dec_t0 & _0058_;
assign _0376_ = illegal_insn_dec_t0 & illegal_csr_insn_i_t0;
assign _0379_ = _0797_ & illegal_dret_insn_t0;
assign _0382_ = _0799_ & illegal_umode_insn_t0;
assign _0385_ = lsu_load_resp_intg_err_i_t0 & lsu_store_resp_intg_err_i_t0;
assign _0388_ = mult_en_dec_t0 & div_en_dec_t0;
assign _0391_ = branch_set_raw_t0 & jump_set_raw_t0;
assign _0394_ = _0803_ & branch_jump_set_done_q_t0;
assign _0397_ = data_ind_timing_i_t0 & \g_sec_branch_taken.branch_taken_q_t0 ;
assign _0400_ = stall_mem_t0 & stall_multdiv_t0;
assign _0403_ = _0807_ & stall_jump_t0;
assign _0406_ = _0809_ & stall_branch_t0;
assign _0409_ = _0811_ & stall_alu_t0;
assign _0412_ = lsu_resp_valid_i_t0 & instr_first_cycle_id_o_t0;
assign _0572_ = _0279_ | _0280_;
assign _0573_ = _0282_ | _0283_;
assign _0619_ = _0371_ | _0372_;
assign _0620_ = _0374_ | _0375_;
assign _0621_ = _0377_ | _0378_;
assign _0622_ = _0380_ | _0381_;
assign _0623_ = _0383_ | _0384_;
assign _0624_ = _0386_ | _0387_;
assign _0625_ = _0389_ | _0390_;
assign _0626_ = _0392_ | _0393_;
assign _0627_ = _0395_ | _0396_;
assign _0628_ = _0398_ | _0399_;
assign _0629_ = _0401_ | _0402_;
assign _0630_ = _0404_ | _0405_;
assign _0631_ = _0407_ | _0408_;
assign _0632_ = _0410_ | _0411_;
assign _0525_ = _0572_ | _0281_;
assign _0527_ = _0573_ | _0284_;
assign _0795_ = _0619_ | _0373_;
assign _0797_ = _0620_ | _0376_;
assign _0799_ = _0621_ | _0379_;
assign _0801_ = _0622_ | _0382_;
assign mem_resp_intg_err_t0 = _0623_ | _0385_;
assign multdiv_en_dec_t0 = _0624_ | _0388_;
assign _0803_ = _0625_ | _0391_;
assign _0805_ = _0626_ | _0394_;
assign branch_taken_t0 = _0627_ | _0397_;
assign _0807_ = _0628_ | _0400_;
assign _0809_ = _0629_ | _0403_;
assign _0811_ = _0630_ | _0406_;
assign stall_id_t0 = _0631_ | _0409_;
assign _0813_ = _0632_ | _0412_;
assign _0524_ = _0822_ | _0820_;
assign _0526_ = _0854_ | _0852_;
assign _0172_ = | { _0818_, _0816_, _0814_ };
assign _0729_ = _0816_ ? imm_j_type : imm_u_type;
assign _0731_ = _0814_ ? _0858_ : _0729_;
assign _0733_ = _0820_ ? imm_b_type : imm_s_type;
assign _0735_ = _0824_ ? imm_i_type : 32'd4;
assign _0737_ = _0524_ ? _0733_ : _0735_;
assign imm_b = _0172_ ? _0731_ : _0737_;
assign id_fsm_d = id_fsm_q ? _0049_ : _0022_;
assign _0010_ = id_fsm_q ? 1'h0 : _0030_;
assign _0008_ = id_fsm_q ? _0045_ : _0028_;
assign _0014_ = id_fsm_q ? _0042_ : _0032_;
assign _0012_ = id_fsm_q ? _0040_ : _0018_;
assign _0016_ = id_fsm_q ? _0047_ : _0034_;
assign _0004_ = id_fsm_q ? 1'h0 : _0024_;
assign _0000_ = id_fsm_q ? 1'h0 : _0018_;
assign _0006_ = id_fsm_q ? 1'h0 : _0026_;
assign rf_wdata_id_o = rf_wdata_sel ? csr_rdata_i : result_ex_i;
assign _0739_ = _0852_ ? imm_a : pc_id_i;
assign _0741_ = _0856_ ? lsu_addr_last_i : rf_rdata_a_i;
assign alu_operand_a_ex_o = _0526_ ? _0739_ : _0741_;
assign _0743_ = csr_op_o == /* src = "generated/sv2v_out.v:17476.34-17476.50" */ 2'h1;
assign _0745_ = csr_op_o == /* src = "generated/sv2v_out.v:17476.56-17476.72" */ 2'h2;
assign _0747_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17477.11-17477.42" */ 12'h300;
assign _0749_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17477.48-17477.79" */ 12'h304;
assign _0751_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17477.86-17477.117" */ 12'h747;
assign _0753_ = instr_rdata_i[31:25] == /* src = "generated/sv2v_out.v:17477.124-17477.153" */ 7'h1d;
assign _0755_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17481.11-17481.42" */ 12'h7b0;
assign _0757_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17481.48-17481.79" */ 12'h7b1;
assign _0759_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17481.86-17481.117" */ 12'h7b2;
assign _0761_ = instr_rdata_i[31:20] == /* src = "generated/sv2v_out.v:17481.124-17481.155" */ 12'h7b3;
assign _0763_ = csr_op_en_o && /* src = "generated/sv2v_out.v:17476.7-17476.74" */ _0767_;
assign _0765_ = csr_op_en_o && /* src = "generated/sv2v_out.v:17480.12-17480.55" */ _0781_;
assign _0767_ = _0743_ || /* src = "generated/sv2v_out.v:17476.33-17476.73" */ _0745_;
assign _0769_ = _0747_ || /* src = "generated/sv2v_out.v:17477.10-17477.80" */ _0749_;
assign _0771_ = _0769_ || /* src = "generated/sv2v_out.v:17477.9-17477.118" */ _0751_;
assign _0773_ = _0771_ || /* src = "generated/sv2v_out.v:17477.8-17477.154" */ _0753_;
assign _0774_ = _0755_ || /* src = "generated/sv2v_out.v:17481.10-17481.80" */ _0757_;
assign _0776_ = _0774_ || /* src = "generated/sv2v_out.v:17481.9-17481.118" */ _0759_;
assign _0778_ = _0776_ || /* src = "generated/sv2v_out.v:17481.8-17481.156" */ _0761_;
assign _0779_ = data_ind_timing_i || /* src = "generated/sv2v_out.v:17655.20-17655.80" */ branch_decision_i;
assign _0781_ = | /* src = "generated/sv2v_out.v:17480.38-17480.54" */ csr_op_o;
assign _0783_ = priv_mode_i != /* src = "generated/sv2v_out.v:17485.31-17485.51" */ 2'h3;
assign _0786_ = ~ /* src = "generated/sv2v_out.v:17295.60-17295.75" */ illegal_insn_o;
assign _0787_ = ~ /* src = "generated/sv2v_out.v:17484.45-17484.58" */ debug_mode_o;
assign _0788_ = ~ /* src = "generated/sv2v_out.v:17592.95-17592.115" */ instr_valid_clear_o;
assign _0789_ = ~ /* src = "generated/sv2v_out.v:17690.23-17690.32" */ stall_id;
assign _0790_ = ~ /* src = "generated/sv2v_out.v:17690.35-17690.44" */ flush_id;
assign _0785_ = ~ /* src = "generated/sv2v_out.v:17727.51-17727.69" */ instr_fetch_err_i;
assign _0791_ = ~ /* src = "generated/sv2v_out.v:17751.65-17751.82" */ lsu_resp_valid_i;
assign _0792_ = ~ /* src = "generated/sv2v_out.v:17755.36-17755.46" */ ebrk_insn;
assign _0793_ = ~ /* src = "generated/sv2v_out.v:17755.49-17755.64" */ ecall_insn_dec;
assign _0794_ = mret_insn_dec | /* src = "generated/sv2v_out.v:17485.56-17485.105" */ _0057_;
assign _0796_ = illegal_insn_dec | /* src = "generated/sv2v_out.v:17486.45-17486.82" */ illegal_csr_insn_i;
assign _0798_ = _0796_ | /* src = "generated/sv2v_out.v:17486.44-17486.103" */ illegal_dret_insn;
assign _0800_ = _0798_ | /* src = "generated/sv2v_out.v:17486.43-17486.125" */ illegal_umode_insn;
assign mem_resp_intg_err = lsu_load_resp_intg_err_i | /* src = "generated/sv2v_out.v:17487.29-17487.81" */ lsu_store_resp_intg_err_i;
assign multdiv_en_dec = mult_en_dec | /* src = "generated/sv2v_out.v:17559.26-17559.50" */ div_en_dec;
assign _0802_ = branch_set_raw | /* src = "generated/sv2v_out.v:17592.36-17592.65" */ jump_set_raw;
assign _0804_ = _0802_ | /* src = "generated/sv2v_out.v:17592.35-17592.91" */ branch_jump_set_done_q;
assign branch_taken = _0105_ | /* src = "generated/sv2v_out.v:17608.26-17608.61" */ \g_sec_branch_taken.branch_taken_q ;
assign _0697_ = branch_decision_i | /* src = "generated/sv2v_out.v:17657.27-17657.64" */ data_ind_timing_i;
assign _0806_ = stall_mem | /* src = "generated/sv2v_out.v:17689.23-17689.64" */ stall_multdiv;
assign _0808_ = _0806_ | /* src = "generated/sv2v_out.v:17689.22-17689.78" */ stall_jump;
assign _0810_ = _0808_ | /* src = "generated/sv2v_out.v:17689.21-17689.94" */ stall_branch;
assign stall_id = _0810_ | /* src = "generated/sv2v_out.v:17689.20-17689.107" */ stall_alu;
assign _0812_ = _0791_ | /* src = "generated/sv2v_out.v:17725.55-17725.92" */ instr_first_cycle_id_o;
/* src = "generated/sv2v_out.v:17603.4-17607.42" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME \g_sec_branch_taken.branch_taken_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_sec_branch_taken.branch_taken_q  <= 1'h0;
else \g_sec_branch_taken.branch_taken_q  <= branch_decision_i;
/* src = "generated/sv2v_out.v:17584.4-17588.43" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME branch_set_raw */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_set_raw <= 1'h0;
else branch_set_raw <= branch_set_raw_d;
/* src = "generated/sv2v_out.v:17593.2-17597.53" */
/* PC_TAINT_INFO MODULE_NAME \$paramod$f727fb3fc3020e3d8c2544b0dd6ded81f558314e\ibex_id_stage  */
/* PC_TAINT_INFO STATE_NAME branch_jump_set_done_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_jump_set_done_q <= 1'h0;
else branch_jump_set_done_q <= branch_jump_set_done_d;
assign _0814_ = imm_b_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17383.5-17392.12" */ 3'h5;
assign _0816_ = imm_b_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17383.5-17392.12" */ 3'h4;
assign _0818_ = imm_b_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17383.5-17392.12" */ 3'h3;
assign _0820_ = imm_b_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17383.5-17392.12" */ 3'h2;
assign _0822_ = imm_b_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17383.5-17392.12" */ 3'h1;
assign _0824_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17383.5-17392.12" */ imm_b_mux_sel;
assign _0049_ = _0065_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17677.10-17677.38|generated/sv2v_out.v:17677.6-17683.9" */ 1'h0 : 1'h1;
assign _0042_ = _0065_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17677.10-17677.38|generated/sv2v_out.v:17677.6-17683.9" */ 1'h0 : jump_in_dec;
assign _0040_ = _0065_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17677.10-17677.38|generated/sv2v_out.v:17677.6-17683.9" */ 1'h0 : branch_in_dec;
assign _0047_ = _0065_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17677.10-17677.38|generated/sv2v_out.v:17677.6-17683.9" */ 1'h0 : multdiv_en_dec;
assign _0045_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17675.10-17675.24|generated/sv2v_out.v:17675.6-17676.42" */ _0063_ : rf_we_dec;
assign _0038_ = ex_valid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17649.12-17649.23|generated/sv2v_out.v:17649.8-17653.11" */ rf_we_dec : 1'h0;
assign _0044_ = ex_valid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17649.12-17649.23|generated/sv2v_out.v:17649.8-17653.11" */ 1'h0 : 1'h1;
assign _0686_ = alu_multicycle_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h1 : 1'h0;
assign _0826_ = jump_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h1 : _0686_;
assign _0828_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ _0859_ : _0826_;
assign _0830_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ _0044_ : _0828_;
assign _0022_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h1 : _0830_;
assign _0687_ = jump_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h0 : _0686_;
assign _0688_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h0 : _0687_;
assign _0689_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h0 : _0688_;
assign _0030_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h0 : _0689_;
assign _0835_ = alu_multicycle_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h0 : rf_we_dec;
assign _0837_ = jump_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ rf_we_dec : _0835_;
assign _0839_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ rf_we_dec : _0837_;
assign _0841_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ _0038_ : _0839_;
assign _0028_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ rf_we_dec : _0841_;
assign _0694_ = jump_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h1 : 1'h0;
assign _0695_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h0 : _0694_;
assign _0696_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h0 : _0695_;
assign _0032_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h0 : _0696_;
assign _0698_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ _0697_ : 1'h0;
assign _0699_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h0 : _0698_;
assign _0018_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h0 : _0699_;
assign _0700_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ _0044_ : 1'h0;
assign _0034_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h0 : _0700_;
assign _0701_ = jump_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ jump_set_dec : 1'h0;
assign _0702_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h0 : _0701_;
assign _0703_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h0 : _0702_;
assign _0024_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h0 : _0703_;
assign _0704_ = branch_in_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h1 : 1'h0;
assign _0705_ = multdiv_en_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h0 : _0704_;
assign _0026_ = lsu_req_dec ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17642.6-17673.13" */ 1'h0 : _0705_;
assign stall_alu = instr_executing ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17639.7-17639.27|generated/sv2v_out.v:17639.3-17686.11" */ _0010_ : 1'h0;
assign rf_we_raw = instr_executing ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17639.7-17639.27|generated/sv2v_out.v:17639.3-17686.11" */ _0008_ : rf_we_dec;
assign stall_jump = instr_executing ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17639.7-17639.27|generated/sv2v_out.v:17639.3-17686.11" */ _0014_ : 1'h0;
assign stall_branch = instr_executing ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17639.7-17639.27|generated/sv2v_out.v:17639.3-17686.11" */ _0012_ : 1'h0;
assign stall_multdiv = instr_executing ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17639.7-17639.27|generated/sv2v_out.v:17639.3-17686.11" */ _0016_ : 1'h0;
assign jump_set_raw = instr_executing ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17639.7-17639.27|generated/sv2v_out.v:17639.3-17686.11" */ _0004_ : 1'h0;
assign branch_set_raw_d = instr_executing ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17639.7-17639.27|generated/sv2v_out.v:17639.3-17686.11" */ _0000_ : 1'h0;
assign perf_branch_o = instr_executing ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17639.7-17639.27|generated/sv2v_out.v:17639.3-17686.11" */ _0006_ : 1'h0;
assign _0036_ = _0778_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17481.8-17481.156|generated/sv2v_out.v:17481.4-17482.27" */ 1'h1 : 1'h0;
assign _0020_ = _0765_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17480.12-17480.55|generated/sv2v_out.v:17480.8-17482.27" */ _0036_ : 1'h0;
assign _0002_ = _0773_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17477.8-17477.154|generated/sv2v_out.v:17477.4-17478.27" */ 1'h1 : 1'h0;
assign csr_pipe_flush = _0763_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:17476.7-17476.74|generated/sv2v_out.v:17476.3-17482.27" */ _0002_ : _0020_;
assign _0852_ = alu_op_a_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17334.3-17340.10" */ 2'h3;
assign _0854_ = alu_op_a_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17334.3-17340.10" */ 2'h2;
assign _0856_ = alu_op_a_mux_sel == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:17334.3-17340.10" */ 2'h1;
assign alu_op_a_mux_sel = lsu_addr_incr_req_i ? /* src = "generated/sv2v_out.v:17329.29-17329.78" */ 2'h1 : alu_op_a_mux_sel_dec;
assign alu_op_b_mux_sel = lsu_addr_incr_req_i ? /* src = "generated/sv2v_out.v:17330.29-17330.78" */ 1'h1 : alu_op_b_mux_sel_dec;
assign imm_b_mux_sel = lsu_addr_incr_req_i ? /* src = "generated/sv2v_out.v:17331.26-17331.72" */ 3'h6 : imm_b_mux_sel_dec;
assign imm_a = imm_a_mux_sel ? /* src = "generated/sv2v_out.v:17332.18-17332.70" */ 32'd0 : zimm_rs1_type;
assign _0858_ = instr_is_compressed_i ? /* src = "generated/sv2v_out.v:17389.21-17389.72" */ 32'd2 : 32'd4;
assign alu_operand_b_ex_o = alu_op_b_mux_sel ? /* src = "generated/sv2v_out.v:17396.26-17396.75" */ imm_b : rf_rdata_b_i;
assign lsu_req_o = instr_executing ? /* src = "generated/sv2v_out.v:17560.20-17560.75" */ _0059_ : 1'h0;
assign mult_en_ex_o = instr_executing ? /* src = "generated/sv2v_out.v:17561.23-17561.59" */ mult_en_dec : 1'h0;
assign div_en_ex_o = instr_executing ? /* src = "generated/sv2v_out.v:17562.22-17562.57" */ div_en_dec : 1'h0;
assign _0859_ = _0779_ ? /* src = "generated/sv2v_out.v:17655.20-17655.94" */ 1'h1 : 1'h0;
assign multicycle_done = lsu_req_dec ? /* src = "generated/sv2v_out.v:17723.30-17723.73" */ lsu_resp_valid_i : ex_valid_i;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:17492.4-17558.3" */
\$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  controller_i (
.branch_not_set_i(1'h0),
.branch_not_set_i_t0(1'h0),
.branch_set_i(branch_set),
.branch_set_i_t0(branch_set_t0),
.clk_i(clk_i),
.controller_run_o(controller_run),
.controller_run_o_t0(controller_run_t0),
.csr_mstatus_mie_i(csr_mstatus_mie_i),
.csr_mstatus_mie_i_t0(csr_mstatus_mie_i_t0),
.csr_mtval_o(csr_mtval_o),
.csr_mtval_o_t0(csr_mtval_o_t0),
.csr_pipe_flush_i(csr_pipe_flush),
.csr_pipe_flush_i_t0(csr_pipe_flush_t0),
.csr_restore_dret_id_o(csr_restore_dret_id_o),
.csr_restore_dret_id_o_t0(csr_restore_dret_id_o_t0),
.csr_restore_mret_id_o(csr_restore_mret_id_o),
.csr_restore_mret_id_o_t0(csr_restore_mret_id_o_t0),
.csr_save_cause_o(csr_save_cause_o),
.csr_save_cause_o_t0(csr_save_cause_o_t0),
.csr_save_id_o(csr_save_id_o),
.csr_save_id_o_t0(csr_save_id_o_t0),
.csr_save_if_o(csr_save_if_o),
.csr_save_if_o_t0(csr_save_if_o_t0),
.csr_save_wb_o(csr_save_wb_o),
.csr_save_wb_o_t0(csr_save_wb_o_t0),
.ctrl_busy_o(ctrl_busy_o),
.ctrl_busy_o_t0(ctrl_busy_o_t0),
.debug_cause_o(debug_cause_o),
.debug_cause_o_t0(debug_cause_o_t0),
.debug_csr_save_o(debug_csr_save_o),
.debug_csr_save_o_t0(debug_csr_save_o_t0),
.debug_ebreakm_i(debug_ebreakm_i),
.debug_ebreakm_i_t0(debug_ebreakm_i_t0),
.debug_ebreaku_i(debug_ebreaku_i),
.debug_ebreaku_i_t0(debug_ebreaku_i_t0),
.debug_mode_entering_o(debug_mode_entering_o),
.debug_mode_entering_o_t0(debug_mode_entering_o_t0),
.debug_mode_o(debug_mode_o),
.debug_mode_o_t0(debug_mode_o_t0),
.debug_req_i(debug_req_i),
.debug_req_i_t0(debug_req_i_t0),
.debug_single_step_i(debug_single_step_i),
.debug_single_step_i_t0(debug_single_step_i_t0),
.dret_insn_i(dret_insn_dec),
.dret_insn_i_t0(dret_insn_dec_t0),
.ebrk_insn_i(ebrk_insn),
.ebrk_insn_i_t0(ebrk_insn_t0),
.ecall_insn_i(ecall_insn_dec),
.ecall_insn_i_t0(ecall_insn_dec_t0),
.exc_cause_o(exc_cause_o),
.exc_cause_o_t0(exc_cause_o_t0),
.exc_pc_mux_o(exc_pc_mux_o),
.exc_pc_mux_o_t0(exc_pc_mux_o_t0),
.flush_id_o(flush_id),
.flush_id_o_t0(flush_id_t0),
.id_exception_o(\gen_no_stall_mem.unused_id_exception ),
.id_exception_o_t0(\gen_no_stall_mem.unused_id_exception_t0 ),
.id_in_ready_o(id_in_ready_o),
.id_in_ready_o_t0(id_in_ready_o_t0),
.illegal_insn_i(illegal_insn_o),
.illegal_insn_i_t0(illegal_insn_o_t0),
.instr_bp_taken_i(instr_bp_taken_i),
.instr_bp_taken_i_t0(instr_bp_taken_i_t0),
.instr_compressed_i(instr_rdata_c_i),
.instr_compressed_i_t0(instr_rdata_c_i_t0),
.instr_exec_i(instr_exec_i),
.instr_exec_i_t0(instr_exec_i_t0),
.instr_fetch_err_i(instr_fetch_err_i),
.instr_fetch_err_i_t0(instr_fetch_err_i_t0),
.instr_fetch_err_plus2_i(instr_fetch_err_plus2_i),
.instr_fetch_err_plus2_i_t0(instr_fetch_err_plus2_i_t0),
.instr_i(instr_rdata_i),
.instr_i_t0(instr_rdata_i_t0),
.instr_is_compressed_i(instr_is_compressed_i),
.instr_is_compressed_i_t0(instr_is_compressed_i_t0),
.instr_req_o(instr_req_o),
.instr_req_o_t0(instr_req_o_t0),
.instr_valid_clear_o(instr_valid_clear_o),
.instr_valid_clear_o_t0(instr_valid_clear_o_t0),
.instr_valid_i(instr_valid_i),
.instr_valid_i_t0(instr_valid_i_t0),
.irq_nm_ext_i(irq_nm_i),
.irq_nm_ext_i_t0(irq_nm_i_t0),
.irq_pending_i(irq_pending_i),
.irq_pending_i_t0(irq_pending_i_t0),
.irqs_i(irqs_i),
.irqs_i_t0(irqs_i_t0),
.jump_set_i(jump_set),
.jump_set_i_t0(jump_set_t0),
.load_err_i(lsu_load_err_i),
.load_err_i_t0(lsu_load_err_i_t0),
.lsu_addr_last_i(lsu_addr_last_i),
.lsu_addr_last_i_t0(lsu_addr_last_i_t0),
.mem_resp_intg_err_i(mem_resp_intg_err),
.mem_resp_intg_err_i_t0(mem_resp_intg_err_t0),
.mret_insn_i(mret_insn_dec),
.mret_insn_i_t0(mret_insn_dec_t0),
.nmi_mode_o(nmi_mode_o),
.nmi_mode_o_t0(nmi_mode_o_t0),
.nt_branch_mispredict_o(nt_branch_mispredict_o),
.nt_branch_mispredict_o_t0(nt_branch_mispredict_o_t0),
.pc_id_i(pc_id_i),
.pc_id_i_t0(pc_id_i_t0),
.pc_mux_o(pc_mux_o),
.pc_mux_o_t0(pc_mux_o_t0),
.pc_set_o(pc_set_o),
.pc_set_o_t0(pc_set_o_t0),
.perf_jump_o(perf_jump_o),
.perf_jump_o_t0(perf_jump_o_t0),
.perf_tbranch_o(perf_tbranch_o),
.perf_tbranch_o_t0(perf_tbranch_o_t0),
.priv_mode_i(priv_mode_i),
.priv_mode_i_t0(priv_mode_i_t0),
.ready_wb_i(ready_wb_i),
.ready_wb_i_t0(ready_wb_i_t0),
.rst_ni(rst_ni),
.stall_id_i(stall_id),
.stall_id_i_t0(stall_id_t0),
.stall_wb_i(1'h0),
.stall_wb_i_t0(1'h0),
.store_err_i(lsu_store_err_i),
.store_err_i_t0(lsu_store_err_i_t0),
.trigger_match_i(trigger_match_i),
.trigger_match_i_t0(trigger_match_i_t0),
.wb_exception_o(\gen_no_stall_mem.unused_wb_exception ),
.wb_exception_o_t0(\gen_no_stall_mem.unused_wb_exception_t0 ),
.wfi_insn_i(wfi_insn_dec),
.wfi_insn_i_t0(wfi_insn_dec_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:17422.4-17473.3" */
\$paramod$5ffe4cc9ba21eb548f33468a0c4a93d38de3dae5\ibex_decoder  decoder_i (
.alu_multicycle_o(alu_multicycle_dec),
.alu_multicycle_o_t0(alu_multicycle_dec_t0),
.alu_op_a_mux_sel_o(alu_op_a_mux_sel_dec),
.alu_op_a_mux_sel_o_t0(alu_op_a_mux_sel_dec_t0),
.alu_op_b_mux_sel_o(alu_op_b_mux_sel_dec),
.alu_op_b_mux_sel_o_t0(alu_op_b_mux_sel_dec_t0),
.alu_operator_o(alu_operator_ex_o),
.alu_operator_o_t0(alu_operator_ex_o_t0),
.branch_in_dec_o(branch_in_dec),
.branch_in_dec_o_t0(branch_in_dec_t0),
.branch_taken_i(branch_taken),
.branch_taken_i_t0(branch_taken_t0),
.bt_a_mux_sel_o(bt_a_mux_sel),
.bt_a_mux_sel_o_t0(bt_a_mux_sel_t0),
.bt_b_mux_sel_o(bt_b_mux_sel),
.bt_b_mux_sel_o_t0(bt_b_mux_sel_t0),
.clk_i(clk_i),
.csr_access_o(csr_access_o),
.csr_access_o_t0(csr_access_o_t0),
.csr_op_o(csr_op_o),
.csr_op_o_t0(csr_op_o_t0),
.data_req_o(lsu_req_dec),
.data_req_o_t0(lsu_req_dec_t0),
.data_sign_extension_o(lsu_sign_ext_o),
.data_sign_extension_o_t0(lsu_sign_ext_o_t0),
.data_type_o(lsu_type_o),
.data_type_o_t0(lsu_type_o_t0),
.data_we_o(lsu_we_o),
.data_we_o_t0(lsu_we_o_t0),
.div_en_o(div_en_dec),
.div_en_o_t0(div_en_dec_t0),
.div_sel_o(div_sel_ex_o),
.div_sel_o_t0(div_sel_ex_o_t0),
.dret_insn_o(dret_insn_dec),
.dret_insn_o_t0(dret_insn_dec_t0),
.ebrk_insn_o(ebrk_insn),
.ebrk_insn_o_t0(ebrk_insn_t0),
.ecall_insn_o(ecall_insn_dec),
.ecall_insn_o_t0(ecall_insn_dec_t0),
.icache_inval_o(icache_inval_o),
.icache_inval_o_t0(icache_inval_o_t0),
.illegal_c_insn_i(illegal_c_insn_i),
.illegal_c_insn_i_t0(illegal_c_insn_i_t0),
.illegal_insn_o(illegal_insn_dec),
.illegal_insn_o_t0(illegal_insn_dec_t0),
.imm_a_mux_sel_o(imm_a_mux_sel),
.imm_a_mux_sel_o_t0(imm_a_mux_sel_t0),
.imm_b_mux_sel_o(imm_b_mux_sel_dec),
.imm_b_mux_sel_o_t0(imm_b_mux_sel_dec_t0),
.imm_b_type_o(imm_b_type),
.imm_b_type_o_t0(imm_b_type_t0),
.imm_i_type_o(imm_i_type),
.imm_i_type_o_t0(imm_i_type_t0),
.imm_j_type_o(imm_j_type),
.imm_j_type_o_t0(imm_j_type_t0),
.imm_s_type_o(imm_s_type),
.imm_s_type_o_t0(imm_s_type_t0),
.imm_u_type_o(imm_u_type),
.imm_u_type_o_t0(imm_u_type_t0),
.instr_first_cycle_i(instr_first_cycle_id_o),
.instr_first_cycle_i_t0(instr_first_cycle_id_o_t0),
.instr_rdata_alu_i(instr_rdata_alu_i),
.instr_rdata_alu_i_t0(instr_rdata_alu_i_t0),
.instr_rdata_i(instr_rdata_i),
.instr_rdata_i_t0(instr_rdata_i_t0),
.jump_in_dec_o(jump_in_dec),
.jump_in_dec_o_t0(jump_in_dec_t0),
.jump_set_o(jump_set_dec),
.jump_set_o_t0(jump_set_dec_t0),
.mret_insn_o(mret_insn_dec),
.mret_insn_o_t0(mret_insn_dec_t0),
.mult_en_o(mult_en_dec),
.mult_en_o_t0(mult_en_dec_t0),
.mult_sel_o(mult_sel_ex_o),
.mult_sel_o_t0(mult_sel_ex_o_t0),
.multdiv_operator_o(multdiv_operator_ex_o),
.multdiv_operator_o_t0(multdiv_operator_ex_o_t0),
.multdiv_signed_mode_o(multdiv_signed_mode_ex_o),
.multdiv_signed_mode_o_t0(multdiv_signed_mode_ex_o_t0),
.rf_raddr_a_o(rf_raddr_a_o),
.rf_raddr_a_o_t0(rf_raddr_a_o_t0),
.rf_raddr_b_o(rf_raddr_b_o),
.rf_raddr_b_o_t0(rf_raddr_b_o_t0),
.rf_ren_a_o(rf_ren_a_dec),
.rf_ren_a_o_t0(rf_ren_a_dec_t0),
.rf_ren_b_o(rf_ren_b_dec),
.rf_ren_b_o_t0(rf_ren_b_dec_t0),
.rf_waddr_o(rf_waddr_id_o),
.rf_waddr_o_t0(rf_waddr_id_o_t0),
.rf_wdata_sel_o(rf_wdata_sel),
.rf_wdata_sel_o_t0(rf_wdata_sel_t0),
.rf_we_o(rf_we_dec),
.rf_we_o_t0(rf_we_dec_t0),
.rst_ni(rst_ni),
.wfi_insn_o(wfi_insn_dec),
.wfi_insn_o_t0(wfi_insn_dec_t0),
.zimm_rs1_type_o(zimm_rs1_type),
.zimm_rs1_type_o_t0(zimm_rs1_type_t0)
);
assign bt_a_operand_o = 32'd0;
assign bt_a_operand_o_t0 = 32'd0;
assign bt_b_operand_o = 32'd0;
assign bt_b_operand_o_t0 = 32'd0;
assign instr_id_done_o = en_wb_o;
assign instr_id_done_o_t0 = en_wb_o_t0;
assign instr_type_wb_o = 2'h2;
assign instr_type_wb_o_t0 = 2'h0;
assign lsu_wdata_o = rf_rdata_b_i;
assign lsu_wdata_o_t0 = rf_rdata_b_i_t0;
assign multdiv_operand_a_ex_o = rf_rdata_a_i;
assign multdiv_operand_a_ex_o_t0 = rf_rdata_a_i_t0;
assign multdiv_operand_b_ex_o = rf_rdata_b_i;
assign multdiv_operand_b_ex_o_t0 = rf_rdata_b_i_t0;
assign multdiv_ready_id_o = ready_wb_i;
assign multdiv_ready_id_o_t0 = ready_wb_i_t0;
assign nt_branch_addr_o = 32'd0;
assign nt_branch_addr_o_t0 = 32'd0;
assign rf_rd_a_wb_match_o = 1'h0;
assign rf_rd_a_wb_match_o_t0 = 1'h0;
assign rf_rd_b_wb_match_o = 1'h0;
assign rf_rd_b_wb_match_o_t0 = 1'h0;
endmodule

module \$paramod\ibex_alu\RV32B=s32'00000000000000000000000000000000 (operator_i, operand_a_i, operand_b_i, instr_first_cycle_i, multdiv_operand_a_i, multdiv_operand_b_i, multdiv_sel_i, imd_val_q_i, imd_val_d_o, imd_val_we_o, adder_result_o, adder_result_ext_o, result_o, comparison_result_o, is_equal_result_o, instr_first_cycle_i_t0, imd_val_d_o_t0, imd_val_q_i_t0, imd_val_we_o_t0, operator_i_t0, adder_result_ext_o_t0
, adder_result_o_t0, comparison_result_o_t0, is_equal_result_o_t0, multdiv_operand_a_i_t0, multdiv_operand_b_i_t0, multdiv_sel_i_t0, operand_a_i_t0, operand_b_i_t0, result_o_t0);
/* src = "generated/sv2v_out.v:11397.52-11397.83" */
wire _0000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11397.52-11397.83" */
wire _0001_;
wire [33:0] _0002_;
wire [33:0] _0003_;
wire _0004_;
wire [6:0] _0005_;
wire _0006_;
wire _0007_;
wire _0008_;
wire _0009_;
wire _0010_;
wire _0011_;
wire _0012_;
wire _0013_;
wire [31:0] _0014_;
wire [7:0] _0015_;
wire [4:0] _0016_;
wire [4:0] _0017_;
wire [5:0] _0018_;
wire [5:0] _0019_;
wire [3:0] _0020_;
wire [4:0] _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire _0026_;
wire _0027_;
wire _0028_;
wire _0029_;
wire _0030_;
wire [31:0] _0031_;
wire [31:0] _0032_;
wire [31:0] _0033_;
wire _0034_;
wire _0035_;
wire _0036_;
wire _0037_;
wire _0038_;
wire _0039_;
wire _0040_;
wire _0041_;
wire [31:0] _0042_;
wire [31:0] _0043_;
wire _0044_;
wire [32:0] _0045_;
wire [32:0] _0046_;
wire _0047_;
wire [4:0] _0048_;
wire [31:0] _0049_;
wire _0050_;
wire _0051_;
wire _0052_;
wire _0053_;
wire [31:0] _0054_;
wire _0055_;
wire _0056_;
wire _0057_;
wire [31:0] _0058_;
wire _0059_;
wire _0060_;
wire [5:0] _0061_;
wire [31:0] _0062_;
wire _0063_;
/* cellift = 32'd1 */
wire _0064_;
wire [33:0] _0065_;
wire [33:0] _0066_;
wire _0067_;
wire _0068_;
wire _0069_;
wire [31:0] _0070_;
wire [31:0] _0071_;
wire [31:0] _0072_;
wire _0073_;
wire _0074_;
wire _0075_;
wire _0076_;
wire _0077_;
wire _0078_;
wire [31:0] _0079_;
wire [31:0] _0080_;
wire [31:0] _0081_;
wire [31:0] _0082_;
wire [31:0] _0083_;
wire [31:0] _0084_;
wire [31:0] _0085_;
wire [31:0] _0086_;
wire [31:0] _0087_;
wire [31:0] _0088_;
wire [31:0] _0089_;
wire _0090_;
wire _0091_;
wire _0092_;
wire _0093_;
wire _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire [31:0] _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire _0109_;
wire _0110_;
wire _0111_;
wire _0112_;
wire _0113_;
wire _0114_;
wire _0115_;
wire _0116_;
wire _0117_;
wire _0118_;
wire _0119_;
wire _0120_;
wire _0121_;
wire _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire [31:0] _0130_;
wire [31:0] _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire [7:0] _0138_;
wire [6:0] _0139_;
wire [4:0] _0140_;
wire [4:0] _0141_;
wire [5:0] _0142_;
wire [31:0] _0143_;
wire [31:0] _0144_;
wire [31:0] _0145_;
wire [31:0] _0146_;
wire [31:0] _0147_;
wire [31:0] _0148_;
wire [5:0] _0149_;
wire [3:0] _0150_;
wire _0151_;
wire _0152_;
wire _0153_;
wire [4:0] _0154_;
wire [32:0] _0155_;
wire [32:0] _0156_;
wire [32:0] _0157_;
wire [32:0] _0158_;
wire [32:0] _0159_;
wire [32:0] _0160_;
wire [32:0] _0161_;
wire [32:0] _0162_;
wire [32:0] _0163_;
wire _0164_;
wire _0165_;
wire [5:0] _0166_;
wire [527:0] _0167_;
/* unused_bits = "32" */
wire [32:0] _0168_;
wire [31:0] _0169_;
wire [4:0] _0170_;
wire [4:0] _0171_;
wire [4:0] _0172_;
wire [31:0] _0173_;
wire [31:0] _0174_;
wire [31:0] _0175_;
wire [31:0] _0176_;
wire [31:0] _0177_;
wire [31:0] _0178_;
wire _0179_;
/* cellift = 32'd1 */
wire _0180_;
wire _0181_;
/* cellift = 32'd1 */
wire _0182_;
wire [33:0] _0183_;
wire [33:0] _0184_;
wire [33:0] _0185_;
wire _0186_;
wire [31:0] _0187_;
wire _0188_;
wire _0189_;
wire [31:0] _0190_;
wire [31:0] _0191_;
wire [31:0] _0192_;
wire [31:0] _0193_;
wire [31:0] _0194_;
wire [31:0] _0195_;
wire [31:0] _0196_;
wire [31:0] _0197_;
wire [31:0] _0198_;
wire [31:0] _0199_;
wire _0200_;
wire _0201_;
wire _0202_;
wire _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
wire _0221_;
wire _0222_;
wire [31:0] _0223_;
wire _0224_;
wire _0225_;
wire [31:0] _0226_;
wire [31:0] _0227_;
wire [31:0] _0228_;
wire [31:0] _0229_;
wire [31:0] _0230_;
wire [31:0] _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire [32:0] _0235_;
wire [32:0] _0236_;
wire [32:0] _0237_;
wire [32:0] _0238_;
wire [32:0] _0239_;
wire [32:0] _0240_;
wire [32:0] _0241_;
wire _0242_;
wire [527:0] _0243_;
wire [527:0] _0244_;
wire [32:0] _0245_;
wire [31:0] _0246_;
wire [31:0] _0247_;
wire [4:0] _0248_;
wire [4:0] _0249_;
wire [4:0] _0250_;
wire [31:0] _0251_;
wire [31:0] _0252_;
wire [31:0] _0253_;
wire [31:0] _0254_;
wire [33:0] _0255_;
wire [31:0] _0256_;
wire [31:0] _0257_;
wire [31:0] _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire _0271_;
wire _0272_;
wire [31:0] _0273_;
wire [31:0] _0274_;
wire _0275_;
wire [32:0] _0276_;
wire [32:0] _0277_;
wire [32:0] _0278_;
wire [527:0] _0279_;
wire [32:0] _0280_;
wire [4:0] _0281_;
wire [31:0] _0282_;
wire [31:0] _0283_;
wire _0284_;
wire _0285_;
wire _0286_;
wire _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire _0294_;
wire _0295_;
wire _0296_;
wire _0297_;
wire _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire _0302_;
wire _0303_;
wire _0304_;
wire _0305_;
wire _0306_;
wire _0307_;
wire _0308_;
wire _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire _0313_;
wire _0314_;
wire _0315_;
wire _0316_;
wire _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire _0322_;
wire _0323_;
wire _0324_;
wire _0325_;
wire _0326_;
wire _0327_;
wire _0328_;
wire _0329_;
wire _0330_;
wire _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire _0335_;
wire _0336_;
wire _0337_;
wire _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire _0344_;
wire _0345_;
wire _0346_;
wire _0347_;
wire _0348_;
wire _0349_;
wire _0350_;
wire _0351_;
wire _0352_;
wire _0353_;
wire _0354_;
wire _0355_;
wire _0356_;
wire _0357_;
wire _0358_;
wire _0359_;
wire _0360_;
wire _0361_;
wire _0362_;
wire _0363_;
wire _0364_;
wire _0365_;
wire _0366_;
wire _0367_;
wire _0368_;
wire _0369_;
wire [33:0] _0370_;
wire [33:0] _0371_;
wire [31:0] _0372_;
wire [31:0] _0373_;
wire [31:0] _0374_;
/* cellift = 32'd1 */
wire [31:0] _0375_;
wire [31:0] _0376_;
/* cellift = 32'd1 */
wire [31:0] _0377_;
wire [31:0] _0378_;
/* cellift = 32'd1 */
wire [31:0] _0379_;
wire _0380_;
/* cellift = 32'd1 */
wire _0381_;
wire _0382_;
/* cellift = 32'd1 */
wire _0383_;
wire [32:0] _0384_;
wire [32:0] _0385_;
/* src = "generated/sv2v_out.v:11318.23-11318.47" */
wire _0386_;
/* src = "generated/sv2v_out.v:11426.23-11426.41" */
wire _0387_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11426.23-11426.41" */
wire _0388_;
/* src = "generated/sv2v_out.v:11426.46-11426.64" */
wire _0389_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11426.46-11426.64" */
wire _0390_;
/* src = "generated/sv2v_out.v:11427.24-11427.42" */
wire _0391_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11427.24-11427.42" */
wire _0392_;
/* src = "generated/sv2v_out.v:11427.47-11427.65" */
wire _0393_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11427.47-11427.65" */
wire _0394_;
wire _0395_;
/* cellift = 32'd1 */
wire _0396_;
wire _0397_;
/* cellift = 32'd1 */
wire _0398_;
wire _0399_;
/* cellift = 32'd1 */
wire _0400_;
wire _0401_;
/* cellift = 32'd1 */
wire _0402_;
/* cellift = 32'd1 */
wire _0403_;
/* cellift = 32'd1 */
wire _0404_;
/* cellift = 32'd1 */
wire _0405_;
wire _0406_;
/* cellift = 32'd1 */
wire _0407_;
wire _0408_;
/* cellift = 32'd1 */
wire _0409_;
/* cellift = 32'd1 */
wire _0410_;
wire _0411_;
/* cellift = 32'd1 */
wire _0412_;
/* cellift = 32'd1 */
wire _0413_;
wire _0414_;
/* cellift = 32'd1 */
wire _0415_;
wire _0416_;
/* cellift = 32'd1 */
wire _0417_;
/* src = "generated/sv2v_out.v:11325.24-11325.33" */
wire _0418_;
/* src = "generated/sv2v_out.v:11327.59-11327.76" */
wire _0419_;
wire [7:0] _0420_;
/* cellift = 32'd1 */
wire [7:0] _0421_;
wire _0422_;
/* cellift = 32'd1 */
wire _0423_;
wire [4:0] _0424_;
/* cellift = 32'd1 */
wire [4:0] _0425_;
wire _0426_;
/* cellift = 32'd1 */
wire _0427_;
wire [4:0] _0428_;
/* cellift = 32'd1 */
wire [4:0] _0429_;
wire _0430_;
/* cellift = 32'd1 */
wire _0431_;
wire [5:0] _0432_;
/* cellift = 32'd1 */
wire [5:0] _0433_;
wire _0434_;
/* cellift = 32'd1 */
wire _0435_;
wire [31:0] _0436_;
/* cellift = 32'd1 */
wire [31:0] _0437_;
wire [5:0] _0438_;
/* cellift = 32'd1 */
wire [5:0] _0439_;
wire _0440_;
/* cellift = 32'd1 */
wire _0441_;
wire [3:0] _0442_;
/* cellift = 32'd1 */
wire [3:0] _0443_;
wire _0444_;
/* cellift = 32'd1 */
wire _0445_;
wire _0446_;
wire [32:0] _0447_;
/* cellift = 32'd1 */
wire [32:0] _0448_;
/* src = "generated/sv2v_out.v:11364.27-11364.48" */
/* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] _0449_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11364.27-11364.48" */
/* unused_bits = "5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" */
wire [31:0] _0450_;
/* src = "generated/sv2v_out.v:11317.8-11317.41" */
wire _0451_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11317.8-11317.41" */
wire _0452_;
/* src = "generated/sv2v_out.v:11320.23-11320.51" */
wire _0453_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11320.23-11320.51" */
wire _0454_;
/* src = "generated/sv2v_out.v:11265.13-11265.23" */
wire [32:0] adder_in_a;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11265.13-11265.23" */
wire [32:0] adder_in_a_t0;
/* src = "generated/sv2v_out.v:11266.13-11266.23" */
wire [32:0] adder_in_b;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11266.13-11266.23" */
wire [32:0] adder_in_b_t0;
/* src = "generated/sv2v_out.v:11264.6-11264.23" */
wire adder_op_b_negate;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11264.6-11264.23" */
wire adder_op_b_negate_t0;
/* src = "generated/sv2v_out.v:11249.21-11249.39" */
output [33:0] adder_result_ext_o;
wire [33:0] adder_result_ext_o;
/* cellift = 32'd1 */
output [33:0] adder_result_ext_o_t0;
wire [33:0] adder_result_ext_o_t0;
/* src = "generated/sv2v_out.v:11248.21-11248.35" */
output [31:0] adder_result_o;
wire [31:0] adder_result_o;
/* cellift = 32'd1 */
output [31:0] adder_result_o_t0;
wire [31:0] adder_result_o_t0;
/* src = "generated/sv2v_out.v:11409.7-11409.18" */
wire bwlogic_and;
/* src = "generated/sv2v_out.v:11412.14-11412.32" */
wire [31:0] bwlogic_and_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11412.14-11412.32" */
wire [31:0] bwlogic_and_result_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11409.7-11409.18" */
wire bwlogic_and_t0;
/* src = "generated/sv2v_out.v:11408.7-11408.17" */
wire bwlogic_or;
/* src = "generated/sv2v_out.v:11411.14-11411.31" */
wire [31:0] bwlogic_or_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11411.14-11411.31" */
wire [31:0] bwlogic_or_result_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11408.7-11408.17" */
wire bwlogic_or_t0;
/* src = "generated/sv2v_out.v:11414.13-11414.27" */
wire [31:0] bwlogic_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11414.13-11414.27" */
wire [31:0] bwlogic_result_t0;
/* src = "generated/sv2v_out.v:11413.14-11413.32" */
wire [31:0] bwlogic_xor_result;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11413.14-11413.32" */
wire [31:0] bwlogic_xor_result_t0;
/* src = "generated/sv2v_out.v:11308.6-11308.16" */
wire cmp_signed;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11308.6-11308.16" */
wire cmp_signed_t0;
/* src = "generated/sv2v_out.v:11251.14-11251.33" */
output comparison_result_o;
wire comparison_result_o;
/* cellift = 32'd1 */
output comparison_result_o_t0;
wire comparison_result_o_t0;
/* src = "generated/sv2v_out.v:11246.20-11246.31" */
output [63:0] imd_val_d_o;
wire [63:0] imd_val_d_o;
/* cellift = 32'd1 */
output [63:0] imd_val_d_o_t0;
wire [63:0] imd_val_d_o_t0;
/* src = "generated/sv2v_out.v:11245.20-11245.31" */
input [63:0] imd_val_q_i;
wire [63:0] imd_val_q_i;
/* cellift = 32'd1 */
input [63:0] imd_val_q_i_t0;
wire [63:0] imd_val_q_i_t0;
/* src = "generated/sv2v_out.v:11247.19-11247.31" */
output [1:0] imd_val_we_o;
wire [1:0] imd_val_we_o;
/* cellift = 32'd1 */
output [1:0] imd_val_we_o_t0;
wire [1:0] imd_val_we_o_t0;
/* src = "generated/sv2v_out.v:11241.13-11241.32" */
input instr_first_cycle_i;
wire instr_first_cycle_i;
/* cellift = 32'd1 */
input instr_first_cycle_i_t0;
wire instr_first_cycle_i_t0;
/* src = "generated/sv2v_out.v:11252.14-11252.31" */
output is_equal_result_o;
wire is_equal_result_o;
/* cellift = 32'd1 */
output is_equal_result_o_t0;
wire is_equal_result_o_t0;
/* src = "generated/sv2v_out.v:11307.6-11307.22" */
wire is_greater_equal;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11307.6-11307.22" */
wire is_greater_equal_t0;
/* src = "generated/sv2v_out.v:11242.20-11242.39" */
input [32:0] multdiv_operand_a_i;
wire [32:0] multdiv_operand_a_i;
/* cellift = 32'd1 */
input [32:0] multdiv_operand_a_i_t0;
wire [32:0] multdiv_operand_a_i_t0;
/* src = "generated/sv2v_out.v:11243.20-11243.39" */
input [32:0] multdiv_operand_b_i;
wire [32:0] multdiv_operand_b_i;
/* cellift = 32'd1 */
input [32:0] multdiv_operand_b_i_t0;
wire [32:0] multdiv_operand_b_i_t0;
/* src = "generated/sv2v_out.v:11244.13-11244.26" */
input multdiv_sel_i;
wire multdiv_sel_i;
/* cellift = 32'd1 */
input multdiv_sel_i_t0;
wire multdiv_sel_i_t0;
/* src = "generated/sv2v_out.v:11239.20-11239.31" */
input [31:0] operand_a_i;
wire [31:0] operand_a_i;
/* cellift = 32'd1 */
input [31:0] operand_a_i_t0;
wire [31:0] operand_a_i_t0;
/* src = "generated/sv2v_out.v:11240.20-11240.31" */
input [31:0] operand_b_i;
wire [31:0] operand_b_i;
/* cellift = 32'd1 */
input [31:0] operand_b_i_t0;
wire [31:0] operand_b_i_t0;
/* src = "generated/sv2v_out.v:11254.14-11254.27" */
wire [32:0] operand_b_neg;
/* src = "generated/sv2v_out.v:11238.19-11238.29" */
input [6:0] operator_i;
wire [6:0] operator_i;
/* cellift = 32'd1 */
input [6:0] operator_i_t0;
wire [6:0] operator_i_t0;
/* src = "generated/sv2v_out.v:11250.20-11250.28" */
output [31:0] result_o;
wire [31:0] result_o;
/* cellift = 32'd1 */
output [31:0] result_o_t0;
wire [31:0] result_o_t0;
/* src = "generated/sv2v_out.v:11336.12-11336.21" */
wire [5:0] shift_amt;
/* src = "generated/sv2v_out.v:11337.13-11337.28" */
/* unused_bits = "5" */
wire [5:0] shift_amt_compl;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11337.13-11337.28" */
/* unused_bits = "5" */
wire [5:0] shift_amt_compl_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11336.12-11336.21" */
wire [5:0] shift_amt_t0;
/* src = "generated/sv2v_out.v:11333.7-11333.18" */
wire shift_arith;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11333.7-11333.18" */
wire shift_arith_t0;
/* src = "generated/sv2v_out.v:11331.6-11331.16" */
wire shift_left;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11331.6-11331.16" */
wire shift_left_t0;
/* src = "generated/sv2v_out.v:11338.13-11338.26" */
wire [31:0] shift_operand;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11338.13-11338.26" */
wire [31:0] shift_operand_t0;
/* src = "generated/sv2v_out.v:11342.13-11342.25" */
wire [31:0] shift_result;
/* src = "generated/sv2v_out.v:11340.13-11340.29" */
/* unused_bits = "32" */
wire [32:0] shift_result_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11340.13-11340.29" */
/* unused_bits = "32" */
wire [32:0] shift_result_ext_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:11342.13-11342.25" */
wire [31:0] shift_result_t0;
assign adder_result_ext_o = { 1'h0, adder_in_a } + /* src = "generated/sv2v_out.v:11303.30-11303.75" */ { 1'h0, adder_in_b };
assign _0000_ = shift_arith & /* src = "generated/sv2v_out.v:11397.52-11397.83" */ shift_operand[31];
assign bwlogic_and_result = operand_a_i & /* src = "generated/sv2v_out.v:11424.30-11424.61" */ operand_b_i;
assign _0002_ = ~ { 1'h0, adder_in_a_t0 };
assign _0003_ = ~ { 1'h0, adder_in_b_t0 };
assign _0065_ = { 1'h0, adder_in_a } & _0002_;
assign _0066_ = { 1'h0, adder_in_b } & _0003_;
assign _0370_ = _0065_ + _0066_;
assign _0183_ = { 1'h0, adder_in_a } | { 1'h0, adder_in_a_t0 };
assign _0184_ = { 1'h0, adder_in_b } | { 1'h0, adder_in_b_t0 };
assign _0371_ = _0183_ + _0184_;
assign _0255_ = _0370_ ^ _0371_;
assign _0185_ = _0255_ | { 1'h0, adder_in_a_t0 };
assign adder_result_ext_o_t0 = _0185_ | { 1'h0, adder_in_b_t0 };
assign _0067_ = shift_arith_t0 & shift_operand[31];
assign _0070_ = operand_a_i_t0 & operand_b_i;
assign _0068_ = shift_operand_t0[31] & shift_arith;
assign _0071_ = operand_b_i_t0 & operand_a_i;
assign _0069_ = shift_arith_t0 & shift_operand_t0[31];
assign _0072_ = operand_a_i_t0 & operand_b_i_t0;
assign _0186_ = _0067_ | _0068_;
assign _0187_ = _0070_ | _0071_;
assign _0001_ = _0186_ | _0069_;
assign bwlogic_and_result_t0 = _0187_ | _0072_;
assign _0005_ = ~ operator_i_t0;
assign _0139_ = operator_i & _0005_;
assign _0284_ = _0139_ == { 2'h0, _0005_[4:2], 1'h0, _0005_[0] };
assign _0285_ = _0139_ == { 3'h0, _0005_[3], 2'h0, _0005_[0] };
assign _0286_ = _0139_ == { 3'h0, _0005_[3], 3'h0 };
assign _0287_ = _0139_ == { 3'h0, _0005_[3:2], 2'h0 };
assign _0288_ = _0139_ == { 3'h0, _0005_[3], 1'h0, _0005_[1:0] };
assign _0289_ = _0139_ == { 6'h00, _0005_[0] };
assign _0290_ = _0139_ == { 2'h0, _0005_[4], 1'h0, _0005_[2:1], 1'h0 };
assign _0291_ = _0139_ == { 2'h0, _0005_[4], 1'h0, _0005_[2:0] };
assign _0292_ = _0139_ == { 2'h0, _0005_[4:3], 3'h0 };
assign _0293_ = _0139_ == { 5'h00, _0005_[1], 1'h0 };
assign _0294_ = _0139_ == { 4'h0, _0005_[2], 1'h0, _0005_[0] };
assign _0295_ = _0139_ == { 5'h00, _0005_[1:0] };
assign _0296_ = _0139_ == { 4'h0, _0005_[2:1], 1'h0 };
assign _0297_ = _0139_ == { 4'h0, _0005_[2], 2'h0 };
assign _0298_ = _0139_ == { 4'h0, _0005_[2:0] };
assign _0299_ = _0139_ == { 3'h0, _0005_[3], 1'h0, _0005_[1], 1'h0 };
assign _0300_ = _0139_ == { 2'h0, _0005_[4:3], 2'h0, _0005_[0] };
assign _0301_ = _0139_ == { 2'h0, _0005_[4:3], 1'h0, _0005_[1], 1'h0 };
assign _0302_ = _0139_ == { 2'h0, _0005_[4:0] };
assign _0303_ = _0139_ == { 1'h0, _0005_[5], 5'h00 };
assign _0304_ = _0139_ == { 1'h0, _0005_[5], 1'h0, _0005_[3], 1'h0, _0005_[1:0] };
assign _0305_ = _0139_ == { 1'h0, _0005_[5], 1'h0, _0005_[3:2], 2'h0 };
assign _0306_ = _0139_ == { 2'h0, _0005_[4:2], 2'h0 };
assign _0307_ = _0139_ == { 1'h0, _0005_[5], 4'h0, _0005_[0] };
assign _0308_ = _0139_ == { 1'h0, _0005_[5], 3'h0, _0005_[1], 1'h0 };
assign _0309_ = _0139_ == { 2'h0, _0005_[4:1], 1'h0 };
assign _0310_ = _0139_ == { 2'h0, _0005_[4:3], 1'h0, _0005_[1:0] };
assign _0421_[0] = _0284_ & _0004_;
assign _0425_[1] = _0285_ & _0004_;
assign shift_arith_t0 = _0286_ & _0004_;
assign _0425_[3] = _0287_ & _0004_;
assign _0425_[4] = _0288_ & _0004_;
assign _0429_[1] = _0289_ & _0004_;
assign _0429_[2] = _0290_ & _0004_;
assign _0429_[3] = _0291_ & _0004_;
assign _0429_[4] = _0292_ & _0004_;
assign _0433_[0] = _0293_ & _0004_;
assign _0433_[1] = _0294_ & _0004_;
assign _0388_ = _0295_ & _0004_;
assign _0390_ = _0296_ & _0004_;
assign _0392_ = _0297_ & _0004_;
assign _0394_ = _0298_ & _0004_;
assign shift_left_t0 = _0299_ & _0004_;
assign _0421_[4] = _0300_ & _0004_;
assign _0421_[5] = _0301_ & _0004_;
assign _0439_[2] = _0302_ & _0004_;
assign _0439_[3] = _0303_ & _0004_;
assign _0421_[6] = _0304_ & _0004_;
assign _0421_[7] = _0305_ & _0004_;
assign _0421_[3] = _0306_ & _0004_;
assign _0443_[2] = _0307_ & _0004_;
assign _0443_[3] = _0308_ & _0004_;
assign _0421_[1] = _0309_ & _0004_;
assign _0421_[2] = _0310_ & _0004_;
assign _0006_ = | adder_result_ext_o_t0[32:1];
assign _0007_ = | _0421_;
assign _0008_ = | { shift_left_t0, _0425_[4:3], _0425_[1], shift_arith_t0 };
assign _0009_ = | _0429_;
assign _0004_ = | operator_i_t0;
assign _0010_ = | { _0433_[1:0], _0394_, _0392_, _0390_, _0388_ };
assign _0011_ = | { _0439_[3:2], _0421_[7:4] };
assign _0012_ = | { _0443_[3:2], _0421_[3:2] };
assign _0013_ = | { _0443_[2], _0439_[2], _0421_[6], _0421_[4], _0421_[2] };
assign _0014_ = ~ adder_result_ext_o_t0[32:1];
assign _0015_ = ~ _0421_;
assign _0016_ = ~ { _0425_[4:3], _0425_[1], shift_left_t0, shift_arith_t0 };
assign _0017_ = ~ _0429_;
assign _0018_ = ~ { _0433_[1:0], _0394_, _0392_, _0390_, _0388_ };
assign _0019_ = ~ { _0439_[3:2], _0421_[7:4] };
assign _0020_ = ~ { _0443_[3:2], _0421_[3:2] };
assign _0021_ = ~ { _0443_[2], _0439_[2], _0421_[6], _0421_[4], _0421_[2] };
assign _0099_ = adder_result_ext_o[32:1] & _0014_;
assign _0138_ = _0420_ & _0015_;
assign _0140_ = { _0424_[4:3], _0424_[1:0], shift_arith } & _0016_;
assign _0141_ = _0428_ & _0017_;
assign _0142_ = { _0432_[1:0], _0393_, _0391_, _0389_, _0387_ } & _0018_;
assign _0149_ = { _0438_[3:2], _0420_[7:4] } & _0019_;
assign _0150_ = { _0442_[3:2], _0420_[3:2] } & _0020_;
assign _0154_ = { _0442_[2], _0438_[2], _0420_[6], _0420_[4], _0420_[2] } & _0021_;
assign _0022_ = ! _0099_;
assign _0023_ = ! _0138_;
assign _0024_ = ! _0140_;
assign _0025_ = ! _0141_;
assign _0026_ = ! _0139_;
assign _0027_ = ! _0142_;
assign _0028_ = ! _0149_;
assign _0029_ = ! _0150_;
assign _0030_ = ! _0154_;
assign is_equal_result_o_t0 = _0022_ & _0006_;
assign _0423_ = _0023_ & _0007_;
assign _0427_ = _0024_ & _0008_;
assign _0431_ = _0025_ & _0009_;
assign _0429_[0] = _0026_ & _0004_;
assign _0435_ = _0027_ & _0010_;
assign _0441_ = _0028_ & _0011_;
assign _0445_ = _0029_ & _0012_;
assign cmp_signed_t0 = _0030_ & _0013_;
assign _0031_ = ~ { _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_ };
assign _0032_ = ~ { _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_ };
assign _0033_ = ~ { _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_ };
assign _0034_ = ~ _0440_;
assign _0035_ = ~ _0420_[1];
assign _0036_ = ~ _0181_;
assign _0037_ = ~ operator_i[5];
assign _0038_ = ~ operator_i[4];
assign _0039_ = ~ operator_i[3];
assign _0040_ = ~ operator_i[2];
assign _0041_ = ~ operator_i[1];
assign _0042_ = ~ { bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and };
assign _0043_ = ~ { bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or };
assign _0044_ = ~ _0451_;
assign _0045_ = ~ { adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate };
assign _0046_ = ~ { multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i };
assign _0047_ = ~ operator_i[6];
assign _0048_ = ~ { instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i };
assign _0049_ = ~ { shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left };
assign _0190_ = { _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_ } | _0031_;
assign _0194_ = { _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_ } | _0032_;
assign _0197_ = { _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_ } | _0033_;
assign _0200_ = _0441_ | _0034_;
assign _0203_ = _0421_[1] | _0035_;
assign _0206_ = _0182_ | _0036_;
assign _0209_ = operator_i_t0[5] | _0037_;
assign _0212_ = operator_i_t0[4] | _0038_;
assign _0215_ = operator_i_t0[3] | _0039_;
assign _0218_ = operator_i_t0[2] | _0040_;
assign _0221_ = operator_i_t0[1] | _0041_;
assign _0226_ = { bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0 } | _0042_;
assign _0229_ = { bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0 } | _0043_;
assign _0232_ = _0452_ | _0044_;
assign _0235_ = { adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0 } | _0045_;
assign _0238_ = { multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0 } | _0046_;
assign _0242_ = operator_i_t0[6] | _0047_;
assign _0248_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0 } | _0048_;
assign _0251_ = { shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0 } | _0049_;
assign _0191_ = { _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_ } | { _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_, _0422_ };
assign _0193_ = { _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_ } | { _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_, _0434_ };
assign _0195_ = { _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_ } | { _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_, _0430_ };
assign _0198_ = { _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_ } | { _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_, _0179_ };
assign _0201_ = _0441_ | _0440_;
assign _0204_ = _0421_[1] | _0420_[1];
assign _0207_ = _0182_ | _0181_;
assign _0210_ = operator_i_t0[5] | operator_i[5];
assign _0213_ = operator_i_t0[4] | operator_i[4];
assign _0216_ = operator_i_t0[3] | operator_i[3];
assign _0219_ = operator_i_t0[2] | operator_i[2];
assign _0222_ = operator_i_t0[1] | operator_i[1];
assign _0227_ = { bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0 } | { bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and, bwlogic_and };
assign _0230_ = { bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0 } | { bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or, bwlogic_or };
assign _0233_ = _0452_ | _0451_;
assign _0236_ = { adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0 } | { adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate, adder_op_b_negate };
assign _0239_ = { multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0 } | { multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i, multdiv_sel_i };
assign _0249_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0 } | { instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i, instr_first_cycle_i };
assign _0252_ = { shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0 } | { shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left, shift_left };
assign _0079_ = shift_result_t0 & _0190_;
assign _0084_ = _0377_ & _0194_;
assign _0087_ = _0379_ & _0197_;
assign _0090_ = is_greater_equal_t0 & _0200_;
assign _0093_ = is_equal_result_o_t0 & _0203_;
assign _0096_ = _0383_ & _0206_;
assign _0100_ = _0396_ & _0209_;
assign _0103_ = _0400_ & _0212_;
assign _0106_ = _0403_ & _0212_;
assign _0108_ = _0404_ & _0215_;
assign _0112_ = _0407_ & _0215_;
assign _0115_ = _0410_ & _0218_;
assign _0117_ = _0412_ & _0218_;
assign _0119_ = _0413_ & _0218_;
assign _0121_ = _0415_ & _0218_;
assign _0124_ = operator_i_t0[0] & _0221_;
assign _0143_ = bwlogic_xor_result_t0 & _0226_;
assign _0146_ = _0437_ & _0229_;
assign _0151_ = adder_result_ext_o_t0[32] & _0232_;
assign _0155_ = { operand_b_i_t0, 1'h0 } & _0235_;
assign _0158_ = _0448_ & _0238_;
assign _0161_ = { operand_a_i_t0, 1'h0 } & _0238_;
assign _0164_ = _0064_ & _0242_;
assign _0170_ = shift_amt_compl_t0[4:0] & _0248_;
assign _0173_ = operand_a_i_t0 & _0251_;
assign _0176_ = shift_result_ext_t0[31:0] & _0251_;
assign _0080_ = { 31'h00000000, comparison_result_o_t0 } & _0191_;
assign _0082_ = bwlogic_result_t0 & _0193_;
assign _0085_ = adder_result_ext_o_t0[32:1] & _0195_;
assign _0088_ = _0375_ & _0198_;
assign _0091_ = is_greater_equal_t0 & _0201_;
assign _0094_ = is_equal_result_o_t0 & _0204_;
assign _0097_ = _0381_ & _0207_;
assign _0101_ = _0398_ & _0210_;
assign _0104_ = _0402_ & _0213_;
assign _0110_ = _0405_ & _0216_;
assign _0113_ = _0409_ & _0216_;
assign _0122_ = _0417_ & _0219_;
assign _0126_ = operator_i_t0[0] & _0222_;
assign _0144_ = bwlogic_and_result_t0 & _0227_;
assign _0147_ = bwlogic_or_result_t0 & _0230_;
assign _0152_ = _0454_ & _0233_;
assign _0156_ = { operand_b_i_t0, 1'h0 } & _0236_;
assign _0159_ = multdiv_operand_b_i_t0 & _0239_;
assign _0162_ = multdiv_operand_a_i_t0 & _0239_;
assign _0171_ = operand_b_i_t0[4:0] & _0249_;
assign _0174_ = { operand_a_i_t0[0], operand_a_i_t0[1], operand_a_i_t0[2], operand_a_i_t0[3], operand_a_i_t0[4], operand_a_i_t0[5], operand_a_i_t0[6], operand_a_i_t0[7], operand_a_i_t0[8], operand_a_i_t0[9], operand_a_i_t0[10], operand_a_i_t0[11], operand_a_i_t0[12], operand_a_i_t0[13], operand_a_i_t0[14], operand_a_i_t0[15], operand_a_i_t0[16], operand_a_i_t0[17], operand_a_i_t0[18], operand_a_i_t0[19], operand_a_i_t0[20], operand_a_i_t0[21], operand_a_i_t0[22], operand_a_i_t0[23], operand_a_i_t0[24], operand_a_i_t0[25], operand_a_i_t0[26], operand_a_i_t0[27], operand_a_i_t0[28], operand_a_i_t0[29], operand_a_i_t0[30], operand_a_i_t0[31] } & _0252_;
assign _0177_ = { shift_result_ext_t0[0], shift_result_ext_t0[1], shift_result_ext_t0[2], shift_result_ext_t0[3], shift_result_ext_t0[4], shift_result_ext_t0[5], shift_result_ext_t0[6], shift_result_ext_t0[7], shift_result_ext_t0[8], shift_result_ext_t0[9], shift_result_ext_t0[10], shift_result_ext_t0[11], shift_result_ext_t0[12], shift_result_ext_t0[13], shift_result_ext_t0[14], shift_result_ext_t0[15], shift_result_ext_t0[16], shift_result_ext_t0[17], shift_result_ext_t0[18], shift_result_ext_t0[19], shift_result_ext_t0[20], shift_result_ext_t0[21], shift_result_ext_t0[22], shift_result_ext_t0[23], shift_result_ext_t0[24], shift_result_ext_t0[25], shift_result_ext_t0[26], shift_result_ext_t0[27], shift_result_ext_t0[28], shift_result_ext_t0[29], shift_result_ext_t0[30], shift_result_ext_t0[31] } & _0252_;
assign _0192_ = _0079_ | _0080_;
assign _0196_ = _0084_ | _0085_;
assign _0199_ = _0087_ | _0088_;
assign _0202_ = _0090_ | _0091_;
assign _0205_ = _0093_ | _0094_;
assign _0208_ = _0096_ | _0097_;
assign _0211_ = _0100_ | _0101_;
assign _0214_ = _0103_ | _0104_;
assign _0217_ = _0112_ | _0113_;
assign _0220_ = _0121_ | _0122_;
assign _0228_ = _0143_ | _0144_;
assign _0231_ = _0146_ | _0147_;
assign _0234_ = _0151_ | _0152_;
assign _0237_ = _0155_ | _0156_;
assign _0240_ = _0158_ | _0159_;
assign _0241_ = _0161_ | _0162_;
assign _0250_ = _0170_ | _0171_;
assign _0253_ = _0173_ | _0174_;
assign _0254_ = _0176_ | _0177_;
assign _0256_ = shift_result ^ { 31'h00000000, comparison_result_o };
assign _0257_ = _0376_ ^ adder_result_ext_o[32:1];
assign _0258_ = _0378_ ^ _0374_;
assign _0259_ = is_greater_equal ^ _0419_;
assign _0260_ = is_equal_result_o ^ _0418_;
assign _0261_ = _0382_ ^ _0380_;
assign _0262_ = _0395_ ^ _0397_;
assign _0263_ = _0399_ ^ _0401_;
assign _0267_ = _0406_ ^ _0408_;
assign _0270_ = _0414_ ^ _0416_;
assign _0273_ = bwlogic_xor_result ^ bwlogic_and_result;
assign _0274_ = _0436_ ^ bwlogic_or_result;
assign _0275_ = _0386_ ^ _0453_;
assign _0276_ = { operand_b_i, 1'h0 } ^ operand_b_neg;
assign _0277_ = _0447_ ^ multdiv_operand_b_i;
assign _0278_ = { operand_a_i, 1'h1 } ^ multdiv_operand_a_i;
assign _0281_ = shift_amt_compl[4:0] ^ operand_b_i[4:0];
assign _0282_ = operand_a_i ^ { operand_a_i[0], operand_a_i[1], operand_a_i[2], operand_a_i[3], operand_a_i[4], operand_a_i[5], operand_a_i[6], operand_a_i[7], operand_a_i[8], operand_a_i[9], operand_a_i[10], operand_a_i[11], operand_a_i[12], operand_a_i[13], operand_a_i[14], operand_a_i[15], operand_a_i[16], operand_a_i[17], operand_a_i[18], operand_a_i[19], operand_a_i[20], operand_a_i[21], operand_a_i[22], operand_a_i[23], operand_a_i[24], operand_a_i[25], operand_a_i[26], operand_a_i[27], operand_a_i[28], operand_a_i[29], operand_a_i[30], operand_a_i[31] };
assign _0283_ = shift_result_ext[31:0] ^ { shift_result_ext[0], shift_result_ext[1], shift_result_ext[2], shift_result_ext[3], shift_result_ext[4], shift_result_ext[5], shift_result_ext[6], shift_result_ext[7], shift_result_ext[8], shift_result_ext[9], shift_result_ext[10], shift_result_ext[11], shift_result_ext[12], shift_result_ext[13], shift_result_ext[14], shift_result_ext[15], shift_result_ext[16], shift_result_ext[17], shift_result_ext[18], shift_result_ext[19], shift_result_ext[20], shift_result_ext[21], shift_result_ext[22], shift_result_ext[23], shift_result_ext[24], shift_result_ext[25], shift_result_ext[26], shift_result_ext[27], shift_result_ext[28], shift_result_ext[29], shift_result_ext[30], shift_result_ext[31] };
assign _0081_ = { _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_, _0423_ } & _0256_;
assign _0083_ = { _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_, _0435_ } & bwlogic_result;
assign _0086_ = { _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_, _0431_ } & _0257_;
assign _0089_ = { _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_, _0180_ } & _0258_;
assign _0092_ = _0441_ & _0259_;
assign _0095_ = _0421_[1] & _0260_;
assign _0098_ = _0182_ & _0261_;
assign _0102_ = operator_i_t0[5] & _0262_;
assign _0105_ = operator_i_t0[4] & _0263_;
assign _0107_ = operator_i_t0[4] & _0264_;
assign _0109_ = operator_i_t0[3] & _0265_;
assign _0111_ = operator_i_t0[3] & _0266_;
assign _0114_ = operator_i_t0[3] & _0267_;
assign _0116_ = operator_i_t0[2] & _0268_;
assign _0118_ = operator_i_t0[2] & _0051_;
assign _0120_ = operator_i_t0[2] & _0269_;
assign _0123_ = operator_i_t0[2] & _0270_;
assign _0125_ = operator_i_t0[1] & _0271_;
assign _0127_ = operator_i_t0[1] & _0272_;
assign _0128_ = operator_i_t0[1] & _0050_;
assign _0129_ = operator_i_t0[1] & operator_i[0];
assign _0145_ = { bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0, bwlogic_and_t0 } & _0273_;
assign _0148_ = { bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0, bwlogic_or_t0 } & _0274_;
assign _0153_ = _0452_ & _0275_;
assign _0157_ = { adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0, adder_op_b_negate_t0 } & _0276_;
assign _0160_ = { multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0 } & _0277_;
assign _0163_ = { multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0, multdiv_sel_i_t0 } & _0278_;
assign _0165_ = operator_i_t0[6] & _0063_;
assign _0172_ = { instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0, instr_first_cycle_i_t0 } & _0281_;
assign _0175_ = { shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0 } & _0282_;
assign _0178_ = { shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0, shift_left_t0 } & _0283_;
assign _0375_ = _0081_ | _0192_;
assign _0377_ = _0083_ | _0082_;
assign _0379_ = _0086_ | _0196_;
assign result_o_t0 = _0089_ | _0199_;
assign _0381_ = _0092_ | _0202_;
assign _0383_ = _0095_ | _0205_;
assign comparison_result_o_t0 = _0098_ | _0208_;
assign _0064_ = _0102_ | _0211_;
assign _0396_ = _0105_ | _0214_;
assign _0398_ = _0107_ | _0106_;
assign _0400_ = _0109_ | _0108_;
assign _0402_ = _0111_ | _0110_;
assign _0403_ = _0114_ | _0217_;
assign _0404_ = _0116_ | _0115_;
assign _0405_ = _0118_ | _0117_;
assign _0407_ = _0120_ | _0119_;
assign _0409_ = _0123_ | _0220_;
assign _0410_ = _0125_ | _0124_;
assign _0415_ = _0125_ | _0126_;
assign _0417_ = _0127_ | _0124_;
assign _0412_ = _0128_ | _0124_;
assign _0413_ = _0129_ | _0126_;
assign _0437_ = _0145_ | _0228_;
assign bwlogic_result_t0 = _0148_ | _0231_;
assign is_greater_equal_t0 = _0153_ | _0234_;
assign _0448_ = _0157_ | _0237_;
assign adder_in_b_t0 = _0160_ | _0240_;
assign adder_in_a_t0 = _0163_ | _0241_;
assign adder_op_b_negate_t0 = _0165_ | _0164_;
assign shift_amt_t0[4:0] = _0172_ | _0250_;
assign shift_operand_t0 = _0175_ | _0253_;
assign shift_result_t0 = _0178_ | _0254_;
assign _0050_ = ~ _0271_;
assign _0051_ = ~ _0411_;
assign operand_b_neg = ~ { operand_b_i, 1'h0 };
assign _0052_ = ~ _0426_;
assign _0053_ = ~ _0444_;
assign _0054_ = ~ operand_a_i;
assign _0055_ = ~ _0387_;
assign _0056_ = ~ _0391_;
assign _0057_ = ~ _0422_;
assign _0058_ = ~ operand_b_i;
assign _0059_ = ~ _0389_;
assign _0060_ = ~ _0393_;
assign _0073_ = _0427_ & _0057_;
assign _0076_ = _0445_ & _0034_;
assign _0130_ = operand_a_i_t0 & _0058_;
assign _0132_ = _0388_ & _0059_;
assign _0135_ = _0392_ & _0060_;
assign _0074_ = _0423_ & _0052_;
assign _0077_ = _0441_ & _0053_;
assign _0131_ = operand_b_i_t0 & _0054_;
assign _0133_ = _0390_ & _0055_;
assign _0136_ = _0394_ & _0056_;
assign _0075_ = _0427_ & _0423_;
assign _0078_ = _0445_ & _0441_;
assign _0134_ = _0388_ & _0390_;
assign _0137_ = _0392_ & _0394_;
assign _0188_ = _0073_ | _0074_;
assign _0189_ = _0076_ | _0077_;
assign _0223_ = _0130_ | _0131_;
assign _0224_ = _0132_ | _0133_;
assign _0225_ = _0135_ | _0136_;
assign _0180_ = _0188_ | _0075_;
assign _0182_ = _0189_ | _0078_;
assign bwlogic_or_result_t0 = _0223_ | _0072_;
assign bwlogic_or_t0 = _0224_ | _0134_;
assign bwlogic_and_t0 = _0225_ | _0137_;
assign _0179_ = _0426_ | _0422_;
assign _0181_ = _0444_ | _0440_;
assign _0374_ = _0422_ ? { 31'h00000000, comparison_result_o } : shift_result;
assign _0376_ = _0434_ ? bwlogic_result : 32'd0;
assign _0378_ = _0430_ ? adder_result_ext_o[32:1] : _0376_;
assign result_o = _0179_ ? _0374_ : _0378_;
assign _0380_ = _0440_ ? _0419_ : is_greater_equal;
assign _0382_ = _0420_[1] ? _0418_ : is_equal_result_o;
assign comparison_result_o = _0181_ ? _0380_ : _0382_;
assign _0311_ = shift_amt_t0[1:0] == 2'h3;
assign _0312_ = { shift_amt_t0[2], shift_amt_t0[0] } == 2'h3;
assign _0313_ = shift_amt_t0[2:1] == 2'h3;
assign _0314_ = shift_amt_t0[2:0] == 3'h7;
assign _0315_ = { shift_amt_t0[3], shift_amt_t0[0] } == 2'h3;
assign _0316_ = { shift_amt_t0[3], shift_amt_t0[1] } == 2'h3;
assign _0317_ = { shift_amt_t0[3], shift_amt_t0[1:0] } == 3'h7;
assign _0318_ = shift_amt_t0[3:2] == 2'h3;
assign _0319_ = { shift_amt_t0[3:2], shift_amt_t0[0] } == 3'h7;
assign _0320_ = shift_amt_t0[3:1] == 3'h7;
assign _0321_ = shift_amt_t0[3:0] == 4'hf;
assign _0322_ = { shift_amt_t0[4], shift_amt_t0[0] } == 2'h3;
assign _0323_ = { shift_amt_t0[4], shift_amt_t0[1] } == 2'h3;
assign _0324_ = { shift_amt_t0[4], shift_amt_t0[1:0] } == 3'h7;
assign _0325_ = { shift_amt_t0[4], shift_amt_t0[2] } == 2'h3;
assign _0326_ = { shift_amt_t0[4], shift_amt_t0[2], shift_amt_t0[0] } == 3'h7;
assign _0327_ = { shift_amt_t0[4], shift_amt_t0[2:1] } == 3'h7;
assign _0328_ = { shift_amt_t0[4], shift_amt_t0[2:0] } == 4'hf;
assign _0329_ = shift_amt_t0[4:3] == 2'h3;
assign _0330_ = { shift_amt_t0[4:3], shift_amt_t0[0] } == 3'h7;
assign _0331_ = { shift_amt_t0[4:3], shift_amt_t0[1] } == 3'h7;
assign _0332_ = { shift_amt_t0[4:3], shift_amt_t0[1:0] } == 4'hf;
assign _0333_ = shift_amt_t0[4:2] == 3'h7;
assign _0334_ = { shift_amt_t0[4:2], shift_amt_t0[0] } == 4'hf;
assign _0335_ = shift_amt_t0[4:1] == 4'hf;
assign _0336_ = shift_amt_t0[4:0] == 5'h1f;
assign _0279_ = { _0384_[31:30], _0384_[30:29], _0384_[29], _0384_[29:28], _0384_[28], _0384_[28], _0384_[28:27], _0384_[27], _0384_[27], _0384_[27], _0384_[27:26], _0384_[26], _0384_[26], _0384_[26], _0384_[26], _0384_[26:25], _0384_[25], _0384_[25], _0384_[25], _0384_[25], _0384_[25], _0384_[25:24], _0384_[24], _0384_[24], _0384_[24], _0384_[24], _0384_[24], _0384_[24], _0384_[24:23], _0384_[23], _0384_[23], _0384_[23], _0384_[23], _0384_[23], _0384_[23], _0384_[23], _0384_[23:22], _0384_[22], _0384_[22], _0384_[22], _0384_[22], _0384_[22], _0384_[22], _0384_[22], _0384_[22], _0384_[22:21], _0384_[21], _0384_[21], _0384_[21], _0384_[21], _0384_[21], _0384_[21], _0384_[21], _0384_[21], _0384_[21], _0384_[21:20], _0384_[20], _0384_[20], _0384_[20], _0384_[20], _0384_[20], _0384_[20], _0384_[20], _0384_[20], _0384_[20], _0384_[20], _0384_[20:19], _0384_[19], _0384_[19], _0384_[19], _0384_[19], _0384_[19], _0384_[19], _0384_[19], _0384_[19], _0384_[19], _0384_[19], _0384_[19], _0384_[19:18], _0384_[18], _0384_[18], _0384_[18], _0384_[18], _0384_[18], _0384_[18], _0384_[18], _0384_[18], _0384_[18], _0384_[18], _0384_[18], _0384_[18], _0384_[18:17], _0384_[17], _0384_[17], _0384_[17], _0384_[17], _0384_[17], _0384_[17], _0384_[17], _0384_[17], _0384_[17], _0384_[17], _0384_[17], _0384_[17], _0384_[17], _0384_[17:16], _0384_[16], _0384_[16], _0384_[16], _0384_[16], _0384_[16], _0384_[16], _0384_[16], _0384_[16], _0384_[16], _0384_[16], _0384_[16], _0384_[16], _0384_[16], _0384_[16], _0384_[16:15], _0384_[15], _0384_[15], _0384_[15], _0384_[15], _0384_[15], _0384_[15], _0384_[15], _0384_[15], _0384_[15], _0384_[15], _0384_[15], _0384_[15], _0384_[15], _0384_[15], _0384_[15], _0384_[15:14], _0384_[14], _0384_[14], _0384_[14], _0384_[14], _0384_[14], _0384_[14], _0384_[14], _0384_[14], _0384_[14], _0384_[14], _0384_[14], _0384_[14], _0384_[14], _0384_[14], _0384_[14], _0384_[14], _0384_[14:13], _0384_[13], _0384_[13], _0384_[13], _0384_[13], _0384_[13], _0384_[13], _0384_[13], _0384_[13], _0384_[13], _0384_[13], _0384_[13], _0384_[13], _0384_[13], _0384_[13], _0384_[13], _0384_[13], _0384_[13], _0384_[13:12], _0384_[12], _0384_[12], _0384_[12], _0384_[12], _0384_[12], _0384_[12], _0384_[12], _0384_[12], _0384_[12], _0384_[12], _0384_[12], _0384_[12], _0384_[12], _0384_[12], _0384_[12], _0384_[12], _0384_[12], _0384_[12], _0384_[12:11], _0384_[11], _0384_[11], _0384_[11], _0384_[11], _0384_[11], _0384_[11], _0384_[11], _0384_[11], _0384_[11], _0384_[11], _0384_[11], _0384_[11], _0384_[11], _0384_[11], _0384_[11], _0384_[11], _0384_[11], _0384_[11], _0384_[11], _0384_[11:10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10], _0384_[10:9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9], _0384_[9:8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8], _0384_[8:7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7], _0384_[7:6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6], _0384_[6:5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5], _0384_[5:4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4], _0384_[4:3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3], _0384_[3:2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2], _0384_[2:1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1], _0384_[1:0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0], _0384_[0] } ^ { _0384_[32], _0384_[32:31], _0384_[32:30], _0384_[32:29], _0384_[32:28], _0384_[32:27], _0384_[32:26], _0384_[32:25], _0384_[32:24], _0384_[32:23], _0384_[32:22], _0384_[32:21], _0384_[32:20], _0384_[32:19], _0384_[32:18], _0384_[32:17], _0384_[32:16], _0384_[32:15], _0384_[32:14], _0384_[32:13], _0384_[32:12], _0384_[32:11], _0384_[32:10], _0384_[32:9], _0384_[32:8], _0384_[32:7], _0384_[32:6], _0384_[32:5], _0384_[32:4], _0384_[32:3], _0384_[32:2], _0384_[32:1] };
assign _0243_ = { _0385_[31:30], _0385_[30:29], _0385_[29], _0385_[29:28], _0385_[28], _0385_[28], _0385_[28:27], _0385_[27], _0385_[27], _0385_[27], _0385_[27:26], _0385_[26], _0385_[26], _0385_[26], _0385_[26], _0385_[26:25], _0385_[25], _0385_[25], _0385_[25], _0385_[25], _0385_[25], _0385_[25:24], _0385_[24], _0385_[24], _0385_[24], _0385_[24], _0385_[24], _0385_[24], _0385_[24:23], _0385_[23], _0385_[23], _0385_[23], _0385_[23], _0385_[23], _0385_[23], _0385_[23], _0385_[23:22], _0385_[22], _0385_[22], _0385_[22], _0385_[22], _0385_[22], _0385_[22], _0385_[22], _0385_[22], _0385_[22:21], _0385_[21], _0385_[21], _0385_[21], _0385_[21], _0385_[21], _0385_[21], _0385_[21], _0385_[21], _0385_[21], _0385_[21:20], _0385_[20], _0385_[20], _0385_[20], _0385_[20], _0385_[20], _0385_[20], _0385_[20], _0385_[20], _0385_[20], _0385_[20], _0385_[20:19], _0385_[19], _0385_[19], _0385_[19], _0385_[19], _0385_[19], _0385_[19], _0385_[19], _0385_[19], _0385_[19], _0385_[19], _0385_[19], _0385_[19:18], _0385_[18], _0385_[18], _0385_[18], _0385_[18], _0385_[18], _0385_[18], _0385_[18], _0385_[18], _0385_[18], _0385_[18], _0385_[18], _0385_[18], _0385_[18:17], _0385_[17], _0385_[17], _0385_[17], _0385_[17], _0385_[17], _0385_[17], _0385_[17], _0385_[17], _0385_[17], _0385_[17], _0385_[17], _0385_[17], _0385_[17], _0385_[17:16], _0385_[16], _0385_[16], _0385_[16], _0385_[16], _0385_[16], _0385_[16], _0385_[16], _0385_[16], _0385_[16], _0385_[16], _0385_[16], _0385_[16], _0385_[16], _0385_[16], _0385_[16:15], _0385_[15], _0385_[15], _0385_[15], _0385_[15], _0385_[15], _0385_[15], _0385_[15], _0385_[15], _0385_[15], _0385_[15], _0385_[15], _0385_[15], _0385_[15], _0385_[15], _0385_[15], _0385_[15:14], _0385_[14], _0385_[14], _0385_[14], _0385_[14], _0385_[14], _0385_[14], _0385_[14], _0385_[14], _0385_[14], _0385_[14], _0385_[14], _0385_[14], _0385_[14], _0385_[14], _0385_[14], _0385_[14], _0385_[14:13], _0385_[13], _0385_[13], _0385_[13], _0385_[13], _0385_[13], _0385_[13], _0385_[13], _0385_[13], _0385_[13], _0385_[13], _0385_[13], _0385_[13], _0385_[13], _0385_[13], _0385_[13], _0385_[13], _0385_[13], _0385_[13:12], _0385_[12], _0385_[12], _0385_[12], _0385_[12], _0385_[12], _0385_[12], _0385_[12], _0385_[12], _0385_[12], _0385_[12], _0385_[12], _0385_[12], _0385_[12], _0385_[12], _0385_[12], _0385_[12], _0385_[12], _0385_[12], _0385_[12:11], _0385_[11], _0385_[11], _0385_[11], _0385_[11], _0385_[11], _0385_[11], _0385_[11], _0385_[11], _0385_[11], _0385_[11], _0385_[11], _0385_[11], _0385_[11], _0385_[11], _0385_[11], _0385_[11], _0385_[11], _0385_[11], _0385_[11], _0385_[11:10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10], _0385_[10:9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9], _0385_[9:8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8], _0385_[8:7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7], _0385_[7:6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6], _0385_[6:5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5], _0385_[5:4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4], _0385_[4:3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3], _0385_[3:2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2], _0385_[2:1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1], _0385_[1:0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0], _0385_[0] } | { _0385_[32], _0385_[32:31], _0385_[32:30], _0385_[32:29], _0385_[32:28], _0385_[32:27], _0385_[32:26], _0385_[32:25], _0385_[32:24], _0385_[32:23], _0385_[32:22], _0385_[32:21], _0385_[32:20], _0385_[32:19], _0385_[32:18], _0385_[32:17], _0385_[32:16], _0385_[32:15], _0385_[32:14], _0385_[32:13], _0385_[32:12], _0385_[32:11], _0385_[32:10], _0385_[32:9], _0385_[32:8], _0385_[32:7], _0385_[32:6], _0385_[32:5], _0385_[32:4], _0385_[32:3], _0385_[32:2], _0385_[32:1] };
assign _0244_ = _0279_ | _0243_;
assign _0167_ = _0244_ & { shift_amt_t0[0], shift_amt_t0[1:0], _0311_, shift_amt_t0[1:0], shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0322_, shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0323_, _0322_, shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0324_, _0323_, _0322_, shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0325_, _0324_, _0323_, _0322_, shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0326_, _0325_, _0324_, _0323_, _0322_, shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0328_, _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0329_, _0328_, _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0330_, _0329_, _0328_, _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0331_, _0330_, _0329_, _0328_, _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0332_, _0331_, _0330_, _0329_, _0328_, _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0333_, _0332_, _0331_, _0330_, _0329_, _0328_, _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0334_, _0333_, _0332_, _0331_, _0330_, _0329_, _0328_, _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0335_, _0334_, _0333_, _0332_, _0331_, _0330_, _0329_, _0328_, _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], _0336_, _0335_, _0334_, _0333_, _0332_, _0331_, _0330_, _0329_, _0328_, _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0], 1'h0, _0336_, _0335_, _0334_, _0333_, _0332_, _0331_, _0330_, _0329_, _0328_, _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, shift_amt_t0[4], _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, shift_amt_t0[3], _0314_, _0313_, _0312_, shift_amt_t0[2], _0311_, shift_amt_t0[1:0] };
assign _0337_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd33;
assign _0338_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd32;
assign _0339_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd31;
assign _0340_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd30;
assign _0341_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd29;
assign _0342_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd28;
assign _0343_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd27;
assign _0344_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd26;
assign _0345_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd25;
assign _0346_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd24;
assign _0347_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd23;
assign _0348_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd22;
assign _0349_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd21;
assign _0350_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd20;
assign _0351_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd19;
assign _0352_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd18;
assign _0353_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd17;
assign _0354_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd16;
assign _0355_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd15;
assign _0356_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd14;
assign _0357_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd13;
assign _0358_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd12;
assign _0359_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd11;
assign _0360_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd10;
assign _0361_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd9;
assign _0362_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd8;
assign _0363_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd7;
assign _0364_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd6;
assign _0365_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd5;
assign _0366_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd4;
assign _0367_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd3;
assign _0368_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd2;
assign _0369_ = { 1'h0, shift_amt_t0[4:0] } >= 32'd1;
assign _0280_ = _0384_ ^ { _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32], _0384_[32] };
assign _0245_ = _0385_ | _0280_;
assign _0168_ = _0245_ & { _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0358_, _0357_, _0356_, _0355_, _0354_, _0353_, _0352_, _0351_, _0350_, _0349_, _0348_, _0347_, _0346_, _0345_, _0344_, _0343_, _0342_, _0341_, _0340_, _0339_, _0338_, _0337_ };
assign shift_result_ext_t0[0] = | { _0168_[0], _0167_[31:0], _0385_[0] };
assign shift_result_ext_t0[1] = | { _0168_[1], _0167_[62:32], _0385_[1] };
assign shift_result_ext_t0[2] = | { _0168_[2], _0167_[92:63], _0385_[2] };
assign shift_result_ext_t0[3] = | { _0168_[3], _0167_[121:93], _0385_[3] };
assign shift_result_ext_t0[4] = | { _0168_[4], _0167_[149:122], _0385_[4] };
assign shift_result_ext_t0[5] = | { _0168_[5], _0167_[176:150], _0385_[5] };
assign shift_result_ext_t0[6] = | { _0168_[6], _0167_[202:177], _0385_[6] };
assign shift_result_ext_t0[7] = | { _0168_[7], _0167_[227:203], _0385_[7] };
assign shift_result_ext_t0[8] = | { _0168_[8], _0167_[251:228], _0385_[8] };
assign shift_result_ext_t0[9] = | { _0168_[9], _0167_[274:252], _0385_[9] };
assign shift_result_ext_t0[10] = | { _0168_[10], _0167_[296:275], _0385_[10] };
assign shift_result_ext_t0[11] = | { _0168_[11], _0167_[317:297], _0385_[11] };
assign shift_result_ext_t0[12] = | { _0168_[12], _0167_[337:318], _0385_[12] };
assign shift_result_ext_t0[13] = | { _0168_[13], _0167_[356:338], _0385_[13] };
assign shift_result_ext_t0[14] = | { _0168_[14], _0167_[374:357], _0385_[14] };
assign shift_result_ext_t0[15] = | { _0168_[15], _0167_[391:375], _0385_[15] };
assign shift_result_ext_t0[16] = | { _0168_[16], _0167_[407:392], _0385_[16] };
assign shift_result_ext_t0[17] = | { _0168_[17], _0167_[422:408], _0385_[17] };
assign shift_result_ext_t0[18] = | { _0168_[18], _0167_[436:423], _0385_[18] };
assign shift_result_ext_t0[19] = | { _0168_[19], _0167_[449:437], _0385_[19] };
assign shift_result_ext_t0[20] = | { _0168_[20], _0167_[461:450], _0385_[20] };
assign shift_result_ext_t0[21] = | { _0168_[21], _0167_[472:462], _0385_[21] };
assign shift_result_ext_t0[22] = | { _0168_[22], _0167_[482:473], _0385_[22] };
assign shift_result_ext_t0[23] = | { _0168_[23], _0167_[491:483], _0385_[23] };
assign shift_result_ext_t0[24] = | { _0168_[24], _0167_[499:492], _0385_[24] };
assign shift_result_ext_t0[25] = | { _0168_[25], _0167_[506:500], _0385_[25] };
assign shift_result_ext_t0[26] = | { _0168_[26], _0167_[512:507], _0385_[26] };
assign shift_result_ext_t0[27] = | { _0168_[27], _0167_[517:513], _0385_[27] };
assign shift_result_ext_t0[28] = | { _0168_[28], _0167_[521:518], _0385_[28] };
assign shift_result_ext_t0[29] = | { _0168_[29], _0167_[524:522], _0385_[29] };
assign shift_result_ext_t0[30] = | { _0168_[30], _0167_[526:525], _0385_[30] };
assign shift_result_ext_t0[31] = | { _0168_[31], _0167_[527], _0385_[31] };
assign _0061_ = ~ { 1'h0, shift_amt_t0[4:0] };
assign _0166_ = { 1'h0, shift_amt[4:0] } & _0061_;
assign _0384_ = $signed({ _0000_, shift_operand }) >>> _0166_;
assign _0385_ = $signed({ _0001_, shift_operand_t0 }) >>> _0166_;
assign _0062_ = ~ { 27'h0000000, operand_b_i_t0[4:0] };
assign _0169_ = { 27'h0000000, operand_b_i[4:0] } & _0062_;
assign _0246_ = { 27'h0000000, operand_b_i[4:0] } | { 27'h0000000, operand_b_i_t0[4:0] };
assign _0372_ = 32'd32 - _0169_;
assign _0373_ = 32'd32 - _0246_;
assign _0247_ = _0372_ ^ _0373_;
assign { _0450_[31:6], shift_amt_compl_t0 } = _0247_ | { 27'h0000000, operand_b_i_t0[4:0] };
assign _0452_ = operand_a_i_t0[31] | operand_b_i_t0[31];
assign _0454_ = operand_a_i_t0[31] | cmp_signed_t0;
assign bwlogic_xor_result_t0 = operand_a_i_t0 | operand_b_i_t0;
assign is_equal_result_o = ! /* src = "generated/sv2v_out.v:11314.20-11314.72" */ adder_result_ext_o[32:1];
assign _0386_ = ~ /* src = "generated/sv2v_out.v:11318.23-11318.47" */ adder_result_ext_o[32];
assign _0063_ = operator_i[5] ? _0397_ : _0395_;
assign _0395_ = operator_i[4] ? _0401_ : _0399_;
assign _0397_ = operator_i[4] ? 1'h0 : _0264_;
assign _0399_ = operator_i[3] ? 1'h0 : _0265_;
assign _0401_ = operator_i[3] ? _0266_ : 1'h0;
assign _0264_ = operator_i[3] ? _0408_ : _0406_;
assign _0265_ = operator_i[2] ? 1'h0 : _0268_;
assign _0266_ = operator_i[2] ? 1'h1 : _0411_;
assign _0406_ = operator_i[2] ? 1'h0 : _0269_;
assign _0408_ = operator_i[2] ? _0416_ : _0414_;
assign _0268_ = operator_i[1] ? 1'h0 : _0271_;
assign _0414_ = operator_i[1] ? _0271_ : 1'h0;
assign _0416_ = operator_i[1] ? 1'h0 : _0272_;
assign _0411_ = operator_i[1] ? 1'h1 : _0271_;
assign _0269_ = operator_i[1] ? _0272_ : 1'h1;
assign _0271_ = operator_i[0] ? 1'h1 : 1'h0;
assign _0272_ = operator_i[0] ? 1'h0 : 1'h1;
assign _0418_ = ~ /* src = "generated/sv2v_out.v:11325.24-11325.33" */ is_equal_result_o;
assign _0419_ = ~ /* src = "generated/sv2v_out.v:11327.59-11327.76" */ is_greater_equal;
assign bwlogic_or_result = operand_a_i | /* src = "generated/sv2v_out.v:11423.29-11423.60" */ operand_b_i;
assign bwlogic_or = _0387_ | /* src = "generated/sv2v_out.v:11426.22-11426.65" */ _0389_;
assign bwlogic_and = _0391_ | /* src = "generated/sv2v_out.v:11427.23-11427.66" */ _0393_;
assign _0422_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ _0420_;
assign _0420_[0] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h1d;
assign _0426_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ { _0424_[4:3], _0424_[1:0], shift_arith };
assign _0424_[1] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h09;
assign shift_arith = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h08;
assign _0424_[3] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h0c;
assign _0424_[4] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h0b;
assign _0430_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ _0428_;
assign _0428_[0] = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ operator_i;
assign _0428_[1] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h01;
assign _0428_[2] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h16;
assign _0428_[3] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h17;
assign _0428_[4] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h18;
assign _0434_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ { _0432_[1:0], _0393_, _0391_, _0389_, _0387_ };
assign _0432_[0] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h02;
assign _0432_[1] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h05;
assign _0387_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h03;
assign _0389_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h06;
assign _0391_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h04;
assign _0393_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11958.3-11976.10" */ 7'h07;
assign _0436_ = bwlogic_and ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11429.3-11433.10" */ bwlogic_and_result : bwlogic_xor_result;
assign bwlogic_result = bwlogic_or ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11429.3-11433.10" */ bwlogic_or_result : _0436_;
assign shift_left = _0424_[0] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11372.3-11381.10" */ 1'h1 : 1'h0;
assign _0424_[0] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11372.3-11381.10" */ 7'h0a;
assign _0440_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ { _0438_[3:2], _0420_[7:4] };
assign _0420_[4] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h19;
assign _0420_[5] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h1a;
assign _0438_[2] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h1f;
assign _0438_[3] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h20;
assign _0420_[6] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h2b;
assign _0420_[7] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h2c;
assign _0444_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ { _0442_[3:2], _0420_[3:2] };
assign _0420_[3] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h1c;
assign _0442_[2] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h21;
assign _0442_[3] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h22;
assign _0420_[1] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11323.3-11329.10" */ 7'h1e;
assign is_greater_equal = _0451_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:11317.7-11317.50|generated/sv2v_out.v:11317.3-11320.52" */ _0453_ : _0386_;
assign cmp_signed = _0446_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11310.3-11313.10" */ 1'h1 : 1'h0;
assign _0446_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11310.3-11313.10" */ { _0442_[2], _0438_[2], _0420_[6], _0420_[4], _0420_[2] };
assign _0420_[2] = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11310.3-11313.10" */ 7'h1b;
assign _0447_ = adder_op_b_negate ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11298.3-11302.10" */ operand_b_neg : { operand_b_i, 1'h0 };
assign adder_in_b = multdiv_sel_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11298.3-11302.10" */ multdiv_operand_b_i : _0447_;
assign adder_in_a = multdiv_sel_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:11289.3-11295.10" */ multdiv_operand_a_i : { operand_a_i, 1'h1 };
assign adder_op_b_negate = operator_i[6] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:11273.3-11286.10" */ 1'h0 : _0063_;
assign shift_result_ext = $signed({ _0000_, shift_operand }) >>> /* src = "generated/sv2v_out.v:11397.29-11397.120" */ shift_amt[4:0];
assign { _0449_[31:6], shift_amt_compl } = 32'd32 - /* src = "generated/sv2v_out.v:11364.27-11364.48" */ operand_b_i[4:0];
assign shift_amt[4:0] = instr_first_cycle_i ? /* src = "generated/sv2v_out.v:11369.22-11369.195" */ operand_b_i[4:0] : shift_amt_compl[4:0];
assign shift_operand = shift_left ? /* src = "generated/sv2v_out.v:11390.21-11390.61" */ { operand_a_i[0], operand_a_i[1], operand_a_i[2], operand_a_i[3], operand_a_i[4], operand_a_i[5], operand_a_i[6], operand_a_i[7], operand_a_i[8], operand_a_i[9], operand_a_i[10], operand_a_i[11], operand_a_i[12], operand_a_i[13], operand_a_i[14], operand_a_i[15], operand_a_i[16], operand_a_i[17], operand_a_i[18], operand_a_i[19], operand_a_i[20], operand_a_i[21], operand_a_i[22], operand_a_i[23], operand_a_i[24], operand_a_i[25], operand_a_i[26], operand_a_i[27], operand_a_i[28], operand_a_i[29], operand_a_i[30], operand_a_i[31] } : operand_a_i;
assign shift_result = shift_left ? /* src = "generated/sv2v_out.v:11406.19-11406.63" */ { shift_result_ext[0], shift_result_ext[1], shift_result_ext[2], shift_result_ext[3], shift_result_ext[4], shift_result_ext[5], shift_result_ext[6], shift_result_ext[7], shift_result_ext[8], shift_result_ext[9], shift_result_ext[10], shift_result_ext[11], shift_result_ext[12], shift_result_ext[13], shift_result_ext[14], shift_result_ext[15], shift_result_ext[16], shift_result_ext[17], shift_result_ext[18], shift_result_ext[19], shift_result_ext[20], shift_result_ext[21], shift_result_ext[22], shift_result_ext[23], shift_result_ext[24], shift_result_ext[25], shift_result_ext[26], shift_result_ext[27], shift_result_ext[28], shift_result_ext[29], shift_result_ext[30], shift_result_ext[31] } : shift_result_ext[31:0];
assign _0451_ = operand_a_i[31] ^ /* src = "generated/sv2v_out.v:11317.8-11317.41" */ operand_b_i[31];
assign _0453_ = operand_a_i[31] ^ /* src = "generated/sv2v_out.v:11320.23-11320.51" */ cmp_signed;
assign bwlogic_xor_result = operand_a_i ^ /* src = "generated/sv2v_out.v:11425.30-11425.61" */ operand_b_i;
assign _0424_[2] = shift_arith;
assign { _0425_[2], _0425_[0] } = { shift_arith_t0, shift_left_t0 };
assign _0432_[5:2] = { _0393_, _0391_, _0389_, _0387_ };
assign _0433_[5:2] = { _0394_, _0392_, _0390_, _0388_ };
assign { _0438_[5:4], _0438_[1:0] } = _0420_[7:4];
assign { _0439_[5:4], _0439_[1:0] } = _0421_[7:4];
assign _0442_[1:0] = _0420_[3:2];
assign _0443_[1:0] = _0421_[3:2];
assign _0449_[5:0] = shift_amt_compl;
assign _0450_[5:0] = shift_amt_compl_t0;
assign adder_result_o = adder_result_ext_o[32:1];
assign adder_result_o_t0 = adder_result_ext_o_t0[32:1];
assign imd_val_d_o = 64'h0000000000000000;
assign imd_val_d_o_t0 = 64'h0000000000000000;
assign imd_val_we_o = 2'h0;
assign imd_val_we_o_t0 = 2'h0;
assign shift_amt[5] = 1'h0;
assign shift_amt_t0[5] = 1'h0;
endmodule

module \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1 (clk_i, rst_ni, ctrl_busy_o, illegal_insn_i, ecall_insn_i, mret_insn_i, dret_insn_i, wfi_insn_i, ebrk_insn_i, csr_pipe_flush_i, instr_valid_i, instr_i, instr_compressed_i, instr_is_compressed_i, instr_bp_taken_i, instr_fetch_err_i, instr_fetch_err_plus2_i, pc_id_i, instr_valid_clear_o, id_in_ready_o, controller_run_o
, instr_exec_i, instr_req_o, pc_set_o, pc_mux_o, nt_branch_mispredict_o, exc_pc_mux_o, exc_cause_o, lsu_addr_last_i, load_err_i, store_err_i, mem_resp_intg_err_i, wb_exception_o, id_exception_o, branch_set_i, branch_not_set_i, jump_set_i, csr_mstatus_mie_i, irq_pending_i, irqs_i, irq_nm_ext_i, nmi_mode_o
, debug_req_i, debug_cause_o, debug_csr_save_o, debug_mode_o, debug_mode_entering_o, debug_single_step_i, debug_ebreakm_i, debug_ebreaku_i, trigger_match_i, csr_save_if_o, csr_save_id_o, csr_save_wb_o, csr_restore_mret_id_o, csr_restore_dret_id_o, csr_save_cause_o, csr_mtval_o, priv_mode_i, stall_id_i, stall_wb_i, flush_id_o, ready_wb_i
, perf_jump_o, perf_tbranch_o, branch_not_set_i_t0, branch_set_i_t0, controller_run_o_t0, csr_mstatus_mie_i_t0, csr_mtval_o_t0, csr_pipe_flush_i_t0, csr_restore_dret_id_o_t0, instr_i_t0, csr_restore_mret_id_o_t0, csr_save_cause_o_t0, csr_save_id_o_t0, csr_save_if_o_t0, csr_save_wb_o_t0, ctrl_busy_o_t0, debug_cause_o_t0, debug_csr_save_o_t0, debug_ebreakm_i_t0, debug_ebreaku_i_t0, debug_mode_entering_o_t0
, debug_mode_o_t0, debug_req_i_t0, debug_single_step_i_t0, dret_insn_i_t0, ebrk_insn_i_t0, ecall_insn_i_t0, exc_cause_o_t0, exc_pc_mux_o_t0, flush_id_o_t0, id_exception_o_t0, id_in_ready_o_t0, illegal_insn_i_t0, instr_bp_taken_i_t0, instr_compressed_i_t0, instr_exec_i_t0, instr_fetch_err_i_t0, instr_fetch_err_plus2_i_t0, instr_is_compressed_i_t0, instr_valid_clear_o_t0, instr_valid_i_t0, irq_nm_ext_i_t0
, irq_pending_i_t0, irqs_i_t0, jump_set_i_t0, load_err_i_t0, lsu_addr_last_i_t0, mem_resp_intg_err_i_t0, mret_insn_i_t0, nmi_mode_o_t0, nt_branch_mispredict_o_t0, pc_id_i_t0, pc_mux_o_t0, pc_set_o_t0, perf_jump_o_t0, perf_tbranch_o_t0, priv_mode_i_t0, ready_wb_i_t0, stall_id_i_t0, stall_wb_i_t0, store_err_i_t0, trigger_match_i_t0, wb_exception_o_t0
, wfi_insn_i_t0, instr_req_o_t0);
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0001_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0003_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0005_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0007_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0009_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0011_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0013_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0015_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0016_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0017_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0018_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0019_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0021_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0022_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0023_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0024_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0025_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0026_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0027_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _0028_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _0029_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0030_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0031_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0032_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0033_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0034_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0035_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0036_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0037_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0038_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0039_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0040_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0041_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0042_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0043_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0044_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _0045_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _0046_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [1:0] _0047_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [1:0] _0048_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0049_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0050_;
/* src = "generated/sv2v_out.v:12399.4-12411.7" */
wire _0051_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12399.4-12411.7" */
wire _0052_;
/* src = "generated/sv2v_out.v:12399.4-12411.7" */
wire _0053_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0054_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0055_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0056_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0057_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0058_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0059_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0060_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [2:0] _0061_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [2:0] _0062_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0063_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0064_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0065_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0066_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0067_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0068_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0069_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0070_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0071_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _0072_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _0073_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0074_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0075_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0076_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0077_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0078_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0079_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0080_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0081_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _0082_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _0083_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0084_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0085_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0086_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0087_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0088_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0089_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0090_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0091_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0092_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0093_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [2:0] _0094_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [2:0] _0095_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0096_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0097_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _0098_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _0099_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0100_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0101_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0102_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0103_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0104_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0105_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0106_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _0107_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _0108_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0109_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0110_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0111_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0112_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0113_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0114_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0115_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0116_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0117_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [2:0] _0118_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0119_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0120_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0121_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0122_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _0123_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _0124_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0125_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0126_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _0127_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _0128_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0129_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0130_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0131_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0132_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0133_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0134_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0135_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0136_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0137_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _0138_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [31:0] _0139_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0140_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0141_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _0142_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0143_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0144_;
/* src = "generated/sv2v_out.v:12368.4-12387.7" */
wire _0145_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0146_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0147_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0148_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0149_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _0150_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _0151_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0152_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0153_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0154_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0155_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0156_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire _0157_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0158_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0159_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _0160_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _0161_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0162_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0163_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0164_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [3:0] _0165_;
/* src = "generated/sv2v_out.v:12474.2-12692.5" */
wire [6:0] _0166_;
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0167_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12441.2-12449.5" */
wire [3:0] _0168_;
/* src = "generated/sv2v_out.v:12638.49-12638.64" */
wire [31:0] _0169_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12638.49-12638.64" */
wire [31:0] _0170_;
/* src = "generated/sv2v_out.v:12404.10-12404.38" */
wire _0171_;
/* src = "generated/sv2v_out.v:12412.46-12412.108" */
wire _0172_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12412.46-12412.108" */
wire _0173_;
/* src = "generated/sv2v_out.v:12434.45-12434.80" */
wire _0174_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12434.45-12434.80" */
wire _0175_;
/* src = "generated/sv2v_out.v:12436.55-12436.86" */
wire _0176_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12436.55-12436.86" */
wire _0177_;
/* src = "generated/sv2v_out.v:12440.24-12440.60" */
wire _0178_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12440.24-12440.60" */
wire _0179_;
/* src = "generated/sv2v_out.v:12440.23-12440.75" */
wire _0180_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12440.23-12440.75" */
wire _0181_;
/* src = "generated/sv2v_out.v:12440.90-12440.117" */
wire _0182_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12440.90-12440.117" */
wire _0183_;
/* src = "generated/sv2v_out.v:12451.52-12451.86" */
wire _0184_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12451.52-12451.86" */
wire _0185_;
/* src = "generated/sv2v_out.v:12578.11-12578.37" */
wire _0186_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12578.11-12578.37" */
wire _0187_;
/* src = "generated/sv2v_out.v:12697.26-12697.43" */
wire _0188_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12697.26-12697.43" */
wire _0189_;
wire [31:0] _0190_;
wire _0191_;
wire _0192_;
wire _0193_;
wire _0194_;
wire _0195_;
wire _0196_;
wire _0197_;
wire _0198_;
wire _0199_;
wire _0200_;
wire [3:0] _0201_;
wire [2:0] _0202_;
wire [1:0] _0203_;
wire [3:0] _0204_;
wire [1:0] _0205_;
wire [1:0] _0206_;
wire [3:0] _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire [1:0] _0217_;
wire [3:0] _0218_;
wire [2:0] _0219_;
wire [2:0] _0220_;
wire [6:0] _0221_;
wire [3:0] _0222_;
wire [1:0] _0223_;
wire [2:0] _0224_;
wire [14:0] _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire _0241_;
wire _0242_;
wire _0243_;
wire _0244_;
wire _0245_;
wire _0246_;
wire _0247_;
wire _0248_;
wire _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire [3:0] _0255_;
wire [3:0] _0256_;
wire [3:0] _0257_;
wire [3:0] _0258_;
wire [3:0] _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire [2:0] _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire [31:0] _0269_;
wire _0270_;
wire [6:0] _0271_;
wire [1:0] _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire _0276_;
wire _0277_;
wire _0278_;
wire _0279_;
wire [3:0] _0280_;
wire _0281_;
wire [3:0] _0282_;
wire _0283_;
wire [2:0] _0284_;
wire [3:0] _0285_;
wire [31:0] _0286_;
wire [31:0] _0287_;
wire [31:0] _0288_;
wire [31:0] _0289_;
wire [31:0] _0290_;
wire [6:0] _0291_;
wire [6:0] _0292_;
wire [6:0] _0293_;
wire [6:0] _0294_;
wire [6:0] _0295_;
wire [3:0] _0296_;
wire [3:0] _0297_;
wire [3:0] _0298_;
wire _0299_;
wire _0300_;
wire _0301_;
wire [3:0] _0302_;
wire _0303_;
wire [2:0] _0304_;
wire [6:0] _0305_;
wire [6:0] _0306_;
wire _0307_;
wire [6:0] _0308_;
wire [3:0] _0309_;
wire [3:0] _0310_;
wire _0311_;
wire [3:0] _0312_;
wire [3:0] _0313_;
wire [3:0] _0314_;
wire [3:0] _0315_;
wire [3:0] _0316_;
wire [3:0] _0317_;
wire [3:0] _0318_;
wire [3:0] _0319_;
wire [3:0] _0320_;
wire [3:0] _0321_;
wire [3:0] _0322_;
wire [3:0] _0323_;
wire [3:0] _0324_;
wire [3:0] _0325_;
wire [3:0] _0326_;
wire [3:0] _0327_;
wire [3:0] _0328_;
wire _0329_;
wire _0330_;
wire _0331_;
wire [2:0] _0332_;
wire [2:0] _0333_;
wire [2:0] _0334_;
wire [31:0] _0335_;
wire [31:0] _0336_;
wire _0337_;
wire _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire _0343_;
wire _0344_;
wire _0345_;
wire _0346_;
wire _0347_;
wire _0348_;
wire _0349_;
wire _0350_;
wire _0351_;
wire _0352_;
wire [1:0] _0353_;
wire [2:0] _0354_;
wire _0355_;
wire [1:0] _0356_;
wire [2:0] _0357_;
wire _0358_;
wire [1:0] _0359_;
wire [1:0] _0360_;
wire [1:0] _0361_;
wire [1:0] _0362_;
wire [1:0] _0363_;
wire [1:0] _0364_;
wire _0365_;
wire [1:0] _0366_;
wire [1:0] _0367_;
wire _0368_;
wire _0369_;
wire [3:0] _0370_;
wire [2:0] _0371_;
wire [1:0] _0372_;
wire [2:0] _0373_;
wire [1:0] _0374_;
wire [1:0] _0375_;
wire _0376_;
wire [2:0] _0377_;
wire [1:0] _0378_;
wire [1:0] _0379_;
wire _0380_;
wire [1:0] _0381_;
wire _0382_;
wire _0383_;
wire [2:0] _0384_;
wire _0385_;
wire _0386_;
wire _0387_;
wire [1:0] _0388_;
wire _0389_;
wire _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire _0398_;
wire _0399_;
wire _0400_;
wire _0401_;
wire _0402_;
wire _0403_;
wire _0404_;
wire _0405_;
wire _0406_;
wire _0407_;
wire _0408_;
wire _0409_;
wire _0410_;
wire _0411_;
wire _0412_;
wire _0413_;
wire _0414_;
wire _0415_;
wire _0416_;
wire _0417_;
wire _0418_;
wire _0419_;
wire _0420_;
wire _0421_;
wire _0422_;
/* cellift = 32'd1 */
wire _0423_;
wire _0424_;
wire _0425_;
wire _0426_;
wire _0427_;
wire _0428_;
wire _0429_;
wire _0430_;
/* cellift = 32'd1 */
wire _0431_;
wire _0432_;
/* cellift = 32'd1 */
wire _0433_;
wire _0434_;
/* cellift = 32'd1 */
wire _0435_;
wire _0436_;
/* cellift = 32'd1 */
wire _0437_;
wire _0438_;
/* cellift = 32'd1 */
wire _0439_;
wire _0440_;
/* cellift = 32'd1 */
wire _0441_;
wire _0442_;
/* cellift = 32'd1 */
wire _0443_;
wire _0444_;
/* cellift = 32'd1 */
wire _0445_;
wire _0446_;
/* cellift = 32'd1 */
wire _0447_;
wire _0448_;
/* cellift = 32'd1 */
wire _0449_;
wire _0450_;
/* cellift = 32'd1 */
wire _0451_;
wire _0452_;
/* cellift = 32'd1 */
wire _0453_;
wire _0454_;
wire _0455_;
/* cellift = 32'd1 */
wire _0456_;
wire [31:0] _0457_;
wire _0458_;
wire _0459_;
wire _0460_;
wire _0461_;
wire _0462_;
wire _0463_;
wire _0464_;
wire _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire _0469_;
wire _0470_;
wire _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire _0477_;
wire _0478_;
wire _0479_;
wire _0480_;
wire _0481_;
wire _0482_;
wire _0483_;
wire _0484_;
wire _0485_;
wire _0486_;
wire _0487_;
wire _0488_;
wire _0489_;
wire _0490_;
wire _0491_;
wire _0492_;
wire _0493_;
wire _0494_;
wire _0495_;
wire _0496_;
wire _0497_;
wire _0498_;
wire _0499_;
wire _0500_;
wire _0501_;
wire _0502_;
wire _0503_;
wire _0504_;
wire _0505_;
wire _0506_;
wire _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0517_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
wire _0525_;
wire _0526_;
wire _0527_;
wire [3:0] _0528_;
wire [3:0] _0529_;
wire [3:0] _0530_;
wire [31:0] _0531_;
wire [31:0] _0532_;
wire [31:0] _0533_;
wire [3:0] _0534_;
wire [2:0] _0535_;
wire [1:0] _0536_;
wire [1:0] _0537_;
wire [3:0] _0538_;
wire [1:0] _0539_;
wire [3:0] _0540_;
wire [2:0] _0541_;
wire [2:0] _0542_;
wire [6:0] _0543_;
wire [3:0] _0544_;
wire [1:0] _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire _0560_;
wire [2:0] _0561_;
wire [3:0] _0562_;
wire [3:0] _0563_;
wire [3:0] _0564_;
wire [3:0] _0565_;
wire [3:0] _0566_;
wire [3:0] _0567_;
wire [3:0] _0568_;
wire [3:0] _0569_;
wire [3:0] _0570_;
wire [3:0] _0571_;
wire [3:0] _0572_;
wire [3:0] _0573_;
wire [3:0] _0574_;
wire [3:0] _0575_;
wire [3:0] _0576_;
wire [3:0] _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire [2:0] _0588_;
wire [2:0] _0589_;
wire [2:0] _0590_;
wire [2:0] _0591_;
wire [2:0] _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire _0596_;
wire _0597_;
wire _0598_;
wire _0599_;
wire _0600_;
wire _0601_;
wire _0602_;
wire _0603_;
wire _0604_;
wire _0605_;
wire _0606_;
wire _0607_;
wire _0608_;
wire _0609_;
wire _0610_;
wire _0611_;
wire [31:0] _0612_;
wire [31:0] _0613_;
wire [31:0] _0614_;
wire [31:0] _0615_;
wire [31:0] _0616_;
wire _0617_;
wire _0618_;
wire _0619_;
wire _0620_;
wire _0621_;
wire _0622_;
wire _0623_;
wire _0624_;
wire _0625_;
wire [6:0] _0626_;
wire [6:0] _0627_;
wire [6:0] _0628_;
wire [6:0] _0629_;
wire [6:0] _0630_;
wire [1:0] _0631_;
wire [1:0] _0632_;
wire [1:0] _0633_;
wire _0634_;
wire _0635_;
wire _0636_;
wire [1:0] _0637_;
wire _0638_;
wire _0639_;
wire _0640_;
wire _0641_;
wire _0642_;
wire _0643_;
wire _0644_;
wire _0645_;
wire _0646_;
wire _0647_;
wire _0648_;
wire _0649_;
wire _0650_;
wire _0651_;
wire _0652_;
wire _0653_;
wire _0654_;
wire _0655_;
wire _0656_;
wire _0657_;
wire _0658_;
wire _0659_;
wire _0660_;
wire _0661_;
wire _0662_;
wire _0663_;
wire _0664_;
wire _0665_;
wire _0666_;
wire _0667_;
wire _0668_;
wire _0669_;
wire _0670_;
wire _0671_;
wire _0672_;
wire _0673_;
wire _0674_;
wire _0675_;
wire _0676_;
wire _0677_;
wire _0678_;
wire _0679_;
wire _0680_;
wire _0681_;
wire _0682_;
wire [3:0] _0683_;
wire [14:0] _0684_;
wire _0685_;
wire _0686_;
wire _0687_;
wire _0688_;
wire _0689_;
wire _0690_;
wire _0691_;
wire _0692_;
wire _0693_;
wire _0694_;
wire _0695_;
wire _0696_;
wire _0697_;
wire _0698_;
wire _0699_;
wire _0700_;
wire _0701_;
wire _0702_;
wire _0703_;
wire _0704_;
wire _0705_;
wire _0706_;
wire _0707_;
wire _0708_;
wire _0709_;
wire _0710_;
wire _0711_;
wire _0712_;
wire _0713_;
wire _0714_;
wire _0715_;
wire _0716_;
wire _0717_;
wire _0718_;
wire _0719_;
wire _0720_;
wire _0721_;
wire _0722_;
wire _0723_;
wire _0724_;
wire _0725_;
wire _0726_;
wire _0727_;
wire _0728_;
wire _0729_;
wire _0730_;
wire _0731_;
wire _0732_;
wire _0733_;
wire _0734_;
wire _0735_;
wire _0736_;
wire _0737_;
wire _0738_;
wire _0739_;
wire _0740_;
wire _0741_;
wire _0742_;
wire _0743_;
wire _0744_;
wire _0745_;
wire _0746_;
wire _0747_;
wire _0748_;
wire _0749_;
wire _0750_;
wire _0751_;
wire _0752_;
wire _0753_;
wire _0754_;
wire _0755_;
wire _0756_;
wire _0757_;
wire _0758_;
wire _0759_;
wire _0760_;
wire _0761_;
wire _0762_;
wire _0763_;
wire _0764_;
wire _0765_;
wire _0766_;
wire _0767_;
wire _0768_;
wire _0769_;
wire _0770_;
wire _0771_;
wire _0772_;
wire _0773_;
wire _0774_;
wire _0775_;
wire _0776_;
wire _0777_;
wire _0778_;
wire _0779_;
wire _0780_;
wire _0781_;
wire [3:0] _0782_;
wire [3:0] _0783_;
wire [3:0] _0784_;
wire [3:0] _0785_;
wire _0786_;
wire _0787_;
wire _0788_;
wire _0789_;
wire [2:0] _0790_;
wire [2:0] _0791_;
wire [3:0] _0792_;
wire [3:0] _0793_;
wire _0794_;
wire [31:0] _0795_;
wire [31:0] _0796_;
wire [31:0] _0797_;
wire [31:0] _0798_;
wire [31:0] _0799_;
wire [31:0] _0800_;
wire [31:0] _0801_;
wire [31:0] _0802_;
wire [31:0] _0803_;
wire [31:0] _0804_;
wire [31:0] _0805_;
wire [31:0] _0806_;
wire [31:0] _0807_;
wire [31:0] _0808_;
wire [31:0] _0809_;
wire [6:0] _0810_;
wire [6:0] _0811_;
wire [6:0] _0812_;
wire [6:0] _0813_;
wire [6:0] _0814_;
wire [6:0] _0815_;
wire [6:0] _0816_;
wire [6:0] _0817_;
wire [6:0] _0818_;
wire [6:0] _0819_;
wire [6:0] _0820_;
wire [6:0] _0821_;
wire [3:0] _0822_;
wire [3:0] _0823_;
wire [3:0] _0824_;
wire [3:0] _0825_;
wire [3:0] _0826_;
wire [3:0] _0827_;
wire [3:0] _0828_;
wire [3:0] _0829_;
wire _0830_;
wire _0831_;
wire _0832_;
wire _0833_;
wire _0834_;
wire _0835_;
wire _0836_;
wire _0837_;
wire [3:0] _0838_;
wire [3:0] _0839_;
wire [3:0] _0840_;
wire _0841_;
wire _0842_;
wire [31:0] _0843_;
wire [31:0] _0844_;
wire _0845_;
wire [6:0] _0846_;
wire [6:0] _0847_;
wire _0848_;
wire _0849_;
wire [1:0] _0850_;
wire [1:0] _0851_;
wire [2:0] _0852_;
wire [2:0] _0853_;
wire _0854_;
wire _0855_;
wire _0856_;
wire _0857_;
wire _0858_;
wire _0859_;
wire _0860_;
wire [6:0] _0861_;
wire [6:0] _0862_;
wire [6:0] _0863_;
wire [6:0] _0864_;
wire [6:0] _0865_;
wire [31:0] _0866_;
wire [31:0] _0867_;
wire _0868_;
wire _0869_;
wire [31:0] _0870_;
wire [31:0] _0871_;
wire [6:0] _0872_;
wire [6:0] _0873_;
wire [6:0] _0874_;
wire _0875_;
wire _0876_;
wire _0877_;
wire [31:0] _0878_;
wire [31:0] _0879_;
wire [6:0] _0880_;
wire [6:0] _0881_;
wire _0882_;
wire _0883_;
wire [3:0] _0884_;
wire [3:0] _0885_;
wire _0886_;
wire _0887_;
wire [3:0] _0888_;
wire [3:0] _0889_;
wire _0890_;
wire _0891_;
wire _0892_;
wire [3:0] _0893_;
wire [3:0] _0894_;
wire [3:0] _0895_;
wire _0896_;
wire _0897_;
wire _0898_;
wire _0899_;
wire [3:0] _0900_;
wire [3:0] _0901_;
wire [3:0] _0902_;
wire [3:0] _0903_;
wire [3:0] _0904_;
wire _0905_;
wire _0906_;
wire [3:0] _0907_;
wire [3:0] _0908_;
wire _0909_;
wire _0910_;
wire _0911_;
wire _0912_;
wire _0913_;
wire _0914_;
wire _0915_;
wire _0916_;
wire _0917_;
wire _0918_;
wire _0919_;
wire [3:0] _0920_;
wire [3:0] _0921_;
wire [3:0] _0922_;
wire [3:0] _0923_;
wire [3:0] _0924_;
wire [3:0] _0925_;
wire [3:0] _0926_;
wire [3:0] _0927_;
wire [3:0] _0928_;
wire [3:0] _0929_;
wire [3:0] _0930_;
wire [3:0] _0931_;
wire [3:0] _0932_;
wire [3:0] _0933_;
wire [3:0] _0934_;
wire [3:0] _0935_;
wire [3:0] _0936_;
wire [3:0] _0937_;
wire [3:0] _0938_;
wire [3:0] _0939_;
wire [3:0] _0940_;
wire [3:0] _0941_;
wire [3:0] _0942_;
wire [3:0] _0943_;
wire [3:0] _0944_;
wire [3:0] _0945_;
wire [3:0] _0946_;
wire [3:0] _0947_;
wire _0948_;
wire _0949_;
wire _0950_;
wire _0951_;
wire _0952_;
wire _0953_;
wire _0954_;
wire _0955_;
wire [2:0] _0956_;
wire [2:0] _0957_;
wire [2:0] _0958_;
wire [2:0] _0959_;
wire [2:0] _0960_;
wire [2:0] _0961_;
wire [31:0] _0962_;
wire [31:0] _0963_;
wire [31:0] _0964_;
wire [31:0] _0965_;
wire [31:0] _0966_;
wire [31:0] _0967_;
wire _0968_;
/* cellift = 32'd1 */
wire _0969_;
wire _0970_;
/* cellift = 32'd1 */
wire _0971_;
wire _0972_;
/* cellift = 32'd1 */
wire _0973_;
wire _0974_;
/* cellift = 32'd1 */
wire _0975_;
wire _0976_;
/* cellift = 32'd1 */
wire _0977_;
wire [31:0] _0978_;
wire _0979_;
wire _0980_;
wire _0981_;
wire _0982_;
wire _0983_;
wire _0984_;
wire _0985_;
wire _0986_;
wire _0987_;
wire _0988_;
wire _0989_;
wire _0990_;
wire _0991_;
wire _0992_;
wire _0993_;
wire _0994_;
wire _0995_;
wire _0996_;
wire _0997_;
wire _0998_;
wire _0999_;
wire _1000_;
wire _1001_;
wire _1002_;
wire _1003_;
wire _1004_;
wire _1005_;
wire [3:0] _1006_;
wire [3:0] _1007_;
wire [3:0] _1008_;
wire [3:0] _1009_;
wire [31:0] _1010_;
wire [31:0] _1011_;
wire [31:0] _1012_;
wire [31:0] _1013_;
wire [3:0] _1014_;
wire [1:0] _1015_;
wire [1:0] _1016_;
wire _1017_;
wire _1018_;
wire _1019_;
wire _1020_;
wire _1021_;
wire [3:0] _1022_;
wire [3:0] _1023_;
wire [3:0] _1024_;
wire [3:0] _1025_;
wire [3:0] _1026_;
wire [3:0] _1027_;
wire [3:0] _1028_;
wire [3:0] _1029_;
wire [3:0] _1030_;
wire [3:0] _1031_;
wire [3:0] _1032_;
wire [3:0] _1033_;
wire [3:0] _1034_;
wire [3:0] _1035_;
wire _1036_;
wire _1037_;
wire _1038_;
wire _1039_;
wire _1040_;
wire _1041_;
wire _1042_;
wire _1043_;
wire _1044_;
wire [2:0] _1045_;
wire [2:0] _1046_;
wire [2:0] _1047_;
wire [2:0] _1048_;
wire _1049_;
wire _1050_;
wire _1051_;
wire _1052_;
wire _1053_;
wire _1054_;
wire _1055_;
wire _1056_;
wire _1057_;
wire _1058_;
wire _1059_;
wire _1060_;
wire [31:0] _1061_;
wire [31:0] _1062_;
wire [31:0] _1063_;
wire [31:0] _1064_;
wire _1065_;
wire _1066_;
wire _1067_;
wire _1068_;
wire [6:0] _1069_;
wire [6:0] _1070_;
wire [6:0] _1071_;
wire [6:0] _1072_;
wire [1:0] _1073_;
wire [1:0] _1074_;
wire [1:0] _1075_;
wire _1076_;
wire _1077_;
wire _1078_;
wire _1079_;
wire _1080_;
wire _1081_;
wire _1082_;
wire _1083_;
wire _1084_;
wire _1085_;
wire _1086_;
wire _1087_;
wire _1088_;
wire _1089_;
wire _1090_;
wire _1091_;
wire _1092_;
wire _1093_;
wire _1094_;
wire _1095_;
wire _1096_;
wire _1097_;
wire _1098_;
wire _1099_;
wire _1100_;
wire _1101_;
wire _1102_;
wire _1103_;
wire _1104_;
wire _1105_;
wire _1106_;
wire _1107_;
wire _1108_;
wire _1109_;
wire _1110_;
wire _1111_;
wire _1112_;
wire _1113_;
wire _1114_;
wire _1115_;
wire _1116_;
wire _1117_;
wire _1118_;
wire _1119_;
wire _1120_;
wire _1121_;
wire _1122_;
wire [3:0] _1123_;
wire [3:0] _1124_;
wire _1125_;
wire [2:0] _1126_;
wire [3:0] _1127_;
wire [31:0] _1128_;
wire [31:0] _1129_;
wire [31:0] _1130_;
wire [31:0] _1131_;
wire [31:0] _1132_;
wire [31:0] _1133_;
wire [31:0] _1134_;
wire [31:0] _1135_;
wire [31:0] _1136_;
wire [31:0] _1137_;
wire [31:0] _1138_;
wire [31:0] _1139_;
wire [6:0] _1140_;
wire [6:0] _1141_;
wire [6:0] _1142_;
wire [6:0] _1143_;
wire [6:0] _1144_;
wire [6:0] _1145_;
wire [6:0] _1146_;
wire [6:0] _1147_;
wire [6:0] _1148_;
wire [3:0] _1149_;
wire [3:0] _1150_;
wire [3:0] _1151_;
wire [3:0] _1152_;
wire _1153_;
wire _1154_;
wire _1155_;
wire _1156_;
wire [3:0] _1157_;
wire [3:0] _1158_;
wire [3:0] _1159_;
wire _1160_;
wire _1161_;
wire [31:0] _1162_;
wire [6:0] _1163_;
wire _1164_;
wire [1:0] _1165_;
wire [2:0] _1166_;
wire _1167_;
wire [6:0] _1168_;
wire [6:0] _1169_;
wire [6:0] _1170_;
wire [6:0] _1171_;
wire [31:0] _1172_;
wire _1173_;
wire [31:0] _1174_;
wire [6:0] _1175_;
wire [6:0] _1176_;
wire [6:0] _1177_;
wire _1178_;
wire _1179_;
wire _1180_;
wire [31:0] _1181_;
wire [6:0] _1182_;
wire [3:0] _1183_;
wire _1184_;
wire [3:0] _1185_;
wire _1186_;
wire _1187_;
wire _1188_;
wire [3:0] _1189_;
wire [3:0] _1190_;
wire [3:0] _1191_;
wire _1192_;
wire [3:0] _1193_;
wire [3:0] _1194_;
wire [3:0] _1195_;
wire [3:0] _1196_;
wire [3:0] _1197_;
wire [3:0] _1198_;
wire [3:0] _1199_;
wire [3:0] _1200_;
wire [3:0] _1201_;
wire [3:0] _1202_;
wire [3:0] _1203_;
wire [3:0] _1204_;
wire [3:0] _1205_;
wire [3:0] _1206_;
wire [3:0] _1207_;
wire [3:0] _1208_;
wire [3:0] _1209_;
wire [3:0] _1210_;
wire _1211_;
wire _1212_;
wire _1213_;
wire _1214_;
wire _1215_;
wire _1216_;
wire _1217_;
wire [2:0] _1218_;
wire [2:0] _1219_;
wire [2:0] _1220_;
wire [31:0] _1221_;
wire [31:0] _1222_;
wire [31:0] _1223_;
wire [31:0] _1224_;
wire [31:0] _1225_;
wire [31:0] _1226_;
wire [31:0] _1227_;
wire _1228_;
wire [3:0] _1229_;
wire [31:0] _1230_;
wire [3:0] _1231_;
wire [3:0] _1232_;
wire [3:0] _1233_;
wire [3:0] _1234_;
wire [3:0] _1235_;
wire _1236_;
wire _1237_;
wire [2:0] _1238_;
wire _1239_;
wire _1240_;
wire _1241_;
wire _1242_;
wire _1243_;
wire [31:0] _1244_;
wire _1245_;
wire _1246_;
wire [6:0] _1247_;
wire [1:0] _1248_;
wire _1249_;
wire [31:0] _1250_;
wire [31:0] _1251_;
wire [31:0] _1252_;
wire [31:0] _1253_;
wire [31:0] _1254_;
wire [6:0] _1255_;
wire [6:0] _1256_;
wire [6:0] _1257_;
wire [6:0] _1258_;
wire [6:0] _1259_;
wire [3:0] _1260_;
wire [3:0] _1261_;
wire [3:0] _1262_;
wire [3:0] _1263_;
wire _1264_;
wire [1:0] _1265_;
wire _1266_;
wire [6:0] _1267_;
wire [6:0] _1268_;
wire _1269_;
wire _1270_;
wire [3:0] _1271_;
wire [3:0] _1272_;
wire _1273_;
wire _1274_;
wire [2:0] _1275_;
wire [2:0] _1276_;
wire [2:0] _1277_;
wire [31:0] _1278_;
wire [31:0] _1279_;
wire _1280_;
wire _1281_;
wire _1282_;
wire _1283_;
wire _1284_;
wire _1285_;
wire _1286_;
wire _1287_;
wire _1288_;
wire _1289_;
wire _1290_;
wire _1291_;
wire _1292_;
wire _1293_;
wire _1294_;
wire [31:0] _1295_;
wire [31:0] _1296_;
wire [3:0] _1297_;
/* cellift = 32'd1 */
wire [3:0] _1298_;
wire [3:0] _1299_;
/* cellift = 32'd1 */
wire [3:0] _1300_;
wire [3:0] _1301_;
/* cellift = 32'd1 */
wire [3:0] _1302_;
wire [3:0] _1303_;
/* cellift = 32'd1 */
wire [3:0] _1304_;
wire [3:0] _1305_;
/* cellift = 32'd1 */
wire [3:0] _1306_;
wire [3:0] _1307_;
/* cellift = 32'd1 */
wire [3:0] _1308_;
wire [3:0] _1309_;
/* cellift = 32'd1 */
wire [3:0] _1310_;
wire _1311_;
/* cellift = 32'd1 */
wire _1312_;
wire _1313_;
/* cellift = 32'd1 */
wire _1314_;
wire _1315_;
/* cellift = 32'd1 */
wire _1316_;
wire [2:0] _1317_;
/* cellift = 32'd1 */
wire [2:0] _1318_;
wire [2:0] _1319_;
wire _1320_;
/* cellift = 32'd1 */
wire _1321_;
wire _1322_;
/* cellift = 32'd1 */
wire _1323_;
wire _1324_;
/* cellift = 32'd1 */
wire _1325_;
wire _1326_;
wire _1327_;
/* cellift = 32'd1 */
wire _1328_;
wire [31:0] _1329_;
/* cellift = 32'd1 */
wire [31:0] _1330_;
wire _1331_;
/* cellift = 32'd1 */
wire _1332_;
wire _1333_;
/* cellift = 32'd1 */
wire _1334_;
wire [6:0] _1335_;
/* cellift = 32'd1 */
wire [6:0] _1336_;
wire [1:0] _1337_;
wire _1338_;
/* cellift = 32'd1 */
wire _1339_;
/* src = "generated/sv2v_out.v:12437.30-12437.50" */
wire _1340_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12437.30-12437.50" */
wire _1341_;
/* src = "generated/sv2v_out.v:12437.72-12437.92" */
wire _1342_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12437.72-12437.92" */
wire _1343_;
/* src = "generated/sv2v_out.v:12557.9-12557.69" */
wire _1344_;
/* src = "generated/sv2v_out.v:12559.10-12559.32" */
wire _1345_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12559.10-12559.32" */
wire _1346_;
/* src = "generated/sv2v_out.v:12559.9-12559.51" */
wire _1347_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12559.9-12559.51" */
wire _1348_;
/* src = "generated/sv2v_out.v:12576.10-12576.31" */
wire _1349_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12576.10-12576.31" */
wire _1350_;
/* src = "generated/sv2v_out.v:12610.9-12610.43" */
wire _1351_;
/* src = "generated/sv2v_out.v:12682.38-12682.73" */
wire _1352_;
/* src = "generated/sv2v_out.v:12682.9-12682.74" */
wire _1353_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12682.9-12682.74" */
wire _1354_;
/* src = "generated/sv2v_out.v:12404.25-12404.38" */
wire _1355_;
/* src = "generated/sv2v_out.v:12559.10-12559.16" */
wire _1356_;
/* src = "generated/sv2v_out.v:12559.20-12559.32" */
wire _1357_;
/* src = "generated/sv2v_out.v:12559.37-12559.51" */
wire _1358_;
/* src = "generated/sv2v_out.v:12576.20-12576.31" */
wire _1359_;
/* src = "generated/sv2v_out.v:12610.30-12610.43" */
wire _1360_;
/* src = "generated/sv2v_out.v:12682.36-12682.74" */
wire _1361_;
/* src = "generated/sv2v_out.v:12524.12-12524.35" */
wire _1362_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12524.12-12524.35" */
wire _1363_;
/* src = "generated/sv2v_out.v:12524.11-12524.51" */
wire _1364_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12524.11-12524.51" */
wire _1365_;
/* src = "generated/sv2v_out.v:12524.10-12524.68" */
wire _1366_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12524.10-12524.68" */
wire _1367_;
/* src = "generated/sv2v_out.v:12524.9-12524.92" */
wire _1368_;
/* src = "generated/sv2v_out.v:12549.9-12549.35" */
wire _1369_;
/* src = "generated/sv2v_out.v:12557.10-12557.40" */
wire _1370_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12557.10-12557.40" */
wire _1371_;
/* src = "generated/sv2v_out.v:12557.46-12557.68" */
wire _1372_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12557.46-12557.68" */
wire _1373_;
/* src = "generated/sv2v_out.v:12623.10-12623.34" */
wire _1374_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12623.10-12623.34" */
wire _1375_;
/* src = "generated/sv2v_out.v:12623.9-12623.49" */
wire _1376_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12623.9-12623.49" */
wire _1377_;
/* src = "generated/sv2v_out.v:12335.44-12335.63" */
wire _1378_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12335.44-12335.63" */
wire _1379_;
/* src = "generated/sv2v_out.v:12582.15-12582.52" */
wire _1380_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12582.15-12582.52" */
wire _1381_;
/* src = "generated/sv2v_out.v:12342.41-12342.52" */
wire _1382_;
/* src = "generated/sv2v_out.v:12412.80-12412.108" */
wire _1383_;
/* src = "generated/sv2v_out.v:12697.35-12697.43" */
wire _1384_;
/* src = "generated/sv2v_out.v:12698.31-12698.51" */
wire _1385_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12698.31-12698.51" */
wire _1386_;
/* src = "generated/sv2v_out.v:12336.24-12336.46" */
wire _1387_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12336.24-12336.46" */
wire _1388_;
/* src = "generated/sv2v_out.v:12336.23-12336.64" */
wire _1389_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12336.23-12336.64" */
wire _1390_;
/* src = "generated/sv2v_out.v:12336.22-12336.83" */
wire _1391_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12336.22-12336.83" */
wire _1392_;
/* src = "generated/sv2v_out.v:12340.35-12340.56" */
wire _1393_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12340.35-12340.56" */
wire _1394_;
/* src = "generated/sv2v_out.v:12340.34-12340.69" */
wire _1395_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12340.34-12340.69" */
wire _1396_;
/* src = "generated/sv2v_out.v:12435.36-12435.66" */
wire _1397_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12435.36-12435.66" */
wire _1398_;
/* src = "generated/sv2v_out.v:12440.80-12440.118" */
wire _1399_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12440.80-12440.118" */
wire _1400_;
wire _1401_;
wire [31:0] _1402_;
/* cellift = 32'd1 */
wire [31:0] _1403_;
/* cellift = 32'd1 */
wire [31:0] _1404_;
/* cellift = 32'd1 */
wire [31:0] _1405_;
wire [31:0] _1406_;
/* cellift = 32'd1 */
wire [31:0] _1407_;
wire [31:0] _1408_;
/* cellift = 32'd1 */
wire [31:0] _1409_;
wire [6:0] _1410_;
wire [6:0] _1411_;
/* cellift = 32'd1 */
wire [6:0] _1412_;
wire [6:0] _1413_;
/* cellift = 32'd1 */
wire [6:0] _1414_;
wire [6:0] _1415_;
/* cellift = 32'd1 */
wire [6:0] _1416_;
wire [6:0] _1417_;
/* cellift = 32'd1 */
wire [6:0] _1418_;
wire [3:0] _1419_;
/* cellift = 32'd1 */
wire [3:0] _1420_;
wire [3:0] _1421_;
/* cellift = 32'd1 */
wire [3:0] _1422_;
wire [3:0] _1423_;
/* cellift = 32'd1 */
wire [3:0] _1424_;
wire _1425_;
/* cellift = 32'd1 */
wire _1426_;
wire _1427_;
/* cellift = 32'd1 */
wire _1428_;
wire _1429_;
/* cellift = 32'd1 */
wire _1430_;
wire _1431_;
/* cellift = 32'd1 */
wire _1432_;
wire _1433_;
/* cellift = 32'd1 */
wire _1434_;
wire _1435_;
wire _1436_;
/* cellift = 32'd1 */
wire _1437_;
wire _1438_;
/* cellift = 32'd1 */
wire _1439_;
wire _1440_;
wire _1441_;
wire _1442_;
/* cellift = 32'd1 */
wire _1443_;
wire _1444_;
/* src = "generated/sv2v_out.v:12437.72-12437.117" */
wire _1445_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12437.72-12437.117" */
wire _1446_;
/* src = "generated/sv2v_out.v:12451.119-12451.149" */
wire [2:0] _1447_;
/* src = "generated/sv2v_out.v:12451.97-12451.150" */
wire [2:0] _1448_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12451.97-12451.150" */
wire [2:0] _1449_;
/* src = "generated/sv2v_out.v:12451.52-12451.151" */
wire [2:0] _1450_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12451.52-12451.151" */
wire [2:0] _1451_;
/* src = "generated/sv2v_out.v:12577.22-12577.87" */
wire [6:0] _1452_;
/* src = "generated/sv2v_out.v:12626.22-12626.48" */
wire [1:0] _1453_;
/* src = "generated/sv2v_out.v:12638.23-12638.74" */
wire [31:0] _1454_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12638.23-12638.74" */
wire [31:0] _1455_;
/* src = "generated/sv2v_out.v:12642.23-12642.99" */
wire [31:0] _1456_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12642.23-12642.99" */
wire [31:0] _1457_;
/* src = "generated/sv2v_out.v:12644.39-12644.119" */
wire [6:0] _1458_;
/* src = "generated/sv2v_out.v:12244.13-12244.29" */
input branch_not_set_i;
wire branch_not_set_i;
/* cellift = 32'd1 */
input branch_not_set_i_t0;
wire branch_not_set_i_t0;
/* src = "generated/sv2v_out.v:12243.13-12243.25" */
input branch_set_i;
wire branch_set_i;
/* cellift = 32'd1 */
input branch_set_i_t0;
wire branch_set_i_t0;
/* src = "generated/sv2v_out.v:12209.13-12209.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:12229.13-12229.29" */
output controller_run_o;
wire controller_run_o;
/* cellift = 32'd1 */
output controller_run_o_t0;
wire controller_run_o_t0;
/* src = "generated/sv2v_out.v:12246.13-12246.30" */
input csr_mstatus_mie_i;
wire csr_mstatus_mie_i;
/* cellift = 32'd1 */
input csr_mstatus_mie_i_t0;
wire csr_mstatus_mie_i_t0;
/* src = "generated/sv2v_out.v:12266.20-12266.31" */
output [31:0] csr_mtval_o;
wire [31:0] csr_mtval_o;
/* cellift = 32'd1 */
output [31:0] csr_mtval_o_t0;
wire [31:0] csr_mtval_o_t0;
/* src = "generated/sv2v_out.v:12324.7-12324.21" */
wire csr_pipe_flush;
/* src = "generated/sv2v_out.v:12218.13-12218.29" */
input csr_pipe_flush_i;
wire csr_pipe_flush_i;
/* cellift = 32'd1 */
input csr_pipe_flush_i_t0;
wire csr_pipe_flush_i_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12324.7-12324.21" */
wire csr_pipe_flush_t0;
/* src = "generated/sv2v_out.v:12264.13-12264.34" */
output csr_restore_dret_id_o;
wire csr_restore_dret_id_o;
/* cellift = 32'd1 */
output csr_restore_dret_id_o_t0;
wire csr_restore_dret_id_o_t0;
/* src = "generated/sv2v_out.v:12263.13-12263.34" */
output csr_restore_mret_id_o;
wire csr_restore_mret_id_o;
/* cellift = 32'd1 */
output csr_restore_mret_id_o_t0;
wire csr_restore_mret_id_o_t0;
/* src = "generated/sv2v_out.v:12265.13-12265.29" */
output csr_save_cause_o;
wire csr_save_cause_o;
/* cellift = 32'd1 */
output csr_save_cause_o_t0;
wire csr_save_cause_o_t0;
/* src = "generated/sv2v_out.v:12261.13-12261.26" */
output csr_save_id_o;
wire csr_save_id_o;
/* cellift = 32'd1 */
output csr_save_id_o_t0;
wire csr_save_id_o_t0;
/* src = "generated/sv2v_out.v:12260.13-12260.26" */
output csr_save_if_o;
wire csr_save_if_o;
/* cellift = 32'd1 */
output csr_save_if_o_t0;
wire csr_save_if_o_t0;
/* src = "generated/sv2v_out.v:12262.13-12262.26" */
output csr_save_wb_o;
wire csr_save_wb_o;
/* cellift = 32'd1 */
output csr_save_wb_o_t0;
wire csr_save_wb_o_t0;
/* src = "generated/sv2v_out.v:12211.13-12211.24" */
output ctrl_busy_o;
wire ctrl_busy_o;
/* cellift = 32'd1 */
output ctrl_busy_o_t0;
wire ctrl_busy_o_t0;
/* src = "generated/sv2v_out.v:12274.12-12274.23" */
reg [3:0] ctrl_fsm_cs;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12274.12-12274.23" */
reg [3:0] ctrl_fsm_cs_t0;
/* src = "generated/sv2v_out.v:12275.12-12275.23" */
wire [3:0] ctrl_fsm_ns;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12275.12-12275.23" */
wire [3:0] ctrl_fsm_ns_t0;
/* src = "generated/sv2v_out.v:12280.13-12280.26" */
wire [2:0] debug_cause_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12280.13-12280.26" */
wire [2:0] debug_cause_d_t0;
/* src = "generated/sv2v_out.v:12252.20-12252.33" */
output [2:0] debug_cause_o;
reg [2:0] debug_cause_o;
/* cellift = 32'd1 */
output [2:0] debug_cause_o_t0;
reg [2:0] debug_cause_o_t0;
/* src = "generated/sv2v_out.v:12253.13-12253.29" */
output debug_csr_save_o;
wire debug_csr_save_o;
/* cellift = 32'd1 */
output debug_csr_save_o_t0;
wire debug_csr_save_o_t0;
/* src = "generated/sv2v_out.v:12257.13-12257.28" */
input debug_ebreakm_i;
wire debug_ebreakm_i;
/* cellift = 32'd1 */
input debug_ebreakm_i_t0;
wire debug_ebreakm_i_t0;
/* src = "generated/sv2v_out.v:12258.13-12258.28" */
input debug_ebreaku_i;
wire debug_ebreaku_i;
/* cellift = 32'd1 */
input debug_ebreaku_i_t0;
wire debug_ebreaku_i_t0;
/* src = "generated/sv2v_out.v:12279.6-12279.18" */
wire debug_mode_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12279.6-12279.18" */
wire debug_mode_d_t0;
/* src = "generated/sv2v_out.v:12255.13-12255.34" */
output debug_mode_entering_o;
wire debug_mode_entering_o;
/* cellift = 32'd1 */
output debug_mode_entering_o_t0;
wire debug_mode_entering_o_t0;
/* src = "generated/sv2v_out.v:12254.14-12254.26" */
output debug_mode_o;
reg debug_mode_o;
/* cellift = 32'd1 */
output debug_mode_o_t0;
reg debug_mode_o_t0;
/* src = "generated/sv2v_out.v:12251.13-12251.24" */
input debug_req_i;
wire debug_req_i;
/* cellift = 32'd1 */
input debug_req_i_t0;
wire debug_req_i_t0;
/* src = "generated/sv2v_out.v:12256.13-12256.32" */
input debug_single_step_i;
wire debug_single_step_i;
/* cellift = 32'd1 */
input debug_single_step_i_t0;
wire debug_single_step_i_t0;
/* src = "generated/sv2v_out.v:12304.7-12304.23" */
wire do_single_step_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12304.7-12304.23" */
wire do_single_step_d_t0;
/* src = "generated/sv2v_out.v:12305.6-12305.22" */
reg do_single_step_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12305.6-12305.22" */
reg do_single_step_q_t0;
/* src = "generated/sv2v_out.v:12321.7-12321.16" */
wire dret_insn;
/* src = "generated/sv2v_out.v:12215.13-12215.24" */
input dret_insn_i;
wire dret_insn_i;
/* cellift = 32'd1 */
input dret_insn_i_t0;
wire dret_insn_i_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12321.7-12321.16" */
wire dret_insn_t0;
/* src = "generated/sv2v_out.v:12309.7-12309.24" */
wire ebreak_into_debug;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12309.7-12309.24" */
wire ebreak_into_debug_t0;
/* src = "generated/sv2v_out.v:12323.7-12323.16" */
wire ebrk_insn;
/* src = "generated/sv2v_out.v:12217.13-12217.24" */
input ebrk_insn_i;
wire ebrk_insn_i;
/* cellift = 32'd1 */
input ebrk_insn_i_t0;
wire ebrk_insn_i_t0;
/* src = "generated/sv2v_out.v:12293.6-12293.20" */
wire ebrk_insn_prio;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12293.6-12293.20" */
wire ebrk_insn_prio_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12323.7-12323.16" */
wire ebrk_insn_t0;
/* src = "generated/sv2v_out.v:12319.7-12319.17" */
wire ecall_insn;
/* src = "generated/sv2v_out.v:12213.13-12213.25" */
input ecall_insn_i;
wire ecall_insn_i;
/* cellift = 32'd1 */
input ecall_insn_i_t0;
wire ecall_insn_i_t0;
/* src = "generated/sv2v_out.v:12292.6-12292.21" */
wire ecall_insn_prio;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12292.6-12292.21" */
wire ecall_insn_prio_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12319.7-12319.17" */
wire ecall_insn_t0;
/* src = "generated/sv2v_out.v:12308.7-12308.23" */
wire enter_debug_mode;
/* src = "generated/sv2v_out.v:12306.7-12306.30" */
wire enter_debug_mode_prio_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12306.7-12306.30" */
wire enter_debug_mode_prio_d_t0;
/* src = "generated/sv2v_out.v:12307.6-12307.29" */
reg enter_debug_mode_prio_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12307.6-12307.29" */
reg enter_debug_mode_prio_q_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12308.7-12308.23" */
wire enter_debug_mode_t0;
/* src = "generated/sv2v_out.v:12236.19-12236.30" */
output [6:0] exc_cause_o;
wire [6:0] exc_cause_o;
/* cellift = 32'd1 */
output [6:0] exc_cause_o_t0;
wire [6:0] exc_cause_o_t0;
/* src = "generated/sv2v_out.v:12235.19-12235.31" */
output [1:0] exc_pc_mux_o;
wire [1:0] exc_pc_mux_o;
/* cellift = 32'd1 */
output [1:0] exc_pc_mux_o_t0;
wire [1:0] exc_pc_mux_o_t0;
/* src = "generated/sv2v_out.v:12300.7-12300.18" */
wire exc_req_lsu;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12300.7-12300.18" */
wire exc_req_lsu_t0;
/* src = "generated/sv2v_out.v:12286.6-12286.15" */
reg exc_req_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12286.6-12286.15" */
reg exc_req_q_t0;
/* src = "generated/sv2v_out.v:12270.14-12270.24" */
output flush_id_o;
wire flush_id_o;
/* cellift = 32'd1 */
output flush_id_o_t0;
wire flush_id_o_t0;
/* src = "generated/sv2v_out.v:12397.9-12397.21" */
wire \g_intg_irq_int.entering_nmi ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12397.9-12397.21" */
wire \g_intg_irq_int.entering_nmi_t0 ;
/* src = "generated/sv2v_out.v:12393.15-12393.39" */
reg [31:0] \g_intg_irq_int.mem_resp_intg_err_addr_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12393.15-12393.39" */
reg [31:0] \g_intg_irq_int.mem_resp_intg_err_addr_q_t0 ;
/* src = "generated/sv2v_out.v:12396.8-12396.35" */
wire \g_intg_irq_int.mem_resp_intg_err_irq_clear ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12396.8-12396.35" */
wire \g_intg_irq_int.mem_resp_intg_err_irq_clear_t0 ;
/* src = "generated/sv2v_out.v:12392.9-12392.40" */
wire \g_intg_irq_int.mem_resp_intg_err_irq_pending_d ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12392.9-12392.40" */
wire \g_intg_irq_int.mem_resp_intg_err_irq_pending_d_t0 ;
/* src = "generated/sv2v_out.v:12391.8-12391.39" */
reg \g_intg_irq_int.mem_resp_intg_err_irq_pending_q ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12391.8-12391.39" */
reg \g_intg_irq_int.mem_resp_intg_err_irq_pending_q_t0 ;
/* src = "generated/sv2v_out.v:12395.8-12395.33" */
wire \g_intg_irq_int.mem_resp_intg_err_irq_set ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12395.8-12395.33" */
wire \g_intg_irq_int.mem_resp_intg_err_irq_set_t0 ;
/* src = "generated/sv2v_out.v:12297.6-12297.13" */
wire halt_if;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12297.6-12297.13" */
wire halt_if_t0;
/* src = "generated/sv2v_out.v:12311.7-12311.17" */
wire handle_irq;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12311.7-12311.17" */
wire handle_irq_t0;
/* src = "generated/sv2v_out.v:12242.14-12242.28" */
output id_exception_o;
wire id_exception_o;
/* cellift = 32'd1 */
output id_exception_o_t0;
wire id_exception_o_t0;
/* src = "generated/sv2v_out.v:12228.14-12228.27" */
output id_in_ready_o;
wire id_in_ready_o;
/* cellift = 32'd1 */
output id_in_ready_o_t0;
wire id_in_ready_o_t0;
/* src = "generated/sv2v_out.v:12312.7-12312.20" */
wire id_wb_pending;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12312.7-12312.20" */
wire id_wb_pending_t0;
/* src = "generated/sv2v_out.v:12289.7-12289.21" */
wire illegal_insn_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12289.7-12289.21" */
wire illegal_insn_d_t0;
/* src = "generated/sv2v_out.v:12212.13-12212.27" */
input illegal_insn_i;
wire illegal_insn_i;
/* cellift = 32'd1 */
input illegal_insn_i_t0;
wire illegal_insn_i_t0;
/* src = "generated/sv2v_out.v:12291.6-12291.23" */
wire illegal_insn_prio;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12291.6-12291.23" */
wire illegal_insn_prio_t0;
/* src = "generated/sv2v_out.v:12288.6-12288.20" */
reg illegal_insn_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12288.6-12288.20" */
reg illegal_insn_q_t0;
/* src = "generated/sv2v_out.v:12223.13-12223.29" */
input instr_bp_taken_i;
wire instr_bp_taken_i;
/* cellift = 32'd1 */
input instr_bp_taken_i_t0;
wire instr_bp_taken_i_t0;
/* src = "generated/sv2v_out.v:12221.20-12221.38" */
input [15:0] instr_compressed_i;
wire [15:0] instr_compressed_i;
/* cellift = 32'd1 */
input [15:0] instr_compressed_i_t0;
wire [15:0] instr_compressed_i_t0;
/* src = "generated/sv2v_out.v:12230.13-12230.25" */
input instr_exec_i;
wire instr_exec_i;
/* cellift = 32'd1 */
input instr_exec_i_t0;
wire instr_exec_i_t0;
/* src = "generated/sv2v_out.v:12325.7-12325.22" */
wire instr_fetch_err;
/* src = "generated/sv2v_out.v:12224.13-12224.30" */
input instr_fetch_err_i;
wire instr_fetch_err_i;
/* cellift = 32'd1 */
input instr_fetch_err_i_t0;
wire instr_fetch_err_i_t0;
/* src = "generated/sv2v_out.v:12225.13-12225.36" */
input instr_fetch_err_plus2_i;
wire instr_fetch_err_plus2_i;
/* cellift = 32'd1 */
input instr_fetch_err_plus2_i_t0;
wire instr_fetch_err_plus2_i_t0;
/* src = "generated/sv2v_out.v:12290.6-12290.26" */
wire instr_fetch_err_prio;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12290.6-12290.26" */
wire instr_fetch_err_prio_t0;
/* src = "generated/sv2v_out.v:12220.20-12220.27" */
input [31:0] instr_i;
wire [31:0] instr_i;
/* cellift = 32'd1 */
input [31:0] instr_i_t0;
wire [31:0] instr_i_t0;
/* src = "generated/sv2v_out.v:12222.13-12222.34" */
input instr_is_compressed_i;
wire instr_is_compressed_i;
/* cellift = 32'd1 */
input instr_is_compressed_i_t0;
wire instr_is_compressed_i_t0;
/* src = "generated/sv2v_out.v:12231.13-12231.24" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:12227.14-12227.33" */
output instr_valid_clear_o;
wire instr_valid_clear_o;
/* cellift = 32'd1 */
output instr_valid_clear_o_t0;
wire instr_valid_clear_o_t0;
/* src = "generated/sv2v_out.v:12219.13-12219.26" */
input instr_valid_i;
wire instr_valid_i;
/* cellift = 32'd1 */
input instr_valid_i_t0;
wire instr_valid_i_t0;
/* src = "generated/sv2v_out.v:12310.7-12310.18" */
wire irq_enabled;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12310.7-12310.18" */
wire irq_enabled_t0;
/* src = "generated/sv2v_out.v:12313.7-12313.13" */
wire irq_nm;
/* src = "generated/sv2v_out.v:12249.13-12249.25" */
input irq_nm_ext_i;
wire irq_nm_ext_i;
/* cellift = 32'd1 */
input irq_nm_ext_i_t0;
wire irq_nm_ext_i_t0;
/* src = "generated/sv2v_out.v:12314.7-12314.17" */
wire irq_nm_int;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12314.7-12314.17" */
wire irq_nm_int_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12313.7-12313.13" */
wire irq_nm_t0;
/* src = "generated/sv2v_out.v:12247.13-12247.26" */
input irq_pending_i;
wire irq_pending_i;
/* cellift = 32'd1 */
input irq_pending_i_t0;
wire irq_pending_i_t0;
/* src = "generated/sv2v_out.v:12248.20-12248.26" */
input [17:0] irqs_i;
wire [17:0] irqs_i;
/* cellift = 32'd1 */
input [17:0] irqs_i_t0;
wire [17:0] irqs_i_t0;
/* src = "generated/sv2v_out.v:12245.13-12245.23" */
input jump_set_i;
wire jump_set_i;
/* cellift = 32'd1 */
input jump_set_i_t0;
wire jump_set_i_t0;
/* src = "generated/sv2v_out.v:12238.13-12238.23" */
input load_err_i;
wire load_err_i;
/* cellift = 32'd1 */
input load_err_i_t0;
wire load_err_i_t0;
/* src = "generated/sv2v_out.v:12295.6-12295.19" */
wire load_err_prio;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12295.6-12295.19" */
wire load_err_prio_t0;
/* src = "generated/sv2v_out.v:12282.6-12282.16" */
reg load_err_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12282.6-12282.16" */
reg load_err_q_t0;
/* src = "generated/sv2v_out.v:12237.20-12237.35" */
input [31:0] lsu_addr_last_i;
wire [31:0] lsu_addr_last_i;
/* cellift = 32'd1 */
input [31:0] lsu_addr_last_i_t0;
wire [31:0] lsu_addr_last_i_t0;
/* src = "generated/sv2v_out.v:12240.13-12240.32" */
input mem_resp_intg_err_i;
wire mem_resp_intg_err_i;
/* cellift = 32'd1 */
input mem_resp_intg_err_i_t0;
wire mem_resp_intg_err_i_t0;
/* src = "generated/sv2v_out.v:12317.12-12317.19" */
wire [3:0] mfip_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12317.12-12317.19" */
wire [3:0] mfip_id_t0;
/* src = "generated/sv2v_out.v:12320.7-12320.16" */
wire mret_insn;
/* src = "generated/sv2v_out.v:12214.13-12214.24" */
input mret_insn_i;
wire mret_insn_i;
/* cellift = 32'd1 */
input mret_insn_i_t0;
wire mret_insn_i_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12320.7-12320.16" */
wire mret_insn_t0;
/* src = "generated/sv2v_out.v:12277.6-12277.16" */
wire nmi_mode_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12277.6-12277.16" */
wire nmi_mode_d_t0;
/* src = "generated/sv2v_out.v:12250.14-12250.24" */
output nmi_mode_o;
reg nmi_mode_o;
/* cellift = 32'd1 */
output nmi_mode_o_t0;
reg nmi_mode_o_t0;
/* src = "generated/sv2v_out.v:12234.13-12234.35" */
output nt_branch_mispredict_o;
wire nt_branch_mispredict_o;
/* cellift = 32'd1 */
output nt_branch_mispredict_o_t0;
wire nt_branch_mispredict_o_t0;
/* src = "generated/sv2v_out.v:12226.20-12226.27" */
input [31:0] pc_id_i;
wire [31:0] pc_id_i;
/* cellift = 32'd1 */
input [31:0] pc_id_i_t0;
wire [31:0] pc_id_i_t0;
/* src = "generated/sv2v_out.v:12233.19-12233.27" */
output [2:0] pc_mux_o;
wire [2:0] pc_mux_o;
/* cellift = 32'd1 */
output [2:0] pc_mux_o_t0;
wire [2:0] pc_mux_o_t0;
/* src = "generated/sv2v_out.v:12232.13-12232.21" */
output pc_set_o;
wire pc_set_o;
/* cellift = 32'd1 */
output pc_set_o_t0;
wire pc_set_o_t0;
/* src = "generated/sv2v_out.v:12272.13-12272.24" */
output perf_jump_o;
wire perf_jump_o;
/* cellift = 32'd1 */
output perf_jump_o_t0;
wire perf_jump_o_t0;
/* src = "generated/sv2v_out.v:12273.13-12273.27" */
output perf_tbranch_o;
wire perf_tbranch_o;
/* cellift = 32'd1 */
output perf_tbranch_o_t0;
wire perf_tbranch_o_t0;
/* src = "generated/sv2v_out.v:12267.19-12267.30" */
input [1:0] priv_mode_i;
wire [1:0] priv_mode_i;
/* cellift = 32'd1 */
input [1:0] priv_mode_i_t0;
wire [1:0] priv_mode_i_t0;
/* src = "generated/sv2v_out.v:12271.13-12271.23" */
input ready_wb_i;
wire ready_wb_i;
/* cellift = 32'd1 */
input ready_wb_i_t0;
wire ready_wb_i_t0;
/* src = "generated/sv2v_out.v:12298.6-12298.15" */
wire retain_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12298.6-12298.15" */
wire retain_id_t0;
/* src = "generated/sv2v_out.v:12210.13-12210.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:12301.7-12301.18" */
wire special_req;
/* src = "generated/sv2v_out.v:12303.7-12303.29" */
wire special_req_flush_only;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12303.7-12303.29" */
wire special_req_flush_only_t0;
/* src = "generated/sv2v_out.v:12302.7-12302.28" */
wire special_req_pc_change;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12302.7-12302.28" */
wire special_req_pc_change_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12301.7-12301.18" */
wire special_req_t0;
/* src = "generated/sv2v_out.v:12296.7-12296.12" */
wire stall;
/* src = "generated/sv2v_out.v:12268.13-12268.23" */
input stall_id_i;
wire stall_id_i;
/* cellift = 32'd1 */
input stall_id_i_t0;
wire stall_id_i_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12296.7-12296.12" */
wire stall_t0;
/* src = "generated/sv2v_out.v:12269.13-12269.23" */
input stall_wb_i;
wire stall_wb_i;
/* cellift = 32'd1 */
input stall_wb_i_t0;
wire stall_wb_i_t0;
/* src = "generated/sv2v_out.v:12239.13-12239.24" */
input store_err_i;
wire store_err_i;
/* cellift = 32'd1 */
input store_err_i_t0;
wire store_err_i_t0;
/* src = "generated/sv2v_out.v:12294.6-12294.20" */
wire store_err_prio;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12294.6-12294.20" */
wire store_err_prio_t0;
/* src = "generated/sv2v_out.v:12284.6-12284.17" */
reg store_err_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12284.6-12284.17" */
reg store_err_q_t0;
/* src = "generated/sv2v_out.v:12259.13-12259.28" */
input trigger_match_i;
wire trigger_match_i;
/* cellift = 32'd1 */
input trigger_match_i_t0;
wire trigger_match_i_t0;
/* src = "generated/sv2v_out.v:12241.14-12241.28" */
output wb_exception_o;
wire wb_exception_o;
/* cellift = 32'd1 */
output wb_exception_o_t0;
wire wb_exception_o_t0;
/* src = "generated/sv2v_out.v:12322.7-12322.15" */
wire wfi_insn;
/* src = "generated/sv2v_out.v:12216.13-12216.23" */
input wfi_insn_i;
wire wfi_insn_i;
/* cellift = 32'd1 */
input wfi_insn_i_t0;
wire wfi_insn_i_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12322.7-12322.15" */
wire wfi_insn_t0;
assign _0169_ = pc_id_i + /* src = "generated/sv2v_out.v:12638.49-12638.64" */ 32'd2;
assign ecall_insn = ecall_insn_i & /* src = "generated/sv2v_out.v:12328.22-12328.50" */ instr_valid_i;
assign mret_insn = mret_insn_i & /* src = "generated/sv2v_out.v:12329.21-12329.48" */ instr_valid_i;
assign dret_insn = dret_insn_i & /* src = "generated/sv2v_out.v:12330.21-12330.48" */ instr_valid_i;
assign wfi_insn = wfi_insn_i & /* src = "generated/sv2v_out.v:12331.20-12331.46" */ instr_valid_i;
assign ebrk_insn = ebrk_insn_i & /* src = "generated/sv2v_out.v:12332.21-12332.48" */ instr_valid_i;
assign csr_pipe_flush = csr_pipe_flush_i & /* src = "generated/sv2v_out.v:12333.26-12333.58" */ instr_valid_i;
assign instr_fetch_err = instr_fetch_err_i & /* src = "generated/sv2v_out.v:12334.27-12334.60" */ instr_valid_i;
assign illegal_insn_d = illegal_insn_i & /* src = "generated/sv2v_out.v:12335.26-12335.64" */ _1378_;
assign id_exception_o = _1391_ & /* src = "generated/sv2v_out.v:12336.21-12336.108" */ _1378_;
assign \g_intg_irq_int.entering_nmi  = nmi_mode_d & /* src = "generated/sv2v_out.v:12398.26-12398.50" */ _0337_;
assign _0171_ = \g_intg_irq_int.entering_nmi  & /* src = "generated/sv2v_out.v:12404.10-12404.38" */ _1355_;
assign _0172_ = \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  & /* src = "generated/sv2v_out.v:12412.46-12412.108" */ _1383_;
assign _0174_ = _0248_ & /* src = "generated/sv2v_out.v:12434.45-12434.80" */ debug_single_step_i;
assign enter_debug_mode_prio_d = _1397_ & /* src = "generated/sv2v_out.v:12435.35-12435.83" */ _0248_;
assign _0176_ = trigger_match_i & /* src = "generated/sv2v_out.v:12436.55-12436.86" */ _0248_;
assign _0178_ = _0248_ & /* src = "generated/sv2v_out.v:12440.24-12440.60" */ _0249_;
assign _0180_ = _0178_ & /* src = "generated/sv2v_out.v:12440.23-12440.75" */ _0337_;
assign _0182_ = irq_pending_i & /* src = "generated/sv2v_out.v:12440.90-12440.117" */ irq_enabled;
assign handle_irq = _0180_ & /* src = "generated/sv2v_out.v:12440.22-12440.119" */ _1399_;
assign _0184_ = ebrk_insn_prio & /* src = "generated/sv2v_out.v:12451.52-12451.86" */ ebreak_into_debug;
assign _0186_ = irq_nm_int & /* src = "generated/sv2v_out.v:12578.11-12578.37" */ _1355_;
assign _0188_ = _0243_ & /* src = "generated/sv2v_out.v:12697.26-12697.43" */ _1384_;
assign id_in_ready_o = _0188_ & /* src = "generated/sv2v_out.v:12697.25-12697.57" */ _0419_;
assign _0190_ = ~ pc_id_i_t0;
assign _0457_ = pc_id_i & _0190_;
assign _1295_ = _0457_ + 32'd2;
assign _0978_ = pc_id_i | pc_id_i_t0;
assign _1296_ = _0978_ + 32'd2;
assign _1227_ = _1295_ ^ _1296_;
assign _0170_ = _1227_ | pc_id_i_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_intg_irq_int.mem_resp_intg_err_irq_pending_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_intg_irq_int.mem_resp_intg_err_irq_pending_q_t0  <= 1'h0;
else \g_intg_irq_int.mem_resp_intg_err_irq_pending_q_t0  <= \g_intg_irq_int.mem_resp_intg_err_irq_pending_d_t0 ;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME nmi_mode_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) nmi_mode_o_t0 <= 1'h0;
else nmi_mode_o_t0 <= nmi_mode_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME load_err_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) load_err_q_t0 <= 1'h0;
else load_err_q_t0 <= load_err_i_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME store_err_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) store_err_q_t0 <= 1'h0;
else store_err_q_t0 <= store_err_i_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME exc_req_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) exc_req_q_t0 <= 1'h0;
else exc_req_q_t0 <= id_exception_o_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME illegal_insn_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) illegal_insn_q_t0 <= 1'h0;
else illegal_insn_q_t0 <= illegal_insn_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME do_single_step_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) do_single_step_q_t0 <= 1'h0;
else do_single_step_q_t0 <= do_single_step_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME enter_debug_mode_prio_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) enter_debug_mode_prio_q_t0 <= 1'h0;
else enter_debug_mode_prio_q_t0 <= enter_debug_mode_prio_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME debug_cause_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) debug_cause_o_t0 <= 3'h0;
else debug_cause_o_t0 <= debug_cause_d_t0;
assign _0191_ = ~ _0442_;
assign _0192_ = ~ _0444_;
assign _0193_ = ~ _0446_;
assign _1228_ = debug_mode_d ^ debug_mode_o;
assign _1229_ = ctrl_fsm_ns ^ ctrl_fsm_cs;
assign _1230_ = lsu_addr_last_i ^ \g_intg_irq_int.mem_resp_intg_err_addr_q ;
assign _1002_ = debug_mode_d_t0 | debug_mode_o_t0;
assign _1006_ = ctrl_fsm_ns_t0 | ctrl_fsm_cs_t0;
assign _1010_ = lsu_addr_last_i_t0 | \g_intg_irq_int.mem_resp_intg_err_addr_q_t0 ;
assign _1003_ = _1228_ | _1002_;
assign _1007_ = _1229_ | _1006_;
assign _1011_ = _1230_ | _1010_;
assign _0525_ = _0442_ & debug_mode_d_t0;
assign _0528_ = { _0444_, _0444_, _0444_, _0444_ } & ctrl_fsm_ns_t0;
assign _0531_ = { _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_, _0446_ } & lsu_addr_last_i_t0;
assign _0526_ = _0191_ & debug_mode_o_t0;
assign _0529_ = { _0192_, _0192_, _0192_, _0192_ } & ctrl_fsm_cs_t0;
assign _0532_ = { _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_, _0193_ } & \g_intg_irq_int.mem_resp_intg_err_addr_q_t0 ;
assign _0527_ = _1003_ & _0443_;
assign _0530_ = _1007_ & { _0445_, _0445_, _0445_, _0445_ };
assign _0533_ = _1011_ & { _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_, _0447_ };
assign _1004_ = _0525_ | _0526_;
assign _1008_ = _0528_ | _0529_;
assign _1012_ = _0531_ | _0532_;
assign _1005_ = _1004_ | _0527_;
assign _1009_ = _1008_ | _0530_;
assign _1013_ = _1012_ | _0533_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME debug_mode_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) debug_mode_o_t0 <= 1'h0;
else debug_mode_o_t0 <= _1005_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME ctrl_fsm_cs_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) ctrl_fsm_cs_t0 <= 4'h0;
else ctrl_fsm_cs_t0 <= _1009_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_intg_irq_int.mem_resp_intg_err_addr_q_t0  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_intg_irq_int.mem_resp_intg_err_addr_q_t0  <= 32'd0;
else \g_intg_irq_int.mem_resp_intg_err_addr_q_t0  <= _1013_;
assign _0458_ = ecall_insn_i_t0 & instr_valid_i;
assign _0461_ = mret_insn_i_t0 & instr_valid_i;
assign _0464_ = dret_insn_i_t0 & instr_valid_i;
assign _0467_ = wfi_insn_i_t0 & instr_valid_i;
assign _0470_ = ebrk_insn_i_t0 & instr_valid_i;
assign _0473_ = csr_pipe_flush_i_t0 & instr_valid_i;
assign _0476_ = instr_fetch_err_i_t0 & instr_valid_i;
assign _0479_ = illegal_insn_i_t0 & _1378_;
assign _0482_ = _1392_ & _1378_;
assign _0485_ = nmi_mode_d_t0 & _0337_;
assign _0488_ = \g_intg_irq_int.entering_nmi_t0  & _1355_;
assign _0491_ = \g_intg_irq_int.mem_resp_intg_err_irq_pending_q_t0  & _1383_;
assign _0494_ = debug_mode_o_t0 & debug_single_step_i;
assign _0497_ = _1398_ & _0248_;
assign _0500_ = trigger_match_i_t0 & _0248_;
assign _0503_ = debug_mode_o_t0 & _0249_;
assign _0504_ = _0179_ & _0337_;
assign _0507_ = irq_pending_i_t0 & irq_enabled;
assign _0510_ = _0181_ & _1399_;
assign _0516_ = irq_nm_int_t0 & _1355_;
assign _0519_ = stall_t0 & _1384_;
assign _0522_ = _0189_ & _0419_;
assign _0459_ = instr_valid_i_t0 & ecall_insn_i;
assign _0462_ = instr_valid_i_t0 & mret_insn_i;
assign _0465_ = instr_valid_i_t0 & dret_insn_i;
assign _0468_ = instr_valid_i_t0 & wfi_insn_i;
assign _0471_ = instr_valid_i_t0 & ebrk_insn_i;
assign _0474_ = instr_valid_i_t0 & csr_pipe_flush_i;
assign _0477_ = instr_valid_i_t0 & instr_fetch_err_i;
assign _0480_ = _1379_ & illegal_insn_i;
assign _0483_ = _1379_ & _1391_;
assign _0486_ = nmi_mode_o_t0 & nmi_mode_d;
assign _0489_ = irq_nm_ext_i_t0 & \g_intg_irq_int.entering_nmi ;
assign _0492_ = \g_intg_irq_int.mem_resp_intg_err_irq_clear_t0  & \g_intg_irq_int.mem_resp_intg_err_irq_pending_q ;
assign _0495_ = debug_single_step_i_t0 & _0248_;
assign _0498_ = debug_mode_o_t0 & _1397_;
assign _0501_ = debug_mode_o_t0 & trigger_match_i;
assign _0505_ = nmi_mode_o_t0 & _0178_;
assign _0508_ = irq_enabled_t0 & irq_pending_i;
assign _0511_ = _1400_ & _0180_;
assign _0517_ = irq_nm_ext_i_t0 & irq_nm_int;
assign _0520_ = halt_if_t0 & _0243_;
assign _0523_ = retain_id_t0 & _0188_;
assign _0460_ = ecall_insn_i_t0 & instr_valid_i_t0;
assign _0463_ = mret_insn_i_t0 & instr_valid_i_t0;
assign _0466_ = dret_insn_i_t0 & instr_valid_i_t0;
assign _0469_ = wfi_insn_i_t0 & instr_valid_i_t0;
assign _0472_ = ebrk_insn_i_t0 & instr_valid_i_t0;
assign _0475_ = csr_pipe_flush_i_t0 & instr_valid_i_t0;
assign _0478_ = instr_fetch_err_i_t0 & instr_valid_i_t0;
assign _0481_ = illegal_insn_i_t0 & _1379_;
assign _0484_ = _1392_ & _1379_;
assign _0487_ = nmi_mode_d_t0 & nmi_mode_o_t0;
assign _0490_ = \g_intg_irq_int.entering_nmi_t0  & irq_nm_ext_i_t0;
assign _0493_ = \g_intg_irq_int.mem_resp_intg_err_irq_pending_q_t0  & \g_intg_irq_int.mem_resp_intg_err_irq_clear_t0 ;
assign _0499_ = _1398_ & debug_mode_o_t0;
assign _0502_ = trigger_match_i_t0 & debug_mode_o_t0;
assign _0496_ = debug_mode_o_t0 & debug_single_step_i_t0;
assign _0506_ = _0179_ & nmi_mode_o_t0;
assign _0509_ = irq_pending_i_t0 & irq_enabled_t0;
assign _0512_ = _0181_ & _1400_;
assign _0515_ = ebrk_insn_prio_t0 & ebreak_into_debug_t0;
assign _0518_ = irq_nm_int_t0 & irq_nm_ext_i_t0;
assign _0521_ = stall_t0 & halt_if_t0;
assign _0524_ = _0189_ & retain_id_t0;
assign _0979_ = _0458_ | _0459_;
assign _0980_ = _0461_ | _0462_;
assign _0981_ = _0464_ | _0465_;
assign _0982_ = _0467_ | _0468_;
assign _0983_ = _0470_ | _0471_;
assign _0984_ = _0473_ | _0474_;
assign _0985_ = _0476_ | _0477_;
assign _0986_ = _0479_ | _0480_;
assign _0987_ = _0482_ | _0483_;
assign _0988_ = _0485_ | _0486_;
assign _0989_ = _0488_ | _0489_;
assign _0990_ = _0491_ | _0492_;
assign _0991_ = _0494_ | _0495_;
assign _0992_ = _0497_ | _0498_;
assign _0993_ = _0500_ | _0501_;
assign _0994_ = _0503_ | _0495_;
assign _0995_ = _0504_ | _0505_;
assign _0996_ = _0507_ | _0508_;
assign _0997_ = _0510_ | _0511_;
assign _0998_ = _0513_ | _0514_;
assign _0999_ = _0516_ | _0517_;
assign _1000_ = _0519_ | _0520_;
assign _1001_ = _0522_ | _0523_;
assign ecall_insn_t0 = _0979_ | _0460_;
assign mret_insn_t0 = _0980_ | _0463_;
assign dret_insn_t0 = _0981_ | _0466_;
assign wfi_insn_t0 = _0982_ | _0469_;
assign ebrk_insn_t0 = _0983_ | _0472_;
assign csr_pipe_flush_t0 = _0984_ | _0475_;
assign instr_fetch_err_prio_t0 = _0985_ | _0478_;
assign illegal_insn_d_t0 = _0986_ | _0481_;
assign id_exception_o_t0 = _0987_ | _0484_;
assign \g_intg_irq_int.entering_nmi_t0  = _0988_ | _0487_;
assign _0052_ = _0989_ | _0490_;
assign _0173_ = _0990_ | _0493_;
assign _0175_ = _0991_ | _0496_;
assign enter_debug_mode_prio_d_t0 = _0992_ | _0499_;
assign _0177_ = _0993_ | _0502_;
assign _0179_ = _0994_ | _0496_;
assign _0181_ = _0995_ | _0506_;
assign _0183_ = _0996_ | _0509_;
assign handle_irq_t0 = _0997_ | _0512_;
assign _0185_ = _0998_ | _0515_;
assign _0187_ = _0999_ | _0518_;
assign _0189_ = _1000_ | _0521_;
assign id_in_ready_o_t0 = _1001_ | _0524_;
assign _0194_ = | { _1377_, _1379_, mret_insn_t0, dret_insn_t0 };
assign _0195_ = | { _1377_, _1379_, mret_insn_t0 };
assign _0196_ = | { _1377_, _1379_ };
assign _0197_ = | { _1437_, enter_debug_mode_t0, handle_irq_t0, id_in_ready_o_t0 };
assign _0198_ = | { _0038_, _1439_ };
assign _0199_ = | priv_mode_i_t0;
assign _0200_ = | ctrl_fsm_cs_t0;
assign _0201_ = ~ { _1379_, _1377_, dret_insn_t0, mret_insn_t0 };
assign _0202_ = ~ { _1379_, _1377_, mret_insn_t0 };
assign _0203_ = ~ { _1379_, _1377_ };
assign _0204_ = ~ { _1437_, id_in_ready_o_t0, handle_irq_t0, enter_debug_mode_t0 };
assign _0205_ = ~ { _1439_, _0038_ };
assign _0206_ = ~ priv_mode_i_t0;
assign _0534_ = { _1401_, _1376_, dret_insn, mret_insn } & _0201_;
assign _0535_ = { _1401_, _1376_, mret_insn } & _0202_;
assign _0536_ = { _1401_, _1376_ } & _0203_;
assign _0538_ = { _1436_, id_in_ready_o, handle_irq, enter_debug_mode } & _0204_;
assign _0539_ = { _1438_, _1368_ } & _0205_;
assign _0637_ = priv_mode_i & _0206_;
assign _0683_ = ctrl_fsm_cs & _0207_;
assign _1280_ = _0534_ == { _0201_[3], 3'h0 };
assign _1281_ = _0535_ == { _0202_[2], 1'h0, _0202_[0] };
assign _1282_ = _0536_ == _0203_;
assign _1283_ = _0538_ == { _0204_[3], 3'h0 };
assign _1284_ = _0539_ == { _0205_[1], 1'h0 };
assign _1285_ = _0637_ == _0206_;
assign _1286_ = _0683_ == { 1'h0, _0207_[2:1], 1'h0 };
assign _1287_ = _0683_ == { 3'h0, _0207_[0] };
assign _1288_ = _0683_ == { 1'h0, _0207_[2], 2'h0 };
assign _1289_ = _0683_ == { 1'h0, _0207_[2:0] };
assign _1290_ = _0683_ == { _0207_[3], 3'h0 };
assign _1291_ = _0683_ == { 2'h0, _0207_[1:0] };
assign _1292_ = _0683_ == { 2'h0, _0207_[1], 1'h0 };
assign _1293_ = _0683_ == { 1'h0, _0207_[2], 1'h0, _0207_[0] };
assign _1294_ = _0683_ == { _0207_[3], 2'h0, _0207_[0] };
assign _0431_ = _1280_ & _0194_;
assign _0433_ = _1281_ & _0195_;
assign _0435_ = _1282_ & _0196_;
assign _0439_ = _1283_ & _0197_;
assign _0441_ = _1284_ & _0198_;
assign _1341_ = _1285_ & _0199_;
assign _1443_ = _1287_ & _0200_;
assign _1437_ = _1288_ & _0200_;
assign _1434_ = _1289_ & _0200_;
assign _1379_ = _1286_ & _0200_;
assign _1328_ = _1290_ & _0200_;
assign _1439_ = _1291_ & _0200_;
assign _1339_ = _1292_ & _0200_;
assign controller_run_o_t0 = _1293_ & _0200_;
assign _1432_ = _1294_ & _0200_;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME debug_mode_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) debug_mode_o <= 1'h0;
else if (_0442_) debug_mode_o <= debug_mode_d;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME ctrl_fsm_cs */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) ctrl_fsm_cs <= 4'h0;
else if (_0444_) ctrl_fsm_cs <= ctrl_fsm_ns;
/* src = "generated/sv2v_out.v:12413.4-12421.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_intg_irq_int.mem_resp_intg_err_addr_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_intg_irq_int.mem_resp_intg_err_addr_q  <= 32'd0;
else if (_0446_) \g_intg_irq_int.mem_resp_intg_err_addr_q  <= lsu_addr_last_i;
assign _0638_ = _1371_ & _1372_;
assign _0641_ = stall_t0 & _1357_;
assign _0644_ = _1346_ & _1358_;
assign _0647_ = irq_nm_t0 & _1359_;
assign _0650_ = ebreak_into_debug_t0 & _1360_;
assign _0513_ = ebrk_insn_prio_t0 & ebreak_into_debug;
assign _0653_ = enter_debug_mode_prio_q_t0 & _1361_;
assign _0639_ = _1373_ & _1370_;
assign _0642_ = special_req_t0 & _1356_;
assign _0645_ = id_wb_pending_t0 & _1345_;
assign _0648_ = nmi_mode_o_t0 & irq_nm;
assign _0651_ = debug_mode_o_t0 & ebreak_into_debug;
assign _0514_ = ebreak_into_debug_t0 & ebrk_insn_prio;
assign _0654_ = _0185_ & enter_debug_mode_prio_q;
assign _0640_ = _1371_ & _1373_;
assign _0643_ = stall_t0 & special_req_t0;
assign _0646_ = _1346_ & id_wb_pending_t0;
assign _0649_ = irq_nm_t0 & nmi_mode_o_t0;
assign _0652_ = ebreak_into_debug_t0 & debug_mode_o_t0;
assign _0655_ = enter_debug_mode_prio_q_t0 & _0185_;
assign _1079_ = _0638_ | _0639_;
assign _1080_ = _0641_ | _0642_;
assign _1081_ = _0644_ | _0645_;
assign _1082_ = _0647_ | _0648_;
assign _1083_ = _0650_ | _0651_;
assign _1084_ = _0653_ | _0654_;
assign _0111_ = _1079_ | _0640_;
assign _1346_ = _1080_ | _0643_;
assign _1348_ = _1081_ | _0646_;
assign _1350_ = _1082_ | _0649_;
assign _0036_ = _1083_ | _0652_;
assign _1354_ = _1084_ | _0655_;
assign _0208_ = | { _1379_, debug_mode_entering_o_t0 };
assign _0209_ = | { _1328_, _1306_[0], _1443_, _1432_ };
assign _0210_ = | { _1328_, _1434_, _1432_ };
assign _0211_ = | { _1339_, _1439_, _1379_ };
assign _0212_ = | { _1328_, _1434_, _1443_, _1432_, _1437_, _1379_, controller_run_o_t0 };
assign _0213_ = | { _1339_, _1328_, _1432_, _1439_ };
assign _0214_ = | { _1328_, _1432_ };
assign _0215_ = | { _0969_, _1437_, controller_run_o_t0 };
assign _0216_ = | irqs_i_t0[14:0];
assign _0217_ = ~ { debug_mode_entering_o_t0, _1379_ };
assign _0218_ = ~ { _1306_[0], _1443_, _1328_, _1432_ };
assign _0219_ = ~ { _1328_, _1434_, _1432_ };
assign _0220_ = ~ { _1339_, _1439_, _1379_ };
assign _0221_ = ~ { _1443_, _1328_, _1437_, controller_run_o_t0, _1434_, _1432_, _1379_ };
assign _0222_ = ~ { _1339_, _1328_, _1439_, _1432_ };
assign _0223_ = ~ { _1328_, _1432_ };
assign _0224_ = ~ { _0969_, _1437_, controller_run_o_t0 };
assign _0225_ = ~ irqs_i_t0[14:0];
assign _0207_ = ~ ctrl_fsm_cs_t0;
assign _0537_ = { _0421_, _1401_ } & _0217_;
assign _0540_ = { _1444_, _1442_, _1440_, _1431_ } & _0218_;
assign _0541_ = { _1440_, _1433_, _1431_ } & _0219_;
assign _0542_ = { _1441_, _1438_, _1401_ } & _0220_;
assign _0543_ = { _1442_, _1440_, _1436_, _1435_, _1433_, _1431_, _1401_ } & _0221_;
assign _0544_ = { _1441_, _1440_, _1438_, _1431_ } & _0222_;
assign _0545_ = { _1440_, _1431_ } & _0223_;
assign _0561_ = { _0968_, _1436_, _1435_ } & _0224_;
assign _0684_ = irqs_i[14:0] & _0225_;
assign _0226_ = ! _0537_;
assign _0227_ = ! _0540_;
assign _0228_ = ! _0541_;
assign _0229_ = ! _0542_;
assign _0230_ = ! _0543_;
assign _0231_ = ! _0544_;
assign _0232_ = ! _0545_;
assign _0233_ = ! _0561_;
assign _0234_ = ! _0637_;
assign _0235_ = ! _0684_;
assign _0236_ = ! _0683_;
assign _0437_ = _0226_ & _0208_;
assign _0449_ = _0227_ & _0209_;
assign _0451_ = _0228_ & _0210_;
assign _0453_ = _0229_ & _0211_;
assign instr_req_o_t0 = _0230_ & _0212_;
assign _0456_ = _0231_ & _0213_;
assign debug_mode_entering_o_t0 = _0232_ & _0214_;
assign _0423_ = _0233_ & _0215_;
assign _1343_ = _0234_ & _0199_;
assign _1381_ = _0235_ & _0216_;
assign _1306_[0] = _0236_ & _0200_;
assign _0237_ = ~ irq_nm;
assign _0238_ = ~ _1362_;
assign _0239_ = ~ _1364_;
assign _0240_ = ~ _1366_;
assign _0241_ = ~ branch_set_i;
assign _0243_ = ~ stall;
assign _0244_ = ~ exc_req_q;
assign _0245_ = ~ _1374_;
assign _0246_ = ~ irq_pending_i;
assign _0247_ = ~ debug_req_i;
assign _0248_ = ~ debug_mode_o;
assign _0249_ = ~ debug_single_step_i;
assign _0250_ = ~ jump_set_i;
assign _0252_ = ~ id_wb_pending;
assign _0254_ = ~ load_err_q;
assign _0656_ = irq_nm_t0 & _0246_;
assign _0659_ = _1363_ & _0247_;
assign _0662_ = _1365_ & _0248_;
assign _0665_ = _1367_ & _0249_;
assign _0668_ = branch_set_i_t0 & _0250_;
assign _0671_ = enter_debug_mode_t0 & _0251_;
assign _0674_ = stall_t0 & _0252_;
assign _0677_ = exc_req_q_t0 & _0253_;
assign _0680_ = _1375_ & _0254_;
assign _0657_ = irq_pending_i_t0 & _0237_;
assign _0660_ = debug_req_i_t0 & _0238_;
assign _0663_ = debug_mode_o_t0 & _0239_;
assign _0666_ = debug_single_step_i_t0 & _0240_;
assign _0669_ = jump_set_i_t0 & _0241_;
assign _0672_ = handle_irq_t0 & _0242_;
assign _0675_ = id_wb_pending_t0 & _0243_;
assign _0678_ = store_err_q_t0 & _0244_;
assign _0681_ = load_err_q_t0 & _0245_;
assign _0658_ = irq_nm_t0 & irq_pending_i_t0;
assign _0661_ = _1363_ & debug_req_i_t0;
assign _0664_ = _1365_ & debug_mode_o_t0;
assign _0667_ = _1367_ & debug_single_step_i_t0;
assign _0670_ = branch_set_i_t0 & jump_set_i_t0;
assign _0673_ = enter_debug_mode_t0 & handle_irq_t0;
assign _0676_ = stall_t0 & id_wb_pending_t0;
assign _0679_ = exc_req_q_t0 & store_err_q_t0;
assign _0682_ = _1375_ & load_err_q_t0;
assign _1085_ = _0656_ | _0657_;
assign _1086_ = _0659_ | _0660_;
assign _1087_ = _0662_ | _0663_;
assign _1088_ = _0665_ | _0666_;
assign _1089_ = _0668_ | _0669_;
assign _1090_ = _0671_ | _0672_;
assign _1091_ = _0674_ | _0675_;
assign _1092_ = _0677_ | _0678_;
assign _1093_ = _0680_ | _0681_;
assign _1363_ = _1085_ | _0658_;
assign _1365_ = _1086_ | _0661_;
assign _1367_ = _1087_ | _0664_;
assign _0038_ = _1088_ | _0667_;
assign _0064_ = _1089_ | _0670_;
assign _1371_ = _1090_ | _0673_;
assign _1373_ = _1091_ | _0676_;
assign _1375_ = _1092_ | _0679_;
assign _1377_ = _1093_ | _0682_;
assign _0255_ = ~ { _1435_, _1435_, _1435_, _1435_ };
assign _0256_ = ~ { _0968_, _0968_, _0968_, _0968_ };
assign _0257_ = ~ { _1442_, _1442_, _1442_, _1442_ };
assign _0258_ = ~ { _0970_, _0970_, _0970_, _0970_ };
assign _0259_ = ~ { _0422_, _0422_, _0422_, _0422_ };
assign _0263_ = ~ _0972_;
assign _0264_ = ~ { _0968_, _0968_, _0968_ };
assign _0265_ = ~ _0452_;
assign _0266_ = ~ _0974_;
assign _0269_ = ~ { _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_ };
assign _0267_ = ~ _1440_;
assign _0270_ = ~ _0976_;
assign _0262_ = ~ _1433_;
assign _0271_ = ~ { _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_ };
assign _0272_ = ~ { _1401_, _1401_ };
assign _0273_ = ~ _1441_;
assign _0274_ = ~ _1438_;
assign _0275_ = ~ \g_intg_irq_int.mem_resp_intg_err_irq_pending_q ;
assign _0253_ = ~ store_err_q;
assign _0276_ = ~ ebrk_insn;
assign _0277_ = ~ ecall_insn;
assign _0278_ = ~ illegal_insn_q;
assign _0279_ = ~ instr_fetch_err;
assign _0280_ = ~ { _1353_, _1353_, _1353_, _1353_ };
assign _0281_ = ~ dret_insn;
assign _0282_ = ~ { dret_insn, dret_insn, dret_insn, dret_insn };
assign _0283_ = ~ mret_insn;
assign _0284_ = ~ { mret_insn, mret_insn, mret_insn };
assign _0285_ = ~ { mret_insn, mret_insn, mret_insn, mret_insn };
assign _0286_ = ~ { store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio };
assign _0287_ = ~ { ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio };
assign _0288_ = ~ { ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio };
assign _0289_ = ~ { illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio };
assign _0290_ = ~ { instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio };
assign _0291_ = ~ { store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio };
assign _0292_ = ~ { ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio };
assign _0293_ = ~ { ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio };
assign _0294_ = ~ { illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio };
assign _0295_ = ~ { instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio };
assign _0296_ = ~ { ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio };
assign _0297_ = ~ { illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio };
assign _0298_ = ~ { instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio };
assign _0299_ = ~ ecall_insn_prio;
assign _0300_ = ~ illegal_insn_prio;
assign _0301_ = ~ instr_fetch_err_prio;
assign _0302_ = ~ { _1376_, _1376_, _1376_, _1376_ };
assign _0303_ = ~ _1376_;
assign _0304_ = ~ { _1376_, _1376_, _1376_ };
assign _0305_ = ~ { irqs_i[15], irqs_i[15], irqs_i[15], irqs_i[15], irqs_i[15], irqs_i[15], irqs_i[15] };
assign _0306_ = ~ { _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_ };
assign _0307_ = ~ _1349_;
assign _0308_ = ~ { _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_ };
assign _0251_ = ~ handle_irq;
assign _0309_ = ~ { handle_irq, handle_irq, handle_irq, handle_irq };
assign _0242_ = ~ enter_debug_mode;
assign _0310_ = ~ { enter_debug_mode, enter_debug_mode, enter_debug_mode, enter_debug_mode };
assign _0311_ = ~ _1347_;
assign _0312_ = ~ { _1347_, _1347_, _1347_, _1347_ };
assign _0313_ = ~ { ready_wb_i, ready_wb_i, ready_wb_i, ready_wb_i };
assign _0314_ = ~ { special_req, special_req, special_req, special_req };
assign _0261_ = ~ _1435_;
assign _0260_ = ~ _1401_;
assign _0268_ = ~ _1431_;
assign _0315_ = ~ { irqs_i[0], irqs_i[0], irqs_i[0], irqs_i[0] };
assign _0316_ = ~ { irqs_i[1], irqs_i[1], irqs_i[1], irqs_i[1] };
assign _0317_ = ~ { irqs_i[2], irqs_i[2], irqs_i[2], irqs_i[2] };
assign _0318_ = ~ { irqs_i[3], irqs_i[3], irqs_i[3], irqs_i[3] };
assign _0319_ = ~ { irqs_i[4], irqs_i[4], irqs_i[4], irqs_i[4] };
assign _0320_ = ~ { irqs_i[5], irqs_i[5], irqs_i[5], irqs_i[5] };
assign _0321_ = ~ { irqs_i[6], irqs_i[6], irqs_i[6], irqs_i[6] };
assign _0322_ = ~ { irqs_i[7], irqs_i[7], irqs_i[7], irqs_i[7] };
assign _0323_ = ~ { irqs_i[8], irqs_i[8], irqs_i[8], irqs_i[8] };
assign _0324_ = ~ { irqs_i[9], irqs_i[9], irqs_i[9], irqs_i[9] };
assign _0325_ = ~ { irqs_i[10], irqs_i[10], irqs_i[10], irqs_i[10] };
assign _0326_ = ~ { irqs_i[11], irqs_i[11], irqs_i[11], irqs_i[11] };
assign _0327_ = ~ { irqs_i[12], irqs_i[12], irqs_i[12], irqs_i[12] };
assign _0328_ = ~ { irqs_i[13], irqs_i[13], irqs_i[13], irqs_i[13] };
assign _0329_ = ~ instr_valid_i;
assign _0330_ = ~ _1342_;
assign _0331_ = ~ _1340_;
assign _0332_ = ~ { debug_req_i, debug_req_i, debug_req_i };
assign _0333_ = ~ { _0184_, _0184_, _0184_ };
assign _0334_ = ~ { trigger_match_i, trigger_match_i, trigger_match_i };
assign _0335_ = ~ { instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i };
assign _0336_ = ~ { instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i };
assign _1023_ = { controller_run_o_t0, controller_run_o_t0, controller_run_o_t0, controller_run_o_t0 } | _0255_;
assign _1026_ = { _0969_, _0969_, _0969_, _0969_ } | _0256_;
assign _1029_ = { _1443_, _1443_, _1443_, _1443_ } | _0257_;
assign _1030_ = { _0971_, _0971_, _0971_, _0971_ } | _0258_;
assign _1033_ = { _0423_, _0423_, _0423_, _0423_ } | _0259_;
assign _1039_ = _1434_ | _0262_;
assign _1042_ = _0973_ | _0263_;
assign _1046_ = { _0969_, _0969_, _0969_ } | _0264_;
assign _1049_ = _0453_ | _0265_;
assign _1051_ = _0975_ | _0266_;
assign _1057_ = _1328_ | _0267_;
assign _1062_ = { _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_ } | _0269_;
assign _1066_ = _0977_ | _0270_;
assign _1070_ = { _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_ } | _0271_;
assign _1073_ = { _1379_, _1379_ } | _0272_;
assign _1076_ = _1439_ | _0274_;
assign _1115_ = \g_intg_irq_int.mem_resp_intg_err_irq_pending_q_t0  | _0275_;
assign _1117_ = store_err_q_t0 | _0253_;
assign _1118_ = ebrk_insn_t0 | _0276_;
assign _1119_ = ecall_insn_t0 | _0277_;
assign _1120_ = illegal_insn_q_t0 | _0278_;
assign _1121_ = instr_fetch_err_prio_t0 | _0279_;
assign _1123_ = { _1354_, _1354_, _1354_, _1354_ } | _0280_;
assign _1124_ = { dret_insn_t0, dret_insn_t0, dret_insn_t0, dret_insn_t0 } | _0282_;
assign _1125_ = mret_insn_t0 | _0283_;
assign _1126_ = { mret_insn_t0, mret_insn_t0, mret_insn_t0 } | _0284_;
assign _1127_ = { mret_insn_t0, mret_insn_t0, mret_insn_t0, mret_insn_t0 } | _0285_;
assign _1129_ = { store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0 } | _0286_;
assign _1132_ = { ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0 } | _0287_;
assign _1133_ = { ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0 } | _0288_;
assign _1134_ = { illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0 } | _0289_;
assign _1137_ = { instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0 } | _0290_;
assign _1140_ = { store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0 } | _0291_;
assign _1141_ = { ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0 } | _0292_;
assign _1144_ = { ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0 } | _0293_;
assign _1147_ = { illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0 } | _0294_;
assign _1148_ = { instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0 } | _0295_;
assign _1150_ = { ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0 } | _0296_;
assign _1151_ = { illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0 } | _0297_;
assign _1152_ = { instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0 } | _0298_;
assign _1153_ = ecall_insn_prio_t0 | _0299_;
assign _1154_ = illegal_insn_prio_t0 | _0300_;
assign _1155_ = instr_fetch_err_prio_t0 | _0301_;
assign _1157_ = { _1377_, _1377_, _1377_, _1377_ } | _0302_;
assign _1160_ = _1377_ | _0303_;
assign _1166_ = { _1377_, _1377_, _1377_ } | _0304_;
assign _1168_ = { irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15] } | _0305_;
assign _1169_ = { _1381_, _1381_, _1381_, _1381_, _1381_, _1381_, _1381_ } | _0306_;
assign _1173_ = _1350_ | _0307_;
assign _1175_ = { _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_ } | _0308_;
assign _1178_ = handle_irq_t0 | _0251_;
assign _1183_ = { handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0 } | _0309_;
assign _1184_ = enter_debug_mode_t0 | _0242_;
assign _1185_ = { enter_debug_mode_t0, enter_debug_mode_t0, enter_debug_mode_t0, enter_debug_mode_t0 } | _0310_;
assign _1186_ = _1348_ | _0311_;
assign _1189_ = { _1348_, _1348_, _1348_, _1348_ } | _0312_;
assign _1193_ = { ready_wb_i_t0, ready_wb_i_t0, ready_wb_i_t0, ready_wb_i_t0 } | _0313_;
assign _1194_ = { special_req_t0, special_req_t0, special_req_t0, special_req_t0 } | _0314_;
assign _1036_ = _1379_ | _0260_;
assign _1058_ = _1432_ | _0268_;
assign _1197_ = { irqs_i_t0[0], irqs_i_t0[0], irqs_i_t0[0], irqs_i_t0[0] } | _0315_;
assign _1198_ = { irqs_i_t0[1], irqs_i_t0[1], irqs_i_t0[1], irqs_i_t0[1] } | _0316_;
assign _1199_ = { irqs_i_t0[2], irqs_i_t0[2], irqs_i_t0[2], irqs_i_t0[2] } | _0317_;
assign _1200_ = { irqs_i_t0[3], irqs_i_t0[3], irqs_i_t0[3], irqs_i_t0[3] } | _0318_;
assign _1201_ = { irqs_i_t0[4], irqs_i_t0[4], irqs_i_t0[4], irqs_i_t0[4] } | _0319_;
assign _1202_ = { irqs_i_t0[5], irqs_i_t0[5], irqs_i_t0[5], irqs_i_t0[5] } | _0320_;
assign _1203_ = { irqs_i_t0[6], irqs_i_t0[6], irqs_i_t0[6], irqs_i_t0[6] } | _0321_;
assign _1204_ = { irqs_i_t0[7], irqs_i_t0[7], irqs_i_t0[7], irqs_i_t0[7] } | _0322_;
assign _1205_ = { irqs_i_t0[8], irqs_i_t0[8], irqs_i_t0[8], irqs_i_t0[8] } | _0323_;
assign _1206_ = { irqs_i_t0[9], irqs_i_t0[9], irqs_i_t0[9], irqs_i_t0[9] } | _0324_;
assign _1207_ = { irqs_i_t0[10], irqs_i_t0[10], irqs_i_t0[10], irqs_i_t0[10] } | _0325_;
assign _1208_ = { irqs_i_t0[11], irqs_i_t0[11], irqs_i_t0[11], irqs_i_t0[11] } | _0326_;
assign _1209_ = { irqs_i_t0[12], irqs_i_t0[12], irqs_i_t0[12], irqs_i_t0[12] } | _0327_;
assign _1210_ = { irqs_i_t0[13], irqs_i_t0[13], irqs_i_t0[13], irqs_i_t0[13] } | _0328_;
assign _1211_ = instr_valid_i_t0 | _0329_;
assign _1215_ = _1341_ | _0331_;
assign _1218_ = { debug_req_i_t0, debug_req_i_t0, debug_req_i_t0 } | _0332_;
assign _1219_ = { _0185_, _0185_, _0185_ } | _0333_;
assign _1220_ = { trigger_match_i_t0, trigger_match_i_t0, trigger_match_i_t0 } | _0334_;
assign _1221_ = { instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0 } | _0335_;
assign _1224_ = { instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0 } | _0336_;
assign _1022_ = { _1379_, _1379_, _1379_, _1379_ } | { _1401_, _1401_, _1401_, _1401_ };
assign _1024_ = { controller_run_o_t0, controller_run_o_t0, controller_run_o_t0, controller_run_o_t0 } | { _1435_, _1435_, _1435_, _1435_ };
assign _1027_ = { _0969_, _0969_, _0969_, _0969_ } | { _0968_, _0968_, _0968_, _0968_ };
assign _1031_ = { _0971_, _0971_, _0971_, _0971_ } | { _0970_, _0970_, _0970_, _0970_ };
assign _1034_ = { _0423_, _0423_, _0423_, _0423_ } | { _0422_, _0422_, _0422_, _0422_ };
assign _1037_ = _1379_ | _1401_;
assign _1038_ = controller_run_o_t0 | _1435_;
assign _1040_ = _1434_ | _1433_;
assign _1043_ = _0973_ | _0972_;
assign _1045_ = { _1379_, _1379_, _1379_ } | { _1401_, _1401_, _1401_ };
assign _1047_ = { _0969_, _0969_, _0969_ } | { _0968_, _0968_, _0968_ };
assign _1050_ = _1437_ | _1436_;
assign _1052_ = _0975_ | _0974_;
assign _1059_ = _1432_ | _1431_;
assign _1061_ = { _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_ } | { _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_ };
assign _1063_ = { _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_ } | { _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_ };
assign _1067_ = _0977_ | _0976_;
assign _1069_ = { _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_ } | { _1433_, _1433_, _1433_, _1433_, _1433_, _1433_, _1433_ };
assign _1071_ = { _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_ } | { _1401_, _1401_, _1401_, _1401_, _1401_, _1401_, _1401_ };
assign _1074_ = { _1379_, _1379_ } | { _1401_, _1401_ };
assign _1077_ = _1439_ | _1438_;
assign _1116_ = \g_intg_irq_int.mem_resp_intg_err_irq_pending_q_t0  | \g_intg_irq_int.mem_resp_intg_err_irq_pending_q ;
assign _1122_ = instr_exec_i_t0 | instr_exec_i;
assign _1128_ = { load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0 } | { load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio, load_err_prio };
assign _1130_ = { store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0 } | { store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio, store_err_prio };
assign _1135_ = { illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0 } | { illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio, illegal_insn_prio };
assign _1138_ = { instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0 } | { instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio, instr_fetch_err_prio };
assign _1142_ = { ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0 } | { ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio };
assign _1145_ = { ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0 } | { ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio, ecall_insn_prio };
assign _1149_ = { ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0 } | { ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio, ebrk_insn_prio };
assign _1156_ = ebrk_insn_prio_t0 | ebrk_insn_prio;
assign _1158_ = { _1377_, _1377_, _1377_, _1377_ } | { _1376_, _1376_, _1376_, _1376_ };
assign _1161_ = _1377_ | _1376_;
assign _1162_ = { _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_ } | { _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_ };
assign _1163_ = { _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_ } | { _1376_, _1376_, _1376_, _1376_, _1376_, _1376_, _1376_ };
assign _1165_ = { _1377_, _1377_ } | { _1376_, _1376_ };
assign _1170_ = { _1381_, _1381_, _1381_, _1381_, _1381_, _1381_, _1381_ } | { _1380_, _1380_, _1380_, _1380_, _1380_, _1380_, _1380_ };
assign _1172_ = { _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_ } | { _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_, _0186_ };
assign _1174_ = { _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_ } | { _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_ };
assign _1176_ = { _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_ } | { _1349_, _1349_, _1349_, _1349_, _1349_, _1349_, _1349_ };
assign _1179_ = handle_irq_t0 | handle_irq;
assign _1181_ = { handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0 } | { handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq };
assign _1182_ = { handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0 } | { handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq, handle_irq };
assign _1187_ = _1348_ | _1347_;
assign _1190_ = { _1348_, _1348_, _1348_, _1348_ } | { _1347_, _1347_, _1347_, _1347_ };
assign _1192_ = _0064_ | _1369_;
assign _1195_ = { special_req_t0, special_req_t0, special_req_t0, special_req_t0 } | { special_req, special_req, special_req, special_req };
assign _1212_ = instr_valid_i_t0 | instr_valid_i;
assign _1214_ = _1343_ | _1342_;
assign _1216_ = _1341_ | _1340_;
assign _1222_ = { instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0 } | { instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i, instr_fetch_err_plus2_i };
assign _1225_ = { instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0 } | { instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i, instr_is_compressed_i };
assign _0564_ = _0126_ & _1023_;
assign _0567_ = _1300_ & _1026_;
assign _0570_ = { 3'h0, _1306_[0] } & _1029_;
assign _0572_ = _1308_ & _1030_;
assign _0575_ = _1310_ & _1033_;
assign _0582_ = _1314_ & _1039_;
assign _0585_ = _1316_ & _1042_;
assign _0590_ = { 2'h0, controller_run_o_t0 } & _1046_;
assign _0593_ = _0130_ & _1049_;
assign _0597_ = _1323_ & _1051_;
assign _0600_ = nmi_mode_o_t0 & _1039_;
assign _0603_ = _1325_ & _1036_;
assign _0606_ = _0456_ & _1036_;
assign _0609_ = _1328_ & _1058_;
assign _0614_ = _1330_ & _1062_;
assign _0617_ = _0036_ & _1036_;
assign _0620_ = _1334_ & _1057_;
assign _0622_ = csr_save_if_o_t0 & _1066_;
assign _0628_ = _1336_ & _1070_;
assign _0631_ = { debug_mode_entering_o_t0, debug_mode_entering_o_t0 } & _1073_;
assign _0634_ = _1339_ & _1076_;
assign _0748_ = mem_resp_intg_err_i_t0 & _1115_;
assign _0750_ = load_err_q_t0 & _1117_;
assign _0752_ = _0132_ & _1118_;
assign _0754_ = store_err_q_t0 & _1118_;
assign _0756_ = _0113_ & _1119_;
assign _0758_ = _0122_ & _1119_;
assign _0760_ = ebrk_insn_t0 & _1119_;
assign _0762_ = _0089_ & _1120_;
assign _0764_ = _0097_ & _1120_;
assign _0766_ = _0080_ & _1120_;
assign _0768_ = ecall_insn_t0 & _1120_;
assign _0770_ = _0056_ & _1121_;
assign _0772_ = _0071_ & _1121_;
assign _0774_ = _0042_ & _1121_;
assign _0776_ = _0044_ & _1121_;
assign _0778_ = illegal_insn_q_t0 & _1121_;
assign _0782_ = _0005_ & _1123_;
assign _0784_ = { 1'h0, wfi_insn_t0, wfi_insn_t0, wfi_insn_t0 } & _1124_;
assign _0786_ = nmi_mode_o_t0 & _1125_;
assign _0788_ = dret_insn_t0 & _1125_;
assign _0790_ = { dret_insn_t0, 2'h0 } & _1126_;
assign _0792_ = _0021_ & _1127_;
assign _0797_ = _1403_ & _1129_;
assign _0800_ = _1404_ & _1132_;
assign _0802_ = _1405_ & _1133_;
assign _0804_ = _1407_ & _1134_;
assign _0807_ = _1409_ & _1137_;
assign _0810_ = { 4'h0, load_err_prio_t0, 1'h0, load_err_prio_t0 } & _1140_;
assign _0812_ = _1412_ & _1141_;
assign _0815_ = _1414_ & _1144_;
assign _0818_ = _1416_ & _1147_;
assign _0820_ = _1418_ & _1148_;
assign _0824_ = _1420_ & _1150_;
assign _0826_ = _1422_ & _1151_;
assign _0828_ = _1424_ & _1152_;
assign _0830_ = _1426_ & _1153_;
assign _0832_ = _1428_ & _1154_;
assign _0834_ = _1430_ & _1155_;
assign _0838_ = _0017_ & _1157_;
assign _0848_ = _0157_ & _1160_;
assign _0852_ = _0095_ & _1166_;
assign _0854_ = _0136_ & _1160_;
assign _0857_ = _0075_ & _1160_;
assign _0859_ = mret_insn_t0 & _1160_;
assign _0861_ = { 4'h0, irqs_i_t0[17], 2'h0 } & _1168_;
assign _0863_ = _0128_ & _1169_;
assign _0868_ = nmi_mode_o_t0 & _1173_;
assign _0872_ = _0108_ & _1175_;
assign _0875_ = nmi_mode_o_t0 & _1178_;
assign _0882_ = _0111_ & _1178_;
assign _0884_ = _0141_ & _1183_;
assign _0886_ = _0153_ & _1184_;
assign _0888_ = _0001_ & _1185_;
assign _0890_ = _0111_ & _1186_;
assign _0893_ = _0141_ & _1189_;
assign _0900_ = ctrl_fsm_cs_t0 & _1193_;
assign _0902_ = ctrl_fsm_cs_t0 & _1194_;
assign _0905_ = handle_irq_t0 & _1184_;
assign _0907_ = _0104_ & _1185_;
assign _0920_ = _0019_ & _1197_;
assign _0922_ = _0015_ & _1198_;
assign _0924_ = _0011_ & _1199_;
assign _0926_ = _0007_ & _1200_;
assign _0928_ = _0003_ & _1201_;
assign _0930_ = _0168_ & _1202_;
assign _0932_ = _0163_ & _1203_;
assign _0934_ = _0155_ & _1204_;
assign _0936_ = _0147_ & _1205_;
assign _0938_ = _0134_ & _1206_;
assign _0940_ = _0115_ & _1207_;
assign _0942_ = _0091_ & _1208_;
assign _0944_ = _0058_ & _1209_;
assign _0946_ = { irqs_i_t0[14], irqs_i_t0[14], irqs_i_t0[14], 1'h0 } & _1210_;
assign _0948_ = do_single_step_q_t0 & _1211_;
assign _0953_ = _1446_ & _1215_;
assign _0956_ = { do_single_step_d_t0, 2'h0 } & _1218_;
assign _0958_ = _1449_ & _1219_;
assign _0960_ = _1451_ & _1220_;
assign _0962_ = pc_id_i_t0 & _1221_;
assign _0965_ = instr_i_t0 & _1224_;
assign _0562_ = _0024_ & _1022_;
assign _0565_ = _0159_ & _1024_;
assign _0568_ = _1298_ & _1027_;
assign _0573_ = _1304_ & _1031_;
assign _0576_ = _1302_ & _1034_;
assign _0578_ = _0120_ & _1037_;
assign _0580_ = _0064_ & _1038_;
assign _0583_ = handle_irq_t0 & _1040_;
assign _0586_ = _1312_ & _1043_;
assign _0588_ = _0062_ & _1045_;
assign _0591_ = _1318_ & _1047_;
assign _0595_ = _0087_ & _1050_;
assign _0598_ = _1321_ & _1052_;
assign _0601_ = _0060_ & _1040_;
assign _0604_ = _0117_ & _1037_;
assign _0607_ = _0050_ & _1037_;
assign _0610_ = _0036_ & _1059_;
assign _0612_ = _0029_ & _1061_;
assign _0615_ = _0124_ & _1063_;
assign _0618_ = _0102_ & _1037_;
assign _0623_ = _1332_ & _1067_;
assign _0626_ = _0046_ & _1069_;
assign _0629_ = _0151_ & _1071_;
assign _0632_ = _0048_ & _1074_;
assign _0635_ = _0038_ & _1077_;
assign _0746_ = _0052_ & _1116_;
assign _0780_ = _0026_ & _1122_;
assign _0795_ = lsu_addr_last_i_t0 & _1128_;
assign _0798_ = lsu_addr_last_i_t0 & _1130_;
assign _0805_ = _1457_ & _1135_;
assign _0808_ = _1455_ & _1138_;
assign _0813_ = { 5'h00, _0013_[3], _0013_[3] } & _1142_;
assign _0816_ = { 5'h00, _1341_, _1341_ } & _1145_;
assign _0822_ = { _0013_[3], _0013_[3], 2'h0 } & _1149_;
assign _0836_ = _0013_[3] & _1156_;
assign _0839_ = _0009_ & _1158_;
assign _0841_ = _0085_ & _1161_;
assign _0843_ = _0139_ & _1162_;
assign _0846_ = _0161_ & _1163_;
assign _0850_ = { debug_mode_o_t0, debug_mode_o_t0 } & _1165_;
assign _0855_ = nmi_mode_o_t0 & _1161_;
assign _0864_ = { 3'h0, mfip_id_t0 } & _1170_;
assign _0866_ = \g_intg_irq_int.mem_resp_intg_err_addr_q_t0  & _1172_;
assign _0870_ = _0099_ & _1174_;
assign _0873_ = { irq_nm_ext_i_t0, irq_nm_ext_i_t0, irq_nm_ext_i_t0, irq_nm_ext_i_t0, irq_nm_ext_i_t0, irq_nm_ext_i_t0, irq_nm_ext_i_t0 } & _1176_;
assign _0876_ = _0093_ & _1179_;
assign _0878_ = _0073_ & _1181_;
assign _0880_ = _0083_ & _1182_;
assign _0891_ = _0144_ & _1187_;
assign _0894_ = _0165_ & _1190_;
assign _0896_ = jump_set_i_t0 & _1192_;
assign _0898_ = branch_set_i_t0 & _1192_;
assign _0903_ = _0149_ & _1195_;
assign _0909_ = special_req_t0 & _1038_;
assign _0911_ = _0068_ & _1038_;
assign _0913_ = _0066_ & _1038_;
assign _0915_ = _0031_ & _1037_;
assign _0917_ = _0033_ & _1037_;
assign _0949_ = _0175_ & _1212_;
assign _0951_ = debug_ebreaku_i_t0 & _1214_;
assign _0954_ = debug_ebreakm_i_t0 & _1216_;
assign _0963_ = _0170_ & _1222_;
assign _0966_ = { 16'h0000, instr_compressed_i_t0 } & _1225_;
assign _1025_ = _0564_ | _0565_;
assign _1028_ = _0567_ | _0568_;
assign _1032_ = _0572_ | _0573_;
assign _1035_ = _0575_ | _0576_;
assign _1041_ = _0582_ | _0583_;
assign _1044_ = _0585_ | _0586_;
assign _1048_ = _0590_ | _0591_;
assign _1053_ = _0597_ | _0598_;
assign _1054_ = _0600_ | _0601_;
assign _1055_ = _0603_ | _0604_;
assign _1056_ = _0606_ | _0607_;
assign _1060_ = _0609_ | _0610_;
assign _1064_ = _0614_ | _0615_;
assign _1065_ = _0617_ | _0618_;
assign _1068_ = _0622_ | _0623_;
assign _1072_ = _0628_ | _0629_;
assign _1075_ = _0631_ | _0632_;
assign _1078_ = _0634_ | _0635_;
assign _1131_ = _0797_ | _0798_;
assign _1136_ = _0804_ | _0805_;
assign _1139_ = _0807_ | _0808_;
assign _1143_ = _0812_ | _0813_;
assign _1146_ = _0815_ | _0816_;
assign _1159_ = _0838_ | _0839_;
assign _1164_ = _0848_ | _0841_;
assign _1167_ = _0854_ | _0855_;
assign _1171_ = _0863_ | _0864_;
assign _1177_ = _0872_ | _0873_;
assign _1180_ = _0875_ | _0876_;
assign _1188_ = _0890_ | _0891_;
assign _1191_ = _0893_ | _0894_;
assign _1196_ = _0902_ | _0903_;
assign _1213_ = _0948_ | _0949_;
assign _1217_ = _0953_ | _0954_;
assign _1223_ = _0962_ | _0963_;
assign _1226_ = _0965_ | _0966_;
assign _1231_ = _0125_ ^ _0158_;
assign _1232_ = _1299_ ^ _1297_;
assign _1234_ = _1307_ ^ _1303_;
assign _1235_ = _1309_ ^ _1301_;
assign _1236_ = _1313_ ^ _0034_;
assign _1237_ = _1315_ ^ _1311_;
assign _1238_ = _1319_ ^ _1317_;
assign _1239_ = _1322_ ^ _1320_;
assign _1240_ = nmi_mode_o ^ _0059_;
assign _1241_ = _1324_ ^ _0116_;
assign _1242_ = _1326_ ^ _0049_;
assign _1243_ = _1327_ ^ _0035_;
assign _1244_ = _1329_ ^ _0123_;
assign _1245_ = _0035_ ^ _0101_;
assign _1246_ = csr_save_if_o ^ _1331_;
assign _1247_ = _1335_ ^ _0150_;
assign _1248_ = _1337_ ^ _0047_;
assign _1249_ = _1338_ ^ _0037_;
assign _1250_ = _1402_ ^ lsu_addr_last_i;
assign _1253_ = _1406_ ^ _1456_;
assign _1254_ = _1408_ ^ _1454_;
assign _1256_ = _1411_ ^ _0166_;
assign _1257_ = _1413_ ^ _1458_;
assign _1263_ = _0016_ ^ _0008_;
assign _1264_ = _0156_ ^ _0084_;
assign _1266_ = _0135_ ^ nmi_mode_o;
assign _1267_ = _0127_ ^ { 3'h3, mfip_id };
assign _1268_ = _0107_ ^ _1452_;
assign _1269_ = nmi_mode_o ^ _0092_;
assign _1270_ = _0110_ ^ _0143_;
assign _1271_ = _0140_ ^ _0164_;
assign _1272_ = ctrl_fsm_cs ^ _0148_;
assign _1273_ = do_single_step_q ^ _0174_;
assign _1274_ = _1445_ ^ debug_ebreakm_i;
assign _1278_ = pc_id_i ^ _0169_;
assign _1279_ = instr_i ^ { 16'h0000, instr_compressed_i };
assign _0563_ = { _1379_, _1379_, _1379_, _1379_ } & { _0023_[3], _0366_[1], _0023_[1], _0366_[0] };
assign _0566_ = { controller_run_o_t0, controller_run_o_t0, controller_run_o_t0, controller_run_o_t0 } & _1231_;
assign _0569_ = { _0969_, _0969_, _0969_, _0969_ } & _1232_;
assign _1304_ = { _1439_, _1439_, _1439_, _1439_ } & { _0039_[3:2], _0353_ };
assign _0571_ = { _1443_, _1443_, _1443_, _1443_ } & { _1233_[3], _0352_, _1233_[1:0] };
assign _0574_ = { _0971_, _0971_, _0971_, _0971_ } & _1234_;
assign _0577_ = { _0423_, _0423_, _0423_, _0423_ } & _1235_;
assign _0579_ = _1379_ & _0349_;
assign _0581_ = controller_run_o_t0 & _0063_;
assign _0584_ = _1434_ & _1236_;
assign _0587_ = _0973_ & _1237_;
assign _0589_ = { _1379_, _1379_, _1379_ } & { _0061_[2], _0369_, _0061_[0] };
assign _0592_ = { _0969_, _0969_, _0969_ } & _1238_;
assign _0594_ = _0453_ & _0341_;
assign _0596_ = _1437_ & _0086_;
assign _0599_ = _0975_ & _1239_;
assign debug_mode_d_t0 = _1379_ & _0343_;
assign _0602_ = _1434_ & _1240_;
assign _0605_ = _1379_ & _1241_;
assign _0608_ = _1379_ & _1242_;
assign _0611_ = _1432_ & _1243_;
assign _0613_ = { _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_ } & _0028_;
assign _0616_ = { _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_ } & _1244_;
assign _0619_ = _1379_ & _1245_;
assign _0621_ = _1328_ & _0351_;
assign _0624_ = _0977_ & _1246_;
assign _0625_ = _1434_ & _0034_;
assign _0627_ = { _1434_, _1434_, _1434_, _1434_, _1434_, _1434_, _1434_ } & _0045_;
assign _0630_ = { _1379_, _1379_, _1379_, _1379_, _1379_, _1379_, _1379_ } & _1247_;
assign _0633_ = { _1379_, _1379_ } & _1248_;
assign _0636_ = _1439_ & _1249_;
assign _0747_ = \g_intg_irq_int.mem_resp_intg_err_irq_pending_q_t0  & _0051_;
assign _0749_ = \g_intg_irq_int.mem_resp_intg_err_irq_pending_q_t0  & _0053_;
assign _0751_ = store_err_q_t0 & _0145_;
assign _0753_ = ebrk_insn_t0 & _0131_;
assign _0755_ = ebrk_insn_t0 & _0137_;
assign _0757_ = ecall_insn_t0 & _0112_;
assign _0759_ = ecall_insn_t0 & _0121_;
assign _0761_ = ecall_insn_t0 & _0106_;
assign _0763_ = illegal_insn_q_t0 & _0088_;
assign _0765_ = illegal_insn_q_t0 & _0096_;
assign _0767_ = illegal_insn_q_t0 & _0079_;
assign _0769_ = illegal_insn_q_t0 & _0081_;
assign _0771_ = instr_fetch_err_prio_t0 & _0055_;
assign _0773_ = instr_fetch_err_prio_t0 & _0070_;
assign _0775_ = instr_fetch_err_prio_t0 & _0041_;
assign _0777_ = instr_fetch_err_prio_t0 & _0043_;
assign _0779_ = instr_fetch_err_prio_t0 & _0054_;
assign _0781_ = instr_exec_i_t0 & _0342_;
assign _0783_ = { _1354_, _1354_, _1354_, _1354_ } & { _0365_, _0004_[2:0] };
assign _0785_ = { dret_insn_t0, dret_insn_t0, dret_insn_t0, dret_insn_t0 } & { _0022_[3], _0359_[1], _0022_[1], _0359_[0] };
assign _0787_ = mret_insn_t0 & nmi_mode_o;
assign _0789_ = mret_insn_t0 & _0344_;
assign _0791_ = { mret_insn_t0, mret_insn_t0, mret_insn_t0 } & { _0118_[2], _0367_ };
assign _0793_ = { mret_insn_t0, mret_insn_t0, mret_insn_t0, mret_insn_t0 } & { _0020_[3], _0360_[1], _0020_[1], _0360_[0] };
assign _0794_ = mret_insn_t0 & _0100_;
assign _0796_ = { load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0, load_err_prio_t0 } & lsu_addr_last_i;
assign _0799_ = { store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0 } & _1250_;
assign _0801_ = { ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0 } & _1251_;
assign _0803_ = { ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0 } & _1252_;
assign _0806_ = { illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0 } & _1253_;
assign _0809_ = { instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0 } & _1254_;
assign _0811_ = { store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0, store_err_prio_t0 } & { _1255_[6:3], _0384_ };
assign _0814_ = { ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0 } & _1256_;
assign _0817_ = { ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0 } & _1257_;
assign _0819_ = { illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0 } & { _1258_[6:2], _0385_, _1258_[0] };
assign _0821_ = { instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0 } & { _1259_[6:1], _0386_ };
assign _0823_ = { ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0, ebrk_insn_prio_t0 } & { _0012_[3], _0361_[1], _0012_[1], _0361_[0] };
assign _0825_ = { ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0, ecall_insn_prio_t0 } & { _1260_[3], _0362_[1], _1260_[1], _0362_[0] };
assign _0827_ = { illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0, illegal_insn_prio_t0 } & { _1261_[3], _0363_[1], _1261_[1], _0363_[0] };
assign _0829_ = { instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0, instr_fetch_err_prio_t0 } & { _1262_[3], _0364_[1], _1262_[1], _0364_[0] };
assign _0831_ = ecall_insn_prio_t0 & _0346_;
assign _0833_ = illegal_insn_prio_t0 & _0347_;
assign _0835_ = instr_fetch_err_prio_t0 & _0348_;
assign _0837_ = ebrk_insn_prio_t0 & _0345_;
assign _0840_ = { _1377_, _1377_, _1377_, _1377_ } & _1263_;
assign _0842_ = _1377_ & _0350_;
assign _0844_ = { _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_ } & _0138_;
assign _0845_ = _1377_ & _0084_;
assign _0847_ = { _1377_, _1377_, _1377_, _1377_, _1377_, _1377_, _1377_ } & _0160_;
assign _0849_ = _1377_ & _1264_;
assign _0851_ = { _1377_, _1377_ } & { _1265_[1], _0387_ };
assign _0853_ = { _1377_, _1377_, _1377_ } & { _0094_[2], _0368_, _0094_[0] };
assign _0856_ = _1377_ & _1266_;
assign _0858_ = _1377_ & _0074_;
assign _0860_ = _1377_ & _0076_;
assign _0862_ = { irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15], irqs_i_t0[15] } & { _0142_[6], _0370_[3], _0142_[4], _0370_[2], _0142_[2], _0370_[1:0] };
assign _0865_ = { _1381_, _1381_, _1381_, _1381_, _1381_, _1381_, _1381_ } & _1267_;
assign _0867_ = { _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_, _0187_ } & \g_intg_irq_int.mem_resp_intg_err_addr_q ;
assign _0869_ = _1350_ & _0337_;
assign _0871_ = { _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_ } & _0098_;
assign _0874_ = { _1350_, _1350_, _1350_, _1350_, _1350_, _1350_, _1350_ } & _1268_;
assign _0877_ = handle_irq_t0 & _1269_;
assign _0879_ = { handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0 } & _0072_;
assign _0881_ = { handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0 } & _0082_;
assign _0883_ = handle_irq_t0 & _0339_;
assign _0885_ = { handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0 } & { _0140_[3], _0357_ };
assign _0887_ = enter_debug_mode_t0 & _0340_;
assign _0889_ = { enter_debug_mode_t0, enter_debug_mode_t0, enter_debug_mode_t0, enter_debug_mode_t0 } & { _0358_, _0000_[2:0] };
assign _0892_ = _1348_ & _1270_;
assign _0895_ = { _1348_, _1348_, _1348_, _1348_ } & _1271_;
assign _0897_ = _0064_ & jump_set_i;
assign _0899_ = _0064_ & branch_set_i;
assign _0901_ = { ready_wb_i_t0, ready_wb_i_t0, ready_wb_i_t0, ready_wb_i_t0 } & { ctrl_fsm_cs[3], _0356_, ctrl_fsm_cs[0] };
assign _0904_ = { special_req_t0, special_req_t0, special_req_t0, special_req_t0 } & _1272_;
assign _0906_ = enter_debug_mode_t0 & _0338_;
assign _0908_ = { enter_debug_mode_t0, enter_debug_mode_t0, enter_debug_mode_t0, enter_debug_mode_t0 } & { _0355_, _0103_[2:0] };
assign _0104_ = { handle_irq_t0, handle_irq_t0, handle_irq_t0, handle_irq_t0 } & { _0077_[3], _0354_ };
assign _0910_ = controller_run_o_t0 & _0069_;
assign _0912_ = controller_run_o_t0 & _0067_;
assign _0914_ = controller_run_o_t0 & _0065_;
assign _0916_ = _1379_ & _0030_;
assign _0918_ = _1379_ & _0032_;
assign _0919_ = _1432_ & _0035_;
assign _0921_ = { irqs_i_t0[0], irqs_i_t0[0], irqs_i_t0[0], irqs_i_t0[0] } & _0018_;
assign _0923_ = { irqs_i_t0[1], irqs_i_t0[1], irqs_i_t0[1], irqs_i_t0[1] } & { _0014_[3:1], _0383_ };
assign _0925_ = { irqs_i_t0[2], irqs_i_t0[2], irqs_i_t0[2], irqs_i_t0[2] } & { _0010_[3:2], _0382_, _0010_[0] };
assign _0927_ = { irqs_i_t0[3], irqs_i_t0[3], irqs_i_t0[3], irqs_i_t0[3] } & { _0006_[3:2], _0381_ };
assign _0929_ = { irqs_i_t0[4], irqs_i_t0[4], irqs_i_t0[4], irqs_i_t0[4] } & { _0002_[3], _0380_, _0002_[1:0] };
assign _0931_ = { irqs_i_t0[5], irqs_i_t0[5], irqs_i_t0[5], irqs_i_t0[5] } & { _0167_[3], _0379_[1], _0167_[1], _0379_[0] };
assign _0933_ = { irqs_i_t0[6], irqs_i_t0[6], irqs_i_t0[6], irqs_i_t0[6] } & { _0162_[3], _0378_, _0162_[0] };
assign _0935_ = { irqs_i_t0[7], irqs_i_t0[7], irqs_i_t0[7], irqs_i_t0[7] } & { _0154_[3], _0377_ };
assign _0937_ = { irqs_i_t0[8], irqs_i_t0[8], irqs_i_t0[8], irqs_i_t0[8] } & { _0376_, _0146_[2:0] };
assign _0939_ = { irqs_i_t0[9], irqs_i_t0[9], irqs_i_t0[9], irqs_i_t0[9] } & { _0375_[1], _0133_[2:1], _0375_[0] };
assign _0941_ = { irqs_i_t0[10], irqs_i_t0[10], irqs_i_t0[10], irqs_i_t0[10] } & { _0374_[1], _0114_[2], _0374_[0], _0114_[0] };
assign _0943_ = { irqs_i_t0[11], irqs_i_t0[11], irqs_i_t0[11], irqs_i_t0[11] } & { _0373_[2], _0090_[2], _0373_[1:0] };
assign _0945_ = { irqs_i_t0[12], irqs_i_t0[12], irqs_i_t0[12], irqs_i_t0[12] } & { _0372_, _0057_[1:0] };
assign _0947_ = { irqs_i_t0[13], irqs_i_t0[13], irqs_i_t0[13], irqs_i_t0[13] } & { _0371_[2:1], _0027_[1], _0371_[0] };
assign _0950_ = instr_valid_i_t0 & _1273_;
assign _0952_ = _1343_ & debug_ebreaku_i;
assign _0955_ = _1341_ & _1274_;
assign _0957_ = { debug_req_i_t0, debug_req_i_t0, debug_req_i_t0 } & { _1275_[2], _0388_ };
assign _0959_ = { _0185_, _0185_, _0185_ } & { _1276_[2:1], _0389_ };
assign _0961_ = { trigger_match_i_t0, trigger_match_i_t0, trigger_match_i_t0 } & { _1277_[2], _0390_, _1277_[0] };
assign _0964_ = { instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0, instr_fetch_err_plus2_i_t0 } & _1278_;
assign _0967_ = { instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0, instr_is_compressed_i_t0 } & _1279_;
assign _1298_ = _0563_ | _0562_;
assign _1300_ = _0566_ | _1025_;
assign _1302_ = _0569_ | _1028_;
assign _1308_ = _0571_ | _0570_;
assign _1310_ = _0574_ | _1032_;
assign ctrl_fsm_ns_t0 = _0577_ | _1035_;
assign _1312_ = _0579_ | _0578_;
assign _1314_ = _0581_ | _0580_;
assign _1316_ = _0584_ | _1041_;
assign pc_set_o_t0 = _0587_ | _1044_;
assign _1318_ = _0589_ | _0588_;
assign pc_mux_o_t0 = _0592_ | _1048_;
assign _1321_ = _0594_ | _0593_;
assign _1323_ = _0596_ | _0595_;
assign _0026_ = _0599_ | _1053_;
assign _1325_ = _0602_ | _1054_;
assign nmi_mode_d_t0 = _0605_ | _1055_;
assign flush_id_o_t0 = _0608_ | _1056_;
assign debug_csr_save_o_t0 = _0611_ | _1060_;
assign _1330_ = _0613_ | _0612_;
assign csr_mtval_o_t0 = _0616_ | _1064_;
assign _1332_ = _0619_ | _1065_;
assign csr_save_if_o_t0 = _0621_ | _0620_;
assign csr_save_cause_o_t0 = _0624_ | _1068_;
assign _1334_ = _0625_ | _0583_;
assign _1336_ = _0627_ | _0626_;
assign exc_cause_o_t0 = _0630_ | _1072_;
assign exc_pc_mux_o_t0 = _0633_ | _1075_;
assign ctrl_busy_o_t0 = _0636_ | _1078_;
assign \g_intg_irq_int.mem_resp_intg_err_irq_clear_t0  = _0747_ | _0746_;
assign \g_intg_irq_int.mem_resp_intg_err_irq_set_t0  = _0749_ | _0748_;
assign _0132_ = _0751_ | _0750_;
assign _0113_ = _0753_ | _0752_;
assign _0122_ = _0755_ | _0754_;
assign _0089_ = _0757_ | _0756_;
assign _0097_ = _0759_ | _0758_;
assign _0080_ = _0761_ | _0760_;
assign _0056_ = _0763_ | _0762_;
assign _0071_ = _0765_ | _0764_;
assign _0042_ = _0767_ | _0766_;
assign _0044_ = _0769_ | _0768_;
assign load_err_prio_t0 = _0771_ | _0770_;
assign store_err_prio_t0 = _0773_ | _0772_;
assign ebrk_insn_prio_t0 = _0775_ | _0774_;
assign ecall_insn_prio_t0 = _0777_ | _0776_;
assign illegal_insn_prio_t0 = _0779_ | _0778_;
assign halt_if_t0 = _0781_ | _0780_;
assign _0024_ = _0783_ | _0782_;
assign _0021_ = _0785_ | _0784_;
assign _0136_ = _0787_ | _0786_;
assign _0157_ = _0789_ | _0788_;
assign _0095_ = _0791_ | _0790_;
assign _0017_ = _0793_ | _0792_;
assign _0075_ = _0794_ | _0788_;
assign _1403_ = _0796_ | _0795_;
assign _1404_ = _0799_ | _1131_;
assign _1405_ = _0801_ | _0800_;
assign _1407_ = _0803_ | _0802_;
assign _1409_ = _0806_ | _1136_;
assign _0139_ = _0809_ | _1139_;
assign _1412_ = _0811_ | _0810_;
assign _1414_ = _0814_ | _1143_;
assign _1416_ = _0817_ | _1146_;
assign _1418_ = _0819_ | _0818_;
assign _0161_ = _0821_ | _0820_;
assign _1420_ = _0823_ | _0822_;
assign _1422_ = _0825_ | _0824_;
assign _1424_ = _0827_ | _0826_;
assign _0009_ = _0829_ | _0828_;
assign _1428_ = _0831_ | _0830_;
assign _1430_ = _0833_ | _0832_;
assign _0085_ = _0835_ | _0834_;
assign _1426_ = _0837_ | _0836_;
assign _0005_ = _0840_ | _1159_;
assign _0050_ = _0842_ | _0841_;
assign _0124_ = _0844_ | _0843_;
assign _0102_ = _0845_ | _0841_;
assign _0151_ = _0847_ | _0846_;
assign _0120_ = _0849_ | _1164_;
assign _0048_ = _0851_ | _0850_;
assign _0062_ = _0853_ | _0852_;
assign _0117_ = _0856_ | _1167_;
assign _0031_ = _0858_ | _0857_;
assign _0033_ = _0860_ | _0859_;
assign _0128_ = _0862_ | _0861_;
assign _0108_ = _0865_ | _1171_;
assign _0099_ = _0867_ | _0866_;
assign _0093_ = _0869_ | _0868_;
assign _0073_ = _0871_ | _0870_;
assign _0083_ = _0874_ | _1177_;
assign _0060_ = _0877_ | _1180_;
assign _0029_ = _0879_ | _0878_;
assign _0046_ = _0881_ | _0880_;
assign _0153_ = _0883_ | _0882_;
assign _0001_ = _0885_ | _0884_;
assign _0144_ = _0887_ | _0886_;
assign _0165_ = _0889_ | _0888_;
assign _0130_ = _0892_ | _1188_;
assign _0159_ = _0895_ | _1191_;
assign _0066_ = _0897_ | _0896_;
assign _0068_ = _0899_ | _0898_;
assign _0149_ = _0901_ | _0900_;
assign _0141_ = _0904_ | _1196_;
assign _0087_ = _0906_ | _0905_;
assign _0126_ = _0908_ | _0907_;
assign retain_id_t0 = _0910_ | _0909_;
assign perf_tbranch_o_t0 = _0912_ | _0911_;
assign perf_jump_o_t0 = _0914_ | _0913_;
assign csr_restore_dret_id_o_t0 = _0916_ | _0915_;
assign csr_restore_mret_id_o_t0 = _0918_ | _0917_;
assign csr_save_id_o_t0 = _0919_ | _0610_;
assign mfip_id_t0 = _0921_ | _0920_;
assign _0019_ = _0923_ | _0922_;
assign _0015_ = _0925_ | _0924_;
assign _0011_ = _0927_ | _0926_;
assign _0007_ = _0929_ | _0928_;
assign _0003_ = _0931_ | _0930_;
assign _0168_ = _0933_ | _0932_;
assign _0163_ = _0935_ | _0934_;
assign _0155_ = _0937_ | _0936_;
assign _0147_ = _0939_ | _0938_;
assign _0134_ = _0941_ | _0940_;
assign _0115_ = _0943_ | _0942_;
assign _0091_ = _0945_ | _0944_;
assign _0058_ = _0947_ | _0946_;
assign do_single_step_d_t0 = _0950_ | _1213_;
assign _1446_ = _0952_ | _0951_;
assign ebreak_into_debug_t0 = _0955_ | _1217_;
assign _1449_ = _0957_ | _0956_;
assign _1451_ = _0959_ | _0958_;
assign debug_cause_d_t0 = _0961_ | _0960_;
assign _1455_ = _0964_ | _1223_;
assign _1457_ = _0967_ | _1226_;
assign _0430_ = { _1401_, _1376_, dret_insn, mret_insn } != 4'h8;
assign _0432_ = { _1401_, _1376_, mret_insn } != 3'h5;
assign _0434_ = { _1401_, _1376_ } != 2'h3;
assign _0436_ = | { _0421_, _1401_ };
assign _0438_ = { _1436_, id_in_ready_o, handle_irq, enter_debug_mode } != 4'h8;
assign _0440_ = { _1438_, _1368_ } != 2'h2;
assign _0442_ = & { _0436_, _0434_, _0432_, _0430_ };
assign _0444_ = & { _0438_, _0440_ };
assign _0446_ = & { _0275_, mem_resp_intg_err_i };
assign _0337_ = ~ nmi_mode_o;
assign _0338_ = ~ _0034_;
assign _0339_ = ~ _0110_;
assign _0340_ = ~ _0152_;
assign _0341_ = ~ _0129_;
assign _0342_ = ~ _0025_;
assign _0343_ = ~ _0040_;
assign _0344_ = ~ _0100_;
assign _0346_ = ~ _1425_;
assign _0347_ = ~ _1427_;
assign _0348_ = ~ _1429_;
assign _0349_ = ~ _0119_;
assign _0350_ = ~ _0084_;
assign _0351_ = ~ _1333_;
assign _0352_ = ~ _1305_[2];
assign _0353_ = ~ _0039_[1:0];
assign _0354_ = ~ _0077_[2:0];
assign _0355_ = ~ _0103_[3];
assign _0356_ = ~ ctrl_fsm_cs[2:1];
assign _0357_ = ~ _0140_[2:0];
assign _0358_ = ~ _0000_[3];
assign _0359_ = ~ { _0022_[2], _0022_[0] };
assign _0360_ = ~ { _0020_[2], _0020_[0] };
assign _0361_ = ~ { _0012_[2], _0012_[0] };
assign _0362_ = ~ { _1419_[2], _1419_[0] };
assign _0363_ = ~ { _1421_[2], _1421_[0] };
assign _0364_ = ~ { _1423_[2], _1423_[0] };
assign _0365_ = ~ _0004_[3];
assign _0366_ = ~ { _0023_[2], _0023_[0] };
assign _0367_ = ~ _0118_[1:0];
assign _0368_ = ~ _0094_[1];
assign _0369_ = ~ _0061_[1];
assign _0370_ = ~ { _0142_[5], _0142_[3], _0142_[1:0] };
assign _0371_ = ~ { _0027_[3:2], _0027_[0] };
assign _0372_ = ~ _0057_[3:2];
assign _0373_ = ~ { _0090_[3], _0090_[1:0] };
assign _0374_ = ~ { _0114_[3], _0114_[1] };
assign _0375_ = ~ { _0133_[3], _0133_[0] };
assign _0376_ = ~ _0146_[3];
assign _0377_ = ~ _0154_[2:0];
assign _0378_ = ~ _0162_[2:1];
assign _0379_ = ~ { _0167_[2], _0167_[0] };
assign _0380_ = ~ _0002_[2];
assign _0381_ = ~ _0006_[1:0];
assign _0382_ = ~ _0010_[1];
assign _0383_ = ~ _0014_[0];
assign _0384_ = ~ _1410_[2:0];
assign _0385_ = ~ _1415_[1];
assign _0386_ = ~ _1417_[0];
assign _0387_ = ~ _1453_[0];
assign _0388_ = ~ _1447_[1:0];
assign _0389_ = ~ _1448_[0];
assign _0390_ = ~ _1450_[1];
assign _0448_ = | { _1444_, _1442_, _1440_, _1431_ };
assign _0450_ = | { _1440_, _1433_, _1431_ };
assign _0452_ = | { _1441_, _1438_, _1401_ };
assign _0454_ = | { _1442_, _1440_, _1436_, _1435_, _1433_, _1431_, _1401_ };
assign _0455_ = | { _1441_, _1440_, _1438_, _1431_ };
assign _0391_ = ~ _0448_;
assign _0392_ = ~ _0450_;
assign _0393_ = ~ _1387_;
assign _0394_ = ~ _1389_;
assign _0395_ = ~ store_err_i;
assign _0396_ = ~ wfi_insn;
assign _0397_ = ~ _1393_;
assign _0398_ = ~ _1395_;
assign _0399_ = ~ special_req_pc_change;
assign _0400_ = ~ _0172_;
assign _0401_ = ~ \g_intg_irq_int.mem_resp_intg_err_irq_set ;
assign _0402_ = ~ enter_debug_mode_prio_d;
assign _0403_ = ~ irq_nm_ext_i;
assign _0404_ = ~ csr_mstatus_mie_i;
assign _0405_ = ~ stall_id_i;
assign _0407_ = ~ illegal_insn_d;
assign _0408_ = ~ load_err_i;
assign _0409_ = ~ csr_pipe_flush;
assign _0410_ = ~ id_exception_o;
assign _0411_ = ~ exc_req_lsu;
assign _0412_ = ~ special_req_flush_only;
assign _0413_ = ~ do_single_step_d;
assign _0414_ = ~ _0176_;
assign _0415_ = ~ irq_nm_int;
assign _0416_ = ~ _0182_;
assign _0417_ = ~ ebreak_into_debug;
assign _0418_ = ~ stall_wb_i;
assign _0419_ = ~ retain_id;
assign _0420_ = ~ flush_id_o;
assign _0546_ = _1339_ & _0274_;
assign _0549_ = _0449_ & _0260_;
assign _0552_ = _0451_ & _0260_;
assign _0555_ = controller_run_o_t0 & _0265_;
assign _0558_ = _1432_ & _0260_;
assign _0685_ = ecall_insn_t0 & _0276_;
assign _0688_ = _1388_ & _0407_;
assign _0691_ = _1390_ & _0279_;
assign _0694_ = store_err_i_t0 & _0408_;
assign _0697_ = wfi_insn_t0 & _0409_;
assign _0700_ = mret_insn_t0 & _0281_;
assign _0703_ = _1394_ & _0410_;
assign _0706_ = _1396_ & _0411_;
assign _0709_ = special_req_pc_change_t0 & _0412_;
assign _0712_ = instr_valid_i_t0 & ready_wb_i;
assign _0715_ = _0173_ & _0401_;
assign _0718_ = \g_intg_irq_int.mem_resp_intg_err_irq_set_t0  & _0275_;
assign _0721_ = debug_req_i_t0 & _0413_;
assign _0724_ = enter_debug_mode_prio_d_t0 & _0414_;
assign _0727_ = irq_nm_ext_i_t0 & _0415_;
assign _0729_ = csr_mstatus_mie_i_t0 & _0330_;
assign _0732_ = irq_nm_t0 & _0416_;
assign _0735_ = debug_mode_o_t0 & _0417_;
assign _0737_ = stall_id_i_t0 & _0418_;
assign _0740_ = stall_t0 & _0419_;
assign _0743_ = _1386_ & _0420_;
assign _0547_ = _1439_ & _0273_;
assign _0550_ = _1379_ & _0391_;
assign _0553_ = _1379_ & _0392_;
assign _0556_ = _0453_ & _0261_;
assign _0559_ = _1379_ & _0268_;
assign _0686_ = ebrk_insn_t0 & _0277_;
assign _0689_ = illegal_insn_d_t0 & _0393_;
assign _0692_ = instr_fetch_err_prio_t0 & _0394_;
assign _0695_ = load_err_i_t0 & _0395_;
assign _0698_ = csr_pipe_flush_t0 & _0396_;
assign _0701_ = dret_insn_t0 & _0283_;
assign _0704_ = id_exception_o_t0 & _0397_;
assign _0707_ = exc_req_lsu_t0 & _0398_;
assign _0710_ = special_req_flush_only_t0 & _0399_;
assign _0713_ = ready_wb_i_t0 & _0329_;
assign _0716_ = \g_intg_irq_int.mem_resp_intg_err_irq_set_t0  & _0400_;
assign _0719_ = \g_intg_irq_int.mem_resp_intg_err_irq_pending_q_t0  & _0401_;
assign _0722_ = do_single_step_d_t0 & _0247_;
assign _0725_ = _0177_ & _0402_;
assign _0728_ = irq_nm_int_t0 & _0403_;
assign _0730_ = _1343_ & _0404_;
assign _0733_ = _0183_ & _0237_;
assign _0736_ = ebreak_into_debug_t0 & _0248_;
assign _0738_ = stall_wb_i_t0 & _0405_;
assign _0741_ = retain_id_t0 & _0243_;
assign _0744_ = flush_id_o_t0 & _0406_;
assign _0548_ = _1339_ & _1439_;
assign _0551_ = _0449_ & _1379_;
assign _0554_ = _0451_ & _1379_;
assign _0557_ = controller_run_o_t0 & _0453_;
assign _0560_ = _1432_ & _1379_;
assign _0687_ = ecall_insn_t0 & ebrk_insn_t0;
assign _0690_ = _1388_ & illegal_insn_d_t0;
assign _0693_ = _1390_ & instr_fetch_err_prio_t0;
assign _0696_ = store_err_i_t0 & load_err_i_t0;
assign _0699_ = wfi_insn_t0 & csr_pipe_flush_t0;
assign _0702_ = mret_insn_t0 & dret_insn_t0;
assign _0705_ = _1394_ & id_exception_o_t0;
assign _0708_ = _1396_ & exc_req_lsu_t0;
assign _0711_ = special_req_pc_change_t0 & special_req_flush_only_t0;
assign _0714_ = instr_valid_i_t0 & ready_wb_i_t0;
assign _0717_ = _0173_ & \g_intg_irq_int.mem_resp_intg_err_irq_set_t0 ;
assign _0720_ = \g_intg_irq_int.mem_resp_intg_err_irq_set_t0  & \g_intg_irq_int.mem_resp_intg_err_irq_pending_q_t0 ;
assign _0723_ = debug_req_i_t0 & do_single_step_d_t0;
assign _0726_ = enter_debug_mode_prio_d_t0 & _0177_;
assign _0731_ = csr_mstatus_mie_i_t0 & _1343_;
assign _0734_ = irq_nm_t0 & _0183_;
assign _0739_ = stall_id_i_t0 & stall_wb_i_t0;
assign _0742_ = stall_t0 & retain_id_t0;
assign _0745_ = _1386_ & flush_id_o_t0;
assign _1017_ = _0546_ | _0547_;
assign _1018_ = _0549_ | _0550_;
assign _1019_ = _0552_ | _0553_;
assign _1020_ = _0555_ | _0556_;
assign _1021_ = _0558_ | _0559_;
assign _1094_ = _0685_ | _0686_;
assign _1095_ = _0688_ | _0689_;
assign _1096_ = _0691_ | _0692_;
assign _1097_ = _0694_ | _0695_;
assign _1098_ = _0697_ | _0698_;
assign _1099_ = _0700_ | _0701_;
assign _1100_ = _0703_ | _0704_;
assign _1101_ = _0706_ | _0707_;
assign _1102_ = _0709_ | _0710_;
assign _1103_ = _0712_ | _0713_;
assign _1104_ = _0715_ | _0716_;
assign _1105_ = _0718_ | _0719_;
assign _1106_ = _0721_ | _0722_;
assign _1107_ = _0724_ | _0725_;
assign _1108_ = _0727_ | _0728_;
assign _1109_ = _0729_ | _0730_;
assign _1110_ = _0732_ | _0733_;
assign _1111_ = _0735_ | _0736_;
assign _1112_ = _0737_ | _0738_;
assign _1113_ = _0740_ | _0741_;
assign _1114_ = _0743_ | _0744_;
assign _0971_ = _1017_ | _0548_;
assign _0973_ = _1018_ | _0551_;
assign _0969_ = _1019_ | _0554_;
assign _0975_ = _1020_ | _0557_;
assign _0977_ = _1021_ | _0560_;
assign _1388_ = _1094_ | _0687_;
assign _1390_ = _1095_ | _0690_;
assign _1392_ = _1096_ | _0693_;
assign exc_req_lsu_t0 = _1097_ | _0696_;
assign special_req_flush_only_t0 = _1098_ | _0699_;
assign _1394_ = _1099_ | _0702_;
assign _1396_ = _1100_ | _0705_;
assign special_req_pc_change_t0 = _1101_ | _0708_;
assign special_req_t0 = _1102_ | _0711_;
assign id_wb_pending_t0 = _1103_ | _0714_;
assign \g_intg_irq_int.mem_resp_intg_err_irq_pending_d_t0  = _1104_ | _0717_;
assign irq_nm_int_t0 = _1105_ | _0720_;
assign _1398_ = _1106_ | _0723_;
assign enter_debug_mode_t0 = _1107_ | _0726_;
assign irq_nm_t0 = _1108_ | _0518_;
assign irq_enabled_t0 = _1109_ | _0731_;
assign _1400_ = _1110_ | _0734_;
assign _0013_[3] = _1111_ | _0652_;
assign stall_t0 = _1112_ | _0739_;
assign _1386_ = _1113_ | _0742_;
assign instr_valid_clear_o_t0 = _1114_ | _0745_;
assign _0421_ = | { _1440_, _1431_ };
assign _0970_ = _1441_ | _1438_;
assign _0972_ = _0448_ | _1401_;
assign _0968_ = _0450_ | _1401_;
assign _0974_ = _1435_ | _0452_;
assign _0976_ = _1431_ | _1401_;
assign _0422_ = | { _0968_, _1436_, _1435_ };
assign _1297_ = _1401_ ? _0023_ : 4'h5;
assign _1299_ = _1435_ ? _0158_ : _0125_;
assign _1301_ = _0968_ ? _1297_ : _1299_;
assign _1303_ = _1438_ ? _0039_ : 4'h3;
assign { _1233_[3], _1305_[2], _1233_[1:0] } = _1444_ ? 4'h1 : 4'h0;
assign _1307_ = _1442_ ? 4'h4 : { _1233_[3], _1305_[2], _1233_[1:0] };
assign _1309_ = _0970_ ? _1303_ : _1307_;
assign ctrl_fsm_ns = _0422_ ? _1301_ : _1309_;
assign _1311_ = _1401_ ? _0119_ : 1'h1;
assign _1313_ = _1435_ ? _0063_ : 1'h0;
assign _1315_ = _1433_ ? _0034_ : _1313_;
assign pc_set_o = _0972_ ? _1311_ : _1315_;
assign _1317_ = _1401_ ? _0061_ : 3'h2;
assign _1319_ = _1435_ ? 3'h1 : 3'h0;
assign pc_mux_o = _0968_ ? _1317_ : _1319_;
assign _1320_ = _0452_ ? 1'h1 : _0129_;
assign _1322_ = _1436_ ? _0086_ : 1'h0;
assign _0025_ = _0974_ ? _1320_ : _1322_;
assign debug_mode_d = _1401_ ? _0040_ : 1'h1;
assign _1324_ = _1433_ ? _0059_ : nmi_mode_o;
assign nmi_mode_d = _1401_ ? _0116_ : _1324_;
assign _1326_ = _0455_ ? 1'h1 : 1'h0;
assign flush_id_o = _1401_ ? _0049_ : _1326_;
assign _1327_ = _1440_ ? 1'h1 : 1'h0;
assign debug_csr_save_o = _1431_ ? _0035_ : _1327_;
assign _1329_ = _1433_ ? _0028_ : 32'd0;
assign csr_mtval_o = _1401_ ? _0123_ : _1329_;
assign _1331_ = _1401_ ? _0101_ : _0035_;
assign csr_save_if_o = _1440_ ? 1'h1 : _1333_;
assign csr_save_cause_o = _0976_ ? _1331_ : csr_save_if_o;
assign _1333_ = _1433_ ? _0034_ : 1'h0;
assign _1335_ = _1433_ ? _0045_ : 7'h00;
assign exc_cause_o = _1401_ ? _0150_ : _1335_;
assign _1337_ = _0421_ ? 2'h2 : 2'h1;
assign exc_pc_mux_o = _1401_ ? _0047_ : _1337_;
assign _1338_ = _1441_ ? 1'h0 : 1'h1;
assign ctrl_busy_o = _1438_ ? _0037_ : _1338_;
assign _0424_ = | { _0437_, _0435_, _0433_, _0431_ };
assign _0425_ = | { _0441_, _0439_ };
assign _0426_ = | { \g_intg_irq_int.mem_resp_intg_err_irq_pending_q_t0 , mem_resp_intg_err_i_t0 };
assign _1014_ = { _0436_, _0434_, _0432_, _0430_ } | { _0437_, _0435_, _0433_, _0431_ };
assign _1015_ = { _0438_, _0440_ } | { _0439_, _0441_ };
assign _1016_ = { _0275_, mem_resp_intg_err_i } | { \g_intg_irq_int.mem_resp_intg_err_irq_pending_q_t0 , mem_resp_intg_err_i_t0 };
assign _0427_ = & _1014_;
assign _0428_ = & _1015_;
assign _0429_ = & _1016_;
assign _0443_ = _0424_ & _0427_;
assign _0445_ = _0425_ & _0428_;
assign _0447_ = _0426_ & _0429_;
assign _1342_ = ! /* src = "generated/sv2v_out.v:12439.44-12439.64" */ priv_mode_i;
assign _1340_ = priv_mode_i == /* src = "generated/sv2v_out.v:12644.39-12644.59" */ 2'h3;
assign _1344_ = _1370_ && /* src = "generated/sv2v_out.v:12557.9-12557.69" */ _1372_;
assign _1345_ = _1356_ && /* src = "generated/sv2v_out.v:12559.10-12559.32" */ _1357_;
assign _1347_ = _1345_ && /* src = "generated/sv2v_out.v:12559.9-12559.51" */ _1358_;
assign _1349_ = irq_nm && /* src = "generated/sv2v_out.v:12576.10-12576.31" */ _1359_;
assign _1351_ = ebreak_into_debug && /* src = "generated/sv2v_out.v:12610.9-12610.43" */ _1360_;
assign _1352_ = ebrk_insn_prio && /* src = "generated/sv2v_out.v:12682.38-12682.73" */ ebreak_into_debug;
assign _1353_ = enter_debug_mode_prio_q && /* src = "generated/sv2v_out.v:12682.9-12682.74" */ _1361_;
assign _1355_ = ! /* src = "generated/sv2v_out.v:12404.25-12404.38" */ irq_nm_ext_i;
assign _1356_ = ! /* src = "generated/sv2v_out.v:12559.10-12559.16" */ stall;
assign _1357_ = ! /* src = "generated/sv2v_out.v:12559.20-12559.32" */ special_req;
assign _1358_ = ! /* src = "generated/sv2v_out.v:12559.37-12559.51" */ id_wb_pending;
assign _1359_ = ! /* src = "generated/sv2v_out.v:12576.20-12576.31" */ nmi_mode_o;
assign _1360_ = ! /* src = "generated/sv2v_out.v:12610.30-12610.43" */ debug_mode_o;
assign _1361_ = ! /* src = "generated/sv2v_out.v:12682.36-12682.74" */ _1352_;
assign _1362_ = irq_nm || /* src = "generated/sv2v_out.v:12524.12-12524.35" */ irq_pending_i;
assign _1364_ = _1362_ || /* src = "generated/sv2v_out.v:12524.11-12524.51" */ debug_req_i;
assign _1366_ = _1364_ || /* src = "generated/sv2v_out.v:12524.10-12524.68" */ debug_mode_o;
assign _1368_ = _1366_ || /* src = "generated/sv2v_out.v:12524.9-12524.92" */ debug_single_step_i;
assign _1369_ = branch_set_i || /* src = "generated/sv2v_out.v:12549.9-12549.35" */ jump_set_i;
assign _1370_ = enter_debug_mode || /* src = "generated/sv2v_out.v:12557.10-12557.40" */ handle_irq;
assign _1372_ = stall || /* src = "generated/sv2v_out.v:12557.46-12557.68" */ id_wb_pending;
assign _1374_ = exc_req_q || /* src = "generated/sv2v_out.v:12623.10-12623.34" */ store_err_q;
assign _1376_ = _1374_ || /* src = "generated/sv2v_out.v:12623.9-12623.49" */ load_err_q;
assign _1378_ = ctrl_fsm_cs != /* src = "generated/sv2v_out.v:12336.88-12336.107" */ 4'h6;
assign _1380_ = | /* src = "generated/sv2v_out.v:12582.15-12582.52" */ irqs_i[14:0];
assign _1382_ = ~ /* src = "generated/sv2v_out.v:12342.41-12342.52" */ ready_wb_i;
assign _1383_ = ~ /* src = "generated/sv2v_out.v:12412.80-12412.108" */ \g_intg_irq_int.mem_resp_intg_err_irq_clear ;
assign _1384_ = ~ /* src = "generated/sv2v_out.v:12697.35-12697.43" */ halt_if;
assign _1385_ = ~ /* src = "generated/sv2v_out.v:12698.31-12698.51" */ _0406_;
assign _1387_ = ecall_insn | /* src = "generated/sv2v_out.v:12336.24-12336.46" */ ebrk_insn;
assign _1389_ = _1387_ | /* src = "generated/sv2v_out.v:12336.23-12336.64" */ illegal_insn_d;
assign _1391_ = _1389_ | /* src = "generated/sv2v_out.v:12336.22-12336.83" */ instr_fetch_err;
assign exc_req_lsu = store_err_i | /* src = "generated/sv2v_out.v:12337.23-12337.47" */ load_err_i;
assign special_req_flush_only = wfi_insn | /* src = "generated/sv2v_out.v:12339.34-12339.59" */ csr_pipe_flush;
assign _1393_ = mret_insn | /* src = "generated/sv2v_out.v:12340.35-12340.56" */ dret_insn;
assign _1395_ = _1393_ | /* src = "generated/sv2v_out.v:12340.34-12340.69" */ id_exception_o;
assign special_req_pc_change = _1395_ | /* src = "generated/sv2v_out.v:12340.33-12340.84" */ exc_req_lsu;
assign special_req = special_req_pc_change | /* src = "generated/sv2v_out.v:12341.23-12341.69" */ special_req_flush_only;
assign id_wb_pending = instr_valid_i | /* src = "generated/sv2v_out.v:12342.25-12342.52" */ _1382_;
assign \g_intg_irq_int.mem_resp_intg_err_irq_pending_d  = _0172_ | /* src = "generated/sv2v_out.v:12412.45-12412.137" */ \g_intg_irq_int.mem_resp_intg_err_irq_set ;
assign irq_nm_int = \g_intg_irq_int.mem_resp_intg_err_irq_set  | /* src = "generated/sv2v_out.v:12422.24-12422.83" */ \g_intg_irq_int.mem_resp_intg_err_irq_pending_q ;
assign _1397_ = debug_req_i | /* src = "generated/sv2v_out.v:12435.36-12435.66" */ do_single_step_d;
assign enter_debug_mode = enter_debug_mode_prio_d | /* src = "generated/sv2v_out.v:12436.28-12436.87" */ _0176_;
assign irq_nm = irq_nm_ext_i | /* src = "generated/sv2v_out.v:12438.18-12438.43" */ irq_nm_int;
assign irq_enabled = csr_mstatus_mie_i | /* src = "generated/sv2v_out.v:12439.23-12439.65" */ _1342_;
assign _1399_ = irq_nm | /* src = "generated/sv2v_out.v:12440.80-12440.118" */ _0182_;
assign _0345_ = debug_mode_o | /* src = "generated/sv2v_out.v:12646.12-12646.44" */ ebreak_into_debug;
assign stall = stall_id_i | /* src = "generated/sv2v_out.v:12696.17-12696.40" */ stall_wb_i;
assign _0406_ = stall | /* src = "generated/sv2v_out.v:12698.33-12698.50" */ retain_id;
assign instr_valid_clear_o = _1385_ | /* src = "generated/sv2v_out.v:12698.31-12698.62" */ flush_id_o;
/* src = "generated/sv2v_out.v:12413.4-12421.8" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  <= 1'h0;
else \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  <= \g_intg_irq_int.mem_resp_intg_err_irq_pending_d ;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME nmi_mode_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) nmi_mode_o <= 1'h0;
else nmi_mode_o <= nmi_mode_d;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME load_err_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) load_err_q <= 1'h0;
else load_err_q <= load_err_i;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME store_err_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) store_err_q <= 1'h0;
else store_err_q <= store_err_i;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME exc_req_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) exc_req_q <= 1'h0;
else exc_req_q <= id_exception_o;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME illegal_insn_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) illegal_insn_q <= 1'h0;
else illegal_insn_q <= illegal_insn_d;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME do_single_step_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) do_single_step_q <= 1'h0;
else do_single_step_q <= do_single_step_d;
/* src = "generated/sv2v_out.v:12699.2-12722.5" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME enter_debug_mode_prio_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) enter_debug_mode_prio_q <= 1'h0;
else enter_debug_mode_prio_q <= enter_debug_mode_prio_d;
/* src = "generated/sv2v_out.v:12452.2-12456.35" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_controller\WritebackStage=1'0\BranchPredictor=1'0\MemECC=1'1  */
/* PC_TAINT_INFO STATE_NAME debug_cause_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) debug_cause_o <= 3'h0;
else debug_cause_o <= debug_cause_d;
assign _0053_ = mem_resp_intg_err_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12407.14-12407.33|generated/sv2v_out.v:12407.10-12410.8" */ 1'h1 : 1'h0;
assign _0051_ = _0171_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12404.10-12404.38|generated/sv2v_out.v:12404.6-12405.42" */ 1'h1 : 1'h0;
assign \g_intg_irq_int.mem_resp_intg_err_irq_clear  = \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12403.9-12403.40|generated/sv2v_out.v:12403.5-12410.8" */ _0051_ : 1'h0;
assign \g_intg_irq_int.mem_resp_intg_err_irq_set  = \g_intg_irq_int.mem_resp_intg_err_irq_pending_q  ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12403.9-12403.40|generated/sv2v_out.v:12403.5-12410.8" */ 1'h0 : _0053_;
assign _0145_ = load_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12385.14-12385.24|generated/sv2v_out.v:12385.10-12386.27" */ 1'h1 : 1'h0;
assign _0137_ = store_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12383.14-12383.25|generated/sv2v_out.v:12383.10-12386.27" */ 1'h1 : 1'h0;
assign _0131_ = store_err_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12383.14-12383.25|generated/sv2v_out.v:12383.10-12386.27" */ 1'h0 : _0145_;
assign _0106_ = ebrk_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12381.14-12381.23|generated/sv2v_out.v:12381.10-12386.27" */ 1'h1 : 1'h0;
assign _0112_ = ebrk_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12381.14-12381.23|generated/sv2v_out.v:12381.10-12386.27" */ 1'h0 : _0131_;
assign _0121_ = ebrk_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12381.14-12381.23|generated/sv2v_out.v:12381.10-12386.27" */ 1'h0 : _0137_;
assign _0081_ = ecall_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12379.14-12379.24|generated/sv2v_out.v:12379.10-12386.27" */ 1'h1 : 1'h0;
assign _0088_ = ecall_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12379.14-12379.24|generated/sv2v_out.v:12379.10-12386.27" */ 1'h0 : _0112_;
assign _0096_ = ecall_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12379.14-12379.24|generated/sv2v_out.v:12379.10-12386.27" */ 1'h0 : _0121_;
assign _0079_ = ecall_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12379.14-12379.24|generated/sv2v_out.v:12379.10-12386.27" */ 1'h0 : _0106_;
assign _0054_ = illegal_insn_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12377.14-12377.28|generated/sv2v_out.v:12377.10-12386.27" */ 1'h1 : 1'h0;
assign _0055_ = illegal_insn_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12377.14-12377.28|generated/sv2v_out.v:12377.10-12386.27" */ 1'h0 : _0088_;
assign _0070_ = illegal_insn_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12377.14-12377.28|generated/sv2v_out.v:12377.10-12386.27" */ 1'h0 : _0096_;
assign _0041_ = illegal_insn_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12377.14-12377.28|generated/sv2v_out.v:12377.10-12386.27" */ 1'h0 : _0079_;
assign _0043_ = illegal_insn_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12377.14-12377.28|generated/sv2v_out.v:12377.10-12386.27" */ 1'h0 : _0081_;
assign instr_fetch_err_prio = instr_fetch_err ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12375.9-12375.24|generated/sv2v_out.v:12375.5-12386.27" */ 1'h1 : 1'h0;
assign load_err_prio = instr_fetch_err ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12375.9-12375.24|generated/sv2v_out.v:12375.5-12386.27" */ 1'h0 : _0055_;
assign store_err_prio = instr_fetch_err ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12375.9-12375.24|generated/sv2v_out.v:12375.5-12386.27" */ 1'h0 : _0070_;
assign ebrk_insn_prio = instr_fetch_err ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12375.9-12375.24|generated/sv2v_out.v:12375.5-12386.27" */ 1'h0 : _0041_;
assign ecall_insn_prio = instr_fetch_err ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12375.9-12375.24|generated/sv2v_out.v:12375.5-12386.27" */ 1'h0 : _0043_;
assign illegal_insn_prio = instr_fetch_err ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12375.9-12375.24|generated/sv2v_out.v:12375.5-12386.27" */ 1'h0 : _0054_;
assign halt_if = instr_exec_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12690.7-12690.20|generated/sv2v_out.v:12690.3-12691.19" */ _0025_ : 1'h1;
assign _0023_ = _1353_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12682.9-12682.74|generated/sv2v_out.v:12682.5-12683.25" */ 4'h8 : _0004_;
assign _0022_ = wfi_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12680.14-12680.22|generated/sv2v_out.v:12680.10-12681.25" */ 4'h2 : 4'h5;
assign _0105_ = dret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12674.14-12674.23|generated/sv2v_out.v:12674.10-12681.25" */ 1'h0 : 1'hx;
assign _0100_ = dret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12674.14-12674.23|generated/sv2v_out.v:12674.10-12681.25" */ 1'h1 : 1'h0;
assign _0118_ = dret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12674.14-12674.23|generated/sv2v_out.v:12674.10-12681.25" */ 3'h4 : 3'h0;
assign _0020_ = dret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12674.14-12674.23|generated/sv2v_out.v:12674.10-12681.25" */ 4'h5 : _0022_;
assign _0135_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12667.14-12667.23|generated/sv2v_out.v:12667.10-12681.25" */ 1'h0 : nmi_mode_o;
assign _0076_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12667.14-12667.23|generated/sv2v_out.v:12667.10-12681.25" */ 1'h1 : 1'h0;
assign _0156_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12667.14-12667.23|generated/sv2v_out.v:12667.10-12681.25" */ 1'h1 : _0100_;
assign _0094_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12667.14-12667.23|generated/sv2v_out.v:12667.10-12681.25" */ 3'h3 : _0118_;
assign _0078_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12667.14-12667.23|generated/sv2v_out.v:12667.10-12681.25" */ 1'hx : _0105_;
assign _0016_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12667.14-12667.23|generated/sv2v_out.v:12667.10-12681.25" */ 4'h5 : _0020_;
assign _0074_ = mret_insn ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12667.14-12667.23|generated/sv2v_out.v:12667.10-12681.25" */ 1'h0 : _0100_;
assign _0012_ = _0345_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12646.12-12646.44|generated/sv2v_out.v:12646.8-12654.51" */ 4'h9 : 4'h5;
assign _0109_ = _0345_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12646.12-12646.44|generated/sv2v_out.v:12646.8-12654.51" */ 1'h0 : 1'h1;
assign _0166_ = _0345_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12646.12-12646.44|generated/sv2v_out.v:12646.8-12654.51" */ 7'h00 : 7'h03;
assign _1402_ = load_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ lsu_addr_last_i : 32'd0;
assign _1251_ = store_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ lsu_addr_last_i : _1402_;
assign _1252_ = ebrk_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 32'd0 : _1251_;
assign _1406_ = ecall_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 32'd0 : _1252_;
assign _1408_ = illegal_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ _1456_ : _1406_;
assign _0138_ = instr_fetch_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ _1454_ : _1408_;
assign { _1255_[6:3], _1410_[2:0] } = load_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 7'h05 : 7'h00;
assign _1411_ = store_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 7'h07 : { _1255_[6:3], _1410_[2:0] };
assign _1413_ = ebrk_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ _0166_ : _1411_;
assign { _1258_[6:2], _1415_[1], _1258_[0] } = ecall_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ _1458_ : _1413_;
assign { _1259_[6:1], _1417_[0] } = illegal_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 7'h02 : { _1258_[6:2], _1415_[1], _1258_[0] };
assign _0160_ = instr_fetch_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 7'h01 : { _1259_[6:1], _1417_[0] };
assign { _1260_[3], _1419_[2], _1260_[1], _1419_[0] } = ebrk_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ _0012_ : 4'h5;
assign { _1261_[3], _1421_[2], _1261_[1], _1421_[0] } = ecall_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 4'h5 : { _1260_[3], _1419_[2], _1260_[1], _1419_[0] };
assign { _1262_[3], _1423_[2], _1262_[1], _1423_[0] } = illegal_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 4'h5 : { _1261_[3], _1421_[2], _1261_[1], _1421_[0] };
assign _0008_ = instr_fetch_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 4'h5 : { _1262_[3], _1423_[2], _1262_[1], _1423_[0] };
assign _1427_ = ecall_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 1'h1 : _1425_;
assign _1429_ = illegal_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 1'h1 : _1427_;
assign _0084_ = instr_fetch_err_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ 1'h1 : _1429_;
assign _1425_ = ebrk_insn_prio ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12635.6-12665.13" */ _0109_ : 1'h1;
assign _0004_ = _1376_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ _0008_ : _0016_;
assign _0049_ = _1376_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ _0084_ : 1'h1;
assign _0123_ = _1376_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ _0138_ : 32'd0;
assign _0101_ = _1376_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ _0084_ : 1'h0;
assign _0150_ = _1376_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ _0160_ : 7'h00;
assign _0119_ = _1376_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ _0084_ : _0156_;
assign _0047_ = _1376_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ { _1265_[1], _1453_[0] } : 2'h1;
assign _0061_ = _1376_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ 3'h2 : _0094_;
assign _0040_ = _1376_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ 1'hx : _0078_;
assign _0116_ = _1376_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ nmi_mode_o : _0135_;
assign _0030_ = _1376_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ 1'h0 : _0074_;
assign _0032_ = _1376_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12623.9-12623.49|generated/sv2v_out.v:12623.5-12681.25" */ 1'h0 : _0076_;
assign _0035_ = _1351_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12610.9-12610.43|generated/sv2v_out.v:12610.5-12614.8" */ 1'h1 : 1'h0;
assign _0142_ = irqs_i[17] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12586.15-12586.25|generated/sv2v_out.v:12586.11-12589.48" */ 7'h23 : 7'h27;
assign _0127_ = irqs_i[15] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12584.15-12584.25|generated/sv2v_out.v:12584.11-12589.48" */ 7'h2b : _0142_;
assign _0107_ = _1380_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12582.15-12582.52|generated/sv2v_out.v:12582.11-12589.48" */ { 3'h3, mfip_id } : _0127_;
assign _0098_ = _0186_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12578.11-12578.37|generated/sv2v_out.v:12578.7-12579.39" */ \g_intg_irq_int.mem_resp_intg_err_addr_q  : 32'd0;
assign _0092_ = _1349_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12576.10-12576.31|generated/sv2v_out.v:12576.6-12589.48" */ 1'h1 : nmi_mode_o;
assign _0072_ = _1349_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12576.10-12576.31|generated/sv2v_out.v:12576.6-12589.48" */ _0098_ : 32'd0;
assign _0082_ = _1349_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12576.10-12576.31|generated/sv2v_out.v:12576.6-12589.48" */ _1452_ : _0107_;
assign _0059_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12572.9-12572.19|generated/sv2v_out.v:12572.5-12590.8" */ _0092_ : nmi_mode_o;
assign _0028_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12572.9-12572.19|generated/sv2v_out.v:12572.5-12590.8" */ _0072_ : 32'd0;
assign _0045_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12572.9-12572.19|generated/sv2v_out.v:12572.5-12590.8" */ _0082_ : 7'h00;
assign _0034_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12572.9-12572.19|generated/sv2v_out.v:12572.5-12590.8" */ 1'h1 : 1'h0;
assign _0152_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12564.15-12564.25|generated/sv2v_out.v:12564.11-12567.9" */ 1'h1 : _0110_;
assign _0000_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12564.15-12564.25|generated/sv2v_out.v:12564.11-12567.9" */ 4'h7 : _0140_;
assign _0143_ = enter_debug_mode ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12560.10-12560.26|generated/sv2v_out.v:12560.6-12567.9" */ 1'h1 : _0152_;
assign _0164_ = enter_debug_mode ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12560.10-12560.26|generated/sv2v_out.v:12560.6-12567.9" */ 4'h8 : _0000_;
assign _0129_ = _1347_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12559.9-12559.51|generated/sv2v_out.v:12559.5-12567.9" */ _0143_ : _0110_;
assign _0158_ = _1347_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12559.9-12559.51|generated/sv2v_out.v:12559.5-12567.9" */ _0164_ : _0140_;
assign _0110_ = _1344_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12557.9-12557.69|generated/sv2v_out.v:12557.5-12558.21" */ 1'h1 : 1'h0;
assign _0065_ = _1369_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12549.9-12549.35|generated/sv2v_out.v:12549.5-12553.8" */ jump_set_i : 1'h0;
assign _0067_ = _1369_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12549.9-12549.35|generated/sv2v_out.v:12549.5-12553.8" */ branch_set_i : 1'h0;
assign _0063_ = _1369_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12549.9-12549.35|generated/sv2v_out.v:12549.5-12553.8" */ 1'h1 : 1'h0;
assign _0148_ = ready_wb_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12546.10-12546.37|generated/sv2v_out.v:12546.6-12547.26" */ 4'h6 : ctrl_fsm_cs;
assign _0140_ = special_req ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12544.9-12544.20|generated/sv2v_out.v:12544.5-12548.8" */ _0148_ : ctrl_fsm_cs;
assign _0069_ = special_req ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12544.9-12544.20|generated/sv2v_out.v:12544.5-12548.8" */ 1'h1 : 1'h0;
assign _0086_ = enter_debug_mode ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12536.9-12536.25|generated/sv2v_out.v:12536.5-12539.8" */ 1'h1 : _0034_;
assign _0125_ = enter_debug_mode ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12536.9-12536.25|generated/sv2v_out.v:12536.5-12539.8" */ 4'h8 : _0103_;
assign _0103_ = handle_irq ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12532.9-12532.19|generated/sv2v_out.v:12532.5-12535.8" */ 4'h7 : _0077_;
assign _0077_ = id_in_ready_o ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12530.9-12530.22|generated/sv2v_out.v:12530.5-12531.25" */ 4'h5 : 4'hx;
assign _0039_ = _1368_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12524.9-12524.92|generated/sv2v_out.v:12524.5-12527.25" */ 4'h4 : 4'hx;
assign _0037_ = _1368_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12524.9-12524.92|generated/sv2v_out.v:12524.5-12527.25" */ 1'h1 : 1'h0;
assign _1444_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ ctrl_fsm_cs;
assign instr_req_o = _0454_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 1'h1 : 1'h0;
assign _1442_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h1;
assign retain_id = _1435_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ _0069_ : 1'h0;
assign _1436_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h4;
assign _1433_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h7;
assign controller_run_o = _1435_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 1'h1 : 1'h0;
assign _1401_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h6;
assign _1440_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h8;
assign _1438_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h3;
assign _1441_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h2;
assign perf_tbranch_o = _1435_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ _0067_ : 1'h0;
assign perf_jump_o = _1435_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ _0065_ : 1'h0;
assign _1435_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h5;
assign _1431_ = ctrl_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 4'h9;
assign debug_mode_entering_o = _0421_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ 1'h1 : 1'h0;
assign csr_restore_dret_id_o = _1401_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ _0030_ : 1'h0;
assign csr_restore_mret_id_o = _1401_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ _0032_ : 1'h0;
assign csr_save_id_o = _1431_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12500.3-12689.10" */ _0035_ : 1'h0;
assign mfip_id = irqs_i[0] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h0 : _0018_;
assign _0018_ = irqs_i[1] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h1 : _0014_;
assign _0014_ = irqs_i[2] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h2 : _0010_;
assign _0010_ = irqs_i[3] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h3 : _0006_;
assign _0006_ = irqs_i[4] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h4 : _0002_;
assign _0002_ = irqs_i[5] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h5 : _0167_;
assign _0167_ = irqs_i[6] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h6 : _0162_;
assign _0162_ = irqs_i[7] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h7 : _0154_;
assign _0154_ = irqs_i[8] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h8 : _0146_;
assign _0146_ = irqs_i[9] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'h9 : _0133_;
assign _0133_ = irqs_i[10] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'ha : _0114_;
assign _0114_ = irqs_i[11] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'hb : _0090_;
assign _0090_ = irqs_i[12] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'hc : _0057_;
assign _0057_ = irqs_i[13] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'hd : _0027_;
assign _0027_ = irqs_i[14] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12446.9-12446.22|generated/sv2v_out.v:12446.5-12447.23" */ 4'he : 4'h0;
assign do_single_step_d = instr_valid_i ? /* src = "generated/sv2v_out.v:12434.29-12434.99" */ _0174_ : do_single_step_q;
assign _1445_ = _1342_ ? /* src = "generated/sv2v_out.v:12437.72-12437.117" */ debug_ebreaku_i : 1'h0;
assign ebreak_into_debug = _1340_ ? /* src = "generated/sv2v_out.v:12437.30-12437.118" */ debug_ebreakm_i : _1445_;
assign { _1275_[2], _1447_[1:0] } = do_single_step_d ? /* src = "generated/sv2v_out.v:12451.119-12451.149" */ 3'h4 : 3'h0;
assign { _1276_[2:1], _1448_[0] } = debug_req_i ? /* src = "generated/sv2v_out.v:12451.97-12451.150" */ 3'h3 : { _1275_[2], _1447_[1:0] };
assign { _1277_[2], _1450_[1], _1277_[0] } = _0184_ ? /* src = "generated/sv2v_out.v:12451.52-12451.151" */ 3'h1 : { _1276_[2:1], _1448_[0] };
assign debug_cause_d = trigger_match_i ? /* src = "generated/sv2v_out.v:12451.26-12451.152" */ 3'h2 : { _1277_[2], _1450_[1], _1277_[0] };
assign _1452_ = irq_nm_ext_i ? /* src = "generated/sv2v_out.v:12577.22-12577.87" */ 7'h3f : 7'h40;
assign { _1265_[1], _1453_[0] } = debug_mode_o ? /* src = "generated/sv2v_out.v:12626.22-12626.48" */ 2'h3 : 2'h0;
assign _1454_ = instr_fetch_err_plus2_i ? /* src = "generated/sv2v_out.v:12638.23-12638.74" */ _0169_ : pc_id_i;
assign _1456_ = instr_is_compressed_i ? /* src = "generated/sv2v_out.v:12642.23-12642.99" */ { 16'h0000, instr_compressed_i } : instr_i;
assign _1458_ = _1340_ ? /* src = "generated/sv2v_out.v:12644.39-12644.119" */ 7'h0b : 7'h08;
assign _0013_[2:0] = { _0013_[3], 2'h0 };
assign _1233_[2] = _0352_;
assign _1255_[2:0] = _0384_;
assign _1258_[1] = _0385_;
assign _1259_[0] = _0386_;
assign { _1260_[2], _1260_[0] } = _0362_;
assign { _1261_[2], _1261_[0] } = _0363_;
assign { _1262_[2], _1262_[0] } = _0364_;
assign _1265_[0] = _0387_;
assign _1275_[1:0] = _0388_;
assign _1276_[0] = _0389_;
assign _1277_[1] = _0390_;
assign { _1305_[3], _1305_[1:0] } = { _1233_[3], _1233_[1:0] };
assign _1306_[3:1] = 3'h0;
assign _1410_[6:3] = _1255_[6:3];
assign { _1415_[6:2], _1415_[0] } = { _1258_[6:2], _1258_[0] };
assign _1417_[6:1] = _1259_[6:1];
assign { _1419_[3], _1419_[1] } = { _1260_[3], _1260_[1] };
assign { _1421_[3], _1421_[1] } = { _1261_[3], _1261_[1] };
assign { _1423_[3], _1423_[1] } = { _1262_[3], _1262_[1] };
assign _1447_[2] = _1275_[2];
assign _1448_[2:1] = _1276_[2:1];
assign { _1450_[2], _1450_[0] } = { _1277_[2], _1277_[0] };
assign _1453_[1] = _1265_[1];
assign csr_save_wb_o = 1'h0;
assign csr_save_wb_o_t0 = 1'h0;
assign nt_branch_mispredict_o = 1'h0;
assign nt_branch_mispredict_o_t0 = 1'h0;
assign wb_exception_o = 1'h0;
assign wb_exception_o_t0 = 1'h0;
endmodule

module \$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000 (clk_i, rst_ni, counter_inc_i, counterh_we_i, counter_we_i, counter_val_i, counter_val_o, counter_val_upd_o, counter_inc_i_t0, counter_val_i_t0, counter_val_o_t0, counter_val_upd_o_t0, counter_we_i_t0, counterh_we_i_t0);
/* src = "generated/sv2v_out.v:13613.2-13627.5" */
wire [63:0] _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13613.2-13627.5" */
wire [63:0] _001_;
wire [63:0] _002_;
wire _003_;
wire _004_;
wire _005_;
wire [1:0] _006_;
wire _007_;
wire [1:0] _008_;
wire _009_;
wire [63:0] _010_;
wire [31:0] _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
/* cellift = 32'd1 */
wire _019_;
wire _020_;
/* cellift = 32'd1 */
wire _021_;
wire _022_;
/* cellift = 32'd1 */
wire _023_;
wire _024_;
/* cellift = 32'd1 */
wire _025_;
wire _026_;
/* cellift = 32'd1 */
wire _027_;
wire [63:0] _028_;
wire [31:0] _029_;
wire [31:0] _030_;
wire [31:0] _031_;
wire [31:0] _032_;
wire [31:0] _033_;
wire [31:0] _034_;
wire [1:0] _035_;
wire [1:0] _036_;
wire _037_;
wire _038_;
wire _039_;
wire [63:0] _040_;
wire [63:0] _041_;
wire [63:0] _042_;
wire [63:0] _043_;
wire [31:0] _044_;
wire [31:0] _045_;
wire [31:0] _046_;
wire [31:0] _047_;
wire [31:0] _048_;
wire [31:0] _049_;
wire [31:0] _050_;
wire [31:0] _051_;
wire [1:0] _052_;
wire [1:0] _053_;
wire _054_;
wire [63:0] _055_;
wire [63:0] _056_;
wire [63:0] _057_;
wire [63:0] _058_;
wire [31:0] _059_;
wire [31:0] _060_;
wire [63:0] _061_;
wire [31:0] _062_;
wire [31:0] _063_;
wire [63:0] _064_;
wire _065_;
wire _066_;
wire [63:0] _067_;
wire [63:0] _068_;
/* src = "generated/sv2v_out.v:13599.13-13599.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:13611.27-13611.36" */
wire [63:0] counter_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13611.27-13611.36" */
wire [63:0] counter_d_t0;
/* src = "generated/sv2v_out.v:13601.13-13601.26" */
input counter_inc_i;
wire counter_inc_i;
/* cellift = 32'd1 */
input counter_inc_i_t0;
wire counter_inc_i_t0;
/* src = "generated/sv2v_out.v:13609.13-13609.25" */
wire [63:0] counter_load;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13609.13-13609.25" */
wire [63:0] counter_load_t0;
/* src = "generated/sv2v_out.v:13608.28-13608.39" */
wire [63:0] counter_upd;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13608.28-13608.39" */
wire [63:0] counter_upd_t0;
/* src = "generated/sv2v_out.v:13604.20-13604.33" */
input [31:0] counter_val_i;
wire [31:0] counter_val_i;
/* cellift = 32'd1 */
input [31:0] counter_val_i_t0;
wire [31:0] counter_val_i_t0;
/* src = "generated/sv2v_out.v:13605.21-13605.34" */
output [63:0] counter_val_o;
reg [63:0] counter_val_o;
/* cellift = 32'd1 */
output [63:0] counter_val_o_t0;
reg [63:0] counter_val_o_t0;
/* src = "generated/sv2v_out.v:13606.21-13606.38" */
output [63:0] counter_val_upd_o;
wire [63:0] counter_val_upd_o;
/* cellift = 32'd1 */
output [63:0] counter_val_upd_o_t0;
wire [63:0] counter_val_upd_o_t0;
/* src = "generated/sv2v_out.v:13603.13-13603.25" */
input counter_we_i;
wire counter_we_i;
/* cellift = 32'd1 */
input counter_we_i_t0;
wire counter_we_i_t0;
/* src = "generated/sv2v_out.v:13602.13-13602.26" */
input counterh_we_i;
wire counterh_we_i;
/* cellift = 32'd1 */
input counterh_we_i_t0;
wire counterh_we_i_t0;
/* src = "generated/sv2v_out.v:13600.13-13600.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:13610.6-13610.8" */
wire we;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:13610.6-13610.8" */
wire we_t0;
assign counter_upd = counter_val_o + /* src = "generated/sv2v_out.v:13612.23-13612.86" */ 64'h0000000000000001;
assign _002_ = ~ counter_val_o_t0;
assign _028_ = counter_val_o & _002_;
assign _067_ = _028_ + 64'h0000000000000001;
assign _043_ = counter_val_o | counter_val_o_t0;
assign _068_ = _043_ + 64'h0000000000000001;
assign _061_ = _067_ ^ _068_;
assign counter_upd_t0 = _061_ | counter_val_o_t0;
assign _003_ = ~ _024_;
assign _004_ = ~ _026_;
assign _062_ = counter_d[63:32] ^ counter_val_o[63:32];
assign _063_ = counter_d[31:0] ^ counter_val_o[31:0];
assign _044_ = counter_d_t0[63:32] | counter_val_o_t0[63:32];
assign _048_ = counter_d_t0[31:0] | counter_val_o_t0[31:0];
assign _045_ = _062_ | _044_;
assign _049_ = _063_ | _048_;
assign _029_ = { _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_, _024_ } & counter_d_t0[63:32];
assign _032_ = { _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_, _026_ } & counter_d_t0[31:0];
assign _030_ = { _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_, _003_ } & counter_val_o_t0[63:32];
assign _033_ = { _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_, _004_ } & counter_val_o_t0[31:0];
assign _031_ = _045_ & { _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_, _025_ };
assign _034_ = _049_ & { _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_, _027_ };
assign _046_ = _029_ | _030_;
assign _050_ = _032_ | _033_;
assign _047_ = _046_ | _031_;
assign _051_ = _050_ | _034_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000  */
/* PC_TAINT_INFO STATE_NAME counter_val_o_t0[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o_t0[63:32] <= 32'd0;
else counter_val_o_t0[63:32] <= _047_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000  */
/* PC_TAINT_INFO STATE_NAME counter_val_o_t0[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o_t0[31:0] <= 32'd0;
else counter_val_o_t0[31:0] <= _051_;
assign _005_ = | { we_t0, counterh_we_i_t0 };
assign _006_ = ~ { we_t0, counterh_we_i_t0 };
assign _036_ = { we, counterh_we_i } & _006_;
assign _065_ = _036_ == { _006_[1], 1'h0 };
assign _066_ = _036_ == _006_;
assign _021_ = _065_ & _005_;
assign _023_ = _066_ & _005_;
/* src = "generated/sv2v_out.v:13629.2-13633.27" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000  */
/* PC_TAINT_INFO STATE_NAME counter_val_o[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o[63:32] <= 32'd0;
else if (_024_) counter_val_o[63:32] <= counter_d[63:32];
/* src = "generated/sv2v_out.v:13629.2-13633.27" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_counter\CounterWidth=s32'00000000000000000000000001000000  */
/* PC_TAINT_INFO STATE_NAME counter_val_o[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) counter_val_o[31:0] <= 32'd0;
else if (_026_) counter_val_o[31:0] <= counter_d[31:0];
assign _007_ = | { we_t0, counter_inc_i_t0 };
assign _008_ = ~ { we_t0, counter_inc_i_t0 };
assign _035_ = { we, counter_inc_i } & _008_;
assign _009_ = ! _035_;
assign _019_ = _009_ & _007_;
assign _010_ = ~ { we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we };
assign _011_ = ~ { counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i };
assign _056_ = { we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0 } | _010_;
assign _059_ = { counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0 } | _011_;
assign _055_ = { counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0, counter_inc_i_t0 } | { counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i, counter_inc_i };
assign _057_ = { we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0 } | { we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we, we };
assign _060_ = { counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0, counterh_we_i_t0 } | { counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i, counterh_we_i };
assign _040_ = _001_ & _056_;
assign counter_load_t0[31:0] = counter_val_i_t0 & _059_;
assign _001_ = counter_upd_t0 & _055_;
assign _041_ = counter_load_t0 & _057_;
assign counter_load_t0[63:32] = counter_val_i_t0 & _060_;
assign _058_ = _040_ | _041_;
assign _064_ = _000_ ^ counter_load;
assign _042_ = { we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0, we_t0 } & _064_;
assign counter_d_t0 = _042_ | _058_;
assign _018_ = | { we, counter_inc_i };
assign _020_ = { we, counterh_we_i } != 2'h2;
assign _022_ = { we, counterh_we_i } != 2'h3;
assign _024_ = & { _018_, _020_ };
assign _026_ = & { _018_, _022_ };
assign _012_ = ~ counter_we_i;
assign _013_ = ~ counterh_we_i;
assign _037_ = counter_we_i_t0 & _013_;
assign _038_ = counterh_we_i_t0 & _012_;
assign _039_ = counter_we_i_t0 & counterh_we_i_t0;
assign _054_ = _037_ | _038_;
assign we_t0 = _054_ | _039_;
assign _014_ = | { _021_, _019_ };
assign _015_ = | { _023_, _019_ };
assign _052_ = { _018_, _020_ } | { _019_, _021_ };
assign _053_ = { _018_, _022_ } | { _019_, _023_ };
assign _016_ = & _052_;
assign _017_ = & _053_;
assign _025_ = _014_ & _016_;
assign _027_ = _015_ & _017_;
assign we = counter_we_i | /* src = "generated/sv2v_out.v:13614.8-13614.36" */ counterh_we_i;
assign _000_ = counter_inc_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13623.12-13623.25|generated/sv2v_out.v:13623.8-13626.44" */ counter_upd : 64'hxxxxxxxxxxxxxxxx;
assign counter_d = we ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13621.7-13621.9|generated/sv2v_out.v:13621.3-13626.44" */ counter_load : _000_;
assign counter_load[63:32] = counterh_we_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13617.7-13617.20|generated/sv2v_out.v:13617.3-13620.6" */ counter_val_i : 32'hxxxxxxxx;
assign counter_load[31:0] = counterh_we_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:13617.7-13617.20|generated/sv2v_out.v:13617.3-13620.6" */ 32'hxxxxxxxx : counter_val_i;
assign counter_val_upd_o = 64'h0000000000000000;
assign counter_val_upd_o_t0 = 64'h0000000000000000;
endmodule

module \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1 (clk_i, rst_ni, clear_i, busy_o, in_valid_i, in_addr_i, in_rdata_i, in_err_i, out_valid_o, out_ready_i, out_addr_o, out_rdata_o, out_err_o, out_err_plus2_o, out_valid_o_t0, out_ready_i_t0, out_rdata_o_t0, out_err_plus2_o_t0, out_err_o_t0, out_addr_o_t0, in_valid_i_t0
, in_rdata_i_t0, in_err_i_t0, in_addr_i_t0, clear_i_t0, busy_o_t0);
/* src = "generated/sv2v_out.v:16127.2-16142.6" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16127.2-16142.6" */
wire _001_;
/* src = "generated/sv2v_out.v:16122.40-16122.75" */
wire _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16122.40-16122.75" */
wire _003_;
/* src = "generated/sv2v_out.v:16122.91-16122.112" */
wire _004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16122.91-16122.112" */
wire _005_;
/* src = "generated/sv2v_out.v:16122.117-16122.168" */
wire _006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16122.117-16122.168" */
wire _007_;
/* src = "generated/sv2v_out.v:16123.35-16123.55" */
wire _008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16123.35-16123.55" */
wire _009_;
/* src = "generated/sv2v_out.v:16123.59-16123.80" */
wire _010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16123.59-16123.80" */
wire _011_;
/* src = "generated/sv2v_out.v:16123.58-16123.93" */
wire _012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16123.58-16123.93" */
wire _013_;
/* src = "generated/sv2v_out.v:16124.48-16124.71" */
wire _014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16124.48-16124.71" */
wire _015_;
/* src = "generated/sv2v_out.v:16143.36-16143.61" */
wire _016_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16143.36-16143.61" */
wire _017_;
/* src = "generated/sv2v_out.v:16174.30-16174.63" */
wire _018_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16174.30-16174.63" */
wire _019_;
/* src = "generated/sv2v_out.v:16174.30-16174.63" */
wire _020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16174.30-16174.63" */
wire _021_;
/* src = "generated/sv2v_out.v:16177.26-16177.56" */
wire _022_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16177.26-16177.56" */
wire _023_;
/* src = "generated/sv2v_out.v:16177.61-16177.108" */
wire _024_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16177.61-16177.108" */
wire _025_;
/* src = "generated/sv2v_out.v:16177.26-16177.56" */
wire _026_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16177.26-16177.56" */
wire _027_;
/* src = "generated/sv2v_out.v:16177.61-16177.108" */
wire _028_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16177.61-16177.108" */
wire _029_;
wire [30:0] _030_;
wire [30:0] _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire [1:0] _038_;
wire [1:0] _039_;
wire _040_;
wire _041_;
wire [31:0] _042_;
wire [31:0] _043_;
wire [31:0] _044_;
wire _045_;
wire [30:0] _046_;
wire _047_;
wire [31:0] _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire [30:0] _064_;
wire [30:0] _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire [31:0] _136_;
wire [31:0] _137_;
wire [31:0] _138_;
wire _139_;
wire _140_;
wire _141_;
wire [31:0] _142_;
wire [31:0] _143_;
wire [31:0] _144_;
wire _145_;
wire _146_;
wire _147_;
wire [31:0] _148_;
wire [31:0] _149_;
wire [31:0] _150_;
wire [30:0] _151_;
wire [30:0] _152_;
wire [30:0] _153_;
wire [1:0] _154_;
wire [1:0] _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire [31:0] _198_;
wire [31:0] _199_;
wire [31:0] _200_;
wire [31:0] _201_;
wire [31:0] _202_;
wire [31:0] _203_;
wire _204_;
wire _205_;
wire _206_;
wire [31:0] _207_;
wire [31:0] _208_;
wire [31:0] _209_;
wire _210_;
wire _211_;
wire _212_;
wire _213_;
wire _214_;
wire _215_;
wire _216_;
wire _217_;
wire _218_;
wire _219_;
wire _220_;
wire [30:0] _221_;
wire [30:0] _222_;
wire [30:0] _223_;
wire _224_;
wire _225_;
wire _226_;
wire _227_;
wire _228_;
wire _229_;
wire [31:0] _230_;
wire [31:0] _231_;
wire [31:0] _232_;
wire [31:0] _233_;
wire [31:0] _234_;
wire [31:0] _235_;
wire _236_;
wire _237_;
wire _238_;
wire _239_;
wire _240_;
wire _241_;
wire _242_;
wire [30:0] _243_;
wire [30:0] _244_;
wire [30:0] _245_;
wire _246_;
wire _247_;
wire _248_;
wire _249_;
wire _250_;
wire _251_;
wire _252_;
wire _253_;
wire _254_;
wire _255_;
wire _256_;
wire _257_;
wire _258_;
wire _259_;
wire _260_;
wire _261_;
wire _262_;
wire _263_;
wire _264_;
wire _265_;
wire _266_;
wire _267_;
wire _268_;
wire _269_;
wire _270_;
wire _271_;
wire _272_;
wire [31:0] _273_;
wire [31:0] _274_;
wire [31:0] _275_;
wire [31:0] _276_;
wire _277_;
wire _278_;
wire _279_;
wire _280_;
wire [31:0] _281_;
wire [31:0] _282_;
wire [31:0] _283_;
wire [31:0] _284_;
wire _285_;
wire _286_;
wire _287_;
wire _288_;
wire [31:0] _289_;
wire [31:0] _290_;
wire [31:0] _291_;
wire [31:0] _292_;
wire [30:0] _293_;
wire [30:0] _294_;
wire [30:0] _295_;
wire [30:0] _296_;
wire _297_;
wire _298_;
wire _299_;
wire _300_;
wire _301_;
wire _302_;
wire _303_;
wire _304_;
wire _305_;
wire _306_;
wire _307_;
wire _308_;
wire _309_;
wire _310_;
wire _311_;
wire _312_;
wire _313_;
wire _314_;
wire [31:0] _315_;
wire [31:0] _316_;
wire [31:0] _317_;
wire [31:0] _318_;
wire [31:0] _319_;
wire [31:0] _320_;
wire _321_;
wire _322_;
wire _323_;
wire [31:0] _324_;
wire [31:0] _325_;
wire [31:0] _326_;
wire _327_;
wire _328_;
wire _329_;
wire _330_;
wire _331_;
wire [30:0] _332_;
wire [30:0] _333_;
wire [30:0] _334_;
wire _335_;
wire _336_;
wire _337_;
wire _338_;
wire [31:0] _339_;
wire [31:0] _340_;
wire [31:0] _341_;
wire [31:0] _342_;
wire _343_;
wire _344_;
wire _345_;
wire _346_;
wire [30:0] _347_;
wire _348_;
wire [31:0] _349_;
wire _350_;
wire [31:0] _351_;
wire _352_;
wire [31:0] _353_;
wire [30:0] _354_;
wire _355_;
wire _356_;
wire _357_;
wire [31:0] _358_;
wire [31:0] _359_;
wire _360_;
wire [31:0] _361_;
wire _362_;
wire _363_;
wire _364_;
wire [30:0] _365_;
wire _366_;
wire _367_;
wire [31:0] _368_;
wire _369_;
wire _370_;
wire _371_;
wire [30:0] _372_;
wire [30:0] _373_;
/* src = "generated/sv2v_out.v:16125.36-16125.57" */
wire _374_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16125.36-16125.57" */
wire _375_;
/* src = "generated/sv2v_out.v:16126.34-16126.53" */
wire _376_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16126.34-16126.53" */
wire _377_;
/* src = "generated/sv2v_out.v:16125.61-16125.65" */
wire _378_;
/* src = "generated/sv2v_out.v:16145.56-16145.70" */
wire _379_;
/* src = "generated/sv2v_out.v:16164.51-16164.73" */
wire _380_;
/* src = "generated/sv2v_out.v:16122.39-16122.87" */
wire _381_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16122.39-16122.87" */
wire _382_;
/* src = "generated/sv2v_out.v:16122.129-16122.167" */
wire _383_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16122.129-16122.167" */
wire _384_;
/* src = "generated/sv2v_out.v:16122.90-16122.169" */
wire _385_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16122.90-16122.169" */
wire _386_;
/* src = "generated/sv2v_out.v:16164.51-16164.89" */
wire _387_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16164.51-16164.89" */
wire _388_;
/* src = "generated/sv2v_out.v:16112.7-16112.20" */
wire addr_incr_two;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16112.7-16112.20" */
wire addr_incr_two_t0;
/* src = "generated/sv2v_out.v:16110.7-16110.28" */
wire aligned_is_compressed;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16110.7-16110.28" */
wire aligned_is_compressed_t0;
/* src = "generated/sv2v_out.v:16080.31-16080.37" */
output [1:0] busy_o;
wire [1:0] busy_o;
/* cellift = 32'd1 */
output [1:0] busy_o_t0;
wire [1:0] busy_o_t0;
/* src = "generated/sv2v_out.v:16079.13-16079.20" */
input clear_i;
wire clear_i;
/* cellift = 32'd1 */
input clear_i_t0;
wire clear_i_t0;
/* src = "generated/sv2v_out.v:16077.13-16077.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:16101.21-16101.29" */
wire [2:0] entry_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16101.21-16101.29" */
wire [2:0] entry_en_t0;
/* src = "generated/sv2v_out.v:16105.7-16105.10" */
wire err;
/* src = "generated/sv2v_out.v:16094.21-16094.26" */
wire [2:0] err_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16094.21-16094.26" */
wire [2:0] err_d_t0;
/* src = "generated/sv2v_out.v:16107.7-16107.16" */
wire err_plus2;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16107.7-16107.16" */
wire err_plus2_t0;
/* src = "generated/sv2v_out.v:16095.20-16095.25" */
reg [2:0] err_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16095.20-16095.25" */
reg [2:0] err_q_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16105.7-16105.10" */
wire err_t0;
/* src = "generated/sv2v_out.v:16106.7-16106.20" */
wire err_unaligned;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16106.7-16106.20" */
wire err_unaligned_t0;
/* src = "generated/sv2v_out.v:16082.20-16082.29" */
input [31:0] in_addr_i;
wire [31:0] in_addr_i;
/* cellift = 32'd1 */
input [31:0] in_addr_i_t0;
wire [31:0] in_addr_i_t0;
/* src = "generated/sv2v_out.v:16084.13-16084.21" */
input in_err_i;
wire in_err_i;
/* cellift = 32'd1 */
input in_err_i_t0;
wire in_err_i_t0;
/* src = "generated/sv2v_out.v:16083.20-16083.30" */
input [31:0] in_rdata_i;
wire [31:0] in_rdata_i;
/* cellift = 32'd1 */
input [31:0] in_rdata_i_t0;
wire [31:0] in_rdata_i_t0;
/* src = "generated/sv2v_out.v:16081.13-16081.23" */
input in_valid_i;
wire in_valid_i;
/* cellift = 32'd1 */
input in_valid_i_t0;
wire in_valid_i_t0;
/* src = "generated/sv2v_out.v:16114.14-16114.26" */
wire [31:1] instr_addr_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16114.14-16114.26" */
wire [31:1] instr_addr_d_t0;
/* src = "generated/sv2v_out.v:16116.7-16116.20" */
wire instr_addr_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16116.7-16116.20" */
wire instr_addr_en_t0;
/* src = "generated/sv2v_out.v:16113.14-16113.29" */
wire [31:1] instr_addr_next;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16113.14-16113.29" */
wire [31:1] instr_addr_next_t0;
/* src = "generated/sv2v_out.v:16115.13-16115.25" */
reg [31:1] instr_addr_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16115.13-16115.25" */
reg [31:1] instr_addr_q_t0;
/* src = "generated/sv2v_out.v:16098.21-16098.38" */
wire [2:0] lowest_free_entry;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16098.21-16098.38" */
wire [2:0] lowest_free_entry_t0;
/* src = "generated/sv2v_out.v:16087.21-16087.31" */
output [31:0] out_addr_o;
wire [31:0] out_addr_o;
/* cellift = 32'd1 */
output [31:0] out_addr_o_t0;
wire [31:0] out_addr_o_t0;
/* src = "generated/sv2v_out.v:16089.13-16089.22" */
output out_err_o;
wire out_err_o;
/* cellift = 32'd1 */
output out_err_o_t0;
wire out_err_o_t0;
/* src = "generated/sv2v_out.v:16090.13-16090.28" */
output out_err_plus2_o;
wire out_err_plus2_o;
/* cellift = 32'd1 */
output out_err_plus2_o_t0;
wire out_err_plus2_o_t0;
/* src = "generated/sv2v_out.v:16088.20-16088.31" */
output [31:0] out_rdata_o;
wire [31:0] out_rdata_o;
/* cellift = 32'd1 */
output [31:0] out_rdata_o_t0;
wire [31:0] out_rdata_o_t0;
/* src = "generated/sv2v_out.v:16086.13-16086.24" */
input out_ready_i;
wire out_ready_i;
/* cellift = 32'd1 */
input out_ready_i_t0;
wire out_ready_i_t0;
/* src = "generated/sv2v_out.v:16085.13-16085.24" */
output out_valid_o;
wire out_valid_o;
/* cellift = 32'd1 */
output out_valid_o_t0;
wire out_valid_o_t0;
/* src = "generated/sv2v_out.v:16102.7-16102.15" */
wire pop_fifo;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16102.7-16102.15" */
wire pop_fifo_t0;
/* src = "generated/sv2v_out.v:16103.14-16103.19" */
wire [31:0] rdata;
/* src = "generated/sv2v_out.v:16092.28-16092.35" */
wire [95:0] rdata_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16092.28-16092.35" */
wire [95:0] rdata_d_t0;
/* src = "generated/sv2v_out.v:16093.27-16093.34" */
reg [95:0] rdata_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16093.27-16093.34" */
reg [95:0] rdata_q_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16103.14-16103.19" */
wire [31:0] rdata_t0;
/* src = "generated/sv2v_out.v:16104.14-16104.29" */
wire [31:0] rdata_unaligned;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16104.14-16104.29" */
wire [31:0] rdata_unaligned_t0;
/* src = "generated/sv2v_out.v:16078.13-16078.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:16111.7-16111.30" */
wire unaligned_is_compressed;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16111.7-16111.30" */
wire unaligned_is_compressed_t0;
/* src = "generated/sv2v_out.v:16108.7-16108.12" */
wire valid;
/* src = "generated/sv2v_out.v:16096.21-16096.28" */
wire [2:0] valid_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16096.21-16096.28" */
wire [2:0] valid_d_t0;
/* src = "generated/sv2v_out.v:16100.21-16100.33" */
wire [2:0] valid_popped;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16100.21-16100.33" */
wire [2:0] valid_popped_t0;
/* src = "generated/sv2v_out.v:16099.21-16099.33" */
wire [2:0] valid_pushed;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16099.21-16099.33" */
wire [2:0] valid_pushed_t0;
/* src = "generated/sv2v_out.v:16097.20-16097.27" */
reg [2:0] valid_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16097.20-16097.27" */
reg [2:0] valid_q_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16108.7-16108.12" */
wire valid_t0;
/* src = "generated/sv2v_out.v:16109.7-16109.22" */
wire valid_unaligned;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:16109.7-16109.22" */
wire valid_unaligned_t0;
assign instr_addr_next = instr_addr_q + /* src = "generated/sv2v_out.v:16145.27-16145.86" */ { 29'h00000000, _379_, addr_incr_two };
assign _002_ = err_q[1] & /* src = "generated/sv2v_out.v:16122.40-16122.75" */ _040_;
assign _004_ = valid_q[0] & /* src = "generated/sv2v_out.v:16122.91-16122.112" */ err_q[0];
assign _006_ = in_err_i & /* src = "generated/sv2v_out.v:16122.117-16122.168" */ _383_;
assign _008_ = err_q[1] & /* src = "generated/sv2v_out.v:16123.35-16123.55" */ _059_;
assign _010_ = in_err_i & /* src = "generated/sv2v_out.v:16123.59-16123.80" */ valid_q[0];
assign _012_ = _010_ & /* src = "generated/sv2v_out.v:16123.58-16123.93" */ _059_;
assign _014_ = valid_q[0] & /* src = "generated/sv2v_out.v:16124.48-16124.71" */ in_valid_i;
assign unaligned_is_compressed = _374_ & /* src = "generated/sv2v_out.v:16125.35-16125.65" */ _378_;
assign aligned_is_compressed = _376_ & /* src = "generated/sv2v_out.v:16126.33-16126.61" */ _378_;
assign _016_ = out_ready_i & /* src = "generated/sv2v_out.v:16164.21-16164.46" */ out_valid_o;
assign pop_fifo = _016_ & /* src = "generated/sv2v_out.v:16164.20-16164.90" */ _387_;
assign lowest_free_entry[1] = _045_ & /* src = "generated/sv2v_out.v:16172.35-16172.63" */ valid_q[0];
assign valid_d[0] = valid_popped[0] & /* src = "generated/sv2v_out.v:16176.24-16176.50" */ _053_;
assign valid_d[1] = valid_popped[1] & /* src = "generated/sv2v_out.v:16176.24-16176.50" */ _053_;
assign _022_ = valid_pushed[1] & /* src = "generated/sv2v_out.v:16177.26-16177.56" */ pop_fifo;
assign _018_ = in_valid_i & /* src = "generated/sv2v_out.v:16177.62-16177.95" */ lowest_free_entry[0];
assign _024_ = _018_ & /* src = "generated/sv2v_out.v:16177.61-16177.108" */ _047_;
assign _026_ = valid_pushed[2] & /* src = "generated/sv2v_out.v:16177.26-16177.56" */ pop_fifo;
assign _020_ = in_valid_i & /* src = "generated/sv2v_out.v:16177.62-16177.95" */ lowest_free_entry[1];
assign _028_ = _020_ & /* src = "generated/sv2v_out.v:16177.61-16177.108" */ _047_;
assign lowest_free_entry[2] = _049_ & /* src = "generated/sv2v_out.v:16182.40-16182.80" */ valid_q[1];
assign valid_d[2] = valid_popped[2] & /* src = "generated/sv2v_out.v:16185.30-16185.64" */ _053_;
assign entry_en[2] = in_valid_i & /* src = "generated/sv2v_out.v:16186.31-16186.72" */ lowest_free_entry[2];
assign _030_ = ~ instr_addr_q_t0;
assign _031_ = ~ { 29'h00000000, addr_incr_two_t0, addr_incr_two_t0 };
assign _064_ = instr_addr_q & _030_;
assign _065_ = { 29'h00000000, _379_, addr_incr_two } & _031_;
assign _372_ = _064_ + _065_;
assign _243_ = instr_addr_q | instr_addr_q_t0;
assign _244_ = { 29'h00000000, _379_, addr_incr_two } | { 29'h00000000, addr_incr_two_t0, addr_incr_two_t0 };
assign _373_ = _243_ + _244_;
assign _347_ = _372_ ^ _373_;
assign _245_ = _347_ | instr_addr_q_t0;
assign instr_addr_next_t0 = _245_ | { 29'h00000000, addr_incr_two_t0, addr_incr_two_t0 };
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME valid_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) valid_q_t0 <= 3'h0;
else valid_q_t0 <= valid_d_t0;
assign _032_ = ~ entry_en[2];
assign _033_ = ~ entry_en[1];
assign _034_ = ~ entry_en[0];
assign _035_ = ~ instr_addr_en;
assign _348_ = in_err_i ^ err_q[2];
assign _349_ = in_rdata_i ^ rdata_q[95:64];
assign _350_ = err_d[1] ^ err_q[1];
assign _351_ = rdata_d[63:32] ^ rdata_q[63:32];
assign _352_ = err_d[0] ^ err_q[0];
assign _353_ = rdata_d[31:0] ^ rdata_q[31:0];
assign _354_ = instr_addr_d ^ instr_addr_q;
assign _269_ = in_err_i_t0 | err_q_t0[2];
assign _273_ = in_rdata_i_t0 | rdata_q_t0[95:64];
assign _277_ = err_d_t0[1] | err_q_t0[1];
assign _281_ = rdata_d_t0[63:32] | rdata_q_t0[63:32];
assign _285_ = err_d_t0[0] | err_q_t0[0];
assign _289_ = rdata_d_t0[31:0] | rdata_q_t0[31:0];
assign _293_ = instr_addr_d_t0 | instr_addr_q_t0;
assign _270_ = _348_ | _269_;
assign _274_ = _349_ | _273_;
assign _278_ = _350_ | _277_;
assign _282_ = _351_ | _281_;
assign _286_ = _352_ | _285_;
assign _290_ = _353_ | _289_;
assign _294_ = _354_ | _293_;
assign _133_ = entry_en[2] & in_err_i_t0;
assign _136_ = { entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2], entry_en[2] } & in_rdata_i_t0;
assign _139_ = entry_en[1] & err_d_t0[1];
assign _142_ = { entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1], entry_en[1] } & rdata_d_t0[63:32];
assign _145_ = entry_en[0] & err_d_t0[0];
assign _148_ = { entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0], entry_en[0] } & rdata_d_t0[31:0];
assign _151_ = { instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en, instr_addr_en } & instr_addr_d_t0;
assign _134_ = _032_ & err_q_t0[2];
assign _137_ = { _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_, _032_ } & rdata_q_t0[95:64];
assign _140_ = _033_ & err_q_t0[1];
assign _143_ = { _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_, _033_ } & rdata_q_t0[63:32];
assign _146_ = _034_ & err_q_t0[0];
assign _149_ = { _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_, _034_ } & rdata_q_t0[31:0];
assign _152_ = { _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_, _035_ } & instr_addr_q_t0;
assign _135_ = _270_ & entry_en_t0[2];
assign _138_ = _274_ & { entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2], entry_en_t0[2] };
assign _141_ = _278_ & entry_en_t0[1];
assign _144_ = _282_ & { entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1], entry_en_t0[1] };
assign _147_ = _286_ & entry_en_t0[0];
assign _150_ = _290_ & { entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0], entry_en_t0[0] };
assign _153_ = _294_ & { instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0, instr_addr_en_t0 };
assign _271_ = _133_ | _134_;
assign _275_ = _136_ | _137_;
assign _279_ = _139_ | _140_;
assign _283_ = _142_ | _143_;
assign _287_ = _145_ | _146_;
assign _291_ = _148_ | _149_;
assign _295_ = _151_ | _152_;
assign _272_ = _271_ | _135_;
assign _276_ = _275_ | _138_;
assign _280_ = _279_ | _141_;
assign _284_ = _283_ | _144_;
assign _288_ = _287_ | _147_;
assign _292_ = _291_ | _150_;
assign _296_ = _295_ | _153_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q_t0[2] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q_t0[2] <= 1'h0;
else err_q_t0[2] <= _272_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q_t0[95:64] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q_t0[95:64] <= 32'd0;
else rdata_q_t0[95:64] <= _276_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q_t0[1] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q_t0[1] <= 1'h0;
else err_q_t0[1] <= _280_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q_t0[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q_t0[63:32] <= 32'd0;
else rdata_q_t0[63:32] <= _284_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q_t0[0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q_t0[0] <= 1'h0;
else err_q_t0[0] <= _288_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q_t0[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q_t0[31:0] <= 32'd0;
else rdata_q_t0[31:0] <= _292_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME instr_addr_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_addr_q_t0 <= 31'h00000000;
else instr_addr_q_t0 <= _296_;
assign _066_ = err_q_t0[1] & _040_;
assign _069_ = valid_q_t0[0] & err_q[0];
assign _072_ = in_err_i_t0 & _383_;
assign _075_ = err_q_t0[1] & _059_;
assign _078_ = in_err_i_t0 & valid_q[0];
assign _081_ = _011_ & _059_;
assign _084_ = valid_q_t0[0] & in_valid_i;
assign _087_ = _375_ & _378_;
assign _090_ = _377_ & _378_;
assign _093_ = out_ready_i_t0 & out_valid_o;
assign _096_ = _017_ & _387_;
assign _099_ = valid_q_t0[1] & valid_q[0];
assign _102_ = valid_popped_t0[0] & _053_;
assign _105_ = valid_popped_t0[1] & _053_;
assign _108_ = valid_pushed_t0[1] & pop_fifo;
assign _111_ = in_valid_i_t0 & lowest_free_entry[0];
assign _112_ = _019_ & _047_;
assign _115_ = valid_pushed_t0[2] & pop_fifo;
assign _118_ = in_valid_i_t0 & lowest_free_entry[1];
assign _121_ = _021_ & _047_;
assign _124_ = valid_q_t0[2] & valid_q[1];
assign _127_ = valid_popped_t0[2] & _053_;
assign _130_ = in_valid_i_t0 & lowest_free_entry[2];
assign _067_ = unaligned_is_compressed_t0 & err_q[1];
assign _070_ = err_q_t0[0] & valid_q[0];
assign _073_ = _384_ & in_err_i;
assign _076_ = err_q_t0[0] & err_q[1];
assign _079_ = valid_q_t0[0] & in_err_i;
assign _082_ = err_q_t0[0] & _010_;
assign _085_ = in_valid_i_t0 & valid_q[0];
assign _088_ = err_t0 & _374_;
assign _091_ = err_t0 & _376_;
assign _094_ = out_valid_o_t0 & out_ready_i;
assign _097_ = _388_ & _016_;
assign _100_ = valid_q_t0[0] & _045_;
assign _103_ = clear_i_t0 & valid_popped[0];
assign _106_ = clear_i_t0 & valid_popped[1];
assign _109_ = pop_fifo_t0 & valid_pushed[1];
assign _113_ = pop_fifo_t0 & _018_;
assign _116_ = pop_fifo_t0 & valid_pushed[2];
assign _119_ = lowest_free_entry_t0[1] & in_valid_i;
assign _122_ = pop_fifo_t0 & _020_;
assign _125_ = valid_q_t0[1] & _049_;
assign _128_ = clear_i_t0 & valid_popped[2];
assign _131_ = lowest_free_entry_t0[2] & in_valid_i;
assign _068_ = err_q_t0[1] & unaligned_is_compressed_t0;
assign _071_ = valid_q_t0[0] & err_q_t0[0];
assign _074_ = in_err_i_t0 & _384_;
assign _077_ = err_q_t0[1] & err_q_t0[0];
assign _080_ = in_err_i_t0 & valid_q_t0[0];
assign _083_ = _011_ & err_q_t0[0];
assign _086_ = valid_q_t0[0] & in_valid_i_t0;
assign _089_ = _375_ & err_t0;
assign _092_ = _377_ & err_t0;
assign _095_ = out_ready_i_t0 & out_valid_o_t0;
assign _098_ = _017_ & _388_;
assign _101_ = valid_q_t0[1] & valid_q_t0[0];
assign _104_ = valid_popped_t0[0] & clear_i_t0;
assign _107_ = valid_popped_t0[1] & clear_i_t0;
assign _110_ = valid_pushed_t0[1] & pop_fifo_t0;
assign _114_ = _019_ & pop_fifo_t0;
assign _117_ = valid_pushed_t0[2] & pop_fifo_t0;
assign _120_ = in_valid_i_t0 & lowest_free_entry_t0[1];
assign _123_ = _021_ & pop_fifo_t0;
assign _126_ = valid_q_t0[2] & valid_q_t0[1];
assign _129_ = valid_popped_t0[2] & clear_i_t0;
assign _132_ = in_valid_i_t0 & lowest_free_entry_t0[2];
assign _246_ = _066_ | _067_;
assign _247_ = _069_ | _070_;
assign _248_ = _072_ | _073_;
assign _249_ = _075_ | _076_;
assign _250_ = _078_ | _079_;
assign _251_ = _081_ | _082_;
assign _252_ = _084_ | _085_;
assign _253_ = _087_ | _088_;
assign _254_ = _090_ | _091_;
assign _255_ = _093_ | _094_;
assign _256_ = _096_ | _097_;
assign _257_ = _099_ | _100_;
assign _258_ = _102_ | _103_;
assign _259_ = _105_ | _106_;
assign _260_ = _108_ | _109_;
assign _261_ = _111_ | _084_;
assign _262_ = _112_ | _113_;
assign _263_ = _115_ | _116_;
assign _264_ = _118_ | _119_;
assign _265_ = _121_ | _122_;
assign _266_ = _124_ | _125_;
assign _267_ = _127_ | _128_;
assign _268_ = _130_ | _131_;
assign _003_ = _246_ | _068_;
assign _005_ = _247_ | _071_;
assign _007_ = _248_ | _074_;
assign _009_ = _249_ | _077_;
assign _011_ = _250_ | _080_;
assign _013_ = _251_ | _083_;
assign _015_ = _252_ | _086_;
assign unaligned_is_compressed_t0 = _253_ | _089_;
assign aligned_is_compressed_t0 = _254_ | _092_;
assign _017_ = _255_ | _095_;
assign pop_fifo_t0 = _256_ | _098_;
assign lowest_free_entry_t0[1] = _257_ | _101_;
assign valid_d_t0[0] = _258_ | _104_;
assign valid_d_t0[1] = _259_ | _107_;
assign _023_ = _260_ | _110_;
assign _019_ = _261_ | _086_;
assign _025_ = _262_ | _114_;
assign _027_ = _263_ | _117_;
assign _021_ = _264_ | _120_;
assign _029_ = _265_ | _123_;
assign lowest_free_entry_t0[2] = _266_ | _126_;
assign valid_d_t0[2] = _267_ | _129_;
assign entry_en_t0[2] = _268_ | _132_;
assign _036_ = | rdata_t0[17:16];
assign _037_ = | rdata_t0[1:0];
assign _038_ = ~ rdata_t0[17:16];
assign _039_ = ~ rdata_t0[1:0];
assign _154_ = rdata[17:16] & _038_;
assign _155_ = rdata[1:0] & _039_;
assign _370_ = _154_ == _038_;
assign _371_ = _155_ == _039_;
assign _375_ = _370_ & _036_;
assign _377_ = _371_ & _037_;
/* src = "generated/sv2v_out.v:16197.5-16205.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q[2] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q[2] <= 1'h0;
else if (entry_en[2]) err_q[2] <= in_err_i;
/* src = "generated/sv2v_out.v:16197.5-16205.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q[95:64] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q[95:64] <= 32'd0;
else if (entry_en[2]) rdata_q[95:64] <= in_rdata_i;
/* src = "generated/sv2v_out.v:16197.5-16205.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q[1] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q[1] <= 1'h0;
else if (entry_en[1]) err_q[1] <= err_d[1];
/* src = "generated/sv2v_out.v:16197.5-16205.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q[63:32] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q[63:32] <= 32'd0;
else if (entry_en[1]) rdata_q[63:32] <= rdata_d[63:32];
/* src = "generated/sv2v_out.v:16197.5-16205.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME err_q[0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) err_q[0] <= 1'h0;
else if (entry_en[0]) err_q[0] <= err_d[0];
/* src = "generated/sv2v_out.v:16197.5-16205.9" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_q[31:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q[31:0] <= 32'd0;
else if (entry_en[0]) rdata_q[31:0] <= rdata_d[31:0];
/* src = "generated/sv2v_out.v:16149.4-16153.35" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME instr_addr_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) instr_addr_q <= 31'h00000000;
else if (instr_addr_en) instr_addr_q <= instr_addr_d;
assign _040_ = ~ unaligned_is_compressed;
assign _041_ = ~ instr_addr_q[1];
assign _042_ = ~ { instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1] };
assign _043_ = ~ { valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0] };
assign lowest_free_entry[0] = ~ valid_q[0];
assign _044_ = ~ { valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1] };
assign _045_ = ~ valid_q[1];
assign _046_ = ~ { clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i };
assign _047_ = ~ pop_fifo;
assign _048_ = ~ { valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2] };
assign _049_ = ~ valid_q[2];
assign _308_ = unaligned_is_compressed_t0 | _040_;
assign _311_ = instr_addr_q_t0[1] | _041_;
assign _315_ = { instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1] } | _042_;
assign _318_ = { valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0] } | _043_;
assign _321_ = valid_q_t0[0] | lowest_free_entry[0];
assign _324_ = { valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1] } | _044_;
assign _327_ = valid_q_t0[1] | _045_;
assign _332_ = { clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0 } | _046_;
assign _335_ = pop_fifo_t0 | _047_;
assign _340_ = { valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2] } | _048_;
assign _344_ = valid_q_t0[2] | _049_;
assign _309_ = unaligned_is_compressed_t0 | unaligned_is_compressed;
assign _312_ = instr_addr_q_t0[1] | instr_addr_q[1];
assign _316_ = { instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1] } | { instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1], instr_addr_q[1] };
assign _319_ = { valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0] } | { valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0], valid_q[0] };
assign _322_ = valid_q_t0[0] | valid_q[0];
assign _325_ = { valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1] } | { valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1], valid_q[1] };
assign _328_ = valid_q_t0[1] | valid_q[1];
assign _333_ = { clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0 } | { clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i, clear_i };
assign _336_ = pop_fifo_t0 | pop_fifo;
assign _341_ = { valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2] } | { valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2], valid_q[2] };
assign _345_ = valid_q_t0[2] | valid_q[2];
assign _187_ = valid_unaligned_t0 & _308_;
assign _190_ = valid_t0 & _311_;
assign _195_ = err_t0 & _311_;
assign _198_ = rdata_t0 & _315_;
assign _201_ = in_rdata_i_t0 & _318_;
assign _204_ = in_err_i_t0 & _321_;
assign _207_ = { in_rdata_i_t0[15:0], rdata_t0[31:16] } & _324_;
assign _210_ = _386_ & _327_;
assign _213_ = _013_ & _327_;
assign _216_ = _015_ & _327_;
assign _218_ = aligned_is_compressed_t0 & _311_;
assign _221_ = instr_addr_next_t0 & _332_;
assign _224_ = valid_pushed_t0[0] & _335_;
assign _227_ = valid_pushed_t0[1] & _335_;
assign _230_ = in_rdata_i_t0 & _324_;
assign _233_ = in_rdata_i_t0 & _340_;
assign _236_ = in_err_i_t0 & _327_;
assign _239_ = in_err_i_t0 & _344_;
assign _242_ = valid_pushed_t0[2] & _335_;
assign _188_ = valid_t0 & _309_;
assign _191_ = _001_ & _312_;
assign _193_ = err_plus2_t0 & _312_;
assign _196_ = err_unaligned_t0 & _312_;
assign _199_ = rdata_unaligned_t0 & _316_;
assign _202_ = rdata_q_t0[31:0] & _319_;
assign _205_ = err_q_t0[0] & _322_;
assign _208_ = { rdata_q_t0[47:32], rdata_t0[31:16] } & _325_;
assign _211_ = _382_ & _328_;
assign _214_ = _009_ & _328_;
assign _219_ = unaligned_is_compressed_t0 & _312_;
assign _222_ = in_addr_i_t0[31:1] & _333_;
assign _225_ = valid_pushed_t0[1] & _336_;
assign _228_ = valid_pushed_t0[2] & _336_;
assign _231_ = rdata_q_t0[63:32] & _325_;
assign _234_ = rdata_q_t0[95:64] & _341_;
assign _237_ = err_q_t0[1] & _328_;
assign _240_ = err_q_t0[2] & _345_;
assign _310_ = _187_ | _188_;
assign _313_ = _190_ | _191_;
assign _314_ = _195_ | _196_;
assign _317_ = _198_ | _199_;
assign _320_ = _201_ | _202_;
assign _323_ = _204_ | _205_;
assign _326_ = _207_ | _208_;
assign _329_ = _210_ | _211_;
assign _330_ = _213_ | _214_;
assign _331_ = _218_ | _219_;
assign _334_ = _221_ | _222_;
assign _337_ = _224_ | _225_;
assign _338_ = _227_ | _228_;
assign _339_ = _230_ | _231_;
assign _342_ = _233_ | _234_;
assign _343_ = _236_ | _237_;
assign _346_ = _239_ | _240_;
assign _355_ = valid_unaligned ^ valid;
assign _356_ = valid ^ _000_;
assign _357_ = err ^ err_unaligned;
assign _358_ = rdata ^ rdata_unaligned;
assign _359_ = in_rdata_i ^ rdata_q[31:0];
assign _360_ = in_err_i ^ err_q[0];
assign _361_ = { in_rdata_i[15:0], rdata[31:16] } ^ { rdata_q[47:32], rdata[31:16] };
assign _362_ = _385_ ^ _381_;
assign _363_ = _012_ ^ _008_;
assign _364_ = aligned_is_compressed ^ unaligned_is_compressed;
assign _365_ = instr_addr_next ^ in_addr_i[31:1];
assign _366_ = valid_pushed[0] ^ valid_pushed[1];
assign _367_ = valid_pushed[1] ^ valid_pushed[2];
assign _368_ = in_rdata_i ^ rdata_q[63:32];
assign _369_ = in_err_i ^ err_q[1];
assign _189_ = unaligned_is_compressed_t0 & _355_;
assign _192_ = instr_addr_q_t0[1] & _356_;
assign _194_ = instr_addr_q_t0[1] & err_plus2;
assign _197_ = instr_addr_q_t0[1] & _357_;
assign _200_ = { instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1], instr_addr_q_t0[1] } & _358_;
assign _203_ = { valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0], valid_q_t0[0] } & _359_;
assign _206_ = valid_q_t0[0] & _360_;
assign _209_ = { valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1] } & _361_;
assign _212_ = valid_q_t0[1] & _362_;
assign _215_ = valid_q_t0[1] & _363_;
assign _217_ = valid_q_t0[1] & _050_;
assign _220_ = instr_addr_q_t0[1] & _364_;
assign _223_ = { clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0, clear_i_t0 } & _365_;
assign _226_ = pop_fifo_t0 & _366_;
assign _229_ = pop_fifo_t0 & _367_;
assign _232_ = { valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1], valid_q_t0[1] } & _368_;
assign _235_ = { valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2], valid_q_t0[2] } & _349_;
assign _238_ = valid_q_t0[1] & _369_;
assign _241_ = valid_q_t0[2] & _348_;
assign _001_ = _189_ | _310_;
assign out_valid_o_t0 = _192_ | _313_;
assign out_err_plus2_o_t0 = _194_ | _193_;
assign out_err_o_t0 = _197_ | _314_;
assign out_rdata_o_t0 = _200_ | _317_;
assign rdata_t0 = _203_ | _320_;
assign err_t0 = _206_ | _323_;
assign rdata_unaligned_t0 = _209_ | _326_;
assign err_unaligned_t0 = _212_ | _329_;
assign err_plus2_t0 = _215_ | _330_;
assign valid_unaligned_t0 = _217_ | _216_;
assign addr_incr_two_t0 = _220_ | _331_;
assign instr_addr_d_t0 = _223_ | _334_;
assign valid_popped_t0[0] = _226_ | _337_;
assign valid_popped_t0[1] = _229_ | _338_;
assign rdata_d_t0[31:0] = _232_ | _339_;
assign rdata_d_t0[63:32] = _235_ | _342_;
assign err_d_t0[0] = _238_ | _343_;
assign err_d_t0[1] = _241_ | _346_;
assign valid_popped_t0[2] = _116_ | _242_;
assign _050_ = ~ _014_;
assign _051_ = ~ _002_;
assign _052_ = ~ _004_;
assign _053_ = ~ clear_i;
assign _054_ = ~ _018_;
assign _055_ = ~ _020_;
assign _056_ = ~ _022_;
assign _057_ = ~ _026_;
assign _058_ = ~ in_valid_i;
assign _059_ = ~ err_q[0];
assign _060_ = ~ _006_;
assign _061_ = ~ _016_;
assign _062_ = ~ _024_;
assign _063_ = ~ _028_;
assign _156_ = valid_q_t0[0] & _058_;
assign _157_ = _003_ & _059_;
assign _160_ = valid_q_t0[0] & unaligned_is_compressed;
assign _163_ = _005_ & _060_;
assign _166_ = clear_i_t0 & _061_;
assign _169_ = aligned_is_compressed_t0 & _041_;
assign _172_ = _019_ & lowest_free_entry[0];
assign _175_ = _021_ & _045_;
assign _178_ = _023_ & _062_;
assign _181_ = _027_ & _063_;
assign _184_ = valid_q_t0[2] & _032_;
assign _158_ = err_q_t0[0] & _051_;
assign _161_ = unaligned_is_compressed_t0 & valid_q[0];
assign _164_ = _007_ & _052_;
assign _167_ = _017_ & _053_;
assign _170_ = instr_addr_q_t0[1] & aligned_is_compressed;
assign _173_ = valid_q_t0[0] & _054_;
assign _176_ = valid_q_t0[1] & _055_;
assign _179_ = _025_ & _056_;
assign _182_ = _029_ & _057_;
assign _185_ = entry_en_t0[2] & _049_;
assign _159_ = _003_ & err_q_t0[0];
assign _162_ = valid_q_t0[0] & unaligned_is_compressed_t0;
assign _165_ = _005_ & _007_;
assign _168_ = clear_i_t0 & _017_;
assign _171_ = aligned_is_compressed_t0 & instr_addr_q_t0[1];
assign _174_ = _019_ & valid_q_t0[0];
assign _177_ = _021_ & valid_q_t0[1];
assign _180_ = _023_ & _025_;
assign _183_ = _027_ & _029_;
assign _186_ = valid_q_t0[2] & entry_en_t0[2];
assign _297_ = _156_ | _111_;
assign _298_ = _157_ | _158_;
assign _299_ = _160_ | _161_;
assign _300_ = _163_ | _164_;
assign _301_ = _166_ | _167_;
assign _302_ = _169_ | _170_;
assign _303_ = _172_ | _173_;
assign _304_ = _175_ | _176_;
assign _305_ = _178_ | _179_;
assign _306_ = _181_ | _182_;
assign _307_ = _184_ | _185_;
assign valid_t0 = _297_ | _086_;
assign _382_ = _298_ | _159_;
assign _384_ = _299_ | _162_;
assign _386_ = _300_ | _165_;
assign instr_addr_en_t0 = _301_ | _168_;
assign _388_ = _302_ | _171_;
assign valid_pushed_t0[0] = _303_ | _174_;
assign valid_pushed_t0[1] = _304_ | _177_;
assign entry_en_t0[0] = _305_ | _180_;
assign entry_en_t0[1] = _306_ | _183_;
assign valid_pushed_t0[2] = _307_ | _186_;
assign _374_ = rdata[17:16] != /* src = "generated/sv2v_out.v:16125.36-16125.57" */ 2'h3;
assign _376_ = rdata[1:0] != /* src = "generated/sv2v_out.v:16126.34-16126.53" */ 2'h3;
assign _378_ = ~ /* src = "generated/sv2v_out.v:16126.57-16126.61" */ err;
assign _379_ = ~ /* src = "generated/sv2v_out.v:16145.56-16145.70" */ addr_incr_two;
assign _380_ = ~ /* src = "generated/sv2v_out.v:16164.51-16164.73" */ aligned_is_compressed;
assign valid = valid_q[0] | /* src = "generated/sv2v_out.v:16120.17-16120.40" */ in_valid_i;
assign _381_ = _002_ | /* src = "generated/sv2v_out.v:16122.39-16122.87" */ err_q[0];
assign _383_ = lowest_free_entry[0] | /* src = "generated/sv2v_out.v:16122.129-16122.167" */ _040_;
assign _385_ = _004_ | /* src = "generated/sv2v_out.v:16122.90-16122.169" */ _006_;
assign instr_addr_en = clear_i | /* src = "generated/sv2v_out.v:16143.25-16143.62" */ _016_;
assign _387_ = _380_ | /* src = "generated/sv2v_out.v:16164.51-16164.89" */ instr_addr_q[1];
assign valid_pushed[0] = _018_ | /* src = "generated/sv2v_out.v:16174.29-16174.77" */ valid_q[0];
assign valid_pushed[1] = _020_ | /* src = "generated/sv2v_out.v:16174.29-16174.77" */ valid_q[1];
assign entry_en[0] = _022_ | /* src = "generated/sv2v_out.v:16177.25-16177.109" */ _024_;
assign entry_en[1] = _026_ | /* src = "generated/sv2v_out.v:16177.25-16177.109" */ _028_;
assign valid_pushed[2] = valid_q[2] | /* src = "generated/sv2v_out.v:16183.35-16183.99" */ entry_en[2];
/* src = "generated/sv2v_out.v:16189.2-16193.23" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME valid_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) valid_q <= 3'h0;
else valid_q <= valid_d;
assign _000_ = unaligned_is_compressed ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:16132.8-16132.31|generated/sv2v_out.v:16132.4-16135.35" */ valid : valid_unaligned;
assign out_valid_o = instr_addr_q[1] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:16128.7-16128.20|generated/sv2v_out.v:16128.3-16142.6" */ _000_ : valid;
assign out_err_plus2_o = instr_addr_q[1] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:16128.7-16128.20|generated/sv2v_out.v:16128.3-16142.6" */ err_plus2 : 1'h0;
assign out_err_o = instr_addr_q[1] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:16128.7-16128.20|generated/sv2v_out.v:16128.3-16142.6" */ err_unaligned : err;
assign out_rdata_o = instr_addr_q[1] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:16128.7-16128.20|generated/sv2v_out.v:16128.3-16142.6" */ rdata_unaligned : rdata;
assign rdata = valid_q[0] ? /* src = "generated/sv2v_out.v:16118.18-16118.58" */ rdata_q[31:0] : in_rdata_i;
assign err = valid_q[0] ? /* src = "generated/sv2v_out.v:16119.16-16119.48" */ err_q[0] : in_err_i;
assign rdata_unaligned = valid_q[1] ? /* src = "generated/sv2v_out.v:16121.28-16121.107" */ { rdata_q[47:32], rdata[31:16] } : { in_rdata_i[15:0], rdata[31:16] };
assign err_unaligned = valid_q[1] ? /* src = "generated/sv2v_out.v:16122.26-16122.169" */ _381_ : _385_;
assign err_plus2 = valid_q[1] ? /* src = "generated/sv2v_out.v:16123.22-16123.93" */ _008_ : _012_;
assign valid_unaligned = valid_q[1] ? /* src = "generated/sv2v_out.v:16124.28-16124.71" */ 1'h1 : _014_;
assign addr_incr_two = instr_addr_q[1] ? /* src = "generated/sv2v_out.v:16144.26-16144.91" */ unaligned_is_compressed : aligned_is_compressed;
assign instr_addr_d = clear_i ? /* src = "generated/sv2v_out.v:16146.25-16146.68" */ in_addr_i[31:1] : instr_addr_next;
assign valid_popped[0] = pop_fifo ? /* src = "generated/sv2v_out.v:16175.30-16175.78" */ valid_pushed[1] : valid_pushed[0];
assign valid_popped[1] = pop_fifo ? /* src = "generated/sv2v_out.v:16175.30-16175.78" */ valid_pushed[2] : valid_pushed[1];
assign rdata_d[31:0] = valid_q[1] ? /* src = "generated/sv2v_out.v:16178.34-16178.89" */ rdata_q[63:32] : in_rdata_i;
assign rdata_d[63:32] = valid_q[2] ? /* src = "generated/sv2v_out.v:16178.34-16178.89" */ rdata_q[95:64] : in_rdata_i;
assign err_d[0] = valid_q[1] ? /* src = "generated/sv2v_out.v:16179.23-16179.63" */ err_q[1] : in_err_i;
assign err_d[1] = valid_q[2] ? /* src = "generated/sv2v_out.v:16179.23-16179.63" */ err_q[2] : in_err_i;
assign valid_popped[2] = pop_fifo ? /* src = "generated/sv2v_out.v:16184.36-16184.77" */ 1'h0 : valid_pushed[2];
assign busy_o = valid_q[2:1];
assign busy_o_t0 = valid_q_t0[2:1];
assign err_d[2] = in_err_i;
assign err_d_t0[2] = in_err_i_t0;
assign lowest_free_entry_t0[0] = valid_q_t0[0];
assign out_addr_o = { instr_addr_q, 1'h0 };
assign out_addr_o_t0 = { instr_addr_q_t0, 1'h0 };
assign rdata_d[95:64] = in_rdata_i;
assign rdata_d_t0[95:64] = in_rdata_i_t0;
endmodule

module \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111 (clk_i, rst_ni, data_req_o, data_gnt_i, data_rvalid_i, data_bus_err_i, data_pmp_err_i, data_addr_o, data_we_o, data_be_o, data_wdata_o, data_rdata_i, lsu_we_i, lsu_type_i, lsu_wdata_i, lsu_sign_ext_i, lsu_rdata_o, lsu_rdata_valid_o, lsu_req_i, adder_result_ex_i, addr_incr_req_o
, addr_last_o, lsu_req_done_o, lsu_resp_valid_o, load_err_o, load_resp_intg_err_o, store_err_o, store_resp_intg_err_o, busy_o, perf_load_o, perf_store_o, data_we_o_t0, data_req_o_t0, busy_o_t0, adder_result_ex_i_t0, addr_incr_req_o_t0, addr_last_o_t0, data_addr_o_t0, data_be_o_t0, data_bus_err_i_t0, data_gnt_i_t0, data_pmp_err_i_t0
, data_rdata_i_t0, data_rvalid_i_t0, data_wdata_o_t0, load_err_o_t0, load_resp_intg_err_o_t0, lsu_rdata_o_t0, lsu_rdata_valid_o_t0, lsu_req_done_o_t0, lsu_req_i_t0, lsu_resp_valid_o_t0, lsu_sign_ext_i_t0, lsu_type_i_t0, lsu_wdata_i_t0, lsu_we_i_t0, perf_load_o_t0, perf_store_o_t0, store_err_o_t0, store_resp_intg_err_o_t0);
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0001_;
/* src = "generated/sv2v_out.v:18407.2-18446.10" */
wire [3:0] _0002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18407.2-18446.10" */
wire [3:0] _0003_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0004_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0005_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0006_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire [2:0] _0007_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire [2:0] _0008_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0009_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0011_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0013_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0015_;
/* src = "generated/sv2v_out.v:18511.2-18534.10" */
wire [31:0] _0016_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18511.2-18534.10" */
wire [31:0] _0017_;
/* src = "generated/sv2v_out.v:18487.2-18510.10" */
wire [31:0] _0018_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18487.2-18510.10" */
wire [31:0] _0019_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0021_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0022_;
/* src = "generated/sv2v_out.v:18407.2-18446.10" */
wire [3:0] _0023_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18407.2-18446.10" */
wire [3:0] _0024_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0025_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0026_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire [2:0] _0027_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire [2:0] _0028_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0029_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0030_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0031_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0032_;
/* src = "generated/sv2v_out.v:18511.2-18534.10" */
wire [31:0] _0033_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18511.2-18534.10" */
wire [31:0] _0034_;
/* src = "generated/sv2v_out.v:18487.2-18510.10" */
wire [31:0] _0035_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18487.2-18510.10" */
wire [31:0] _0036_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0037_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0038_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0039_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0040_;
/* src = "generated/sv2v_out.v:18407.2-18446.10" */
wire [3:0] _0041_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18407.2-18446.10" */
wire [3:0] _0042_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0043_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire [2:0] _0044_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire [2:0] _0045_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0046_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0047_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0048_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0049_;
/* src = "generated/sv2v_out.v:18511.2-18534.10" */
wire [31:0] _0050_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18511.2-18534.10" */
wire [31:0] _0051_;
/* src = "generated/sv2v_out.v:18487.2-18510.10" */
wire [31:0] _0052_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18487.2-18510.10" */
wire [31:0] _0053_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0054_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0055_;
/* src = "generated/sv2v_out.v:18407.2-18446.10" */
wire [3:0] _0056_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18407.2-18446.10" */
wire [3:0] _0057_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0058_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0059_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire [2:0] _0060_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire [2:0] _0061_;
/* src = "generated/sv2v_out.v:18511.2-18534.10" */
wire [31:0] _0062_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18511.2-18534.10" */
wire [31:0] _0063_;
/* src = "generated/sv2v_out.v:18487.2-18510.10" */
wire [31:0] _0064_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18487.2-18510.10" */
wire [31:0] _0065_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0066_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0067_;
/* src = "generated/sv2v_out.v:18407.2-18446.10" */
wire [3:0] _0068_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18407.2-18446.10" */
wire [3:0] _0069_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0070_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire [2:0] _0071_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire [2:0] _0072_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0073_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0074_;
/* src = "generated/sv2v_out.v:18407.2-18446.10" */
wire [3:0] _0075_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18407.2-18446.10" */
wire [3:0] _0076_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire _0077_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire [2:0] _0078_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire [2:0] _0079_;
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire [2:0] _0080_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18561.2-18639.5" */
wire [2:0] _0081_;
/* src = "generated/sv2v_out.v:18609.20-18609.62" */
wire _0082_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18609.20-18609.62" */
wire _0083_;
/* src = "generated/sv2v_out.v:18656.32-18656.67" */
wire _0084_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18656.32-18656.67" */
wire _0085_;
/* src = "generated/sv2v_out.v:18656.31-18656.87" */
wire _0086_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18656.31-18656.87" */
wire _0087_;
/* src = "generated/sv2v_out.v:18656.30-18656.101" */
wire _0088_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18656.30-18656.101" */
wire _0089_;
/* src = "generated/sv2v_out.v:18674.23-18674.51" */
wire _0090_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18674.23-18674.51" */
wire _0091_;
/* src = "generated/sv2v_out.v:18675.24-18675.51" */
wire _0092_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18675.24-18675.51" */
wire _0093_;
/* src = "generated/sv2v_out.v:18676.33-18676.62" */
wire _0094_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18676.33-18676.62" */
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire _0109_;
wire _0110_;
wire _0111_;
wire _0112_;
wire _0113_;
wire [2:0] _0114_;
wire [2:0] _0115_;
wire [1:0] _0116_;
wire [1:0] _0117_;
wire [1:0] _0118_;
wire [1:0] _0119_;
wire [1:0] _0120_;
wire [2:0] _0121_;
wire [1:0] _0122_;
wire [1:0] _0123_;
wire [1:0] _0124_;
wire [1:0] _0125_;
wire _0126_;
wire _0127_;
wire _0128_;
wire _0129_;
wire _0130_;
wire _0131_;
wire _0132_;
wire _0133_;
wire _0134_;
wire _0135_;
wire [3:0] _0136_;
wire [2:0] _0137_;
wire [2:0] _0138_;
wire [1:0] _0139_;
wire [1:0] _0140_;
wire [2:0] _0141_;
wire [2:0] _0142_;
wire [1:0] _0143_;
wire [1:0] _0144_;
wire [1:0] _0145_;
wire _0146_;
wire _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
wire _0152_;
wire _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire [2:0] _0164_;
wire [2:0] _0165_;
wire [2:0] _0166_;
wire [2:0] _0167_;
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire [31:0] _0177_;
wire [31:0] _0178_;
wire [31:0] _0179_;
wire [31:0] _0180_;
wire [31:0] _0181_;
wire [31:0] _0182_;
wire [31:0] _0183_;
wire [31:0] _0184_;
wire [3:0] _0185_;
wire [3:0] _0186_;
wire [3:0] _0187_;
wire [2:0] _0188_;
wire [2:0] _0189_;
wire [2:0] _0190_;
wire [2:0] _0191_;
wire [2:0] _0192_;
wire _0193_;
wire [31:0] _0194_;
wire [3:0] _0195_;
wire [31:0] _0196_;
wire _0197_;
wire _0198_;
wire _0199_;
wire _0200_;
wire _0201_;
wire _0202_;
wire _0203_;
wire _0204_;
wire _0205_;
wire _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
/* cellift = 32'd1 */
wire _0211_;
wire _0212_;
/* cellift = 32'd1 */
wire _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
/* cellift = 32'd1 */
wire _0221_;
wire _0222_;
/* cellift = 32'd1 */
wire _0223_;
wire _0224_;
/* cellift = 32'd1 */
wire _0225_;
wire _0226_;
/* cellift = 32'd1 */
wire _0227_;
wire _0228_;
/* cellift = 32'd1 */
wire _0229_;
wire _0230_;
/* cellift = 32'd1 */
wire _0231_;
wire _0232_;
/* cellift = 32'd1 */
wire _0233_;
wire _0234_;
/* cellift = 32'd1 */
wire _0235_;
wire _0236_;
/* cellift = 32'd1 */
wire _0237_;
wire _0238_;
/* cellift = 32'd1 */
wire _0239_;
wire _0240_;
/* cellift = 32'd1 */
wire _0241_;
wire _0242_;
/* cellift = 32'd1 */
wire _0243_;
wire _0244_;
/* cellift = 32'd1 */
wire _0245_;
wire _0246_;
/* cellift = 32'd1 */
wire _0247_;
wire _0248_;
wire _0249_;
wire _0250_;
wire _0251_;
wire _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire _0259_;
wire _0260_;
wire _0261_;
wire _0262_;
wire _0263_;
wire _0264_;
wire _0265_;
wire _0266_;
wire _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire _0271_;
wire _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire _0276_;
wire _0277_;
wire _0278_;
wire _0279_;
wire _0280_;
wire _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire _0285_;
wire _0286_;
wire _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire _0294_;
wire _0295_;
wire _0296_;
wire _0297_;
wire [23:0] _0298_;
wire [23:0] _0299_;
wire [23:0] _0300_;
wire [31:0] _0301_;
wire [31:0] _0302_;
wire [31:0] _0303_;
wire [1:0] _0304_;
wire [1:0] _0305_;
wire [1:0] _0306_;
wire [1:0] _0307_;
wire [1:0] _0308_;
wire [1:0] _0309_;
wire _0310_;
wire _0311_;
wire _0312_;
wire [2:0] _0313_;
wire [2:0] _0314_;
wire [1:0] _0315_;
wire [1:0] _0316_;
wire [1:0] _0317_;
wire [3:0] _0318_;
wire [1:0] _0319_;
wire [1:0] _0320_;
wire [2:0] _0321_;
wire [2:0] _0322_;
wire [1:0] _0323_;
wire [1:0] _0324_;
wire [2:0] _0325_;
wire _0326_;
wire _0327_;
wire _0328_;
wire _0329_;
wire _0330_;
wire _0331_;
wire _0332_;
wire _0333_;
wire _0334_;
wire [2:0] _0335_;
wire [2:0] _0336_;
wire [2:0] _0337_;
wire [2:0] _0338_;
wire [2:0] _0339_;
wire [2:0] _0340_;
wire [2:0] _0341_;
wire [2:0] _0342_;
wire [2:0] _0343_;
wire [2:0] _0344_;
wire [2:0] _0345_;
wire [2:0] _0346_;
wire [2:0] _0347_;
wire [2:0] _0348_;
wire _0349_;
wire _0350_;
wire _0351_;
wire _0352_;
wire _0353_;
wire _0354_;
wire _0355_;
wire _0356_;
wire _0357_;
wire _0358_;
wire _0359_;
wire _0360_;
wire _0361_;
wire _0362_;
wire _0363_;
wire _0364_;
wire _0365_;
wire _0366_;
wire _0367_;
wire _0368_;
wire _0369_;
wire _0370_;
wire _0371_;
wire _0372_;
wire _0373_;
wire _0374_;
wire _0375_;
wire _0376_;
wire _0377_;
wire _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire _0382_;
wire _0383_;
wire _0384_;
wire _0385_;
wire _0386_;
wire _0387_;
wire _0388_;
wire _0389_;
wire _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire [31:0] _0397_;
wire [31:0] _0398_;
wire [31:0] _0399_;
wire [31:0] _0400_;
wire [31:0] _0401_;
wire [31:0] _0402_;
wire [31:0] _0403_;
wire [31:0] _0404_;
wire [31:0] _0405_;
wire [31:0] _0406_;
wire [31:0] _0407_;
wire [31:0] _0408_;
wire [31:0] _0409_;
wire [31:0] _0410_;
wire [31:0] _0411_;
wire [31:0] _0412_;
wire [31:0] _0413_;
wire [31:0] _0414_;
wire [31:0] _0415_;
wire [31:0] _0416_;
wire [31:0] _0417_;
wire [31:0] _0418_;
wire [31:0] _0419_;
wire [31:0] _0420_;
wire [31:0] _0421_;
wire [31:0] _0422_;
wire [31:0] _0423_;
wire [31:0] _0424_;
wire [31:0] _0425_;
wire [31:0] _0426_;
wire [31:0] _0427_;
wire [31:0] _0428_;
wire [31:0] _0429_;
wire [31:0] _0430_;
wire [31:0] _0431_;
wire [31:0] _0432_;
wire [31:0] _0433_;
wire [31:0] _0434_;
wire [31:0] _0435_;
wire [31:0] _0436_;
wire [31:0] _0437_;
wire [31:0] _0438_;
wire [3:0] _0439_;
wire [3:0] _0440_;
wire [3:0] _0441_;
wire [3:0] _0442_;
wire [3:0] _0443_;
wire [3:0] _0444_;
wire [3:0] _0445_;
wire [3:0] _0446_;
wire [3:0] _0447_;
wire [3:0] _0448_;
wire [3:0] _0449_;
wire [3:0] _0450_;
wire [3:0] _0451_;
wire [3:0] _0452_;
wire [3:0] _0453_;
wire [2:0] _0454_;
wire _0455_;
wire _0456_;
wire _0457_;
wire _0458_;
wire _0459_;
wire _0460_;
wire _0461_;
wire _0462_;
wire _0463_;
wire _0464_;
wire _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire _0469_;
wire [1:0] _0470_;
wire [2:0] _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire _0477_;
wire _0478_;
wire _0479_;
wire _0480_;
wire _0481_;
wire _0482_;
wire _0483_;
wire [2:0] _0484_;
wire [2:0] _0485_;
wire _0486_;
wire _0487_;
wire _0488_;
wire [2:0] _0489_;
wire [2:0] _0490_;
wire _0491_;
wire _0492_;
wire [2:0] _0493_;
wire [2:0] _0494_;
wire _0495_;
wire _0496_;
wire _0497_;
wire _0498_;
wire [2:0] _0499_;
wire [2:0] _0500_;
wire [2:0] _0501_;
wire _0502_;
wire _0503_;
wire [2:0] _0504_;
wire [2:0] _0505_;
wire [2:0] _0506_;
wire [2:0] _0507_;
wire [2:0] _0508_;
wire [2:0] _0509_;
wire [2:0] _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0517_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire [1:0] _0522_;
wire [1:0] _0523_;
wire [31:0] _0524_;
wire [31:0] _0525_;
wire [31:0] _0526_;
wire [31:0] _0527_;
wire [31:0] _0528_;
wire [31:0] _0529_;
wire [31:0] _0530_;
wire [31:0] _0531_;
wire [31:0] _0532_;
wire [31:0] _0533_;
wire [31:0] _0534_;
wire [31:0] _0535_;
wire [31:0] _0536_;
wire [31:0] _0537_;
wire [31:0] _0538_;
wire [31:0] _0539_;
wire [31:0] _0540_;
wire [31:0] _0541_;
wire [31:0] _0542_;
wire [31:0] _0543_;
wire [31:0] _0544_;
wire [31:0] _0545_;
wire [31:0] _0546_;
wire [31:0] _0547_;
wire [1:0] _0548_;
wire [1:0] _0549_;
wire [3:0] _0550_;
wire [3:0] _0551_;
wire [3:0] _0552_;
wire [3:0] _0553_;
wire [3:0] _0554_;
wire [1:0] _0555_;
wire [1:0] _0556_;
wire [31:0] _0557_;
wire [31:0] _0558_;
wire [31:0] _0559_;
wire _0560_;
/* cellift = 32'd1 */
wire _0561_;
wire _0562_;
/* cellift = 32'd1 */
wire _0563_;
wire _0564_;
/* cellift = 32'd1 */
wire _0565_;
wire _0566_;
wire _0567_;
wire _0568_;
wire _0569_;
wire _0570_;
wire _0571_;
wire _0572_;
wire _0573_;
wire _0574_;
wire _0575_;
wire _0576_;
wire _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire [23:0] _0596_;
wire [23:0] _0597_;
wire [23:0] _0598_;
wire [23:0] _0599_;
wire [31:0] _0600_;
wire [31:0] _0601_;
wire [31:0] _0602_;
wire [31:0] _0603_;
wire [1:0] _0604_;
wire [1:0] _0605_;
wire [1:0] _0606_;
wire [1:0] _0607_;
wire [1:0] _0608_;
wire [1:0] _0609_;
wire [1:0] _0610_;
wire [1:0] _0611_;
wire _0612_;
wire _0613_;
wire _0614_;
wire _0615_;
wire [5:0] _0616_;
wire [2:0] _0617_;
wire [3:0] _0618_;
wire _0619_;
wire _0620_;
wire _0621_;
wire [2:0] _0622_;
wire [2:0] _0623_;
wire [2:0] _0624_;
wire [2:0] _0625_;
wire [2:0] _0626_;
wire [2:0] _0627_;
wire [2:0] _0628_;
wire [2:0] _0629_;
wire [2:0] _0630_;
wire [2:0] _0631_;
wire [2:0] _0632_;
wire [2:0] _0633_;
wire [2:0] _0634_;
wire _0635_;
wire _0636_;
wire _0637_;
wire _0638_;
wire _0639_;
wire _0640_;
wire _0641_;
wire _0642_;
wire _0643_;
wire _0644_;
wire _0645_;
wire _0646_;
wire _0647_;
wire _0648_;
wire _0649_;
wire _0650_;
wire _0651_;
wire _0652_;
wire _0653_;
wire _0654_;
wire _0655_;
wire _0656_;
wire _0657_;
wire _0658_;
wire _0659_;
wire _0660_;
wire _0661_;
wire [31:0] _0662_;
wire [31:0] _0663_;
wire [31:0] _0664_;
wire [31:0] _0665_;
wire [31:0] _0666_;
wire [31:0] _0667_;
wire [31:0] _0668_;
wire [31:0] _0669_;
wire [31:0] _0670_;
wire [31:0] _0671_;
wire [31:0] _0672_;
wire [31:0] _0673_;
wire [31:0] _0674_;
wire [31:0] _0675_;
wire [31:0] _0676_;
wire [31:0] _0677_;
wire [31:0] _0678_;
wire [31:0] _0679_;
wire [31:0] _0680_;
wire [31:0] _0681_;
wire [31:0] _0682_;
wire [31:0] _0683_;
wire [31:0] _0684_;
wire [31:0] _0685_;
wire [31:0] _0686_;
wire [31:0] _0687_;
wire [31:0] _0688_;
wire [31:0] _0689_;
wire [31:0] _0690_;
wire [31:0] _0691_;
wire [3:0] _0692_;
wire [3:0] _0693_;
wire [3:0] _0694_;
wire [3:0] _0695_;
wire [3:0] _0696_;
wire [3:0] _0697_;
wire [3:0] _0698_;
wire [3:0] _0699_;
wire [3:0] _0700_;
wire [3:0] _0701_;
wire [3:0] _0702_;
wire _0703_;
wire _0704_;
wire _0705_;
wire _0706_;
wire _0707_;
wire _0708_;
wire _0709_;
wire _0710_;
wire _0711_;
wire [2:0] _0712_;
wire _0713_;
wire _0714_;
wire [2:0] _0715_;
wire _0716_;
wire [2:0] _0717_;
wire [2:0] _0718_;
wire _0719_;
wire [2:0] _0720_;
wire [2:0] _0721_;
wire [2:0] _0722_;
wire [2:0] _0723_;
wire [2:0] _0724_;
wire [2:0] _0725_;
wire [2:0] _0726_;
wire _0727_;
wire [31:0] _0728_;
wire [31:0] _0729_;
wire [31:0] _0730_;
wire [31:0] _0731_;
wire [31:0] _0732_;
wire [31:0] _0733_;
wire [31:0] _0734_;
wire [31:0] _0735_;
wire [31:0] _0736_;
wire [31:0] _0737_;
wire [3:0] _0738_;
wire [3:0] _0739_;
wire [3:0] _0740_;
wire [31:0] _0741_;
wire [31:0] _0742_;
wire [31:0] _0743_;
wire _0744_;
wire _0745_;
wire _0746_;
wire _0747_;
wire [23:0] _0748_;
wire [31:0] _0749_;
wire [1:0] _0750_;
wire [1:0] _0751_;
wire _0752_;
wire [2:0] _0753_;
wire [2:0] _0754_;
wire [2:0] _0755_;
wire [2:0] _0756_;
wire _0757_;
wire _0758_;
wire _0759_;
wire _0760_;
wire _0761_;
wire _0762_;
wire _0763_;
wire _0764_;
wire _0765_;
wire _0766_;
wire _0767_;
wire _0768_;
wire [31:0] _0769_;
wire [31:0] _0770_;
wire [31:0] _0771_;
wire [31:0] _0772_;
wire [31:0] _0773_;
wire [31:0] _0774_;
wire [31:0] _0775_;
wire [31:0] _0776_;
wire [31:0] _0777_;
wire [31:0] _0778_;
wire [31:0] _0779_;
wire [31:0] _0780_;
wire [31:0] _0781_;
wire [31:0] _0782_;
wire [3:0] _0783_;
wire [3:0] _0784_;
wire [3:0] _0785_;
wire [3:0] _0786_;
wire [3:0] _0787_;
wire [3:0] _0788_;
wire _0789_;
wire _0790_;
wire [2:0] _0791_;
wire [2:0] _0792_;
wire [2:0] _0793_;
wire _0794_;
wire [31:0] _0795_;
wire [31:0] _0796_;
wire [31:0] _0797_;
wire [31:0] _0798_;
wire [31:0] _0799_;
wire [31:0] _0800_;
wire [31:0] _0801_;
wire [31:0] _0802_;
wire [3:0] _0803_;
wire [31:0] _0804_;
wire _0805_;
wire _0806_;
wire _0807_;
wire _0808_;
wire _0809_;
wire _0810_;
wire _0811_;
wire _0812_;
wire _0813_;
wire _0814_;
wire _0815_;
wire _0816_;
wire _0817_;
wire _0818_;
wire _0819_;
wire _0820_;
wire _0821_;
wire _0822_;
wire _0823_;
wire _0824_;
wire _0825_;
wire _0826_;
wire _0827_;
wire [2:0] _0828_;
/* cellift = 32'd1 */
wire [2:0] _0829_;
wire [2:0] _0830_;
/* cellift = 32'd1 */
wire [2:0] _0831_;
wire [2:0] _0832_;
/* cellift = 32'd1 */
wire [2:0] _0833_;
wire [2:0] _0834_;
/* cellift = 32'd1 */
wire [2:0] _0835_;
wire _0836_;
/* cellift = 32'd1 */
wire _0837_;
wire _0838_;
/* cellift = 32'd1 */
wire _0839_;
wire _0840_;
/* cellift = 32'd1 */
wire _0841_;
wire _0842_;
/* cellift = 32'd1 */
wire _0843_;
wire _0844_;
/* cellift = 32'd1 */
wire _0845_;
wire _0846_;
/* cellift = 32'd1 */
wire _0847_;
wire _0848_;
/* cellift = 32'd1 */
wire _0849_;
wire _0850_;
/* cellift = 32'd1 */
wire _0851_;
wire _0852_;
/* cellift = 32'd1 */
wire _0853_;
wire _0854_;
/* cellift = 32'd1 */
wire _0855_;
wire _0856_;
/* cellift = 32'd1 */
wire _0857_;
wire [31:0] _0858_;
/* cellift = 32'd1 */
wire [31:0] _0859_;
wire [31:0] _0860_;
/* cellift = 32'd1 */
wire [31:0] _0861_;
wire [31:0] _0862_;
/* cellift = 32'd1 */
wire [31:0] _0863_;
wire [31:0] _0864_;
/* cellift = 32'd1 */
wire [31:0] _0865_;
wire [31:0] _0866_;
/* cellift = 32'd1 */
wire [31:0] _0867_;
wire [31:0] _0868_;
/* cellift = 32'd1 */
wire [31:0] _0869_;
wire [31:0] _0870_;
/* cellift = 32'd1 */
wire [31:0] _0871_;
wire [31:0] _0872_;
/* cellift = 32'd1 */
wire [31:0] _0873_;
wire [31:0] _0874_;
/* cellift = 32'd1 */
wire [31:0] _0875_;
wire [3:0] _0876_;
/* cellift = 32'd1 */
wire [3:0] _0877_;
wire [3:0] _0878_;
/* cellift = 32'd1 */
wire [3:0] _0879_;
wire [3:0] _0880_;
wire [3:0] _0881_;
wire [3:0] _0882_;
wire [3:0] _0883_;
wire [3:0] _0884_;
wire [3:0] _0885_;
/* cellift = 32'd1 */
wire [3:0] _0886_;
/* src = "generated/sv2v_out.v:18560.37-18560.56" */
wire _0887_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18560.37-18560.56" */
wire _0888_;
/* src = "generated/sv2v_out.v:18560.90-18560.109" */
wire _0889_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18560.90-18560.109" */
wire _0890_;
/* src = "generated/sv2v_out.v:18560.115-18560.135" */
wire _0891_;
/* src = "generated/sv2v_out.v:18640.63-18640.80" */
wire _0892_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18640.63-18640.80" */
wire _0893_;
/* src = "generated/sv2v_out.v:18655.59-18655.76" */
wire _0894_;
/* src = "generated/sv2v_out.v:18560.36-18560.83" */
wire _0895_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18560.36-18560.83" */
wire _0896_;
/* src = "generated/sv2v_out.v:18560.89-18560.136" */
wire _0897_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18560.89-18560.136" */
wire _0898_;
/* src = "generated/sv2v_out.v:18594.9-18594.32" */
wire _0899_;
/* src = "generated/sv2v_out.v:18604.9-18604.35" */
wire _0900_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18604.9-18604.35" */
wire _0901_;
/* src = "generated/sv2v_out.v:18560.62-18560.82" */
wire _0902_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18560.62-18560.82" */
wire _0903_;
/* src = "generated/sv2v_out.v:18609.33-18609.62" */
wire _0904_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18609.33-18609.62" */
wire _0905_;
/* src = "generated/sv2v_out.v:18656.71-18656.87" */
wire _0906_;
/* src = "generated/sv2v_out.v:18656.105-18656.119" */
wire _0907_;
/* src = "generated/sv2v_out.v:18606.18-18606.44" */
wire _0908_;
/* src = "generated/sv2v_out.v:18640.27-18640.58" */
wire _0909_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18640.27-18640.58" */
wire _0910_;
/* src = "generated/sv2v_out.v:18654.28-18654.54" */
wire _0911_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18654.28-18654.54" */
wire _0912_;
/* src = "generated/sv2v_out.v:18655.29-18655.54" */
wire _0913_;
wire _0914_;
/* cellift = 32'd1 */
wire _0915_;
wire _0916_;
/* cellift = 32'd1 */
wire _0917_;
wire _0918_;
/* cellift = 32'd1 */
wire _0919_;
wire _0920_;
/* cellift = 32'd1 */
wire _0921_;
wire [1:0] _0922_;
/* cellift = 32'd1 */
wire [1:0] _0923_;
wire _0924_;
/* cellift = 32'd1 */
wire _0925_;
wire _0926_;
/* cellift = 32'd1 */
wire _0927_;
wire _0928_;
/* cellift = 32'd1 */
wire _0929_;
wire _0930_;
/* cellift = 32'd1 */
wire _0931_;
wire _0932_;
/* cellift = 32'd1 */
wire _0933_;
wire _0934_;
/* cellift = 32'd1 */
wire _0935_;
wire _0936_;
wire [1:0] _0937_;
/* cellift = 32'd1 */
wire [1:0] _0938_;
wire _0939_;
/* cellift = 32'd1 */
wire _0940_;
/* src = "generated/sv2v_out.v:18586.20-18586.57" */
wire [2:0] _0941_;
/* src = "generated/sv2v_out.v:18589.20-18589.57" */
wire [2:0] _0942_;
/* src = "generated/sv2v_out.v:18608.19-18608.43" */
wire [2:0] _0943_;
/* src = "generated/sv2v_out.v:18363.20-18363.37" */
input [31:0] adder_result_ex_i;
wire [31:0] adder_result_ex_i;
/* cellift = 32'd1 */
input [31:0] adder_result_ex_i_t0;
wire [31:0] adder_result_ex_i_t0;
/* src = "generated/sv2v_out.v:18364.13-18364.28" */
output addr_incr_req_o;
wire addr_incr_req_o;
/* cellift = 32'd1 */
output addr_incr_req_o_t0;
wire addr_incr_req_o_t0;
/* src = "generated/sv2v_out.v:18378.14-18378.25" */
wire [31:0] addr_last_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18378.14-18378.25" */
wire [31:0] addr_last_d_t0;
/* src = "generated/sv2v_out.v:18365.21-18365.32" */
output [31:0] addr_last_o;
reg [31:0] addr_last_o;
/* cellift = 32'd1 */
output [31:0] addr_last_o_t0;
reg [31:0] addr_last_o_t0;
/* src = "generated/sv2v_out.v:18379.6-18379.17" */
wire addr_update;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18379.6-18379.17" */
wire addr_update_t0;
/* src = "generated/sv2v_out.v:18372.14-18372.20" */
output busy_o;
wire busy_o;
/* cellift = 32'd1 */
output busy_o_t0;
wire busy_o_t0;
/* src = "generated/sv2v_out.v:18344.13-18344.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:18380.6-18380.17" */
wire ctrl_update;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18380.6-18380.17" */
wire ctrl_update_t0;
/* src = "generated/sv2v_out.v:18351.21-18351.32" */
output [31:0] data_addr_o;
wire [31:0] data_addr_o;
/* cellift = 32'd1 */
output [31:0] data_addr_o_t0;
wire [31:0] data_addr_o_t0;
/* src = "generated/sv2v_out.v:18353.20-18353.29" */
output [3:0] data_be_o;
wire [3:0] data_be_o;
/* cellift = 32'd1 */
output [3:0] data_be_o_t0;
wire [3:0] data_be_o_t0;
/* src = "generated/sv2v_out.v:18349.13-18349.27" */
input data_bus_err_i;
wire data_bus_err_i;
/* cellift = 32'd1 */
input data_bus_err_i_t0;
wire data_bus_err_i_t0;
/* src = "generated/sv2v_out.v:18347.13-18347.23" */
input data_gnt_i;
wire data_gnt_i;
/* cellift = 32'd1 */
input data_gnt_i_t0;
wire data_gnt_i_t0;
/* src = "generated/sv2v_out.v:18401.7-18401.20" */
wire data_intg_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18401.7-18401.20" */
wire data_intg_err_t0;
/* src = "generated/sv2v_out.v:18402.7-18402.22" */
wire data_or_pmp_err;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18402.7-18402.22" */
wire data_or_pmp_err_t0;
/* src = "generated/sv2v_out.v:18350.13-18350.27" */
input data_pmp_err_i;
wire data_pmp_err_i;
/* cellift = 32'd1 */
input data_pmp_err_i_t0;
wire data_pmp_err_i_t0;
/* src = "generated/sv2v_out.v:18355.34-18355.46" */
input [38:0] data_rdata_i;
wire [38:0] data_rdata_i;
/* cellift = 32'd1 */
input [38:0] data_rdata_i_t0;
wire [38:0] data_rdata_i_t0;
/* src = "generated/sv2v_out.v:18346.13-18346.23" */
output data_req_o;
wire data_req_o;
/* cellift = 32'd1 */
output data_req_o_t0;
wire data_req_o_t0;
/* src = "generated/sv2v_out.v:18348.13-18348.26" */
input data_rvalid_i;
wire data_rvalid_i;
/* cellift = 32'd1 */
input data_rvalid_i_t0;
wire data_rvalid_i_t0;
/* src = "generated/sv2v_out.v:18385.6-18385.21" */
reg data_sign_ext_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18385.6-18385.21" */
reg data_sign_ext_q_t0;
/* src = "generated/sv2v_out.v:18384.12-18384.23" */
reg [1:0] data_type_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18384.12-18384.23" */
reg [1:0] data_type_q_t0;
/* src = "generated/sv2v_out.v:18389.13-18389.23" */
wire [31:0] data_wdata;
/* src = "generated/sv2v_out.v:18354.35-18354.47" */
output [38:0] data_wdata_o;
wire [38:0] data_wdata_o;
/* cellift = 32'd1 */
output [38:0] data_wdata_o_t0;
wire [38:0] data_wdata_o_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18389.13-18389.23" */
wire [31:0] data_wdata_t0;
/* src = "generated/sv2v_out.v:18352.14-18352.23" */
output data_we_o;
wire data_we_o;
/* cellift = 32'd1 */
output data_we_o_t0;
wire data_we_o_t0;
/* src = "generated/sv2v_out.v:18386.6-18386.15" */
reg data_we_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18386.6-18386.15" */
reg data_we_q_t0;
/* src = "generated/sv2v_out.v:18545.30-18545.44" */
wire [38:0] \g_mem_rdata_ecc.data_rdata_buf ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18545.30-18545.44" */
wire [38:0] \g_mem_rdata_ecc.data_rdata_buf_t0 ;
/* src = "generated/sv2v_out.v:18544.15-18544.22" */
wire [1:0] \g_mem_rdata_ecc.ecc_err ;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18544.15-18544.22" */
wire [1:0] \g_mem_rdata_ecc.ecc_err_t0 ;
/* src = "generated/sv2v_out.v:18396.6-18396.25" */
wire handle_misaligned_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18396.6-18396.25" */
wire handle_misaligned_d_t0;
/* src = "generated/sv2v_out.v:18395.6-18395.25" */
reg handle_misaligned_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18395.6-18395.25" */
reg handle_misaligned_q_t0;
/* src = "generated/sv2v_out.v:18368.14-18368.24" */
output load_err_o;
wire load_err_o;
/* cellift = 32'd1 */
output load_err_o_t0;
wire load_err_o_t0;
/* src = "generated/sv2v_out.v:18369.14-18369.34" */
output load_resp_intg_err_o;
wire load_resp_intg_err_o;
/* cellift = 32'd1 */
output load_resp_intg_err_o_t0;
wire load_resp_intg_err_o_t0;
/* src = "generated/sv2v_out.v:18403.12-18403.21" */
reg [2:0] ls_fsm_cs;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18403.12-18403.21" */
reg [2:0] ls_fsm_cs_t0;
/* src = "generated/sv2v_out.v:18404.12-18404.21" */
wire [2:0] ls_fsm_ns;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18404.12-18404.21" */
wire [2:0] ls_fsm_ns_t0;
/* src = "generated/sv2v_out.v:18400.6-18400.15" */
wire lsu_err_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18400.6-18400.15" */
wire lsu_err_d_t0;
/* src = "generated/sv2v_out.v:18399.6-18399.15" */
reg lsu_err_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18399.6-18399.15" */
reg lsu_err_q_t0;
/* src = "generated/sv2v_out.v:18360.21-18360.32" */
output [31:0] lsu_rdata_o;
wire [31:0] lsu_rdata_o;
/* cellift = 32'd1 */
output [31:0] lsu_rdata_o_t0;
wire [31:0] lsu_rdata_o_t0;
/* src = "generated/sv2v_out.v:18361.14-18361.31" */
output lsu_rdata_valid_o;
wire lsu_rdata_valid_o;
/* cellift = 32'd1 */
output lsu_rdata_valid_o_t0;
wire lsu_rdata_valid_o_t0;
/* src = "generated/sv2v_out.v:18366.14-18366.28" */
output lsu_req_done_o;
wire lsu_req_done_o;
/* cellift = 32'd1 */
output lsu_req_done_o_t0;
wire lsu_req_done_o_t0;
/* src = "generated/sv2v_out.v:18362.13-18362.22" */
input lsu_req_i;
wire lsu_req_i;
/* cellift = 32'd1 */
input lsu_req_i_t0;
wire lsu_req_i_t0;
/* src = "generated/sv2v_out.v:18367.14-18367.30" */
output lsu_resp_valid_o;
wire lsu_resp_valid_o;
/* cellift = 32'd1 */
output lsu_resp_valid_o_t0;
wire lsu_resp_valid_o_t0;
/* src = "generated/sv2v_out.v:18359.13-18359.27" */
input lsu_sign_ext_i;
wire lsu_sign_ext_i;
/* cellift = 32'd1 */
input lsu_sign_ext_i_t0;
wire lsu_sign_ext_i_t0;
/* src = "generated/sv2v_out.v:18357.19-18357.29" */
input [1:0] lsu_type_i;
wire [1:0] lsu_type_i;
/* cellift = 32'd1 */
input [1:0] lsu_type_i_t0;
wire [1:0] lsu_type_i_t0;
/* src = "generated/sv2v_out.v:18358.20-18358.31" */
input [31:0] lsu_wdata_i;
wire [31:0] lsu_wdata_i;
/* cellift = 32'd1 */
input [31:0] lsu_wdata_i_t0;
wire [31:0] lsu_wdata_i_t0;
/* src = "generated/sv2v_out.v:18356.13-18356.21" */
input lsu_we_i;
wire lsu_we_i;
/* cellift = 32'd1 */
input lsu_we_i_t0;
wire lsu_we_i_t0;
/* src = "generated/sv2v_out.v:18373.13-18373.24" */
output perf_load_o;
wire perf_load_o;
/* cellift = 32'd1 */
output perf_load_o_t0;
wire perf_load_o_t0;
/* src = "generated/sv2v_out.v:18374.13-18374.25" */
output perf_store_o;
wire perf_store_o;
/* cellift = 32'd1 */
output perf_store_o_t0;
wire perf_store_o_t0;
/* src = "generated/sv2v_out.v:18398.6-18398.15" */
wire pmp_err_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18398.6-18398.15" */
wire pmp_err_d_t0;
/* src = "generated/sv2v_out.v:18397.6-18397.15" */
reg pmp_err_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18397.6-18397.15" */
reg pmp_err_q_t0;
/* src = "generated/sv2v_out.v:18393.13-18393.24" */
wire [31:0] rdata_b_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18393.13-18393.24" */
wire [31:0] rdata_b_ext_t0;
/* src = "generated/sv2v_out.v:18392.13-18392.24" */
wire [31:0] rdata_h_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18392.13-18392.24" */
wire [31:0] rdata_h_ext_t0;
/* src = "generated/sv2v_out.v:18383.12-18383.26" */
reg [1:0] rdata_offset_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18383.12-18383.26" */
reg [1:0] rdata_offset_q_t0;
/* src = "generated/sv2v_out.v:18382.13-18382.20" */
reg [31:8] rdata_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18382.13-18382.20" */
reg [31:8] rdata_q_t0;
/* src = "generated/sv2v_out.v:18381.6-18381.18" */
wire rdata_update;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18381.6-18381.18" */
wire rdata_update_t0;
/* src = "generated/sv2v_out.v:18391.13-18391.24" */
wire [31:0] rdata_w_ext;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18391.13-18391.24" */
wire [31:0] rdata_w_ext_t0;
/* src = "generated/sv2v_out.v:18345.13-18345.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:18394.7-18394.30" */
wire split_misaligned_access;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:18394.7-18394.30" */
wire split_misaligned_access_t0;
/* src = "generated/sv2v_out.v:18370.14-18370.25" */
output store_err_o;
wire store_err_o;
/* cellift = 32'd1 */
output store_err_o_t0;
wire store_err_o_t0;
/* src = "generated/sv2v_out.v:18371.14-18371.35" */
output store_resp_intg_err_o;
wire store_resp_intg_err_o;
/* cellift = 32'd1 */
output store_resp_intg_err_o_t0;
wire store_resp_intg_err_o_t0;
assign _0082_ = data_gnt_i & /* src = "generated/sv2v_out.v:18609.20-18609.62" */ _0904_;
assign lsu_req_done_o = _0909_ & /* src = "generated/sv2v_out.v:18640.26-18640.81" */ _0892_;
assign lsu_resp_valid_o = _0913_ & /* src = "generated/sv2v_out.v:18655.28-18655.77" */ _0894_;
assign _0084_ = _0894_ & /* src = "generated/sv2v_out.v:18656.32-18656.67" */ data_rvalid_i;
assign _0086_ = _0084_ & /* src = "generated/sv2v_out.v:18656.31-18656.87" */ _0906_;
assign _0088_ = _0086_ & /* src = "generated/sv2v_out.v:18656.30-18656.101" */ _0789_;
assign lsu_rdata_valid_o = _0088_ & /* src = "generated/sv2v_out.v:18656.29-18656.119" */ _0907_;
assign _0090_ = data_or_pmp_err & /* src = "generated/sv2v_out.v:18674.23-18674.51" */ _0789_;
assign load_err_o = _0090_ & /* src = "generated/sv2v_out.v:18674.22-18674.71" */ lsu_resp_valid_o;
assign _0092_ = data_or_pmp_err & /* src = "generated/sv2v_out.v:18675.24-18675.51" */ data_we_q;
assign store_err_o = _0092_ & /* src = "generated/sv2v_out.v:18675.23-18675.71" */ lsu_resp_valid_o;
assign load_resp_intg_err_o = _0094_ & /* src = "generated/sv2v_out.v:18676.32-18676.76" */ _0789_;
assign _0094_ = data_intg_err & /* src = "generated/sv2v_out.v:18677.34-18677.63" */ data_rvalid_i;
assign store_resp_intg_err_o = _0094_ & /* src = "generated/sv2v_out.v:18677.33-18677.76" */ data_we_q;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME ls_fsm_cs_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) ls_fsm_cs_t0 <= 3'h0;
else ls_fsm_cs_t0 <= ls_fsm_ns_t0;
assign _0096_ = ~ _0238_;
assign _0098_ = ~ _0240_;
assign _0099_ = ~ _0242_;
assign _0100_ = ~ rdata_update;
assign _0101_ = ~ addr_update;
assign _0097_ = ~ ctrl_update;
assign _0744_ = handle_misaligned_d ^ handle_misaligned_q;
assign _0745_ = lsu_we_i ^ data_we_q;
assign _0746_ = pmp_err_d ^ pmp_err_q;
assign _0747_ = lsu_err_d ^ lsu_err_q;
assign _0748_ = data_rdata_i[31:8] ^ rdata_q;
assign _0749_ = addr_last_d ^ addr_last_o;
assign _0750_ = adder_result_ex_i[1:0] ^ rdata_offset_q;
assign _0751_ = lsu_type_i ^ data_type_q;
assign _0752_ = lsu_sign_ext_i ^ data_sign_ext_q;
assign _0580_ = handle_misaligned_d_t0 | handle_misaligned_q_t0;
assign _0584_ = lsu_we_i_t0 | data_we_q_t0;
assign _0588_ = pmp_err_d_t0 | pmp_err_q_t0;
assign _0592_ = lsu_err_d_t0 | lsu_err_q_t0;
assign _0596_ = data_rdata_i_t0[31:8] | rdata_q_t0;
assign _0600_ = addr_last_d_t0 | addr_last_o_t0;
assign _0604_ = adder_result_ex_i_t0[1:0] | rdata_offset_q_t0;
assign _0608_ = lsu_type_i_t0 | data_type_q_t0;
assign _0612_ = lsu_sign_ext_i_t0 | data_sign_ext_q_t0;
assign _0581_ = _0744_ | _0580_;
assign _0585_ = _0745_ | _0584_;
assign _0589_ = _0746_ | _0588_;
assign _0593_ = _0747_ | _0592_;
assign _0597_ = _0748_ | _0596_;
assign _0601_ = _0749_ | _0600_;
assign _0605_ = _0750_ | _0604_;
assign _0609_ = _0751_ | _0608_;
assign _0613_ = _0752_ | _0612_;
assign _0286_ = _0238_ & handle_misaligned_d_t0;
assign _0289_ = ctrl_update & lsu_we_i_t0;
assign _0292_ = _0240_ & pmp_err_d_t0;
assign _0295_ = _0242_ & lsu_err_d_t0;
assign _0298_ = { rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update, rdata_update } & data_rdata_i_t0[31:8];
assign _0301_ = { addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update, addr_update } & addr_last_d_t0;
assign _0304_ = { ctrl_update, ctrl_update } & adder_result_ex_i_t0[1:0];
assign _0307_ = { ctrl_update, ctrl_update } & lsu_type_i_t0;
assign _0310_ = ctrl_update & lsu_sign_ext_i_t0;
assign _0287_ = _0096_ & handle_misaligned_q_t0;
assign _0290_ = _0097_ & data_we_q_t0;
assign _0293_ = _0098_ & pmp_err_q_t0;
assign _0296_ = _0099_ & lsu_err_q_t0;
assign _0299_ = { _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_, _0100_ } & rdata_q_t0;
assign _0302_ = { _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_, _0101_ } & addr_last_o_t0;
assign _0305_ = { _0097_, _0097_ } & rdata_offset_q_t0;
assign _0308_ = { _0097_, _0097_ } & data_type_q_t0;
assign _0311_ = _0097_ & data_sign_ext_q_t0;
assign _0288_ = _0581_ & _0239_;
assign _0291_ = _0585_ & ctrl_update_t0;
assign _0294_ = _0589_ & _0241_;
assign _0297_ = _0593_ & _0243_;
assign _0300_ = _0597_ & { rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0, rdata_update_t0 };
assign _0303_ = _0601_ & { addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0, addr_update_t0 };
assign _0306_ = _0605_ & { ctrl_update_t0, ctrl_update_t0 };
assign _0309_ = _0609_ & { ctrl_update_t0, ctrl_update_t0 };
assign _0312_ = _0613_ & ctrl_update_t0;
assign _0582_ = _0286_ | _0287_;
assign _0586_ = _0289_ | _0290_;
assign _0590_ = _0292_ | _0293_;
assign _0594_ = _0295_ | _0296_;
assign _0598_ = _0298_ | _0299_;
assign _0602_ = _0301_ | _0302_;
assign _0606_ = _0304_ | _0305_;
assign _0610_ = _0307_ | _0308_;
assign _0614_ = _0310_ | _0311_;
assign _0583_ = _0582_ | _0288_;
assign _0587_ = _0586_ | _0291_;
assign _0591_ = _0590_ | _0294_;
assign _0595_ = _0594_ | _0297_;
assign _0599_ = _0598_ | _0300_;
assign _0603_ = _0602_ | _0303_;
assign _0607_ = _0606_ | _0306_;
assign _0611_ = _0610_ | _0309_;
assign _0615_ = _0614_ | _0312_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME handle_misaligned_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) handle_misaligned_q_t0 <= 1'h0;
else handle_misaligned_q_t0 <= _0583_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME data_we_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) data_we_q_t0 <= 1'h0;
else data_we_q_t0 <= _0587_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME pmp_err_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) pmp_err_q_t0 <= 1'h0;
else pmp_err_q_t0 <= _0591_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME lsu_err_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) lsu_err_q_t0 <= 1'h0;
else lsu_err_q_t0 <= _0595_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME rdata_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q_t0 <= 24'h000000;
else rdata_q_t0 <= _0599_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME addr_last_o_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) addr_last_o_t0 <= 32'd0;
else addr_last_o_t0 <= _0603_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME rdata_offset_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_offset_q_t0 <= 2'h0;
else rdata_offset_q_t0 <= _0607_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME data_type_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) data_type_q_t0 <= 2'h0;
else data_type_q_t0 <= _0611_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME data_sign_ext_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) data_sign_ext_q_t0 <= 1'h0;
else data_sign_ext_q_t0 <= _0615_;
assign _0248_ = data_gnt_i_t0 & _0904_;
assign _0251_ = _0910_ & _0892_;
assign _0254_ = _0901_ & _0894_;
assign _0257_ = busy_o_t0 & data_rvalid_i;
assign _0260_ = _0085_ & _0906_;
assign _0263_ = _0087_ & _0789_;
assign _0266_ = _0089_ & _0907_;
assign _0269_ = data_or_pmp_err_t0 & _0789_;
assign _0272_ = _0091_ & lsu_resp_valid_o;
assign _0275_ = data_or_pmp_err_t0 & data_we_q;
assign _0276_ = _0093_ & lsu_resp_valid_o;
assign _0279_ = _0095_ & _0789_;
assign _0282_ = data_intg_err_t0 & data_rvalid_i;
assign _0285_ = _0095_ & data_we_q;
assign _0249_ = _0905_ & data_gnt_i;
assign _0252_ = _0893_ & _0909_;
assign _0255_ = busy_o_t0 & _0913_;
assign _0258_ = data_rvalid_i_t0 & _0894_;
assign _0261_ = data_or_pmp_err_t0 & _0084_;
assign _0264_ = data_we_q_t0 & _0086_;
assign _0267_ = data_intg_err_t0 & _0088_;
assign _0273_ = lsu_resp_valid_o_t0 & _0090_;
assign _0270_ = data_we_q_t0 & data_or_pmp_err;
assign _0277_ = lsu_resp_valid_o_t0 & _0092_;
assign _0280_ = data_we_q_t0 & _0094_;
assign _0283_ = data_rvalid_i_t0 & data_intg_err;
assign _0250_ = data_gnt_i_t0 & _0905_;
assign _0253_ = _0910_ & _0893_;
assign _0256_ = _0901_ & busy_o_t0;
assign _0259_ = busy_o_t0 & data_rvalid_i_t0;
assign _0262_ = _0085_ & data_or_pmp_err_t0;
assign _0265_ = _0087_ & data_we_q_t0;
assign _0268_ = _0089_ & data_intg_err_t0;
assign _0271_ = data_or_pmp_err_t0 & data_we_q_t0;
assign _0274_ = _0091_ & lsu_resp_valid_o_t0;
assign _0278_ = _0093_ & lsu_resp_valid_o_t0;
assign _0284_ = data_intg_err_t0 & data_rvalid_i_t0;
assign _0281_ = _0095_ & data_we_q_t0;
assign _0566_ = _0248_ | _0249_;
assign _0567_ = _0251_ | _0252_;
assign _0568_ = _0254_ | _0255_;
assign _0569_ = _0257_ | _0258_;
assign _0570_ = _0260_ | _0261_;
assign _0571_ = _0263_ | _0264_;
assign _0572_ = _0266_ | _0267_;
assign _0573_ = _0269_ | _0270_;
assign _0574_ = _0272_ | _0273_;
assign _0575_ = _0275_ | _0270_;
assign _0576_ = _0276_ | _0277_;
assign _0577_ = _0279_ | _0280_;
assign _0578_ = _0282_ | _0283_;
assign _0579_ = _0285_ | _0280_;
assign _0083_ = _0566_ | _0250_;
assign lsu_req_done_o_t0 = _0567_ | _0253_;
assign lsu_resp_valid_o_t0 = _0568_ | _0256_;
assign _0085_ = _0569_ | _0259_;
assign _0087_ = _0570_ | _0262_;
assign _0089_ = _0571_ | _0265_;
assign lsu_rdata_valid_o_t0 = _0572_ | _0268_;
assign _0091_ = _0573_ | _0271_;
assign load_err_o_t0 = _0574_ | _0274_;
assign _0093_ = _0575_ | _0271_;
assign store_err_o_t0 = _0576_ | _0278_;
assign load_resp_intg_err_o_t0 = _0577_ | _0281_;
assign _0095_ = _0578_ | _0284_;
assign store_resp_intg_err_o_t0 = _0579_ | _0281_;
assign _0102_ = | { lsu_req_i_t0, data_gnt_i_t0, busy_o_t0 };
assign _0103_ = | { _0919_, _0901_, data_gnt_i_t0 };
assign _0104_ = | { lsu_req_i_t0, busy_o_t0 };
assign _0105_ = | { _0040_, _0921_ };
assign _0106_ = | { _0040_, _0917_ };
assign _0107_ = | { _0915_, data_rvalid_i_t0 };
assign _0108_ = | { _0919_, _0901_ };
assign _0110_ = | data_type_q_t0;
assign _0111_ = | rdata_offset_q_t0;
assign _0114_ = ~ { busy_o_t0, lsu_req_i_t0, data_gnt_i_t0 };
assign _0115_ = ~ { _0919_, _0901_, data_gnt_i_t0 };
assign _0116_ = ~ { busy_o_t0, lsu_req_i_t0 };
assign _0117_ = ~ { _0921_, _0040_ };
assign _0118_ = ~ { _0917_, _0040_ };
assign _0119_ = ~ { _0915_, data_rvalid_i_t0 };
assign _0120_ = ~ { _0919_, _0901_ };
assign _0122_ = ~ data_type_q_t0;
assign _0123_ = ~ rdata_offset_q_t0;
assign _0313_ = { _0894_, lsu_req_i, data_gnt_i } & _0114_;
assign _0314_ = { _0918_, _0900_, data_gnt_i } & _0115_;
assign _0315_ = { _0894_, lsu_req_i } & _0116_;
assign _0316_ = { _0920_, _0899_ } & _0117_;
assign _0317_ = { _0916_, _0899_ } & _0118_;
assign _0319_ = { _0914_, data_rvalid_i } & _0119_;
assign _0320_ = { _0918_, _0900_ } & _0120_;
assign _0471_ = ls_fsm_cs & _0121_;
assign _0523_ = data_type_q & _0122_;
assign _0548_ = rdata_offset_q & _0123_;
assign _0805_ = _0313_ == { _0114_[2:1], 1'h0 };
assign _0806_ = _0314_ == { _0115_[2], 2'h0 };
assign _0807_ = _0315_ == { _0116_[1], 1'h0 };
assign _0808_ = _0316_ == { _0117_[1], 1'h0 };
assign _0809_ = _0317_ == { _0118_[1], 1'h0 };
assign _0810_ = _0319_ == { _0119_[1], 1'h0 };
assign _0811_ = _0320_ == { _0120_[1], 1'h0 };
assign _0812_ = _0471_ == { 2'h0, _0121_[0] };
assign _0813_ = _0471_ == { _0121_[2], 2'h0 };
assign _0814_ = _0471_ == { 1'h0, _0121_[1:0] };
assign _0815_ = _0471_ == { 1'h0, _0121_[1], 1'h0 };
assign _0816_ = _0523_ == { _0122_[1], 1'h0 };
assign _0817_ = _0523_ == _0122_;
assign _0818_ = _0523_ == { 1'h0, _0122_[0] };
assign _0819_ = _0548_ == _0123_;
assign _0820_ = _0548_ == { _0123_[1], 1'h0 };
assign _0821_ = _0548_ == { 1'h0, _0123_[0] };
assign _0822_ = _0470_ == _0124_;
assign _0823_ = _0470_ == { _0124_[1], 1'h0 };
assign _0824_ = _0470_ == { 1'h0, _0124_[0] };
assign _0825_ = _0555_ == { _0125_[1], 1'h0 };
assign _0826_ = _0555_ == _0125_;
assign _0827_ = _0555_ == { 1'h0, _0125_[0] };
assign _0221_ = _0805_ & _0102_;
assign _0223_ = _0806_ & _0103_;
assign _0225_ = _0807_ & _0104_;
assign _0227_ = _0808_ & _0105_;
assign _0229_ = _0809_ & _0106_;
assign _0233_ = _0810_ & _0107_;
assign _0235_ = _0811_ & _0108_;
assign _0921_ = _0812_ & _0109_;
assign _0915_ = _0813_ & _0109_;
assign _0917_ = _0814_ & _0109_;
assign _0919_ = _0815_ & _0109_;
assign _0923_[0] = _0816_ & _0110_;
assign _0923_[1] = _0817_ & _0110_;
assign _0927_ = _0818_ & _0110_;
assign _0929_ = _0819_ & _0111_;
assign _0931_ = _0820_ & _0111_;
assign _0933_ = _0821_ & _0111_;
assign _0877_[3] = _0822_ & _0112_;
assign _0935_ = _0823_ & _0112_;
assign _0879_[1] = _0824_ & _0112_;
assign _0938_[0] = _0825_ & _0113_;
assign _0938_[1] = _0826_ & _0113_;
assign _0890_ = _0827_ & _0113_;
/* src = "generated/sv2v_out.v:18641.2-18653.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME handle_misaligned_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) handle_misaligned_q <= 1'h0;
else if (_0238_) handle_misaligned_q <= handle_misaligned_d;
/* src = "generated/sv2v_out.v:18460.2-18472.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME data_we_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) data_we_q <= 1'h0;
else if (ctrl_update) data_we_q <= lsu_we_i;
/* src = "generated/sv2v_out.v:18641.2-18653.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME pmp_err_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) pmp_err_q <= 1'h0;
else if (_0240_) pmp_err_q <= pmp_err_d;
/* src = "generated/sv2v_out.v:18641.2-18653.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME lsu_err_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) lsu_err_q <= 1'h0;
else if (_0242_) lsu_err_q <= lsu_err_d;
/* src = "generated/sv2v_out.v:18455.2-18459.34" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME rdata_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_q <= 24'h000000;
else if (rdata_update) rdata_q <= data_rdata_i[31:8];
/* src = "generated/sv2v_out.v:18474.2-18478.31" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME addr_last_o */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) addr_last_o <= 32'd0;
else if (addr_update) addr_last_o <= addr_last_d;
/* src = "generated/sv2v_out.v:18460.2-18472.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME rdata_offset_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_offset_q <= 2'h0;
else if (ctrl_update) rdata_offset_q <= adder_result_ex_i[1:0];
/* src = "generated/sv2v_out.v:18460.2-18472.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME data_type_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) data_type_q <= 2'h0;
else if (ctrl_update) data_type_q <= lsu_type_i;
/* src = "generated/sv2v_out.v:18460.2-18472.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME data_sign_ext_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) data_sign_ext_q <= 1'h0;
else if (ctrl_update) data_sign_ext_q <= lsu_sign_ext_i;
assign _0455_ = _0888_ & _0902_;
assign _0458_ = _0890_ & _0891_;
assign _0456_ = _0903_ & _0887_;
assign _0459_ = _0877_[3] & _0889_;
assign _0457_ = _0888_ & _0903_;
assign _0460_ = _0890_ & _0877_[3];
assign _0703_ = _0455_ | _0456_;
assign _0704_ = _0458_ | _0459_;
assign _0896_ = _0703_ | _0457_;
assign _0898_ = _0704_ | _0460_;
assign _0126_ = | { _0917_, _0921_, _0919_, busy_o_t0 };
assign _0127_ = | { _0915_, _0919_, busy_o_t0 };
assign _0128_ = | { _0917_, _0921_, _0919_ };
assign _0129_ = | { _0917_, _0921_ };
assign _0130_ = | { _0915_, _0919_ };
assign _0131_ = | { _0915_, _0917_, _0919_ };
assign _0132_ = | ls_fsm_ns_t0;
assign _0112_ = | adder_result_ex_i_t0[1:0];
assign _0109_ = | ls_fsm_cs_t0;
assign _0133_ = | _0923_;
assign _0134_ = | _0938_;
assign _0113_ = | lsu_type_i_t0;
assign _0135_ = | \g_mem_rdata_ecc.ecc_err_t0 ;
assign _0136_ = ~ { _0919_, _0917_, busy_o_t0, _0921_ };
assign _0137_ = ~ { _0919_, _0915_, busy_o_t0 };
assign _0138_ = ~ { _0921_, _0919_, _0917_ };
assign _0139_ = ~ { _0921_, _0917_ };
assign _0140_ = ~ { _0919_, _0915_ };
assign _0141_ = ~ { _0919_, _0917_, _0915_ };
assign _0142_ = ~ ls_fsm_ns_t0;
assign _0124_ = ~ adder_result_ex_i_t0[1:0];
assign _0121_ = ~ ls_fsm_cs_t0;
assign _0143_ = ~ _0923_;
assign _0144_ = ~ _0938_;
assign _0125_ = ~ lsu_type_i_t0;
assign _0145_ = ~ \g_mem_rdata_ecc.ecc_err_t0 ;
assign _0318_ = { _0918_, _0916_, _0894_, _0920_ } & _0136_;
assign _0321_ = { _0918_, _0914_, _0894_ } & _0137_;
assign _0322_ = { _0920_, _0918_, _0916_ } & _0138_;
assign _0323_ = { _0920_, _0916_ } & _0139_;
assign _0324_ = { _0918_, _0914_ } & _0140_;
assign _0325_ = { _0918_, _0916_, _0914_ } & _0141_;
assign _0454_ = ls_fsm_ns & _0142_;
assign _0470_ = adder_result_ex_i[1:0] & _0124_;
assign _0522_ = _0922_ & _0143_;
assign _0549_ = _0937_ & _0144_;
assign _0555_ = lsu_type_i & _0125_;
assign _0556_ = \g_mem_rdata_ecc.ecc_err  & _0145_;
assign _0146_ = ! _0318_;
assign _0147_ = ! _0321_;
assign _0148_ = ! _0322_;
assign _0149_ = ! _0323_;
assign _0150_ = ! _0324_;
assign _0151_ = ! _0325_;
assign _0152_ = ! _0454_;
assign _0153_ = ! _0470_;
assign _0154_ = ! _0471_;
assign _0155_ = ! _0522_;
assign _0156_ = ! _0549_;
assign _0157_ = ! _0555_;
assign _0158_ = ! _0556_;
assign _0231_ = _0146_ & _0126_;
assign _0237_ = _0147_ & _0127_;
assign _0245_ = _0148_ & _0128_;
assign _0247_ = _0149_ & _0129_;
assign _0211_ = _0150_ & _0130_;
assign _0213_ = _0151_ & _0131_;
assign _0893_ = _0152_ & _0132_;
assign _0903_ = _0153_ & _0112_;
assign busy_o_t0 = _0154_ & _0109_;
assign _0925_ = _0155_ & _0133_;
assign _0940_ = _0156_ & _0134_;
assign _0888_ = _0157_ & _0113_;
assign data_intg_err_t0 = _0158_ & _0135_;
assign _0159_ = ~ _0895_;
assign _0160_ = ~ data_rvalid_i;
assign _0161_ = ~ data_gnt_i;
assign _0162_ = ~ _0897_;
assign _0163_ = ~ pmp_err_q;
assign _0461_ = _0896_ & _0162_;
assign _0464_ = data_rvalid_i_t0 & _0163_;
assign _0467_ = data_gnt_i_t0 & _0163_;
assign _0462_ = _0898_ & _0159_;
assign _0465_ = pmp_err_q_t0 & _0160_;
assign _0468_ = pmp_err_q_t0 & _0161_;
assign _0463_ = _0896_ & _0898_;
assign _0466_ = data_rvalid_i_t0 & pmp_err_q_t0;
assign _0469_ = data_gnt_i_t0 & pmp_err_q_t0;
assign _0705_ = _0461_ | _0462_;
assign _0706_ = _0464_ | _0465_;
assign _0707_ = _0467_ | _0468_;
assign split_misaligned_access_t0 = _0705_ | _0463_;
assign _0901_ = _0706_ | _0466_;
assign _0040_ = _0707_ | _0469_;
assign _0164_ = ~ { _0916_, _0916_, _0916_ };
assign _0165_ = ~ { _0914_, _0914_, _0914_ };
assign _0166_ = ~ { _0920_, _0920_, _0920_ };
assign _0167_ = ~ { _0212_, _0212_, _0212_ };
assign _0168_ = ~ _0918_;
assign _0169_ = ~ _0914_;
assign _0170_ = ~ _0916_;
assign _0171_ = ~ _0920_;
assign _0172_ = ~ _0560_;
assign _0173_ = ~ _0246_;
assign _0174_ = ~ _0212_;
assign _0175_ = ~ _0244_;
assign _0176_ = ~ _0210_;
assign _0177_ = ~ { _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_ };
assign _0178_ = ~ { _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_ };
assign _0179_ = ~ { _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_ };
assign _0180_ = ~ { _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_ };
assign _0181_ = ~ { _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_ };
assign _0182_ = ~ { _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_ };
assign _0183_ = ~ { _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_ };
assign _0184_ = ~ { _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_ };
assign _0185_ = ~ { _0564_, _0564_, _0564_, _0564_ };
assign _0186_ = ~ { _0889_, _0889_, _0889_, _0889_ };
assign _0187_ = ~ { _0939_, _0939_, _0939_, _0939_ };
assign _0188_ = ~ { data_rvalid_i, data_rvalid_i, data_rvalid_i };
assign _0189_ = ~ { _0899_, _0899_, _0899_ };
assign _0190_ = ~ { data_gnt_i, data_gnt_i, data_gnt_i };
assign _0191_ = ~ { _0900_, _0900_, _0900_ };
assign _0192_ = ~ { lsu_req_i, lsu_req_i, lsu_req_i };
assign _0193_ = ~ lsu_req_i;
assign _0194_ = ~ { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q };
assign _0195_ = ~ { handle_misaligned_q, handle_misaligned_q, handle_misaligned_q, handle_misaligned_q };
assign _0196_ = ~ { addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o };
assign _0622_ = { _0917_, _0917_, _0917_ } | _0164_;
assign _0625_ = { _0915_, _0915_, _0915_ } | _0165_;
assign _0629_ = { _0921_, _0921_, _0921_ } | _0166_;
assign _0632_ = { _0213_, _0213_, _0213_ } | _0167_;
assign _0635_ = _0919_ | _0168_;
assign _0637_ = _0915_ | _0169_;
assign _0642_ = _0917_ | _0170_;
assign _0644_ = _0921_ | _0171_;
assign _0646_ = _0561_ | _0172_;
assign _0649_ = _0247_ | _0173_;
assign _0656_ = _0213_ | _0174_;
assign _0659_ = _0245_ | _0175_;
assign _0661_ = _0211_ | _0176_;
assign _0662_ = { _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_ } | _0177_;
assign _0665_ = { _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_ } | _0178_;
assign _0668_ = { _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_ } | _0179_;
assign _0671_ = { _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_ } | _0180_;
assign _0674_ = { _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_ } | _0181_;
assign _0683_ = { _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3] } | _0182_;
assign _0686_ = { _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1] } | _0183_;
assign _0689_ = { _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_ } | _0184_;
assign _0692_ = { _0565_, _0565_, _0565_, _0565_ } | _0185_;
assign _0697_ = { _0890_, _0890_, _0890_, _0890_ } | _0186_;
assign _0700_ = { _0940_, _0940_, _0940_, _0940_ } | _0187_;
assign _0712_ = { data_rvalid_i_t0, data_rvalid_i_t0, data_rvalid_i_t0 } | _0188_;
assign _0715_ = { _0040_, _0040_, _0040_ } | _0189_;
assign _0717_ = { data_gnt_i_t0, data_gnt_i_t0, data_gnt_i_t0 } | _0190_;
assign _0720_ = { _0901_, _0901_, _0901_ } | _0191_;
assign _0724_ = { lsu_req_i_t0, lsu_req_i_t0, lsu_req_i_t0 } | _0192_;
assign _0728_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } | _0194_;
assign _0738_ = { handle_misaligned_q_t0, handle_misaligned_q_t0, handle_misaligned_q_t0, handle_misaligned_q_t0 } | _0195_;
assign _0741_ = { addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0 } | _0196_;
assign _0623_ = { _0917_, _0917_, _0917_ } | { _0916_, _0916_, _0916_ };
assign _0626_ = { _0915_, _0915_, _0915_ } | { _0914_, _0914_, _0914_ };
assign _0628_ = { busy_o_t0, busy_o_t0, busy_o_t0 } | { _0894_, _0894_, _0894_ };
assign _0630_ = { _0921_, _0921_, _0921_ } | { _0920_, _0920_, _0920_ };
assign _0633_ = { _0213_, _0213_, _0213_ } | { _0212_, _0212_, _0212_ };
assign _0636_ = _0919_ | _0918_;
assign _0638_ = _0915_ | _0914_;
assign _0643_ = _0917_ | _0916_;
assign _0645_ = _0921_ | _0920_;
assign _0647_ = _0561_ | _0560_;
assign _0650_ = _0247_ | _0246_;
assign _0654_ = busy_o_t0 | _0894_;
assign _0657_ = _0213_ | _0212_;
assign _0663_ = { _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_ } | { _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_, _0926_ };
assign _0666_ = { _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_ } | { _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_, _0924_ };
assign _0669_ = { _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_ } | { _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_, _0928_ };
assign _0672_ = { _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_ } | { _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_, _0932_ };
assign _0675_ = { _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_ } | { _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_, _0562_ };
assign _0684_ = { _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3] } | { _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_, _0891_ };
assign _0687_ = { _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1] } | { _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_, _0936_ };
assign _0690_ = { _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_ } | { _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_, _0564_ };
assign _0693_ = { _0565_, _0565_, _0565_, _0565_ } | { _0564_, _0564_, _0564_, _0564_ };
assign _0698_ = { _0890_, _0890_, _0890_, _0890_ } | { _0889_, _0889_, _0889_, _0889_ };
assign _0701_ = { _0940_, _0940_, _0940_, _0940_ } | { _0939_, _0939_, _0939_, _0939_ };
assign _0713_ = data_rvalid_i_t0 | data_rvalid_i;
assign _0714_ = _0040_ | _0899_;
assign _0716_ = data_gnt_i_t0 | data_gnt_i;
assign _0718_ = { data_gnt_i_t0, data_gnt_i_t0, data_gnt_i_t0 } | { data_gnt_i, data_gnt_i, data_gnt_i };
assign _0719_ = _0901_ | _0900_;
assign _0721_ = { _0901_, _0901_, _0901_ } | { _0900_, _0900_, _0900_ };
assign _0725_ = { lsu_req_i_t0, lsu_req_i_t0, lsu_req_i_t0 } | { lsu_req_i, lsu_req_i, lsu_req_i };
assign _0727_ = lsu_req_i_t0 | lsu_req_i;
assign _0729_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } | { data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q, data_sign_ext_q };
assign _0739_ = { handle_misaligned_q_t0, handle_misaligned_q_t0, handle_misaligned_q_t0, handle_misaligned_q_t0 } | { handle_misaligned_q, handle_misaligned_q, handle_misaligned_q, handle_misaligned_q };
assign _0742_ = { addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0 } | { addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o, addr_incr_req_o };
assign _0335_ = _0061_ & _0622_;
assign _0338_ = _0829_ & _0625_;
assign _0343_ = _0833_ & _0629_;
assign _0346_ = _0835_ & _0632_;
assign _0351_ = _0837_ & _0637_;
assign _0354_ = _0015_ & _0635_;
assign _0357_ = _0839_ & _0637_;
assign _0360_ = _0059_ & _0642_;
assign _0362_ = _0006_ & _0644_;
assign _0364_ = _0843_ & _0646_;
assign _0367_ = _0845_ & _0649_;
assign _0370_ = _0055_ & _0642_;
assign _0373_ = _0847_ & _0637_;
assign _0378_ = _0845_ & _0644_;
assign _0381_ = _0851_ & _0656_;
assign _0386_ = _0853_ & _0659_;
assign _0390_ = _0855_ & _0637_;
assign _0395_ = _0857_ & _0661_;
assign _0397_ = rdata_w_ext_t0 & _0662_;
assign _0400_ = _0859_ & _0665_;
assign _0403_ = _0051_ & _0668_;
assign _0406_ = _0017_ & _0671_;
assign _0409_ = _0863_ & _0674_;
assign _0412_ = _0053_ & _0668_;
assign _0415_ = _0019_ & _0671_;
assign _0418_ = _0867_ & _0674_;
assign _0421_ = { data_rdata_i_t0[15:0], rdata_q_t0[31:16] } & _0668_;
assign _0424_ = data_rdata_i_t0[31:0] & _0671_;
assign _0427_ = _0871_ & _0674_;
assign _0430_ = { lsu_wdata_i_t0[15:0], lsu_wdata_i_t0[31:16] } & _0683_;
assign _0433_ = lsu_wdata_i_t0 & _0686_;
assign _0436_ = _0875_ & _0689_;
assign _0439_ = { 2'h0, _0879_[1], _0879_[1] } & _0692_;
assign _0442_ = { 1'h0, _0879_[1], 1'h0, _0879_[1] } & _0692_;
assign _0445_ = { 3'h0, _0879_[1] } & _0692_;
assign _0448_ = _0003_ & _0697_;
assign _0451_ = _0886_ & _0700_;
assign _0484_ = ls_fsm_cs_t0 & _0712_;
assign _0489_ = ls_fsm_cs_t0 & _0715_;
assign _0493_ = ls_fsm_cs_t0 & _0717_;
assign _0499_ = _0072_ & _0720_;
assign _0505_ = { 1'h0, split_misaligned_access_t0, 1'h0 } & _0717_;
assign _0508_ = ls_fsm_cs_t0 & _0724_;
assign _0524_ = { 24'h000000, data_rdata_i_t0[31:24] } & _0728_;
assign _0527_ = { 24'h000000, data_rdata_i_t0[23:16] } & _0728_;
assign _0530_ = { 24'h000000, data_rdata_i_t0[15:8] } & _0728_;
assign _0533_ = { 24'h000000, data_rdata_i_t0[7:0] } & _0728_;
assign _0536_ = { 16'h0000, data_rdata_i_t0[7:0], rdata_q_t0[31:24] } & _0728_;
assign _0539_ = { 16'h0000, data_rdata_i_t0[31:16] } & _0728_;
assign _0542_ = { 16'h0000, data_rdata_i_t0[23:8] } & _0728_;
assign _0545_ = { 16'h0000, data_rdata_i_t0[15:0] } & _0728_;
assign _0550_ = _0069_ & _0738_;
assign _0552_ = _0024_ & _0738_;
assign _0557_ = adder_result_ex_i_t0 & _0741_;
assign _0336_ = _0079_ & _0623_;
assign _0339_ = _0081_ & _0626_;
assign _0341_ = _0008_ & _0628_;
assign _0344_ = _0045_ & _0630_;
assign _0347_ = _0831_ & _0633_;
assign _0349_ = _0030_ & _0636_;
assign _0352_ = _0047_ & _0638_;
assign _0355_ = _0032_ & _0636_;
assign _0358_ = _0049_ & _0638_;
assign _0365_ = _0841_ & _0647_;
assign _0368_ = _0040_ & _0650_;
assign _0371_ = _0067_ & _0643_;
assign _0374_ = _0074_ & _0638_;
assign _0376_ = _0001_ & _0654_;
assign _0379_ = _0040_ & _0645_;
assign _0382_ = _0849_ & _0657_;
assign _0384_ = lsu_req_i_t0 & _0654_;
assign _0388_ = _0021_ & _0636_;
assign _0391_ = _0038_ & _0638_;
assign _0393_ = handle_misaligned_q_t0 & _0643_;
assign _0398_ = rdata_h_ext_t0 & _0663_;
assign _0401_ = rdata_b_ext_t0 & _0666_;
assign _0404_ = _0063_ & _0669_;
assign _0407_ = _0034_ & _0672_;
assign _0410_ = _0861_ & _0675_;
assign _0413_ = _0065_ & _0669_;
assign _0416_ = _0036_ & _0672_;
assign _0419_ = _0865_ & _0675_;
assign _0422_ = { data_rdata_i_t0[23:0], rdata_q_t0[31:24] } & _0669_;
assign _0425_ = { data_rdata_i_t0[7:0], rdata_q_t0 } & _0672_;
assign _0428_ = _0869_ & _0675_;
assign _0431_ = { lsu_wdata_i_t0[7:0], lsu_wdata_i_t0[31:8] } & _0684_;
assign _0434_ = { lsu_wdata_i_t0[23:0], lsu_wdata_i_t0[31:24] } & _0687_;
assign _0437_ = _0873_ & _0690_;
assign _0440_ = { _0877_[3], _0877_[3], 2'h0 } & _0693_;
assign _0443_ = { 1'h0, _0877_[3], 2'h0 } & _0693_;
assign _0449_ = _0057_ & _0698_;
assign _0452_ = _0076_ & _0701_;
assign _0486_ = data_we_q_t0 & _0713_;
assign _0047_ = data_bus_err_i_t0 & _0713_;
assign _0049_ = data_pmp_err_i_t0 & _0713_;
assign _0491_ = lsu_err_q_t0 & _0714_;
assign _0495_ = data_gnt_i_t0 & _0719_;
assign _0497_ = _0083_ & _0719_;
assign _0500_ = { 1'h0, data_gnt_i_t0, data_gnt_i_t0 } & _0721_;
assign _0502_ = data_we_q_t0 & _0719_;
assign _0030_ = _0905_ & _0719_;
assign _0032_ = data_pmp_err_i_t0 & _0719_;
assign _0506_ = { 1'h0, split_misaligned_access_t0, 1'h0 } & _0718_;
assign _0026_ = split_misaligned_access_t0 & _0716_;
assign _0509_ = _0028_ & _0725_;
assign _0006_ = _0026_ & _0727_;
assign _0511_ = data_gnt_i_t0 & _0727_;
assign _0513_ = lsu_we_i_t0 & _0727_;
assign _0516_ = data_pmp_err_i_t0 & _0727_;
assign _0518_ = _0013_ & _0654_;
assign _0520_ = _0011_ & _0654_;
assign _0525_ = { data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31:24] } & _0729_;
assign _0528_ = { data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23:16] } & _0729_;
assign _0531_ = { data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15:8] } & _0729_;
assign _0534_ = { data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7:0] } & _0729_;
assign _0537_ = { data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7], data_rdata_i_t0[7:0], rdata_q_t0[31:24] } & _0729_;
assign _0540_ = { data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31], data_rdata_i_t0[31:16] } & _0729_;
assign _0543_ = { data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23], data_rdata_i_t0[23:8] } & _0729_;
assign _0546_ = { data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15], data_rdata_i_t0[15:0] } & _0729_;
assign _0553_ = _0042_ & _0739_;
assign _0558_ = { adder_result_ex_i_t0[31:2], 2'h0 } & _0742_;
assign _0624_ = _0335_ | _0336_;
assign _0627_ = _0338_ | _0339_;
assign _0631_ = _0343_ | _0344_;
assign _0634_ = _0346_ | _0347_;
assign _0639_ = _0351_ | _0352_;
assign _0640_ = _0354_ | _0355_;
assign _0641_ = _0357_ | _0358_;
assign _0648_ = _0364_ | _0365_;
assign _0651_ = _0367_ | _0368_;
assign _0652_ = _0370_ | _0371_;
assign _0653_ = _0373_ | _0374_;
assign _0655_ = _0378_ | _0379_;
assign _0658_ = _0381_ | _0382_;
assign _0660_ = _0390_ | _0391_;
assign _0664_ = _0397_ | _0398_;
assign _0667_ = _0400_ | _0401_;
assign _0670_ = _0403_ | _0404_;
assign _0673_ = _0406_ | _0407_;
assign _0676_ = _0409_ | _0410_;
assign _0677_ = _0412_ | _0413_;
assign _0678_ = _0415_ | _0416_;
assign _0679_ = _0418_ | _0419_;
assign _0680_ = _0421_ | _0422_;
assign _0681_ = _0424_ | _0425_;
assign _0682_ = _0427_ | _0428_;
assign _0685_ = _0430_ | _0431_;
assign _0688_ = _0433_ | _0434_;
assign _0691_ = _0436_ | _0437_;
assign _0694_ = _0439_ | _0440_;
assign _0695_ = _0442_ | _0443_;
assign _0696_ = _0445_ | _0443_;
assign _0699_ = _0448_ | _0449_;
assign _0702_ = _0451_ | _0452_;
assign _0722_ = _0499_ | _0500_;
assign _0723_ = _0505_ | _0506_;
assign _0726_ = _0508_ | _0509_;
assign _0730_ = _0524_ | _0525_;
assign _0731_ = _0527_ | _0528_;
assign _0732_ = _0530_ | _0531_;
assign _0733_ = _0533_ | _0534_;
assign _0734_ = _0536_ | _0537_;
assign _0735_ = _0539_ | _0540_;
assign _0736_ = _0542_ | _0543_;
assign _0737_ = _0545_ | _0546_;
assign _0740_ = _0552_ | _0553_;
assign _0743_ = _0557_ | _0558_;
assign _0753_ = _0060_ ^ _0078_;
assign _0754_ = _0828_ ^ _0080_;
assign _0755_ = _0832_ ^ _0044_;
assign _0756_ = _0834_ ^ _0830_;
assign _0757_ = _0009_ ^ _0029_;
assign _0758_ = _0836_ ^ _0046_;
assign _0759_ = _0014_ ^ _0031_;
assign _0760_ = _0838_ ^ _0048_;
assign _0761_ = _0058_ ^ _0077_;
assign _0762_ = _0005_ ^ _0043_;
assign _0763_ = _0842_ ^ _0840_;
assign _0764_ = _0844_ ^ _0039_;
assign _0765_ = _0054_ ^ _0066_;
assign _0766_ = _0846_ ^ _0073_;
assign _0767_ = _0850_ ^ _0848_;
assign _0768_ = _0854_ ^ _0037_;
assign _0769_ = rdata_w_ext ^ rdata_h_ext;
assign _0770_ = _0858_ ^ rdata_b_ext;
assign _0771_ = _0050_ ^ _0062_;
assign _0772_ = _0016_ ^ _0033_;
assign _0773_ = _0862_ ^ _0860_;
assign _0774_ = _0052_ ^ _0064_;
assign _0775_ = _0018_ ^ _0035_;
assign _0776_ = _0866_ ^ _0864_;
assign _0777_ = { data_rdata_i[15:0], rdata_q[31:16] } ^ { data_rdata_i[23:0], rdata_q[31:24] };
assign _0778_ = data_rdata_i[31:0] ^ { data_rdata_i[7:0], rdata_q };
assign _0779_ = _0870_ ^ _0868_;
assign _0780_ = { lsu_wdata_i[15:0], lsu_wdata_i[31:16] } ^ { lsu_wdata_i[7:0], lsu_wdata_i[31:8] };
assign _0781_ = lsu_wdata_i ^ { lsu_wdata_i[23:0], lsu_wdata_i[31:24] };
assign _0782_ = _0874_ ^ _0872_;
assign _0783_ = _0878_ ^ _0876_;
assign _0784_ = _0881_ ^ _0880_;
assign _0785_ = _0883_ ^ _0882_;
assign _0786_ = _0884_ ^ _0880_;
assign _0787_ = _0002_ ^ _0056_;
assign _0788_ = _0885_ ^ _0075_;
assign _0790_ = _0070_ ^ _0161_;
assign _0791_ = _0071_ ^ _0943_;
assign _0792_ = _0942_ ^ _0941_;
assign _0793_ = ls_fsm_cs ^ _0027_;
assign _0795_ = { 24'h000000, data_rdata_i[31:24] } ^ { data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31:24] };
assign _0796_ = { 24'h000000, data_rdata_i[23:16] } ^ { data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23:16] };
assign _0797_ = { 24'h000000, data_rdata_i[15:8] } ^ { data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15:8] };
assign _0798_ = { 24'h000000, data_rdata_i[7:0] } ^ { data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7:0] };
assign _0799_ = { 16'h0000, data_rdata_i[7:0], rdata_q[31:24] } ^ { data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7:0], rdata_q[31:24] };
assign _0800_ = { 16'h0000, data_rdata_i[31:16] } ^ { data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31:16] };
assign _0801_ = { 16'h0000, data_rdata_i[23:8] } ^ { data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23:8] };
assign _0802_ = { 16'h0000, data_rdata_i[15:0] } ^ { data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15:0] };
assign _0803_ = _0023_ ^ _0041_;
assign _0804_ = adder_result_ex_i ^ { adder_result_ex_i[31:2], 2'h0 };
assign _0337_ = { _0917_, _0917_, _0917_ } & _0753_;
assign _0340_ = { _0915_, _0915_, _0915_ } & _0754_;
assign _0342_ = { busy_o_t0, busy_o_t0, busy_o_t0 } & _0007_;
assign _0345_ = { _0921_, _0921_, _0921_ } & _0755_;
assign _0348_ = { _0213_, _0213_, _0213_ } & _0756_;
assign _0350_ = _0919_ & _0757_;
assign _0353_ = _0915_ & _0758_;
assign _0356_ = _0919_ & _0759_;
assign _0359_ = _0915_ & _0760_;
assign _0361_ = _0917_ & _0761_;
assign _0363_ = _0921_ & _0762_;
assign _0366_ = _0561_ & _0763_;
assign _0369_ = _0247_ & _0764_;
assign _0372_ = _0917_ & _0765_;
assign _0375_ = _0915_ & _0766_;
assign _0377_ = busy_o_t0 & _0000_;
assign _0380_ = _0921_ & _0764_;
assign _0383_ = _0213_ & _0767_;
assign _0385_ = busy_o_t0 & _0004_;
assign _0387_ = _0245_ & _0198_;
assign _0389_ = _0919_ & _0020_;
assign _0392_ = _0915_ & _0768_;
assign _0394_ = _0917_ & handle_misaligned_q;
assign _0396_ = _0211_ & _0197_;
assign _0399_ = { _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_, _0927_ } & _0769_;
assign _0402_ = { _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_, _0925_ } & _0770_;
assign _0405_ = { _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_ } & _0771_;
assign _0408_ = { _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_ } & _0772_;
assign _0411_ = { _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_ } & _0773_;
assign _0414_ = { _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_ } & _0774_;
assign _0417_ = { _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_ } & _0775_;
assign _0420_ = { _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_ } & _0776_;
assign _0423_ = { _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_, _0929_ } & _0777_;
assign _0426_ = { _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_, _0933_ } & _0778_;
assign _0429_ = { _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_, _0563_ } & _0779_;
assign _0432_ = { _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3], _0877_[3] } & _0780_;
assign _0435_ = { _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1], _0879_[1] } & _0781_;
assign _0438_ = { _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_, _0565_ } & _0782_;
assign _0441_ = { _0565_, _0565_, _0565_, _0565_ } & _0783_;
assign _0444_ = { _0565_, _0565_, _0565_, _0565_ } & _0784_;
assign _0446_ = { _0565_, _0565_, _0565_, _0565_ } & _0785_;
assign _0447_ = { _0565_, _0565_, _0565_, _0565_ } & _0786_;
assign _0450_ = { _0890_, _0890_, _0890_, _0890_ } & _0787_;
assign _0453_ = { _0940_, _0940_, _0940_, _0940_ } & _0788_;
assign _0485_ = { data_rvalid_i_t0, data_rvalid_i_t0, data_rvalid_i_t0 } & ls_fsm_cs;
assign _0487_ = data_rvalid_i_t0 & _0789_;
assign _0488_ = data_rvalid_i_t0 & _0204_;
assign _0490_ = { _0040_, _0040_, _0040_ } & ls_fsm_cs;
assign _0492_ = _0040_ & _0205_;
assign _0494_ = { data_gnt_i_t0, data_gnt_i_t0, data_gnt_i_t0 } & { _0200_, ls_fsm_cs[1:0] };
assign _0496_ = _0901_ & _0790_;
assign _0498_ = _0901_ & _0082_;
assign _0501_ = { _0901_, _0901_, _0901_ } & _0791_;
assign _0503_ = _0901_ & _0789_;
assign _0504_ = { _0040_, _0040_, _0040_ } & { ls_fsm_cs[2], _0199_, ls_fsm_cs[0] };
assign _0507_ = { data_gnt_i_t0, data_gnt_i_t0, data_gnt_i_t0 } & _0792_;
assign _0510_ = { lsu_req_i_t0, lsu_req_i_t0, lsu_req_i_t0 } & _0793_;
assign _0512_ = lsu_req_i_t0 & _0022_;
assign _0514_ = lsu_req_i_t0 & lsu_we_i;
assign _0515_ = lsu_req_i_t0 & _0794_;
assign _0517_ = lsu_req_i_t0 & data_pmp_err_i;
assign _0519_ = busy_o_t0 & _0012_;
assign _0521_ = busy_o_t0 & _0010_;
assign _0526_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } & _0795_;
assign _0529_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } & _0796_;
assign _0532_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } & _0797_;
assign _0535_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } & _0798_;
assign _0538_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } & _0799_;
assign _0541_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } & _0800_;
assign _0544_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } & _0801_;
assign _0547_ = { data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0, data_sign_ext_q_t0 } & _0802_;
assign _0551_ = { handle_misaligned_q_t0, handle_misaligned_q_t0, handle_misaligned_q_t0, handle_misaligned_q_t0 } & { _0068_[3:1], _0201_ };
assign _0554_ = { handle_misaligned_q_t0, handle_misaligned_q_t0, handle_misaligned_q_t0, handle_misaligned_q_t0 } & _0803_;
assign _0559_ = { addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0, addr_incr_req_o_t0 } & _0804_;
assign _0829_ = _0337_ | _0624_;
assign _0831_ = _0340_ | _0627_;
assign _0833_ = _0342_ | _0341_;
assign _0835_ = _0345_ | _0631_;
assign ls_fsm_ns_t0 = _0348_ | _0634_;
assign _0837_ = _0350_ | _0349_;
assign lsu_err_d_t0 = _0353_ | _0639_;
assign _0839_ = _0356_ | _0640_;
assign pmp_err_d_t0 = _0359_ | _0641_;
assign _0841_ = _0361_ | _0360_;
assign _0843_ = _0363_ | _0362_;
assign handle_misaligned_d_t0 = _0366_ | _0648_;
assign ctrl_update_t0 = _0369_ | _0651_;
assign _0847_ = _0372_ | _0652_;
assign _0849_ = _0375_ | _0653_;
assign _0845_ = _0377_ | _0376_;
assign _0851_ = _0380_ | _0655_;
assign addr_update_t0 = _0383_ | _0658_;
assign _0853_ = _0385_ | _0384_;
assign data_req_o_t0 = _0387_ | _0386_;
assign _0855_ = _0389_ | _0388_;
assign rdata_update_t0 = _0392_ | _0660_;
assign _0857_ = _0394_ | _0393_;
assign addr_incr_req_o_t0 = _0396_ | _0395_;
assign _0859_ = _0399_ | _0664_;
assign lsu_rdata_o_t0 = _0402_ | _0667_;
assign _0861_ = _0405_ | _0670_;
assign _0863_ = _0408_ | _0673_;
assign rdata_b_ext_t0 = _0411_ | _0676_;
assign _0865_ = _0414_ | _0677_;
assign _0867_ = _0417_ | _0678_;
assign rdata_h_ext_t0 = _0420_ | _0679_;
assign _0869_ = _0423_ | _0680_;
assign _0871_ = _0426_ | _0681_;
assign rdata_w_ext_t0 = _0429_ | _0682_;
assign _0873_ = _0432_ | _0685_;
assign _0875_ = _0435_ | _0688_;
assign data_wdata_t0 = _0438_ | _0691_;
assign _0076_ = _0441_ | _0694_;
assign _0069_ = _0444_ | _0695_;
assign _0042_ = _0446_ | _0696_;
assign _0024_ = _0447_ | _0696_;
assign _0886_ = _0450_ | _0699_;
assign data_be_o_t0 = _0453_ | _0702_;
assign _0081_ = _0485_ | _0484_;
assign _0038_ = _0487_ | _0486_;
assign _0074_ = _0488_ | _0047_;
assign _0079_ = _0490_ | _0489_;
assign _0067_ = _0492_ | _0491_;
assign _0072_ = _0494_ | _0493_;
assign _0059_ = _0496_ | _0495_;
assign _0055_ = _0498_ | _0497_;
assign _0061_ = _0501_ | _0722_;
assign _0021_ = _0503_ | _0502_;
assign _0045_ = _0504_ | _0489_;
assign _0028_ = _0507_ | _0723_;
assign _0008_ = _0510_ | _0726_;
assign _0001_ = _0512_ | _0511_;
assign _0013_ = _0514_ | _0513_;
assign _0011_ = _0515_ | _0513_;
assign _0015_ = _0517_ | _0516_;
assign perf_store_o_t0 = _0519_ | _0518_;
assign perf_load_o_t0 = _0521_ | _0520_;
assign _0063_ = _0526_ | _0730_;
assign _0051_ = _0529_ | _0731_;
assign _0034_ = _0532_ | _0732_;
assign _0017_ = _0535_ | _0733_;
assign _0065_ = _0538_ | _0734_;
assign _0053_ = _0541_ | _0735_;
assign _0036_ = _0544_ | _0736_;
assign _0019_ = _0547_ | _0737_;
assign _0057_ = _0551_ | _0550_;
assign _0003_ = _0554_ | _0740_;
assign addr_last_d_t0 = _0559_ | _0743_;
assign _0220_ = { _0894_, lsu_req_i, data_gnt_i } != 3'h6;
assign _0222_ = { _0918_, _0900_, data_gnt_i } != 3'h4;
assign _0224_ = { _0894_, lsu_req_i } != 2'h2;
assign _0226_ = { _0920_, _0899_ } != 2'h2;
assign _0228_ = { _0916_, _0899_ } != 2'h2;
assign _0230_ = | { _0918_, _0916_, _0894_, _0920_ };
assign _0232_ = { _0914_, data_rvalid_i } != 2'h2;
assign _0234_ = { _0918_, _0900_ } != 2'h2;
assign _0236_ = | { _0918_, _0914_, _0894_ };
assign _0238_ = & { _0220_, _0224_, _0226_, _0230_, _0228_, _0222_ };
assign _0240_ = & { _0232_, _0236_, _0234_ };
assign _0242_ = & { _0224_, _0232_, _0236_, _0234_ };
assign _0197_ = ~ _0856_;
assign _0198_ = ~ _0852_;
assign _0199_ = ~ ls_fsm_cs[1];
assign _0200_ = ~ ls_fsm_cs[2];
assign _0201_ = ~ _0068_[0];
assign _0244_ = | { _0920_, _0918_, _0916_ };
assign _0246_ = | { _0920_, _0916_ };
assign _0202_ = ~ _0930_;
assign _0203_ = ~ _0934_;
assign _0204_ = ~ data_bus_err_i;
assign _0205_ = ~ lsu_err_q;
assign _0206_ = ~ _0911_;
assign _0207_ = ~ _0928_;
assign _0208_ = ~ _0891_;
assign _0209_ = ~ busy_o;
assign _0326_ = _0919_ & _0170_;
assign _0329_ = _0931_ & _0207_;
assign _0332_ = _0935_ & _0208_;
assign _0472_ = data_bus_err_i_t0 & _0163_;
assign _0475_ = lsu_req_i_t0 & _0209_;
assign _0478_ = lsu_err_q_t0 & _0204_;
assign _0481_ = _0912_ & _0163_;
assign _0327_ = _0917_ & _0168_;
assign _0330_ = _0929_ & _0202_;
assign _0333_ = _0877_[3] & _0203_;
assign _0473_ = pmp_err_q_t0 & _0204_;
assign _0476_ = busy_o_t0 & _0193_;
assign _0479_ = data_bus_err_i_t0 & _0205_;
assign _0482_ = pmp_err_q_t0 & _0206_;
assign _0328_ = _0919_ & _0917_;
assign _0331_ = _0931_ & _0929_;
assign _0334_ = _0935_ & _0877_[3];
assign _0474_ = data_bus_err_i_t0 & pmp_err_q_t0;
assign _0477_ = lsu_req_i_t0 & busy_o_t0;
assign _0480_ = lsu_err_q_t0 & data_bus_err_i_t0;
assign _0483_ = _0912_ & pmp_err_q_t0;
assign _0619_ = _0326_ | _0327_;
assign _0620_ = _0329_ | _0330_;
assign _0621_ = _0332_ | _0333_;
assign _0708_ = _0472_ | _0473_;
assign _0709_ = _0475_ | _0476_;
assign _0710_ = _0478_ | _0479_;
assign _0711_ = _0481_ | _0482_;
assign _0561_ = _0619_ | _0328_;
assign _0563_ = _0620_ | _0331_;
assign _0565_ = _0621_ | _0334_;
assign _0905_ = _0708_ | _0474_;
assign _0910_ = _0709_ | _0477_;
assign _0912_ = _0710_ | _0480_;
assign data_or_pmp_err_t0 = _0711_ | _0483_;
assign _0210_ = | { _0918_, _0914_ };
assign _0212_ = | { _0918_, _0916_, _0914_ };
assign _0560_ = _0918_ | _0916_;
assign _0562_ = _0930_ | _0928_;
assign _0564_ = _0934_ | _0891_;
assign _0828_ = _0916_ ? _0078_ : _0060_;
assign _0830_ = _0914_ ? _0080_ : _0828_;
assign _0832_ = _0894_ ? _0007_ : 3'h0;
assign _0834_ = _0920_ ? _0044_ : _0832_;
assign ls_fsm_ns = _0212_ ? _0830_ : _0834_;
assign _0836_ = _0918_ ? _0029_ : _0009_;
assign lsu_err_d = _0914_ ? _0046_ : _0836_;
assign _0838_ = _0918_ ? _0031_ : _0014_;
assign pmp_err_d = _0914_ ? _0048_ : _0838_;
assign _0840_ = _0916_ ? _0077_ : _0058_;
assign _0842_ = _0920_ ? _0043_ : _0005_;
assign handle_misaligned_d = _0560_ ? _0840_ : _0842_;
assign ctrl_update = _0246_ ? _0039_ : _0844_;
assign _0846_ = _0916_ ? _0066_ : _0054_;
assign _0848_ = _0914_ ? _0073_ : _0846_;
assign _0844_ = _0894_ ? _0000_ : 1'h0;
assign _0850_ = _0920_ ? _0039_ : _0844_;
assign addr_update = _0212_ ? _0848_ : _0850_;
assign _0852_ = _0894_ ? _0004_ : 1'h0;
assign data_req_o = _0244_ ? 1'h1 : _0852_;
assign _0854_ = _0918_ ? _0020_ : 1'h0;
assign rdata_update = _0914_ ? _0037_ : _0854_;
assign _0856_ = _0916_ ? handle_misaligned_q : 1'h0;
assign addr_incr_req_o = _0210_ ? 1'h1 : _0856_;
assign _0858_ = _0926_ ? rdata_h_ext : rdata_w_ext;
assign lsu_rdata_o = _0924_ ? rdata_b_ext : _0858_;
assign _0860_ = _0928_ ? _0062_ : _0050_;
assign _0862_ = _0932_ ? _0033_ : _0016_;
assign rdata_b_ext = _0562_ ? _0860_ : _0862_;
assign _0864_ = _0928_ ? _0064_ : _0052_;
assign _0866_ = _0932_ ? _0035_ : _0018_;
assign rdata_h_ext = _0562_ ? _0864_ : _0866_;
assign _0868_ = _0928_ ? { data_rdata_i[23:0], rdata_q[31:24] } : { data_rdata_i[15:0], rdata_q[31:16] };
assign _0870_ = _0932_ ? { data_rdata_i[7:0], rdata_q } : data_rdata_i[31:0];
assign rdata_w_ext = _0562_ ? _0868_ : _0870_;
assign _0872_ = _0891_ ? { lsu_wdata_i[7:0], lsu_wdata_i[31:8] } : { lsu_wdata_i[15:0], lsu_wdata_i[31:16] };
assign _0874_ = _0936_ ? { lsu_wdata_i[23:0], lsu_wdata_i[31:24] } : lsu_wdata_i;
assign data_wdata = _0564_ ? _0872_ : _0874_;
assign _0876_ = _0891_ ? 4'h8 : 4'h4;
assign _0878_ = _0936_ ? 4'h2 : 4'h1;
assign _0075_ = _0564_ ? _0876_ : _0878_;
assign _0881_ = _0936_ ? 4'h6 : 4'h3;
assign _0068_ = _0564_ ? _0880_ : _0881_;
assign _0882_ = _0891_ ? 4'h7 : 4'h3;
assign _0883_ = _0936_ ? 4'h1 : 4'h0;
assign _0041_ = _0564_ ? _0882_ : _0883_;
assign _0880_ = _0891_ ? 4'h8 : 4'hc;
assign _0884_ = _0936_ ? 4'he : 4'hf;
assign _0023_ = _0564_ ? _0880_ : _0884_;
assign _0885_ = _0889_ ? _0056_ : _0002_;
assign data_be_o = _0939_ ? _0075_ : _0885_;
assign _0214_ = | { _0231_, _0229_, _0227_, _0225_, _0223_, _0221_ };
assign _0215_ = | { _0237_, _0235_, _0233_ };
assign _0216_ = | { _0237_, _0235_, _0233_, _0225_ };
assign _0616_ = { _0220_, _0224_, _0226_, _0230_, _0228_, _0222_ } | { _0221_, _0225_, _0227_, _0231_, _0229_, _0223_ };
assign _0617_ = { _0232_, _0236_, _0234_ } | { _0233_, _0237_, _0235_ };
assign _0618_ = { _0224_, _0232_, _0236_, _0234_ } | { _0225_, _0233_, _0237_, _0235_ };
assign _0217_ = & _0616_;
assign _0218_ = & _0617_;
assign _0219_ = & _0618_;
assign _0239_ = _0214_ & _0217_;
assign _0241_ = _0215_ & _0218_;
assign _0243_ = _0216_ & _0219_;
assign _0892_ = ! /* src = "generated/sv2v_out.v:18640.63-18640.80" */ ls_fsm_ns;
assign _0895_ = _0887_ && /* src = "generated/sv2v_out.v:18560.36-18560.83" */ _0902_;
assign _0897_ = _0889_ && /* src = "generated/sv2v_out.v:18560.89-18560.136" */ _0891_;
assign split_misaligned_access = _0895_ || /* src = "generated/sv2v_out.v:18560.35-18560.137" */ _0897_;
assign _0900_ = data_rvalid_i || /* src = "generated/sv2v_out.v:18604.9-18604.35" */ pmp_err_q;
assign _0899_ = data_gnt_i || /* src = "generated/sv2v_out.v:18620.9-18620.32" */ pmp_err_q;
assign _0902_ = | /* src = "generated/sv2v_out.v:18560.62-18560.82" */ adder_result_ex_i[1:0];
assign busy_o = | /* src = "generated/sv2v_out.v:18678.18-18678.35" */ ls_fsm_cs;
assign _0794_ = ~ /* src = "generated/sv2v_out.v:18580.20-18580.29" */ lsu_we_i;
assign _0904_ = ~ /* src = "generated/sv2v_out.v:18609.33-18609.62" */ _0908_;
assign _0906_ = ~ /* src = "generated/sv2v_out.v:18656.71-18656.87" */ data_or_pmp_err;
assign _0907_ = ~ /* src = "generated/sv2v_out.v:18656.105-18656.119" */ data_intg_err;
assign _0789_ = ~ /* src = "generated/sv2v_out.v:18676.66-18676.76" */ data_we_q;
assign _0908_ = data_bus_err_i | /* src = "generated/sv2v_out.v:18609.35-18609.61" */ pmp_err_q;
assign _0909_ = lsu_req_i | /* src = "generated/sv2v_out.v:18640.27-18640.58" */ busy_o;
assign _0911_ = lsu_err_q | /* src = "generated/sv2v_out.v:18654.28-18654.54" */ data_bus_err_i;
assign data_or_pmp_err = _0911_ | /* src = "generated/sv2v_out.v:18654.27-18654.67" */ pmp_err_q;
assign _0913_ = data_rvalid_i | /* src = "generated/sv2v_out.v:18655.29-18655.54" */ pmp_err_q;
/* src = "generated/sv2v_out.v:18641.2-18653.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_load_store_unit\MemECC=1'1\MemDataWidth=32'00000000000000000000000000100111  */
/* PC_TAINT_INFO STATE_NAME ls_fsm_cs */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) ls_fsm_cs <= 3'h0;
else ls_fsm_cs <= ls_fsm_ns;
assign _0080_ = data_rvalid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18629.9-18629.22|generated/sv2v_out.v:18629.5-18635.8" */ 3'h0 : ls_fsm_cs;
assign _0037_ = data_rvalid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18629.9-18629.22|generated/sv2v_out.v:18629.5-18635.8" */ _0789_ : 1'h0;
assign _0073_ = data_rvalid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18629.9-18629.22|generated/sv2v_out.v:18629.5-18635.8" */ _0204_ : 1'h0;
assign _0046_ = data_rvalid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18629.9-18629.22|generated/sv2v_out.v:18629.5-18635.8" */ data_bus_err_i : 1'hx;
assign _0048_ = data_rvalid_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18629.9-18629.22|generated/sv2v_out.v:18629.5-18635.8" */ data_pmp_err_i : 1'hx;
assign _0077_ = _0899_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18620.9-18620.32|generated/sv2v_out.v:18620.5-18625.8" */ 1'h0 : 1'hx;
assign _0078_ = _0899_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18620.9-18620.32|generated/sv2v_out.v:18620.5-18625.8" */ 3'h0 : ls_fsm_cs;
assign _0066_ = _0899_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18620.9-18620.32|generated/sv2v_out.v:18620.5-18625.8" */ _0205_ : 1'h0;
assign _0070_ = data_gnt_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18612.14-18612.24|generated/sv2v_out.v:18612.10-18615.8" */ 1'h0 : 1'hx;
assign _0071_ = data_gnt_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18612.14-18612.24|generated/sv2v_out.v:18612.10-18615.8" */ 3'h4 : ls_fsm_cs;
assign _0058_ = _0900_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18604.9-18604.35|generated/sv2v_out.v:18604.5-18615.8" */ _0161_ : _0070_;
assign _0054_ = _0900_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18604.9-18604.35|generated/sv2v_out.v:18604.5-18615.8" */ _0082_ : 1'h0;
assign _0060_ = _0900_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18604.9-18604.35|generated/sv2v_out.v:18604.5-18615.8" */ _0943_ : _0071_;
assign _0020_ = _0900_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18604.9-18604.35|generated/sv2v_out.v:18604.5-18615.8" */ _0789_ : 1'h0;
assign _0029_ = _0900_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18604.9-18604.35|generated/sv2v_out.v:18604.5-18615.8" */ _0908_ : 1'hx;
assign _0031_ = _0900_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18604.9-18604.35|generated/sv2v_out.v:18604.5-18615.8" */ data_pmp_err_i : 1'hx;
assign _0044_ = _0899_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18594.9-18594.32|generated/sv2v_out.v:18594.5-18599.8" */ 3'h2 : ls_fsm_cs;
assign _0043_ = _0899_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18594.9-18594.32|generated/sv2v_out.v:18594.5-18599.8" */ 1'h1 : 1'hx;
assign _0039_ = _0899_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18594.9-18594.32|generated/sv2v_out.v:18594.5-18599.8" */ 1'h1 : 1'h0;
assign _0027_ = data_gnt_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18582.10-18582.20|generated/sv2v_out.v:18582.6-18589.59" */ _0941_ : _0942_;
assign _0025_ = data_gnt_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18582.10-18582.20|generated/sv2v_out.v:18582.6-18589.59" */ split_misaligned_access : 1'hx;
assign _0022_ = data_gnt_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18582.10-18582.20|generated/sv2v_out.v:18582.6-18589.59" */ 1'h1 : 1'h0;
assign _0007_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18576.9-18576.18|generated/sv2v_out.v:18576.5-18590.8" */ _0027_ : ls_fsm_cs;
assign _0005_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18576.9-18576.18|generated/sv2v_out.v:18576.5-18590.8" */ _0025_ : 1'hx;
assign _0000_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18576.9-18576.18|generated/sv2v_out.v:18576.5-18590.8" */ _0022_ : 1'h0;
assign _0012_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18576.9-18576.18|generated/sv2v_out.v:18576.5-18590.8" */ lsu_we_i : 1'h0;
assign _0010_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18576.9-18576.18|generated/sv2v_out.v:18576.5-18590.8" */ _0794_ : 1'h0;
assign _0009_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18576.9-18576.18|generated/sv2v_out.v:18576.5-18590.8" */ 1'h0 : 1'hx;
assign _0014_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18576.9-18576.18|generated/sv2v_out.v:18576.5-18590.8" */ data_pmp_err_i : 1'h0;
assign _0004_ = lsu_req_i ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18576.9-18576.18|generated/sv2v_out.v:18576.5-18590.8" */ 1'h1 : 1'h0;
assign perf_store_o = _0894_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18573.3-18638.10" */ _0012_ : 1'h0;
assign perf_load_o = _0894_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18573.3-18638.10" */ _0010_ : 1'h0;
assign _0920_ = ls_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18573.3-18638.10" */ 3'h1;
assign _0894_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18573.3-18638.10" */ ls_fsm_cs;
assign _0914_ = ls_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18573.3-18638.10" */ 3'h4;
assign _0916_ = ls_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18573.3-18638.10" */ 3'h3;
assign _0918_ = ls_fsm_cs == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18573.3-18638.10" */ 3'h2;
assign _0924_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18536.3-18541.10" */ _0922_;
assign _0922_[0] = data_type_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18536.3-18541.10" */ 2'h2;
assign _0922_[1] = data_type_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18536.3-18541.10" */ 2'h3;
assign _0926_ = data_type_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18536.3-18541.10" */ 2'h1;
assign _0062_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18529.9-18529.25|generated/sv2v_out.v:18529.5-18532.67" */ { data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31:24] } : { 24'h000000, data_rdata_i[31:24] };
assign _0050_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18524.9-18524.25|generated/sv2v_out.v:18524.5-18527.67" */ { data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23:16] } : { 24'h000000, data_rdata_i[23:16] };
assign _0033_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18519.9-18519.25|generated/sv2v_out.v:18519.5-18522.66" */ { data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15:8] } : { 24'h000000, data_rdata_i[15:8] };
assign _0016_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18514.9-18514.25|generated/sv2v_out.v:18514.5-18517.64" */ { data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7:0] } : { 24'h000000, data_rdata_i[7:0] };
assign _0064_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18505.9-18505.25|generated/sv2v_out.v:18505.5-18508.80" */ { data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7], data_rdata_i[7:0], rdata_q[31:24] } : { 16'h0000, data_rdata_i[7:0], rdata_q[31:24] };
assign _0052_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18500.9-18500.25|generated/sv2v_out.v:18500.5-18503.67" */ { data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31], data_rdata_i[31:16] } : { 16'h0000, data_rdata_i[31:16] };
assign _0035_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18495.9-18495.25|generated/sv2v_out.v:18495.5-18498.66" */ { data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23], data_rdata_i[23:8] } : { 16'h0000, data_rdata_i[23:8] };
assign _0018_ = data_sign_ext_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18490.9-18490.25|generated/sv2v_out.v:18490.5-18493.66" */ { data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15], data_rdata_i[15:0] } : { 16'h0000, data_rdata_i[15:0] };
assign _0928_ = rdata_offset_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18480.3-18486.10" */ 2'h3;
assign _0930_ = rdata_offset_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18480.3-18486.10" */ 2'h2;
assign _0932_ = rdata_offset_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18480.3-18486.10" */ 2'h1;
assign _0939_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18408.3-18446.10" */ _0937_;
assign _0056_ = handle_misaligned_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18427.9-18427.29|generated/sv2v_out.v:18427.5-18436.24" */ 4'h1 : _0068_;
assign _0891_ = adder_result_ex_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18411.6-18417.13" */ 2'h3;
assign _0934_ = adder_result_ex_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18411.6-18417.13" */ 2'h2;
assign _0936_ = adder_result_ex_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18411.6-18417.13" */ 2'h1;
assign _0002_ = handle_misaligned_q ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:18410.9-18410.29|generated/sv2v_out.v:18410.5-18425.13" */ _0041_ : _0023_;
assign _0937_[0] = lsu_type_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18408.3-18446.10" */ 2'h2;
assign _0937_[1] = lsu_type_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18408.3-18446.10" */ 2'h3;
assign _0889_ = lsu_type_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18408.3-18446.10" */ 2'h1;
assign _0887_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:18408.3-18446.10" */ lsu_type_i;
assign data_intg_err = | /* src = "generated/sv2v_out.v:18554.27-18554.35" */ \g_mem_rdata_ecc.ecc_err ;
assign addr_last_d = addr_incr_req_o ? /* src = "generated/sv2v_out.v:18473.24-18473.73" */ { adder_result_ex_i[31:2], 2'h0 } : adder_result_ex_i;
assign _0941_ = split_misaligned_access ? /* src = "generated/sv2v_out.v:18586.20-18586.57" */ 3'h2 : 3'h0;
assign _0942_ = split_misaligned_access ? /* src = "generated/sv2v_out.v:18589.20-18589.57" */ 3'h1 : 3'h3;
assign _0943_ = data_gnt_i ? /* src = "generated/sv2v_out.v:18608.19-18608.43" */ 3'h0 : 3'h3;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18550.30-18553.5" */
prim_secded_inv_39_32_dec \g_mem_rdata_ecc.u_data_intg_dec  (
.data_i(\g_mem_rdata_ecc.data_rdata_buf ),
.data_i_t0(\g_mem_rdata_ecc.data_rdata_buf_t0 ),
.err_o(\g_mem_rdata_ecc.ecc_err ),
.err_o_t0(\g_mem_rdata_ecc.ecc_err_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18546.37-18549.5" */
\$paramod\prim_buf\Width=32'00000000000000000000000000100111  \g_mem_rdata_ecc.u_prim_buf_instr_rdata  (
.in_i(data_rdata_i),
.in_i_t0(data_rdata_i_t0),
.out_o(\g_mem_rdata_ecc.data_rdata_buf ),
.out_o_t0(\g_mem_rdata_ecc.data_rdata_buf_t0 )
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:18664.30-18667.5" */
prim_secded_inv_39_32_enc \g_mem_wdata_ecc.u_data_gen  (
.data_i(data_wdata),
.data_i_t0(data_wdata_t0),
.data_o(data_wdata_o),
.data_o_t0(data_wdata_o_t0)
);
assign _0877_[2:0] = { _0877_[3], 2'h0 };
assign { _0879_[3:2], _0879_[0] } = { 2'h0, _0879_[1] };
assign data_addr_o = { adder_result_ex_i[31:2], 2'h0 };
assign data_addr_o_t0 = { adder_result_ex_i_t0[31:2], 2'h0 };
assign data_we_o = lsu_we_i;
assign data_we_o_t0 = lsu_we_i_t0;
endmodule

module \$paramod\ibex_prefetch_buffer\ResetAll=1'1 (clk_i, rst_ni, req_i, branch_i, addr_i, ready_i, valid_o, rdata_o, addr_o, err_o, err_plus2_o, instr_req_o, instr_gnt_i, instr_addr_o, instr_rdata_i, instr_err_i, instr_rvalid_i, busy_o, valid_o_t0, req_i_t0, ready_i_t0
, rdata_o_t0, instr_rvalid_i_t0, instr_req_o_t0, instr_rdata_i_t0, instr_gnt_i_t0, instr_err_i_t0, instr_addr_o_t0, err_plus2_o_t0, branch_i_t0, addr_o_t0, addr_i_t0, busy_o_t0, err_o_t0);
/* src = "generated/sv2v_out.v:19959.26-19959.57" */
wire _000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19959.26-19959.57" */
wire _001_;
/* src = "generated/sv2v_out.v:19963.27-19963.55" */
wire _002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19963.27-19963.55" */
wire _003_;
/* src = "generated/sv2v_out.v:20000.38-20000.61" */
wire _004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20000.38-20000.61" */
wire _005_;
/* src = "generated/sv2v_out.v:20001.36-20001.77" */
wire _006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20001.36-20001.77" */
wire _007_;
/* src = "generated/sv2v_out.v:20001.82-20001.115" */
wire _008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20001.82-20001.115" */
wire _009_;
/* src = "generated/sv2v_out.v:20004.38-20004.92" */
wire _010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20004.38-20004.92" */
wire _011_;
/* src = "generated/sv2v_out.v:20005.36-20005.108" */
wire _012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20005.36-20005.108" */
wire _013_;
/* src = "generated/sv2v_out.v:20005.113-20005.146" */
wire _014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20005.113-20005.146" */
wire _015_;
wire [31:0] _016_;
wire [31:0] _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire [1:0] _022_;
wire _023_;
wire [31:0] _024_;
wire [31:0] _025_;
wire [1:0] _026_;
wire _027_;
wire _028_;
wire [1:0] _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire [1:0] _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
/* cellift = 32'd1 */
wire _054_;
wire [31:0] _055_;
wire [31:0] _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire [31:0] _094_;
wire [31:0] _095_;
wire [31:0] _096_;
wire [1:0] _097_;
wire [1:0] _098_;
wire [1:0] _099_;
wire [29:0] _100_;
wire [29:0] _101_;
wire [29:0] _102_;
wire _103_;
wire _104_;
wire _105_;
wire [1:0] _106_;
wire [1:0] _107_;
wire [1:0] _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire [1:0] _136_;
wire [31:0] _137_;
wire [31:0] _138_;
wire [31:0] _139_;
wire [31:0] _140_;
wire [31:0] _141_;
wire [31:0] _142_;
wire [31:0] _143_;
wire [31:0] _144_;
wire [1:0] _145_;
wire [1:0] _146_;
wire [1:0] _147_;
wire [1:0] _148_;
wire [1:0] _149_;
wire [1:0] _150_;
wire [31:0] _151_;
wire [31:0] _152_;
wire [31:0] _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire [31:0] _167_;
wire [31:0] _168_;
wire [31:0] _169_;
wire [31:0] _170_;
wire [1:0] _171_;
wire [1:0] _172_;
wire [1:0] _173_;
wire [1:0] _174_;
wire [29:0] _175_;
wire [29:0] _176_;
wire [29:0] _177_;
wire [29:0] _178_;
wire [1:0] _179_;
wire _180_;
wire [1:0] _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire [1:0] _192_;
wire [31:0] _193_;
wire [31:0] _194_;
wire [31:0] _195_;
wire [31:0] _196_;
wire [31:0] _197_;
wire [31:0] _198_;
wire [31:0] _199_;
wire [1:0] _200_;
wire [1:0] _201_;
wire [1:0] _202_;
wire [1:0] _203_;
wire [31:0] _204_;
wire [31:0] _205_;
wire [1:0] _206_;
wire [29:0] _207_;
wire [31:0] _208_;
wire [31:0] _209_;
wire [31:0] _210_;
wire [1:0] _211_;
wire [1:0] _212_;
wire [31:0] _213_;
wire [31:0] _214_;
/* src = "generated/sv2v_out.v:19961.35-19961.47" */
wire _215_;
/* src = "generated/sv2v_out.v:19939.25-19939.58" */
wire [1:0] _216_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19939.25-19939.58" */
wire [1:0] _217_;
/* src = "generated/sv2v_out.v:19959.35-19959.56" */
wire _218_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19959.35-19959.56" */
wire _219_;
/* src = "generated/sv2v_out.v:19962.40-19962.64" */
wire _220_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19962.40-19962.64" */
wire _221_;
/* src = "generated/sv2v_out.v:20001.35-20001.116" */
wire _222_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20001.35-20001.116" */
wire _223_;
/* src = "generated/sv2v_out.v:20005.35-20005.147" */
wire _224_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20005.35-20005.147" */
wire _225_;
/* src = "generated/sv2v_out.v:19931.18-19931.38" */
wire _226_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19931.18-19931.38" */
wire _227_;
/* src = "generated/sv2v_out.v:19980.25-19980.72" */
wire [31:0] _228_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19980.25-19980.72" */
wire [31:0] _229_;
/* src = "generated/sv2v_out.v:19995.54-19995.86" */
wire [31:0] _230_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19995.54-19995.86" */
wire [31:0] _231_;
/* src = "generated/sv2v_out.v:19890.20-19890.26" */
input [31:0] addr_i;
wire [31:0] addr_i;
/* cellift = 32'd1 */
input [31:0] addr_i_t0;
wire [31:0] addr_i_t0;
/* src = "generated/sv2v_out.v:19894.21-19894.27" */
output [31:0] addr_o;
wire [31:0] addr_o;
/* cellift = 32'd1 */
output [31:0] addr_o_t0;
wire [31:0] addr_o_t0;
/* src = "generated/sv2v_out.v:19914.13-19914.29" */
wire [1:0] branch_discard_n;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19914.13-19914.29" */
wire [1:0] branch_discard_n_t0;
/* src = "generated/sv2v_out.v:19916.12-19916.28" */
reg [1:0] branch_discard_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19916.12-19916.28" */
reg [1:0] branch_discard_q_t0;
/* src = "generated/sv2v_out.v:19915.13-19915.29" */
wire [1:0] branch_discard_s;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19915.13-19915.29" */
wire [1:0] branch_discard_s_t0;
/* src = "generated/sv2v_out.v:19889.13-19889.21" */
input branch_i;
wire branch_i;
/* cellift = 32'd1 */
input branch_i_t0;
wire branch_i_t0;
/* src = "generated/sv2v_out.v:19903.14-19903.20" */
output busy_o;
wire busy_o;
/* cellift = 32'd1 */
output busy_o_t0;
wire busy_o_t0;
/* src = "generated/sv2v_out.v:19886.13-19886.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:19909.7-19909.20" */
wire discard_req_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19909.7-19909.20" */
wire discard_req_d_t0;
/* src = "generated/sv2v_out.v:19910.6-19910.19" */
reg discard_req_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19910.6-19910.19" */
reg discard_req_q_t0;
/* src = "generated/sv2v_out.v:19895.14-19895.19" */
output err_o;
wire err_o;
/* cellift = 32'd1 */
output err_o_t0;
wire err_o_t0;
/* src = "generated/sv2v_out.v:19896.14-19896.25" */
output err_plus2_o;
wire err_plus2_o;
/* cellift = 32'd1 */
output err_plus2_o_t0;
wire err_plus2_o_t0;
/* src = "generated/sv2v_out.v:19921.14-19921.26" */
wire [31:0] fetch_addr_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19921.14-19921.26" */
wire [31:0] fetch_addr_d_t0;
/* src = "generated/sv2v_out.v:19923.7-19923.20" */
wire fetch_addr_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19923.7-19923.20" */
wire fetch_addr_en_t0;
/* src = "generated/sv2v_out.v:19922.13-19922.25" */
reg [31:0] fetch_addr_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19922.13-19922.25" */
reg [31:0] fetch_addr_q_t0;
/* src = "generated/sv2v_out.v:19930.13-19930.22" */
wire [1:0] fifo_busy;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19930.13-19930.22" */
wire [1:0] fifo_busy_t0;
/* src = "generated/sv2v_out.v:19928.7-19928.17" */
wire fifo_ready;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19928.7-19928.17" */
wire fifo_ready_t0;
/* src = "generated/sv2v_out.v:19926.7-19926.17" */
wire fifo_valid;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19926.7-19926.17" */
wire fifo_valid_t0;
/* src = "generated/sv2v_out.v:19924.14-19924.24" */
/* unused_bits = "0 1" */
wire [31:0] instr_addr;
/* src = "generated/sv2v_out.v:19899.21-19899.33" */
output [31:0] instr_addr_o;
wire [31:0] instr_addr_o;
/* cellift = 32'd1 */
output [31:0] instr_addr_o_t0;
wire [31:0] instr_addr_o_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19924.14-19924.24" */
/* unused_bits = "0 1" */
wire [31:0] instr_addr_t0;
/* src = "generated/sv2v_out.v:19901.13-19901.24" */
input instr_err_i;
wire instr_err_i;
/* cellift = 32'd1 */
input instr_err_i_t0;
wire instr_err_i_t0;
/* src = "generated/sv2v_out.v:19898.13-19898.24" */
input instr_gnt_i;
wire instr_gnt_i;
/* cellift = 32'd1 */
input instr_gnt_i_t0;
wire instr_gnt_i_t0;
/* src = "generated/sv2v_out.v:19900.20-19900.33" */
input [31:0] instr_rdata_i;
wire [31:0] instr_rdata_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_i_t0;
wire [31:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:19897.14-19897.25" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:19902.13-19902.27" */
input instr_rvalid_i;
wire instr_rvalid_i;
/* cellift = 32'd1 */
input instr_rvalid_i_t0;
wire instr_rvalid_i_t0;
/* src = "generated/sv2v_out.v:19893.21-19893.28" */
output [31:0] rdata_o;
wire [31:0] rdata_o;
/* cellift = 32'd1 */
output [31:0] rdata_o_t0;
wire [31:0] rdata_o_t0;
/* src = "generated/sv2v_out.v:19911.13-19911.32" */
wire [1:0] rdata_outstanding_n;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19911.13-19911.32" */
wire [1:0] rdata_outstanding_n_t0;
/* src = "generated/sv2v_out.v:19913.12-19913.31" */
reg [1:0] rdata_outstanding_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19913.12-19913.31" */
reg [1:0] rdata_outstanding_q_t0;
/* src = "generated/sv2v_out.v:19912.13-19912.32" */
wire [1:0] rdata_outstanding_s;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19912.13-19912.32" */
wire [1:0] rdata_outstanding_s_t0;
/* src = "generated/sv2v_out.v:19891.13-19891.20" */
input ready_i;
wire ready_i;
/* cellift = 32'd1 */
input ready_i_t0;
wire ready_i_t0;
/* src = "generated/sv2v_out.v:19888.13-19888.18" */
input req_i;
wire req_i;
/* cellift = 32'd1 */
input req_i_t0;
wire req_i_t0;
/* src = "generated/sv2v_out.v:19887.13-19887.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:19920.7-19920.21" */
wire stored_addr_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19920.7-19920.21" */
wire stored_addr_en_t0;
/* src = "generated/sv2v_out.v:19919.13-19919.26" */
reg [31:0] stored_addr_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19919.13-19919.26" */
reg [31:0] stored_addr_q_t0;
/* src = "generated/sv2v_out.v:19905.7-19905.20" */
wire valid_new_req;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19905.7-19905.20" */
wire valid_new_req_t0;
/* src = "generated/sv2v_out.v:19892.14-19892.21" */
output valid_o;
wire valid_o;
/* cellift = 32'd1 */
output valid_o_t0;
wire valid_o_t0;
/* src = "generated/sv2v_out.v:19907.7-19907.18" */
wire valid_req_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19907.7-19907.18" */
wire valid_req_d_t0;
/* src = "generated/sv2v_out.v:19908.6-19908.17" */
reg valid_req_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19908.6-19908.17" */
reg valid_req_q_t0;
assign fetch_addr_d = _228_ + /* src = "generated/sv2v_out.v:19980.24-19980.126" */ { 29'h00000000, _002_, 2'h0 };
assign _000_ = req_i & /* src = "generated/sv2v_out.v:19959.26-19959.57" */ _218_;
assign valid_new_req = _000_ & /* src = "generated/sv2v_out.v:19959.25-19959.84" */ _046_;
assign valid_req_d = instr_req_o & /* src = "generated/sv2v_out.v:19961.23-19961.47" */ _215_;
assign discard_req_d = valid_req_q & /* src = "generated/sv2v_out.v:19962.25-19962.65" */ _220_;
assign stored_addr_en = _002_ & /* src = "generated/sv2v_out.v:19963.26-19963.71" */ _215_;
assign _002_ = valid_new_req & /* src = "generated/sv2v_out.v:19980.90-19980.118" */ _027_;
assign _008_ = branch_i & /* src = "generated/sv2v_out.v:20001.82-20001.115" */ rdata_outstanding_q[0];
assign _010_ = _004_ & /* src = "generated/sv2v_out.v:20004.38-20004.92" */ rdata_outstanding_q[0];
assign _004_ = instr_req_o & /* src = "generated/sv2v_out.v:20005.38-20005.61" */ instr_gnt_i;
assign _006_ = _004_ & /* src = "generated/sv2v_out.v:20005.37-20005.78" */ discard_req_d;
assign _012_ = _006_ & /* src = "generated/sv2v_out.v:20005.36-20005.108" */ rdata_outstanding_q[0];
assign _014_ = branch_i & /* src = "generated/sv2v_out.v:20005.113-20005.146" */ rdata_outstanding_q[1];
assign fifo_valid = instr_rvalid_i & /* src = "generated/sv2v_out.v:20011.22-20011.59" */ _045_;
assign _016_ = ~ _229_;
assign _017_ = ~ { 29'h00000000, _003_, 2'h0 };
assign _055_ = _228_ & _016_;
assign _056_ = { 29'h00000000, _002_, 2'h0 } & _017_;
assign _213_ = _055_ + _056_;
assign _151_ = _228_ | _229_;
assign _152_ = { 29'h00000000, _002_, 2'h0 } | { 29'h00000000, _003_, 2'h0 };
assign _214_ = _151_ + _152_;
assign _204_ = _213_ ^ _214_;
assign _153_ = _204_ | _229_;
assign fetch_addr_d_t0 = _153_ | { 29'h00000000, _003_, 2'h0 };
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME valid_req_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) valid_req_q_t0 <= 1'h0;
else valid_req_q_t0 <= valid_req_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME discard_req_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) discard_req_q_t0 <= 1'h0;
else discard_req_q_t0 <= discard_req_d_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_outstanding_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_outstanding_q_t0 <= 2'h0;
else rdata_outstanding_q_t0 <= rdata_outstanding_s_t0;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME branch_discard_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_discard_q_t0 <= 2'h0;
else branch_discard_q_t0 <= branch_discard_s_t0;
assign _018_ = ~ fetch_addr_en;
assign _019_ = ~ _053_;
assign _020_ = ~ stored_addr_en;
assign _205_ = fetch_addr_d ^ fetch_addr_q;
assign _206_ = _230_[1:0] ^ stored_addr_q[1:0];
assign _207_ = instr_addr[31:2] ^ stored_addr_q[31:2];
assign _167_ = fetch_addr_d_t0 | fetch_addr_q_t0;
assign _171_ = _231_[1:0] | stored_addr_q_t0[1:0];
assign _175_ = instr_addr_t0[31:2] | stored_addr_q_t0[31:2];
assign _168_ = _205_ | _167_;
assign _172_ = _206_ | _171_;
assign _176_ = _207_ | _175_;
assign _094_ = { fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en, fetch_addr_en } & fetch_addr_d_t0;
assign _097_ = { _053_, _053_ } & _231_[1:0];
assign _100_ = { stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en, stored_addr_en } & instr_addr_t0[31:2];
assign _095_ = { _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_, _018_ } & fetch_addr_q_t0;
assign _098_ = { _019_, _019_ } & stored_addr_q_t0[1:0];
assign _101_ = { _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_, _020_ } & stored_addr_q_t0[31:2];
assign _096_ = _168_ & { fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0, fetch_addr_en_t0 };
assign _099_ = _172_ & { _054_, _054_ };
assign _102_ = _176_ & { stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0, stored_addr_en_t0 };
assign _169_ = _094_ | _095_;
assign _173_ = _097_ | _098_;
assign _177_ = _100_ | _101_;
assign _170_ = _169_ | _096_;
assign _174_ = _173_ | _099_;
assign _178_ = _177_ | _102_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME fetch_addr_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) fetch_addr_q_t0 <= 32'd0;
else fetch_addr_q_t0 <= _170_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME stored_addr_q_t0[1:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) stored_addr_q_t0[1:0] <= 2'h0;
else stored_addr_q_t0[1:0] <= _174_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME stored_addr_q_t0[31:2] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) stored_addr_q_t0[31:2] <= 30'h00000000;
else stored_addr_q_t0[31:2] <= _178_;
assign _057_ = req_i_t0 & _218_;
assign _060_ = _001_ & _046_;
assign _063_ = instr_req_o_t0 & _215_;
assign _066_ = valid_req_q_t0 & _220_;
assign _069_ = _003_ & _215_;
assign _072_ = valid_new_req_t0 & _027_;
assign _075_ = branch_i_t0 & rdata_outstanding_q[0];
assign _078_ = _005_ & rdata_outstanding_q[0];
assign _081_ = instr_req_o_t0 & instr_gnt_i;
assign _082_ = _005_ & discard_req_d;
assign _085_ = _007_ & rdata_outstanding_q[0];
assign _088_ = branch_i_t0 & rdata_outstanding_q[1];
assign _091_ = instr_rvalid_i_t0 & _045_;
assign _058_ = _219_ & req_i;
assign _061_ = rdata_outstanding_q_t0[1] & _000_;
assign _064_ = instr_gnt_i_t0 & instr_req_o;
assign _067_ = _221_ & valid_req_q;
assign _070_ = instr_gnt_i_t0 & _002_;
assign _073_ = valid_req_q_t0 & valid_new_req;
assign _076_ = rdata_outstanding_q_t0[0] & branch_i;
assign _079_ = rdata_outstanding_q_t0[0] & _004_;
assign _083_ = discard_req_d_t0 & _004_;
assign _086_ = rdata_outstanding_q_t0[0] & _006_;
assign _089_ = rdata_outstanding_q_t0[1] & branch_i;
assign _092_ = branch_discard_q_t0[0] & instr_rvalid_i;
assign _059_ = req_i_t0 & _219_;
assign _062_ = _001_ & rdata_outstanding_q_t0[1];
assign _065_ = instr_req_o_t0 & instr_gnt_i_t0;
assign _068_ = valid_req_q_t0 & _221_;
assign _071_ = _003_ & instr_gnt_i_t0;
assign _074_ = valid_new_req_t0 & valid_req_q_t0;
assign _077_ = branch_i_t0 & rdata_outstanding_q_t0[0];
assign _080_ = _005_ & rdata_outstanding_q_t0[0];
assign _084_ = _005_ & discard_req_d_t0;
assign _087_ = _007_ & rdata_outstanding_q_t0[0];
assign _090_ = branch_i_t0 & rdata_outstanding_q_t0[1];
assign _093_ = instr_rvalid_i_t0 & branch_discard_q_t0[0];
assign _154_ = _057_ | _058_;
assign _155_ = _060_ | _061_;
assign _156_ = _063_ | _064_;
assign _157_ = _066_ | _067_;
assign _158_ = _069_ | _070_;
assign _159_ = _072_ | _073_;
assign _160_ = _075_ | _076_;
assign _161_ = _078_ | _079_;
assign _162_ = _081_ | _064_;
assign _163_ = _082_ | _083_;
assign _164_ = _085_ | _086_;
assign _165_ = _088_ | _089_;
assign _166_ = _091_ | _092_;
assign _001_ = _154_ | _059_;
assign valid_new_req_t0 = _155_ | _062_;
assign valid_req_d_t0 = _156_ | _065_;
assign discard_req_d_t0 = _157_ | _068_;
assign stored_addr_en_t0 = _158_ | _071_;
assign _003_ = _159_ | _074_;
assign _009_ = _160_ | _077_;
assign _011_ = _161_ | _080_;
assign _005_ = _162_ | _065_;
assign _007_ = _163_ | _084_;
assign _013_ = _164_ | _087_;
assign _015_ = _165_ | _090_;
assign fifo_valid_t0 = _166_ | _093_;
/* src = "generated/sv2v_out.v:19983.4-19987.35" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME fetch_addr_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) fetch_addr_q <= 32'd0;
else if (fetch_addr_en) fetch_addr_q <= fetch_addr_d;
/* src = "generated/sv2v_out.v:19967.4-19971.37" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME stored_addr_q[1:0] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) stored_addr_q[1:0] <= 2'h0;
else if (_053_) stored_addr_q[1:0] <= _230_[1:0];
/* src = "generated/sv2v_out.v:19967.4-19971.37" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME stored_addr_q[31:2] */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) stored_addr_q[31:2] <= 30'h00000000;
else if (stored_addr_en) stored_addr_q[31:2] <= instr_addr[31:2];
assign _021_ = | rdata_outstanding_q_t0;
assign _022_ = ~ rdata_outstanding_q_t0;
assign _136_ = rdata_outstanding_q & _022_;
assign _023_ = ! _136_;
assign _227_ = _023_ & _021_;
assign _024_ = ~ { branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i };
assign _025_ = ~ { valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q };
assign _026_ = ~ { instr_rvalid_i, instr_rvalid_i };
assign _193_ = { branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0 } | _024_;
assign _197_ = { valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0 } | _025_;
assign _200_ = { instr_rvalid_i_t0, instr_rvalid_i_t0 } | _026_;
assign _194_ = { branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0 } | { branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i, branch_i };
assign _198_ = { valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0 } | { valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q, valid_req_q };
assign _201_ = { instr_rvalid_i_t0, instr_rvalid_i_t0 } | { instr_rvalid_i, instr_rvalid_i };
assign _137_ = { fetch_addr_q_t0[31:2], 2'h0 } & _193_;
assign _140_ = fetch_addr_q_t0 & _193_;
assign _142_ = _231_ & _197_;
assign _145_ = rdata_outstanding_n_t0 & _200_;
assign _148_ = branch_discard_n_t0 & _200_;
assign _138_ = addr_i_t0 & _194_;
assign _143_ = stored_addr_q_t0 & _198_;
assign _146_ = { 1'h0, rdata_outstanding_n_t0[1] } & _201_;
assign _149_ = { 1'h0, branch_discard_n_t0[1] } & _201_;
assign _195_ = _137_ | _138_;
assign _196_ = _140_ | _138_;
assign _199_ = _142_ | _143_;
assign _202_ = _145_ | _146_;
assign _203_ = _148_ | _149_;
assign _208_ = { fetch_addr_q[31:2], 2'h0 } ^ addr_i;
assign _209_ = fetch_addr_q ^ addr_i;
assign _210_ = _230_ ^ stored_addr_q;
assign _211_ = rdata_outstanding_n ^ { 1'h0, rdata_outstanding_n[1] };
assign _212_ = branch_discard_n ^ { 1'h0, branch_discard_n[1] };
assign _139_ = { branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0 } & _208_;
assign _141_ = { branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0, branch_i_t0 } & _209_;
assign _144_ = { valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0, valid_req_q_t0 } & _210_;
assign _147_ = { instr_rvalid_i_t0, instr_rvalid_i_t0 } & _211_;
assign _150_ = { instr_rvalid_i_t0, instr_rvalid_i_t0 } & _212_;
assign _229_ = _139_ | _195_;
assign _231_ = _141_ | _196_;
assign instr_addr_t0 = _144_ | _199_;
assign rdata_outstanding_s_t0 = _147_ | _202_;
assign branch_discard_s_t0 = _150_ | _203_;
assign _027_ = ~ valid_req_q;
assign _053_ = & { _027_, stored_addr_en };
assign _028_ = ~ _226_;
assign _029_ = ~ fifo_busy;
assign _031_ = ~ branch_i;
assign _032_ = ~ _004_;
assign _033_ = ~ _006_;
assign _034_ = ~ _222_;
assign _035_ = ~ _010_;
assign _036_ = ~ _012_;
assign _037_ = ~ _224_;
assign _038_ = ~ instr_req_o;
assign _039_ = ~ { rdata_outstanding_q[0], rdata_outstanding_q[1] };
assign _040_ = ~ valid_new_req;
assign _041_ = ~ discard_req_q;
assign _042_ = ~ _002_;
assign _043_ = ~ rdata_outstanding_q[0];
assign _044_ = ~ _008_;
assign _045_ = ~ branch_discard_q[0];
assign _046_ = ~ rdata_outstanding_q[1];
assign _047_ = ~ _014_;
assign _048_ = ~ branch_discard_q[1];
assign _103_ = _227_ & _038_;
assign _106_ = fifo_busy_t0 & _039_;
assign _109_ = fifo_ready_t0 & _031_;
assign _112_ = valid_req_q_t0 & _040_;
assign _113_ = branch_i_t0 & _041_;
assign _116_ = branch_i_t0 & _042_;
assign _119_ = _005_ & _043_;
assign _121_ = _007_ & _044_;
assign _124_ = _223_ & _045_;
assign _127_ = _011_ & _046_;
assign _130_ = _013_ & _047_;
assign _133_ = _225_ & _048_;
assign _104_ = instr_req_o_t0 & _028_;
assign _107_ = { rdata_outstanding_q_t0[0], rdata_outstanding_q_t0[1] } & _029_;
assign _110_ = branch_i_t0 & _030_;
assign _114_ = discard_req_q_t0 & _031_;
assign _117_ = _003_ & _031_;
assign _120_ = rdata_outstanding_q_t0[0] & _032_;
assign _122_ = _009_ & _033_;
assign _125_ = branch_discard_q_t0[0] & _034_;
assign _128_ = rdata_outstanding_q_t0[1] & _035_;
assign _131_ = _015_ & _036_;
assign _134_ = branch_discard_q_t0[1] & _037_;
assign _105_ = _227_ & instr_req_o_t0;
assign _108_ = fifo_busy_t0 & { rdata_outstanding_q_t0[0], rdata_outstanding_q_t0[1] };
assign _111_ = fifo_ready_t0 & branch_i_t0;
assign _115_ = branch_i_t0 & discard_req_q_t0;
assign _118_ = branch_i_t0 & _003_;
assign _123_ = _007_ & _009_;
assign _126_ = _223_ & branch_discard_q_t0[0];
assign _129_ = _011_ & rdata_outstanding_q_t0[1];
assign _132_ = _013_ & _015_;
assign _135_ = _225_ & branch_discard_q_t0[1];
assign _180_ = _103_ | _104_;
assign _181_ = _106_ | _107_;
assign _182_ = _109_ | _110_;
assign _183_ = _112_ | _072_;
assign _184_ = _113_ | _114_;
assign _185_ = _116_ | _117_;
assign _186_ = _119_ | _120_;
assign _187_ = _121_ | _122_;
assign _188_ = _124_ | _125_;
assign _189_ = _127_ | _128_;
assign _190_ = _130_ | _131_;
assign _191_ = _133_ | _134_;
assign busy_o_t0 = _180_ | _105_;
assign _217_ = _181_ | _108_;
assign _219_ = _182_ | _111_;
assign instr_req_o_t0 = _183_ | _074_;
assign _221_ = _184_ | _115_;
assign fetch_addr_en_t0 = _185_ | _118_;
assign rdata_outstanding_n_t0[0] = _186_ | _080_;
assign _223_ = _187_ | _123_;
assign branch_discard_n_t0[0] = _188_ | _126_;
assign rdata_outstanding_n_t0[1] = _189_ | _129_;
assign _225_ = _190_ | _132_;
assign branch_discard_n_t0[1] = _191_ | _135_;
assign _049_ = | { valid_req_q_t0, stored_addr_en_t0 };
assign _050_ = | _217_;
assign _179_ = { _027_, stored_addr_en } | { valid_req_q_t0, stored_addr_en_t0 };
assign _192_ = _216_ | _217_;
assign _051_ = & _179_;
assign _052_ = & _192_;
assign _054_ = _049_ & _051_;
assign fifo_ready_t0 = _050_ & _052_;
assign fifo_ready = ! /* src = "generated/sv2v_out.v:0.0-0.0" */ _030_;
assign _215_ = ~ /* src = "generated/sv2v_out.v:19963.59-19963.71" */ instr_gnt_i;
assign busy_o = _226_ | /* src = "generated/sv2v_out.v:19931.18-19931.52" */ instr_req_o;
assign _216_ = fifo_busy | /* src = "generated/sv2v_out.v:19939.25-19939.58" */ { rdata_outstanding_q[0], rdata_outstanding_q[1] };
assign _218_ = fifo_ready | /* src = "generated/sv2v_out.v:19959.35-19959.56" */ branch_i;
assign instr_req_o = valid_req_q | /* src = "generated/sv2v_out.v:19960.21-19960.48" */ valid_new_req;
assign _220_ = branch_i | /* src = "generated/sv2v_out.v:19962.40-19962.64" */ discard_req_q;
assign fetch_addr_en = branch_i | /* src = "generated/sv2v_out.v:19979.25-19979.66" */ _002_;
assign rdata_outstanding_n[0] = _004_ | /* src = "generated/sv2v_out.v:20000.37-20000.87" */ rdata_outstanding_q[0];
assign _222_ = _006_ | /* src = "generated/sv2v_out.v:20001.35-20001.116" */ _008_;
assign branch_discard_n[0] = _222_ | /* src = "generated/sv2v_out.v:20001.34-20001.139" */ branch_discard_q[0];
assign rdata_outstanding_n[1] = _010_ | /* src = "generated/sv2v_out.v:20004.37-20004.118" */ rdata_outstanding_q[1];
assign _224_ = _012_ | /* src = "generated/sv2v_out.v:20005.35-20005.147" */ _014_;
assign branch_discard_n[1] = _224_ | /* src = "generated/sv2v_out.v:20005.34-20005.170" */ branch_discard_q[1];
/* src = "generated/sv2v_out.v:20013.2-20025.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME valid_req_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) valid_req_q <= 1'h0;
else valid_req_q <= valid_req_d;
/* src = "generated/sv2v_out.v:20013.2-20025.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME discard_req_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) discard_req_q <= 1'h0;
else discard_req_q <= discard_req_d;
/* src = "generated/sv2v_out.v:20013.2-20025.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME rdata_outstanding_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) rdata_outstanding_q <= 2'h0;
else rdata_outstanding_q <= rdata_outstanding_s;
/* src = "generated/sv2v_out.v:20013.2-20025.6" */
/* PC_TAINT_INFO MODULE_NAME \$paramod\ibex_prefetch_buffer\ResetAll=1'1  */
/* PC_TAINT_INFO STATE_NAME branch_discard_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) branch_discard_q <= 2'h0;
else branch_discard_q <= branch_discard_s;
assign _030_ = & /* src = "generated/sv2v_out.v:19939.22-19939.59" */ _216_;
assign _226_ = | /* src = "generated/sv2v_out.v:19931.18-19931.38" */ rdata_outstanding_q;
assign _228_ = branch_i ? /* src = "generated/sv2v_out.v:19980.25-19980.72" */ addr_i : { fetch_addr_q[31:2], 2'h0 };
assign _230_ = branch_i ? /* src = "generated/sv2v_out.v:19995.54-19995.86" */ addr_i : fetch_addr_q;
assign instr_addr = valid_req_q ? /* src = "generated/sv2v_out.v:19995.23-19995.87" */ stored_addr_q : _230_;
assign rdata_outstanding_s = instr_rvalid_i ? /* src = "generated/sv2v_out.v:20009.32-20009.103" */ { 1'h0, rdata_outstanding_n[1] } : rdata_outstanding_n;
assign branch_discard_s = instr_rvalid_i ? /* src = "generated/sv2v_out.v:20010.29-20010.94" */ { 1'h0, branch_discard_n[1] } : branch_discard_n;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:19943.4-19958.3" */
\$paramod\ibex_fetch_fifo\NUM_REQS=32'00000000000000000000000000000010\ResetAll=1'1  fifo_i (
.busy_o(fifo_busy),
.busy_o_t0(fifo_busy_t0),
.clear_i(branch_i),
.clear_i_t0(branch_i_t0),
.clk_i(clk_i),
.in_addr_i(addr_i),
.in_addr_i_t0(addr_i_t0),
.in_err_i(instr_err_i),
.in_err_i_t0(instr_err_i_t0),
.in_rdata_i(instr_rdata_i),
.in_rdata_i_t0(instr_rdata_i_t0),
.in_valid_i(fifo_valid),
.in_valid_i_t0(fifo_valid_t0),
.out_addr_o(addr_o),
.out_addr_o_t0(addr_o_t0),
.out_err_o(err_o),
.out_err_o_t0(err_o_t0),
.out_err_plus2_o(err_plus2_o),
.out_err_plus2_o_t0(err_plus2_o_t0),
.out_rdata_o(rdata_o),
.out_rdata_o_t0(rdata_o_t0),
.out_ready_i(ready_i),
.out_ready_i_t0(ready_i_t0),
.out_valid_o(valid_o),
.out_valid_o_t0(valid_o_t0),
.rst_ni(rst_ni)
);
assign instr_addr_o = { instr_addr[31:2], 2'h0 };
assign instr_addr_o_t0 = { instr_addr_t0[31:2], 2'h0 };
endmodule

module \$paramod\ibex_wb_stage\ResetAll=1'1\WritebackStage=1'0\DummyInstructions=1'1 (clk_i, rst_ni, en_wb_i, instr_type_wb_i, pc_id_i, instr_is_compressed_id_i, instr_perf_count_id_i, ready_wb_o, rf_write_wb_o, outstanding_load_wb_o, outstanding_store_wb_o, pc_wb_o, perf_instr_ret_wb_o, perf_instr_ret_compressed_wb_o, perf_instr_ret_wb_spec_o, perf_instr_ret_compressed_wb_spec_o, rf_waddr_id_i, rf_wdata_id_i, rf_we_id_i, dummy_instr_id_i, rf_wdata_lsu_i
, rf_we_lsu_i, rf_wdata_fwd_wb_o, rf_waddr_wb_o, rf_wdata_wb_o, rf_we_wb_o, dummy_instr_wb_o, lsu_resp_valid_i, lsu_resp_err_i, instr_done_wb_o, pc_id_i_t0, lsu_resp_valid_i_t0, dummy_instr_id_i_t0, dummy_instr_wb_o_t0, en_wb_i_t0, instr_done_wb_o_t0, instr_is_compressed_id_i_t0, instr_perf_count_id_i_t0, instr_type_wb_i_t0, lsu_resp_err_i_t0, outstanding_load_wb_o_t0, outstanding_store_wb_o_t0
, pc_wb_o_t0, perf_instr_ret_compressed_wb_o_t0, perf_instr_ret_compressed_wb_spec_o_t0, perf_instr_ret_wb_o_t0, perf_instr_ret_wb_spec_o_t0, ready_wb_o_t0, rf_waddr_id_i_t0, rf_waddr_wb_o_t0, rf_wdata_fwd_wb_o_t0, rf_wdata_id_i_t0, rf_wdata_lsu_i_t0, rf_wdata_wb_o_t0, rf_we_id_i_t0, rf_we_lsu_i_t0, rf_we_wb_o_t0, rf_write_wb_o_t0);
/* src = "generated/sv2v_out.v:21045.34-21045.65" */
wire _00_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21045.34-21045.65" */
wire _01_;
/* src = "generated/sv2v_out.v:21045.71-21045.104" */
wire _02_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21045.71-21045.104" */
wire _03_;
/* src = "generated/sv2v_out.v:21067.26-21067.75" */
wire [31:0] _04_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21067.26-21067.75" */
wire [31:0] _05_;
/* src = "generated/sv2v_out.v:21067.80-21067.129" */
wire [31:0] _06_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:21067.80-21067.129" */
wire [31:0] _07_;
wire _08_;
wire [1:0] _09_;
wire _10_;
wire [31:0] _11_;
wire [31:0] _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire [31:0] _25_;
wire [31:0] _26_;
wire [31:0] _27_;
wire [31:0] _28_;
wire [31:0] _29_;
wire [31:0] _30_;
wire [31:0] _31_;
wire [31:0] _32_;
wire [31:0] _33_;
wire [1:0] _34_;
wire _35_;
wire _36_;
wire _37_;
wire _38_;
wire [31:0] _39_;
wire [31:0] _40_;
wire [31:0] _41_;
/* src = "generated/sv2v_out.v:21045.69-21045.105" */
wire _42_;
/* src = "generated/sv2v_out.v:20916.13-20916.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:20935.13-20935.29" */
input dummy_instr_id_i;
wire dummy_instr_id_i;
/* cellift = 32'd1 */
input dummy_instr_id_i_t0;
wire dummy_instr_id_i_t0;
/* src = "generated/sv2v_out.v:20942.14-20942.30" */
output dummy_instr_wb_o;
wire dummy_instr_wb_o;
/* cellift = 32'd1 */
output dummy_instr_wb_o_t0;
wire dummy_instr_wb_o_t0;
/* src = "generated/sv2v_out.v:20918.13-20918.20" */
input en_wb_i;
wire en_wb_i;
/* cellift = 32'd1 */
input en_wb_i_t0;
wire en_wb_i_t0;
/* src = "generated/sv2v_out.v:20945.14-20945.29" */
output instr_done_wb_o;
wire instr_done_wb_o;
/* cellift = 32'd1 */
output instr_done_wb_o_t0;
wire instr_done_wb_o_t0;
/* src = "generated/sv2v_out.v:20921.13-20921.37" */
input instr_is_compressed_id_i;
wire instr_is_compressed_id_i;
/* cellift = 32'd1 */
input instr_is_compressed_id_i_t0;
wire instr_is_compressed_id_i_t0;
/* src = "generated/sv2v_out.v:20922.13-20922.34" */
input instr_perf_count_id_i;
wire instr_perf_count_id_i;
/* cellift = 32'd1 */
input instr_perf_count_id_i_t0;
wire instr_perf_count_id_i_t0;
/* src = "generated/sv2v_out.v:20919.19-20919.34" */
input [1:0] instr_type_wb_i;
wire [1:0] instr_type_wb_i;
/* cellift = 32'd1 */
input [1:0] instr_type_wb_i_t0;
wire [1:0] instr_type_wb_i_t0;
/* src = "generated/sv2v_out.v:20944.13-20944.27" */
input lsu_resp_err_i;
wire lsu_resp_err_i;
/* cellift = 32'd1 */
input lsu_resp_err_i_t0;
wire lsu_resp_err_i_t0;
/* src = "generated/sv2v_out.v:20943.13-20943.29" */
input lsu_resp_valid_i;
wire lsu_resp_valid_i;
/* cellift = 32'd1 */
input lsu_resp_valid_i_t0;
wire lsu_resp_valid_i_t0;
/* src = "generated/sv2v_out.v:20925.14-20925.35" */
output outstanding_load_wb_o;
wire outstanding_load_wb_o;
/* cellift = 32'd1 */
output outstanding_load_wb_o_t0;
wire outstanding_load_wb_o_t0;
/* src = "generated/sv2v_out.v:20926.14-20926.36" */
output outstanding_store_wb_o;
wire outstanding_store_wb_o;
/* cellift = 32'd1 */
output outstanding_store_wb_o_t0;
wire outstanding_store_wb_o_t0;
/* src = "generated/sv2v_out.v:20920.20-20920.27" */
input [31:0] pc_id_i;
wire [31:0] pc_id_i;
/* cellift = 32'd1 */
input [31:0] pc_id_i_t0;
wire [31:0] pc_id_i_t0;
/* src = "generated/sv2v_out.v:20927.21-20927.28" */
output [31:0] pc_wb_o;
wire [31:0] pc_wb_o;
/* cellift = 32'd1 */
output [31:0] pc_wb_o_t0;
wire [31:0] pc_wb_o_t0;
/* src = "generated/sv2v_out.v:20929.14-20929.44" */
output perf_instr_ret_compressed_wb_o;
wire perf_instr_ret_compressed_wb_o;
/* cellift = 32'd1 */
output perf_instr_ret_compressed_wb_o_t0;
wire perf_instr_ret_compressed_wb_o_t0;
/* src = "generated/sv2v_out.v:20931.14-20931.49" */
output perf_instr_ret_compressed_wb_spec_o;
wire perf_instr_ret_compressed_wb_spec_o;
/* cellift = 32'd1 */
output perf_instr_ret_compressed_wb_spec_o_t0;
wire perf_instr_ret_compressed_wb_spec_o_t0;
/* src = "generated/sv2v_out.v:20928.14-20928.33" */
output perf_instr_ret_wb_o;
wire perf_instr_ret_wb_o;
/* cellift = 32'd1 */
output perf_instr_ret_wb_o_t0;
wire perf_instr_ret_wb_o_t0;
/* src = "generated/sv2v_out.v:20930.14-20930.38" */
output perf_instr_ret_wb_spec_o;
wire perf_instr_ret_wb_spec_o;
/* cellift = 32'd1 */
output perf_instr_ret_wb_spec_o_t0;
wire perf_instr_ret_wb_spec_o_t0;
/* src = "generated/sv2v_out.v:20923.14-20923.24" */
output ready_wb_o;
wire ready_wb_o;
/* cellift = 32'd1 */
output ready_wb_o_t0;
wire ready_wb_o_t0;
/* src = "generated/sv2v_out.v:20932.19-20932.32" */
input [4:0] rf_waddr_id_i;
wire [4:0] rf_waddr_id_i;
/* cellift = 32'd1 */
input [4:0] rf_waddr_id_i_t0;
wire [4:0] rf_waddr_id_i_t0;
/* src = "generated/sv2v_out.v:20939.20-20939.33" */
output [4:0] rf_waddr_wb_o;
wire [4:0] rf_waddr_wb_o;
/* cellift = 32'd1 */
output [4:0] rf_waddr_wb_o_t0;
wire [4:0] rf_waddr_wb_o_t0;
/* src = "generated/sv2v_out.v:20938.21-20938.38" */
output [31:0] rf_wdata_fwd_wb_o;
wire [31:0] rf_wdata_fwd_wb_o;
/* cellift = 32'd1 */
output [31:0] rf_wdata_fwd_wb_o_t0;
wire [31:0] rf_wdata_fwd_wb_o_t0;
/* src = "generated/sv2v_out.v:20933.20-20933.33" */
input [31:0] rf_wdata_id_i;
wire [31:0] rf_wdata_id_i;
/* cellift = 32'd1 */
input [31:0] rf_wdata_id_i_t0;
wire [31:0] rf_wdata_id_i_t0;
/* src = "generated/sv2v_out.v:20936.20-20936.34" */
input [31:0] rf_wdata_lsu_i;
wire [31:0] rf_wdata_lsu_i;
/* cellift = 32'd1 */
input [31:0] rf_wdata_lsu_i_t0;
wire [31:0] rf_wdata_lsu_i_t0;
/* src = "generated/sv2v_out.v:20940.21-20940.34" */
output [31:0] rf_wdata_wb_o;
wire [31:0] rf_wdata_wb_o;
/* cellift = 32'd1 */
output [31:0] rf_wdata_wb_o_t0;
wire [31:0] rf_wdata_wb_o_t0;
/* src = "generated/sv2v_out.v:20934.13-20934.23" */
input rf_we_id_i;
wire rf_we_id_i;
/* cellift = 32'd1 */
input rf_we_id_i_t0;
wire rf_we_id_i_t0;
/* src = "generated/sv2v_out.v:20937.13-20937.24" */
input rf_we_lsu_i;
wire rf_we_lsu_i;
/* cellift = 32'd1 */
input rf_we_lsu_i_t0;
wire rf_we_lsu_i_t0;
/* src = "generated/sv2v_out.v:20941.14-20941.24" */
output rf_we_wb_o;
wire rf_we_wb_o;
/* cellift = 32'd1 */
output rf_we_wb_o_t0;
wire rf_we_wb_o_t0;
/* src = "generated/sv2v_out.v:20924.14-20924.27" */
output rf_write_wb_o;
wire rf_write_wb_o;
/* cellift = 32'd1 */
output rf_write_wb_o_t0;
wire rf_write_wb_o_t0;
/* src = "generated/sv2v_out.v:20917.13-20917.19" */
input rst_ni;
wire rst_ni;
assign _00_ = instr_perf_count_id_i & /* src = "generated/sv2v_out.v:21045.34-21045.65" */ en_wb_i;
assign _02_ = lsu_resp_valid_i & /* src = "generated/sv2v_out.v:21045.71-21045.104" */ lsu_resp_err_i;
assign perf_instr_ret_wb_o = _00_ & /* src = "generated/sv2v_out.v:21045.33-21045.105" */ _42_;
assign perf_instr_ret_compressed_wb_o = perf_instr_ret_wb_o & /* src = "generated/sv2v_out.v:21046.44-21046.90" */ instr_is_compressed_id_i;
assign _04_ = { rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i } & /* src = "generated/sv2v_out.v:21067.26-21067.75" */ rf_wdata_id_i;
assign _06_ = { rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i } & /* src = "generated/sv2v_out.v:21067.80-21067.129" */ rf_wdata_lsu_i;
assign _13_ = instr_perf_count_id_i_t0 & en_wb_i;
assign _16_ = lsu_resp_valid_i_t0 & lsu_resp_err_i;
assign _19_ = _01_ & _42_;
assign _22_ = perf_instr_ret_wb_o_t0 & instr_is_compressed_id_i;
assign _25_ = { rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0 } & rf_wdata_id_i;
assign _28_ = { rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0 } & rf_wdata_lsu_i;
assign _14_ = en_wb_i_t0 & instr_perf_count_id_i;
assign _17_ = lsu_resp_err_i_t0 & lsu_resp_valid_i;
assign _20_ = _03_ & _00_;
assign _23_ = instr_is_compressed_id_i_t0 & perf_instr_ret_wb_o;
assign _26_ = rf_wdata_id_i_t0 & { rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i, rf_we_id_i };
assign _29_ = rf_wdata_lsu_i_t0 & { rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i, rf_we_lsu_i };
assign _15_ = instr_perf_count_id_i_t0 & en_wb_i_t0;
assign _18_ = lsu_resp_valid_i_t0 & lsu_resp_err_i_t0;
assign _21_ = _01_ & _03_;
assign _24_ = perf_instr_ret_wb_o_t0 & instr_is_compressed_id_i_t0;
assign _27_ = { rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0, rf_we_id_i_t0 } & rf_wdata_id_i_t0;
assign _30_ = { rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0, rf_we_lsu_i_t0 } & rf_wdata_lsu_i_t0;
assign _35_ = _13_ | _14_;
assign _36_ = _16_ | _17_;
assign _37_ = _19_ | _20_;
assign _38_ = _22_ | _23_;
assign _39_ = _25_ | _26_;
assign _40_ = _28_ | _29_;
assign _01_ = _35_ | _15_;
assign _03_ = _36_ | _18_;
assign perf_instr_ret_wb_o_t0 = _37_ | _21_;
assign perf_instr_ret_compressed_wb_o_t0 = _38_ | _24_;
assign _05_ = _39_ | _27_;
assign _07_ = _40_ | _30_;
assign _08_ = | { rf_we_lsu_i_t0, rf_we_id_i_t0 };
assign _09_ = ~ { rf_we_lsu_i_t0, rf_we_id_i_t0 };
assign _34_ = { rf_we_lsu_i, rf_we_id_i } & _09_;
assign _10_ = ! _34_;
assign rf_we_wb_o_t0 = _10_ & _08_;
assign _11_ = ~ _04_;
assign _12_ = ~ _06_;
assign _31_ = _05_ & _12_;
assign _32_ = _07_ & _11_;
assign _33_ = _05_ & _07_;
assign _41_ = _31_ | _32_;
assign rf_wdata_wb_o_t0 = _41_ | _33_;
assign _42_ = ~ /* src = "generated/sv2v_out.v:21045.69-21045.105" */ _02_;
assign rf_wdata_wb_o = _04_ | /* src = "generated/sv2v_out.v:21067.25-21067.130" */ _06_;
assign rf_we_wb_o = | /* src = "generated/sv2v_out.v:21068.22-21068.41" */ { rf_we_lsu_i, rf_we_id_i };
assign dummy_instr_wb_o = dummy_instr_id_i;
assign dummy_instr_wb_o_t0 = dummy_instr_id_i_t0;
assign instr_done_wb_o = 1'h0;
assign instr_done_wb_o_t0 = 1'h0;
assign outstanding_load_wb_o = 1'h0;
assign outstanding_load_wb_o_t0 = 1'h0;
assign outstanding_store_wb_o = 1'h0;
assign outstanding_store_wb_o_t0 = 1'h0;
assign pc_wb_o = 32'd0;
assign pc_wb_o_t0 = 32'd0;
assign perf_instr_ret_compressed_wb_spec_o = 1'h0;
assign perf_instr_ret_compressed_wb_spec_o_t0 = 1'h0;
assign perf_instr_ret_wb_spec_o = 1'h0;
assign perf_instr_ret_wb_spec_o_t0 = 1'h0;
assign ready_wb_o = 1'h1;
assign ready_wb_o_t0 = 1'h0;
assign rf_waddr_wb_o = rf_waddr_id_i;
assign rf_waddr_wb_o_t0 = rf_waddr_id_i_t0;
assign rf_wdata_fwd_wb_o = 32'd0;
assign rf_wdata_fwd_wb_o_t0 = 32'd0;
assign rf_write_wb_o = 1'h0;
assign rf_write_wb_o_t0 = 1'h0;
endmodule

module \$paramod\prim_buf\Width=32'00000000000000000000000000001100 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23015.22-23015.26" */
input [11:0] in_i;
wire [11:0] in_i;
/* cellift = 32'd1 */
input [11:0] in_i_t0;
wire [11:0] in_i_t0;
/* src = "generated/sv2v_out.v:23016.28-23016.33" */
output [11:0] out_o;
wire [11:0] out_o;
/* cellift = 32'd1 */
output [11:0] out_o_t0;
wire [11:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23026.38-23029.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000001100  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_buf\Width=32'00000000000000000000000000100000 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23015.22-23015.26" */
input [31:0] in_i;
wire [31:0] in_i;
/* cellift = 32'd1 */
input [31:0] in_i_t0;
wire [31:0] in_i_t0;
/* src = "generated/sv2v_out.v:23016.28-23016.33" */
output [31:0] out_o;
wire [31:0] out_o;
/* cellift = 32'd1 */
output [31:0] out_o_t0;
wire [31:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23026.38-23029.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000100000  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_buf\Width=32'00000000000000000000000000100111 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23015.22-23015.26" */
input [38:0] in_i;
wire [38:0] in_i;
/* cellift = 32'd1 */
input [38:0] in_i_t0;
wire [38:0] in_i_t0;
/* src = "generated/sv2v_out.v:23016.28-23016.33" */
output [38:0] out_o;
wire [38:0] out_o;
/* cellift = 32'd1 */
output [38:0] out_o_t0;
wire [38:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23026.38-23029.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000100111  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_buf\Width=s32'00000000000000000000000000000100 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23015.22-23015.26" */
input [3:0] in_i;
wire [3:0] in_i;
/* cellift = 32'd1 */
input [3:0] in_i_t0;
wire [3:0] in_i_t0;
/* src = "generated/sv2v_out.v:23016.28-23016.33" */
output [3:0] out_o;
wire [3:0] out_o;
/* cellift = 32'd1 */
output [3:0] out_o_t0;
wire [3:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23026.38-23029.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000000100  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_buf\Width=s32'00000000000000000000000000000111 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23015.22-23015.26" */
input [6:0] in_i;
wire [6:0] in_i;
/* cellift = 32'd1 */
input [6:0] in_i_t0;
wire [6:0] in_i_t0;
/* src = "generated/sv2v_out.v:23016.28-23016.33" */
output [6:0] out_o;
wire [6:0] out_o;
/* cellift = 32'd1 */
output [6:0] out_o_t0;
wire [6:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23026.38-23029.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000000111  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_buf\Width=s32'00000000000000000000000000100000 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:23015.22-23015.26" */
input [31:0] in_i;
wire [31:0] in_i;
/* cellift = 32'd1 */
input [31:0] in_i_t0;
wire [31:0] in_i_t0;
/* src = "generated/sv2v_out.v:23016.28-23016.33" */
output [31:0] out_o;
wire [31:0] out_o;
/* cellift = 32'd1 */
output [31:0] out_o_t0;
wire [31:0] out_o_t0;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:23026.38-23029.5" */
\$paramod\prim_generic_buf\Width=s32'00000000000000000000000000100000  \gen_generic.u_impl_generic  (
.in_i(in_i),
.in_i_t0(in_i_t0),
.out_o(out_o),
.out_o_t0(out_o_t0)
);
endmodule

module \$paramod\prim_generic_buf\Width=s32'00000000000000000000000000000100 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:24862.22-24862.26" */
input [3:0] in_i;
wire [3:0] in_i;
/* cellift = 32'd1 */
input [3:0] in_i_t0;
wire [3:0] in_i_t0;
/* src = "generated/sv2v_out.v:24864.21-24864.24" */
wire [3:0] inv;
/* src = "generated/sv2v_out.v:24863.28-24863.33" */
output [3:0] out_o;
wire [3:0] out_o;
/* cellift = 32'd1 */
output [3:0] out_o_t0;
wire [3:0] out_o_t0;
assign inv = ~ /* src = "generated/sv2v_out.v:24865.15-24865.20" */ in_i;
assign out_o = ~ /* src = "generated/sv2v_out.v:24866.17-24866.21" */ inv;
assign out_o_t0 = in_i_t0;
endmodule

module \$paramod\prim_generic_buf\Width=s32'00000000000000000000000000000111 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:24862.22-24862.26" */
input [6:0] in_i;
wire [6:0] in_i;
/* cellift = 32'd1 */
input [6:0] in_i_t0;
wire [6:0] in_i_t0;
/* src = "generated/sv2v_out.v:24864.21-24864.24" */
wire [6:0] inv;
/* src = "generated/sv2v_out.v:24863.28-24863.33" */
output [6:0] out_o;
wire [6:0] out_o;
/* cellift = 32'd1 */
output [6:0] out_o_t0;
wire [6:0] out_o_t0;
assign inv = ~ /* src = "generated/sv2v_out.v:24865.15-24865.20" */ in_i;
assign out_o = ~ /* src = "generated/sv2v_out.v:24866.17-24866.21" */ inv;
assign out_o_t0 = in_i_t0;
endmodule

module \$paramod\prim_generic_buf\Width=s32'00000000000000000000000000001100 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:24862.22-24862.26" */
input [11:0] in_i;
wire [11:0] in_i;
/* cellift = 32'd1 */
input [11:0] in_i_t0;
wire [11:0] in_i_t0;
/* src = "generated/sv2v_out.v:24864.21-24864.24" */
wire [11:0] inv;
/* src = "generated/sv2v_out.v:24863.28-24863.33" */
output [11:0] out_o;
wire [11:0] out_o;
/* cellift = 32'd1 */
output [11:0] out_o_t0;
wire [11:0] out_o_t0;
assign inv = ~ /* src = "generated/sv2v_out.v:24865.15-24865.20" */ in_i;
assign out_o = ~ /* src = "generated/sv2v_out.v:24866.17-24866.21" */ inv;
assign out_o_t0 = in_i_t0;
endmodule

module \$paramod\prim_generic_buf\Width=s32'00000000000000000000000000100000 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:24862.22-24862.26" */
input [31:0] in_i;
wire [31:0] in_i;
/* cellift = 32'd1 */
input [31:0] in_i_t0;
wire [31:0] in_i_t0;
/* src = "generated/sv2v_out.v:24864.21-24864.24" */
wire [31:0] inv;
/* src = "generated/sv2v_out.v:24863.28-24863.33" */
output [31:0] out_o;
wire [31:0] out_o;
/* cellift = 32'd1 */
output [31:0] out_o_t0;
wire [31:0] out_o_t0;
assign inv = ~ /* src = "generated/sv2v_out.v:24865.15-24865.20" */ in_i;
assign out_o = ~ /* src = "generated/sv2v_out.v:24866.17-24866.21" */ inv;
assign out_o_t0 = in_i_t0;
endmodule

module \$paramod\prim_generic_buf\Width=s32'00000000000000000000000000100111 (in_i, out_o, out_o_t0, in_i_t0);
/* src = "generated/sv2v_out.v:24862.22-24862.26" */
input [38:0] in_i;
wire [38:0] in_i;
/* cellift = 32'd1 */
input [38:0] in_i_t0;
wire [38:0] in_i_t0;
/* src = "generated/sv2v_out.v:24864.21-24864.24" */
wire [38:0] inv;
/* src = "generated/sv2v_out.v:24863.28-24863.33" */
output [38:0] out_o;
wire [38:0] out_o;
/* cellift = 32'd1 */
output [38:0] out_o_t0;
wire [38:0] out_o_t0;
assign inv = ~ /* src = "generated/sv2v_out.v:24865.15-24865.20" */ in_i;
assign out_o = ~ /* src = "generated/sv2v_out.v:24866.17-24866.21" */ inv;
assign out_o_t0 = in_i_t0;
endmodule

module ibex_compressed_decoder(clk_i, rst_ni, valid_i, instr_i, instr_o, is_compressed_o, illegal_instr_o, valid_i_t0, is_compressed_o_t0, instr_o_t0, instr_i_t0, illegal_instr_o_t0);
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0000_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0001_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0002_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0003_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0004_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0005_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0006_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0007_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0008_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0009_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0010_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0011_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0012_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0013_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0014_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0015_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0016_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0017_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0018_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0019_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0020_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0021_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0022_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0023_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0024_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0025_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0026_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0027_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0028_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0029_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0030_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0031_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0032_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0033_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0034_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0035_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0036_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0037_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire _0038_;
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0039_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12050.2-12136.5" */
wire [31:0] _0040_;
wire _0041_;
wire _0042_;
wire _0043_;
wire _0044_;
wire _0045_;
wire [4:0] _0046_;
wire [1:0] _0047_;
wire [2:0] _0048_;
wire [1:0] _0049_;
wire [2:0] _0050_;
wire _0051_;
wire _0052_;
wire _0053_;
wire _0054_;
wire _0055_;
wire _0056_;
wire _0057_;
wire _0058_;
wire _0059_;
wire _0060_;
wire _0061_;
wire [1:0] _0062_;
wire [5:0] _0063_;
wire [3:0] _0064_;
wire [7:0] _0065_;
wire [5:0] _0066_;
wire [4:0] _0067_;
wire [3:0] _0068_;
wire [3:0] _0069_;
wire [1:0] _0070_;
wire [1:0] _0071_;
wire [4:0] _0072_;
wire _0073_;
wire _0074_;
wire _0075_;
wire _0076_;
wire _0077_;
wire _0078_;
wire _0079_;
wire _0080_;
wire _0081_;
wire _0082_;
wire _0083_;
wire _0084_;
wire _0085_;
wire _0086_;
wire _0087_;
wire _0088_;
wire _0089_;
wire [31:0] _0090_;
wire [31:0] _0091_;
wire [31:0] _0092_;
wire [31:0] _0093_;
wire [31:0] _0094_;
wire [31:0] _0095_;
wire [31:0] _0096_;
wire [31:0] _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire [31:0] _0101_;
wire [31:0] _0102_;
wire [31:0] _0103_;
wire [31:0] _0104_;
wire [31:0] _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire [31:0] _0109_;
wire [31:0] _0110_;
wire _0111_;
wire _0112_;
wire _0113_;
wire [31:0] _0114_;
wire [31:0] _0115_;
wire [31:0] _0116_;
wire [31:0] _0117_;
wire [31:0] _0118_;
wire _0119_;
wire _0120_;
wire [31:0] _0121_;
wire [31:0] _0122_;
wire _0123_;
wire _0124_;
wire _0125_;
wire _0126_;
wire _0127_;
/* cellift = 32'd1 */
wire _0128_;
wire _0129_;
/* cellift = 32'd1 */
wire _0130_;
wire _0131_;
/* cellift = 32'd1 */
wire _0132_;
wire [1:0] _0133_;
wire [5:0] _0134_;
wire _0135_;
wire _0136_;
wire _0137_;
wire _0138_;
wire _0139_;
wire _0140_;
wire _0141_;
wire _0142_;
wire _0143_;
wire _0144_;
wire _0145_;
wire _0146_;
wire [3:0] _0147_;
wire _0148_;
wire _0149_;
wire _0150_;
wire _0151_;
wire _0152_;
wire _0153_;
wire _0154_;
wire _0155_;
wire _0156_;
wire [31:0] _0157_;
wire [31:0] _0158_;
wire [31:0] _0159_;
wire [31:0] _0160_;
wire [31:0] _0161_;
wire [31:0] _0162_;
wire [31:0] _0163_;
wire [31:0] _0164_;
wire [31:0] _0165_;
wire [31:0] _0166_;
wire [31:0] _0167_;
wire [31:0] _0168_;
wire [31:0] _0169_;
wire [31:0] _0170_;
wire [31:0] _0171_;
wire [31:0] _0172_;
wire [31:0] _0173_;
wire [31:0] _0174_;
wire [31:0] _0175_;
wire [31:0] _0176_;
wire [31:0] _0177_;
wire [31:0] _0178_;
wire [31:0] _0179_;
wire [31:0] _0180_;
wire _0181_;
wire _0182_;
wire _0183_;
wire _0184_;
wire _0185_;
wire [31:0] _0186_;
wire [31:0] _0187_;
wire [31:0] _0188_;
wire [31:0] _0189_;
wire [31:0] _0190_;
wire [31:0] _0191_;
wire [31:0] _0192_;
wire [31:0] _0193_;
wire [31:0] _0194_;
wire [31:0] _0195_;
wire [31:0] _0196_;
wire [31:0] _0197_;
wire [31:0] _0198_;
wire [31:0] _0199_;
wire [31:0] _0200_;
wire [31:0] _0201_;
wire [31:0] _0202_;
wire [31:0] _0203_;
wire [31:0] _0204_;
wire [31:0] _0205_;
wire [31:0] _0206_;
wire _0207_;
wire _0208_;
wire _0209_;
wire _0210_;
wire _0211_;
wire _0212_;
wire _0213_;
wire _0214_;
wire _0215_;
wire [31:0] _0216_;
wire [31:0] _0217_;
wire [31:0] _0218_;
wire [31:0] _0219_;
wire [31:0] _0220_;
wire [31:0] _0221_;
wire [31:0] _0222_;
wire [31:0] _0223_;
wire [31:0] _0224_;
wire _0225_;
wire _0226_;
wire _0227_;
wire _0228_;
wire _0229_;
wire _0230_;
wire _0231_;
wire _0232_;
wire [31:0] _0233_;
wire [31:0] _0234_;
wire [31:0] _0235_;
wire [31:0] _0236_;
wire [31:0] _0237_;
wire [31:0] _0238_;
wire [31:0] _0239_;
wire [31:0] _0240_;
wire [31:0] _0241_;
wire [7:0] _0242_;
wire [4:0] _0243_;
wire [5:0] _0244_;
wire [4:0] _0245_;
wire [1:0] _0246_;
wire [31:0] _0247_;
wire [31:0] _0248_;
wire [31:0] _0249_;
wire [31:0] _0250_;
wire [31:0] _0251_;
wire [31:0] _0252_;
wire [31:0] _0253_;
wire [31:0] _0254_;
wire _0255_;
wire _0256_;
wire _0257_;
wire _0258_;
wire [31:0] _0259_;
wire [31:0] _0260_;
wire [31:0] _0261_;
wire [3:0] _0262_;
wire [3:0] _0263_;
wire [2:0] _0264_;
wire [1:0] _0265_;
wire [31:0] _0266_;
wire [31:0] _0267_;
wire [31:0] _0268_;
wire [1:0] _0269_;
wire [1:0] _0270_;
wire [4:0] _0271_;
wire [2:0] _0272_;
wire _0273_;
/* cellift = 32'd1 */
wire _0274_;
wire _0275_;
/* cellift = 32'd1 */
wire _0276_;
wire _0277_;
/* cellift = 32'd1 */
wire _0278_;
wire _0279_;
/* cellift = 32'd1 */
wire _0280_;
wire _0281_;
wire _0282_;
wire _0283_;
wire _0284_;
wire _0285_;
wire _0286_;
wire _0287_;
wire _0288_;
wire _0289_;
wire _0290_;
wire _0291_;
wire _0292_;
wire _0293_;
wire [31:0] _0294_;
wire [31:0] _0295_;
wire [31:0] _0296_;
wire [31:0] _0297_;
wire [31:0] _0298_;
wire [31:0] _0299_;
wire [31:0] _0300_;
wire [31:0] _0301_;
wire [31:0] _0302_;
wire [31:0] _0303_;
wire [31:0] _0304_;
wire [31:0] _0305_;
wire [31:0] _0306_;
wire [31:0] _0307_;
wire [31:0] _0308_;
wire [31:0] _0309_;
wire [31:0] _0310_;
wire [31:0] _0311_;
wire [31:0] _0312_;
wire [31:0] _0313_;
wire [31:0] _0314_;
wire [31:0] _0315_;
wire [31:0] _0316_;
wire [31:0] _0317_;
wire _0318_;
wire _0319_;
wire _0320_;
wire _0321_;
wire [31:0] _0322_;
wire [31:0] _0323_;
wire [31:0] _0324_;
wire [31:0] _0325_;
wire [31:0] _0326_;
wire [31:0] _0327_;
wire [31:0] _0328_;
wire [31:0] _0329_;
wire [31:0] _0330_;
wire [31:0] _0331_;
wire [31:0] _0332_;
wire [31:0] _0333_;
wire [31:0] _0334_;
wire [31:0] _0335_;
wire [31:0] _0336_;
wire [31:0] _0337_;
wire [31:0] _0338_;
wire _0339_;
wire _0340_;
wire _0341_;
wire _0342_;
wire [31:0] _0343_;
wire [31:0] _0344_;
wire [31:0] _0345_;
wire [31:0] _0346_;
wire [31:0] _0347_;
wire [31:0] _0348_;
wire [31:0] _0349_;
wire _0350_;
wire _0351_;
wire _0352_;
wire _0353_;
wire _0354_;
wire _0355_;
wire _0356_;
wire [31:0] _0357_;
wire [31:0] _0358_;
wire [31:0] _0359_;
wire [31:0] _0360_;
wire [31:0] _0361_;
wire [31:0] _0362_;
wire [31:0] _0363_;
wire [31:0] _0364_;
wire [31:0] _0365_;
wire [31:0] _0366_;
wire [31:0] _0367_;
wire [31:0] _0368_;
wire [31:0] _0369_;
wire [31:0] _0370_;
wire _0371_;
wire _0372_;
wire [31:0] _0373_;
wire [31:0] _0374_;
wire [31:0] _0375_;
wire [31:0] _0376_;
wire [31:0] _0377_;
wire [31:0] _0378_;
wire _0379_;
wire _0380_;
wire _0381_;
wire [31:0] _0382_;
wire [31:0] _0383_;
wire [31:0] _0384_;
wire [31:0] _0385_;
wire [31:0] _0386_;
wire [31:0] _0387_;
wire [31:0] _0388_;
wire [31:0] _0389_;
wire _0390_;
wire [31:0] _0391_;
wire [31:0] _0392_;
wire [31:0] _0393_;
wire [31:0] _0394_;
wire [31:0] _0395_;
wire [31:0] _0396_;
wire [31:0] _0397_;
wire _0398_;
wire _0399_;
wire [31:0] _0400_;
wire [31:0] _0401_;
wire [31:0] _0402_;
wire _0403_;
wire _0404_;
wire [31:0] _0405_;
wire [31:0] _0406_;
wire [31:0] _0407_;
wire [31:0] _0408_;
wire [31:0] _0409_;
wire [31:0] _0410_;
wire [31:0] _0411_;
wire _0412_;
wire _0413_;
wire _0414_;
wire _0415_;
wire _0416_;
wire _0417_;
wire _0418_;
wire _0419_;
wire _0420_;
wire _0421_;
wire _0422_;
wire _0423_;
wire _0424_;
wire _0425_;
wire _0426_;
wire _0427_;
wire _0428_;
wire _0429_;
wire _0430_;
wire _0431_;
wire _0432_;
/* cellift = 32'd1 */
wire _0433_;
wire _0434_;
/* cellift = 32'd1 */
wire _0435_;
wire _0436_;
/* cellift = 32'd1 */
wire _0437_;
wire [31:0] _0438_;
/* cellift = 32'd1 */
wire [31:0] _0439_;
wire [31:0] _0440_;
/* cellift = 32'd1 */
wire [31:0] _0441_;
wire [31:0] _0442_;
/* cellift = 32'd1 */
wire [31:0] _0443_;
wire [31:0] _0444_;
/* cellift = 32'd1 */
wire [31:0] _0445_;
wire [31:0] _0446_;
/* cellift = 32'd1 */
wire [31:0] _0447_;
wire [31:0] _0448_;
/* cellift = 32'd1 */
wire [31:0] _0449_;
wire _0450_;
/* cellift = 32'd1 */
wire _0451_;
wire [31:0] _0452_;
/* cellift = 32'd1 */
wire [31:0] _0453_;
wire [31:0] _0454_;
/* cellift = 32'd1 */
wire [31:0] _0455_;
wire [31:0] _0456_;
/* cellift = 32'd1 */
wire [31:0] _0457_;
wire [31:0] _0458_;
/* cellift = 32'd1 */
wire [31:0] _0459_;
wire [31:0] _0460_;
/* cellift = 32'd1 */
wire [31:0] _0461_;
/* cellift = 32'd1 */
wire _0462_;
wire _0463_;
/* cellift = 32'd1 */
wire _0464_;
wire [31:0] _0465_;
/* cellift = 32'd1 */
wire [31:0] _0466_;
wire [31:0] _0467_;
/* cellift = 32'd1 */
wire [31:0] _0468_;
wire _0469_;
/* cellift = 32'd1 */
wire _0470_;
wire _0471_;
/* cellift = 32'd1 */
wire _0472_;
wire [31:0] _0473_;
/* cellift = 32'd1 */
wire [31:0] _0474_;
wire [31:0] _0475_;
/* cellift = 32'd1 */
wire [31:0] _0476_;
/* src = "generated/sv2v_out.v:12058.11-12058.39" */
wire _0477_;
/* src = "generated/sv2v_out.v:12073.11-12073.33" */
wire _0478_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12073.11-12073.33" */
wire _0479_;
/* src = "generated/sv2v_out.v:12075.11-12075.51" */
wire _0480_;
/* src = "generated/sv2v_out.v:12109.11-12109.36" */
wire _0481_;
/* src = "generated/sv2v_out.v:12114.12-12114.36" */
wire _0482_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:12114.12-12114.36" */
wire _0483_;
/* src = "generated/sv2v_out.v:12069.164-12069.176" */
wire _0484_;
wire _0485_;
/* cellift = 32'd1 */
wire _0486_;
wire _0487_;
/* cellift = 32'd1 */
wire _0488_;
wire _0489_;
/* cellift = 32'd1 */
wire _0490_;
wire _0491_;
/* cellift = 32'd1 */
wire _0492_;
wire [3:0] _0493_;
/* cellift = 32'd1 */
wire [3:0] _0494_;
wire _0495_;
wire _0496_;
/* cellift = 32'd1 */
wire _0497_;
wire [3:0] _0498_;
/* cellift = 32'd1 */
wire [3:0] _0499_;
wire _0500_;
wire _0501_;
/* cellift = 32'd1 */
wire _0502_;
wire _0503_;
/* cellift = 32'd1 */
wire _0504_;
wire _0505_;
/* cellift = 32'd1 */
wire _0506_;
wire _0507_;
/* cellift = 32'd1 */
wire _0508_;
wire _0509_;
/* cellift = 32'd1 */
wire _0510_;
wire _0511_;
/* cellift = 32'd1 */
wire _0512_;
wire _0513_;
/* cellift = 32'd1 */
wire _0514_;
wire _0515_;
/* cellift = 32'd1 */
wire _0516_;
wire _0517_;
/* cellift = 32'd1 */
wire _0518_;
wire _0519_;
/* src = "generated/sv2v_out.v:12041.13-12041.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:12047.13-12047.28" */
output illegal_instr_o;
wire illegal_instr_o;
/* cellift = 32'd1 */
output illegal_instr_o_t0;
wire illegal_instr_o_t0;
/* src = "generated/sv2v_out.v:12044.20-12044.27" */
input [31:0] instr_i;
wire [31:0] instr_i;
/* cellift = 32'd1 */
input [31:0] instr_i_t0;
wire [31:0] instr_i_t0;
/* src = "generated/sv2v_out.v:12045.20-12045.27" */
output [31:0] instr_o;
wire [31:0] instr_o;
/* cellift = 32'd1 */
output [31:0] instr_o_t0;
wire [31:0] instr_o_t0;
/* src = "generated/sv2v_out.v:12046.14-12046.29" */
output is_compressed_o;
wire is_compressed_o;
/* cellift = 32'd1 */
output is_compressed_o_t0;
wire is_compressed_o_t0;
/* src = "generated/sv2v_out.v:12042.13-12042.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:12043.13-12043.20" */
input valid_i;
wire valid_i;
/* cellift = 32'd1 */
input valid_i_t0;
wire valid_i_t0;
assign _0041_ = | instr_i_t0[11:7];
assign _0042_ = | instr_i_t0[1:0];
assign _0043_ = | { instr_i_t0[12], instr_i_t0[6:5] };
assign _0044_ = | instr_i_t0[11:10];
assign _0045_ = | instr_i_t0[15:13];
assign _0047_ = ~ instr_i_t0[1:0];
assign _0048_ = ~ { instr_i_t0[12], instr_i_t0[6:5] };
assign _0049_ = ~ instr_i_t0[11:10];
assign _0264_ = { instr_i[12], instr_i[6:5] } & _0048_;
assign _0265_ = instr_i[11:10] & _0049_;
assign _0246_ = instr_i[1:0] & _0047_;
assign _0412_ = _0243_ == { 3'h0, _0046_[1], 1'h0 };
assign _0413_ = _0246_ == _0047_;
assign _0414_ = _0264_ == { _0048_[2], 2'h0 };
assign _0415_ = _0264_ == { _0048_[2], 1'h0, _0048_[0] };
assign _0416_ = _0264_ == { _0048_[2:1], 1'h0 };
assign _0417_ = _0264_ == _0048_;
assign _0418_ = _0264_ == { 1'h0, _0048_[1:0] };
assign _0419_ = _0264_ == { 1'h0, _0048_[1], 1'h0 };
assign _0420_ = _0264_ == { 2'h0, _0048_[0] };
assign _0421_ = _0265_ == _0049_;
assign _0422_ = _0265_ == { _0049_[1], 1'h0 };
assign _0423_ = _0272_ == { 2'h0, _0050_[0] };
assign _0424_ = _0272_ == { 1'h0, _0050_[1:0] };
assign _0425_ = _0272_ == { _0050_[2], 2'h0 };
assign _0426_ = _0272_ == { _0050_[2], 1'h0, _0050_[0] };
assign _0427_ = _0272_ == _0050_;
assign _0428_ = _0272_ == { _0050_[2:1], 1'h0 };
assign _0429_ = _0272_ == { 1'h0, _0050_[1], 1'h0 };
assign _0430_ = _0246_ == { 1'h0, _0047_[0] };
assign _0431_ = _0246_ == { _0047_[1], 1'h0 };
assign _0479_ = _0412_ & _0041_;
assign is_compressed_o_t0 = _0413_ & _0042_;
assign _0499_[0] = _0414_ & _0043_;
assign _0499_[1] = _0415_ & _0043_;
assign _0499_[2] = _0416_ & _0043_;
assign _0499_[3] = _0417_ & _0043_;
assign _0502_ = _0418_ & _0043_;
assign _0504_ = _0419_ & _0043_;
assign _0506_ = _0420_ & _0043_;
assign _0508_ = _0421_ & _0044_;
assign _0512_ = _0422_ & _0044_;
assign _0494_[0] = _0423_ & _0045_;
assign _0494_[1] = _0424_ & _0045_;
assign _0486_ = _0425_ & _0045_;
assign _0494_[2] = _0426_ & _0045_;
assign _0494_[3] = _0427_ & _0045_;
assign _0497_ = _0428_ & _0045_;
assign _0490_ = _0429_ & _0045_;
assign _0510_ = _0430_ & _0042_;
assign _0488_ = _0431_ & _0042_;
assign _0051_ = | { _0497_, _0490_ };
assign _0052_ = | { _0497_, _0494_[3:2], _0494_[0], _0492_, _0490_ };
assign _0053_ = | { _0497_, _0494_[3], _0494_[1], _0486_ };
assign _0054_ = | instr_i_t0[12:5];
assign _0055_ = | { instr_i_t0[12], instr_i_t0[6:2] };
assign _0056_ = | instr_i_t0[6:2];
assign _0057_ = | _0494_;
assign _0058_ = | _0499_;
assign _0059_ = | { _0497_, _0494_[3] };
assign _0060_ = | { _0494_[2], _0494_[0] };
assign _0061_ = | { _0494_, _0486_ };
assign _0062_ = ~ { _0497_, _0490_ };
assign _0063_ = ~ { _0497_, _0494_[3:2], _0494_[0], _0492_, _0490_ };
assign _0064_ = ~ { _0497_, _0494_[3], _0494_[1], _0486_ };
assign _0065_ = ~ instr_i_t0[12:5];
assign _0066_ = ~ { instr_i_t0[12], instr_i_t0[6:2] };
assign _0046_ = ~ instr_i_t0[11:7];
assign _0067_ = ~ instr_i_t0[6:2];
assign _0068_ = ~ _0494_;
assign _0069_ = ~ _0499_;
assign _0070_ = ~ { _0497_, _0494_[3] };
assign _0071_ = ~ { _0494_[2], _0494_[0] };
assign _0072_ = ~ { _0494_, _0486_ };
assign _0050_ = ~ instr_i_t0[15:13];
assign _0133_ = { _0496_, _0489_ } & _0062_;
assign _0134_ = { _0496_, _0493_[3:2], _0493_[0], _0491_, _0489_ } & _0063_;
assign _0147_ = { _0496_, _0493_[3], _0493_[1], _0485_ } & _0064_;
assign _0242_ = instr_i[12:5] & _0065_;
assign _0244_ = { instr_i[12], instr_i[6:2] } & _0066_;
assign _0243_ = instr_i[11:7] & _0046_;
assign _0245_ = instr_i[6:2] & _0067_;
assign _0262_ = _0493_ & _0068_;
assign _0263_ = _0498_ & _0069_;
assign _0269_ = { _0496_, _0493_[3] } & _0070_;
assign _0270_ = { _0493_[2], _0493_[0] } & _0071_;
assign _0271_ = { _0493_, _0485_ } & _0072_;
assign _0272_ = instr_i[15:13] & _0050_;
assign _0073_ = ! _0133_;
assign _0074_ = ! _0134_;
assign _0075_ = ! _0147_;
assign _0076_ = ! _0242_;
assign _0077_ = ! _0244_;
assign _0078_ = ! _0243_;
assign _0079_ = ! _0245_;
assign _0080_ = ! _0262_;
assign _0081_ = ! _0263_;
assign _0082_ = ! _0269_;
assign _0083_ = ! _0270_;
assign _0084_ = ! _0271_;
assign _0085_ = ! _0272_;
assign _0130_ = _0073_ & _0051_;
assign _0132_ = _0074_ & _0052_;
assign _0128_ = _0075_ & _0053_;
assign _0016_ = _0076_ & _0054_;
assign _0024_ = _0077_ & _0055_;
assign _0004_ = _0078_ & _0041_;
assign _0483_ = _0079_ & _0056_;
assign _0433_ = _0080_ & _0057_;
assign _0034_ = _0081_ & _0058_;
assign _0514_ = _0082_ & _0059_;
assign _0516_ = _0083_ & _0060_;
assign _0518_ = _0084_ & _0061_;
assign _0492_ = _0085_ & _0045_;
assign _0086_ = ~ _0495_;
assign _0087_ = ~ _0489_;
assign _0088_ = ~ _0485_;
assign _0089_ = ~ _0273_;
assign _0090_ = ~ { _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_ };
assign _0091_ = ~ { _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_ };
assign _0092_ = ~ { _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_ };
assign _0093_ = ~ { _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_ };
assign _0094_ = ~ { _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_ };
assign _0095_ = ~ { _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_ };
assign _0096_ = ~ { _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_ };
assign _0097_ = ~ { _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_ };
assign _0098_ = ~ _0500_;
assign _0099_ = ~ _0511_;
assign _0100_ = ~ _0507_;
assign _0101_ = ~ { _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_ };
assign _0102_ = ~ { _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_ };
assign _0103_ = ~ { _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_ };
assign _0104_ = ~ { _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_ };
assign _0105_ = ~ { _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_ };
assign _0106_ = ~ _0131_;
assign _0107_ = ~ _0129_;
assign _0108_ = ~ _0517_;
assign _0109_ = ~ { _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_ };
assign _0110_ = ~ { _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_ };
assign _0111_ = ~ _0519_;
assign _0112_ = ~ _0509_;
assign _0113_ = ~ _0279_;
assign _0114_ = ~ { _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_ };
assign _0115_ = ~ { _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_ };
assign _0116_ = ~ { _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_ };
assign _0117_ = ~ { _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_, _0481_ };
assign _0118_ = ~ { _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_ };
assign _0119_ = ~ _0482_;
assign _0120_ = ~ instr_i[12];
assign _0121_ = ~ { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12] };
assign _0122_ = ~ { _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_ };
assign _0285_ = _0490_ | _0087_;
assign _0288_ = _0486_ | _0088_;
assign _0291_ = _0274_ | _0089_;
assign _0294_ = { _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_ } | _0090_;
assign _0297_ = { _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_ } | _0091_;
assign _0300_ = { _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_ } | _0092_;
assign _0303_ = { _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_ } | _0093_;
assign _0306_ = { _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_ } | _0094_;
assign _0309_ = { _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_ } | _0095_;
assign _0312_ = { _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_ } | _0096_;
assign _0315_ = { _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_ } | _0097_;
assign _0318_ = _0512_ | _0099_;
assign _0319_ = _0508_ | _0100_;
assign _0322_ = { _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_ } | _0101_;
assign _0325_ = { _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_ } | _0102_;
assign _0329_ = { _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_ } | _0103_;
assign _0332_ = { _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_ } | _0104_;
assign _0336_ = { _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_ } | _0105_;
assign _0340_ = _0132_ | _0106_;
assign _0341_ = _0130_ | _0107_;
assign _0342_ = _0518_ | _0108_;
assign _0343_ = { _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_ } | _0109_;
assign _0347_ = { _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_ } | _0110_;
assign _0350_ = is_compressed_o_t0 | _0111_;
assign _0351_ = _0510_ | _0112_;
assign _0354_ = _0280_ | _0113_;
assign _0357_ = { is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0 } | _0114_;
assign _0360_ = { _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_ } | _0115_;
assign _0363_ = { _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_ } | _0116_;
assign _0366_ = { _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_ } | _0117_;
assign _0367_ = { _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_ } | _0118_;
assign _0371_ = _0483_ | _0119_;
assign _0372_ = instr_i_t0[12] | _0120_;
assign _0373_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12] } | _0121_;
assign _0376_ = { _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_ } | _0122_;
assign _0286_ = _0490_ | _0489_;
assign _0289_ = _0486_ | _0485_;
assign _0292_ = _0274_ | _0273_;
assign _0295_ = { _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_ } | { _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_, _0495_ };
assign _0298_ = { _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_ } | { _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_, _0489_ };
assign _0301_ = { _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_ } | { _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_, _0485_ };
assign _0304_ = { _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_ } | { _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_, _0273_ };
assign _0307_ = { _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_ } | { _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_, _0500_ };
assign _0310_ = { _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_ } | { _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_, _0505_ };
assign _0313_ = { _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_ } | { _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_, _0503_ };
assign _0316_ = { _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_ } | { _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_, _0275_ };
assign _0320_ = _0508_ | _0507_;
assign _0323_ = { _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_ } | { _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_, _0511_ };
assign _0326_ = { _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_ } | { _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_, _0507_ };
assign _0330_ = { _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_ } | { _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_, _0513_ };
assign _0333_ = { _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_ } | { _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_, _0515_ };
assign _0337_ = { _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_ } | { _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_, _0127_ };
assign _0344_ = { _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_ } | { _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_, _0517_ };
assign _0348_ = { _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_ } | { _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_, _0277_ };
assign _0352_ = _0510_ | _0509_;
assign _0355_ = _0280_ | _0279_;
assign _0358_ = { is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0 } | { _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_, _0519_ };
assign _0361_ = { _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_ } | { _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_, _0509_ };
assign _0364_ = { _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_ } | { _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_, _0279_ };
assign _0368_ = { _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_ } | { _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_, _0482_ };
assign _0374_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12] } | { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12] };
assign _0377_ = { _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_ } | { _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_, _0478_ };
assign _0148_ = instr_i_t0[12] & _0285_;
assign _0151_ = _0435_ & _0288_;
assign _0154_ = _0437_ & _0291_;
assign _0157_ = { 4'h0, instr_i_t0[8:7], instr_i_t0[12], instr_i_t0[6:2], 8'h00, instr_i_t0[11:9], 9'h000 } & _0294_;
assign _0160_ = { 7'h00, instr_i_t0[6:2], instr_i_t0[11:7], 3'h0, instr_i_t0[11:7], 7'h00 } & _0297_;
assign _0163_ = _0441_ & _0300_;
assign _0166_ = _0443_ & _0303_;
assign _0169_ = { 9'h000, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 } & _0306_;
assign _0172_ = { 9'h000, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 } & _0309_;
assign _0175_ = _0447_ & _0312_;
assign _0178_ = _0449_ & _0315_;
assign _0181_ = instr_i_t0[12] & _0318_;
assign _0183_ = _0451_ & _0319_;
assign _0186_ = { 1'h0, instr_i_t0[10], 5'h00, instr_i_t0[6:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 } & _0322_;
assign _0189_ = _0453_ & _0325_;
assign _0192_ = _0022_ & _0300_;
assign _0195_ = _0455_ & _0329_;
assign _0198_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:2], instr_i_t0[11:7], 3'h0, instr_i_t0[11:7], 7'h00 } & _0332_;
assign _0201_ = _0459_ & _0297_;
assign _0204_ = _0461_ & _0336_;
assign _0207_ = _0024_ & _0288_;
assign _0210_ = _0462_ & _0340_;
assign _0212_ = _0016_ & _0341_;
assign _0214_ = _0464_ & _0342_;
assign _0216_ = { 5'h00, instr_i_t0[5], instr_i_t0[12], 2'h0, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 3'h0, instr_i_t0[11:10], instr_i_t0[6], 9'h000 } & _0343_;
assign _0219_ = { 2'h0, instr_i_t0[10:7], instr_i_t0[12:11], instr_i_t0[5], instr_i_t0[6], 12'h000, instr_i_t0[4:2], 7'h00 } & _0297_;
assign _0222_ = _0468_ & _0347_;
assign _0225_ = _0038_ & _0350_;
assign _0227_ = _0012_ & _0351_;
assign _0230_ = _0472_ & _0354_;
assign _0233_ = _0032_ & _0357_;
assign _0236_ = _0014_ & _0360_;
assign _0239_ = _0476_ & _0363_;
assign _0247_ = { 12'h000, instr_i_t0[11:7], 15'h0000 } & _0366_;
assign _0249_ = _0006_ & _0367_;
assign _0252_ = { 12'h000, instr_i_t0[11:7], 15'h0000 } & _0367_;
assign _0255_ = _0004_ & _0371_;
assign _0257_ = _0010_ & _0372_;
assign _0259_ = _0040_ & _0373_;
assign _0266_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:2], instr_i_t0[11:7], 7'h00 } & _0376_;
assign _0149_ = _0004_ & _0286_;
assign _0152_ = _0008_ & _0289_;
assign _0155_ = _0433_ & _0292_;
assign _0158_ = instr_i_t0 & _0295_;
assign _0161_ = { 4'h0, instr_i_t0[3:2], instr_i_t0[12], instr_i_t0[6:4], 10'h000, instr_i_t0[11:7], 7'h00 } & _0298_;
assign _0164_ = _0036_ & _0301_;
assign _0167_ = _0439_ & _0304_;
assign _0170_ = instr_i_t0 & _0307_;
assign _0173_ = { 9'h000, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 } & _0310_;
assign _0176_ = { 9'h000, instr_i_t0[4:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 } & _0313_;
assign _0179_ = _0445_ & _0316_;
assign _0184_ = _0034_ & _0320_;
assign _0187_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:2], 2'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[9:7], 7'h00 } & _0323_;
assign _0190_ = _0030_ & _0326_;
assign _0193_ = _0026_ & _0301_;
assign _0196_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:5], instr_i_t0[2], 7'h00, instr_i_t0[9:7], 2'h0, instr_i_t0[13], instr_i_t0[11:10], instr_i_t0[4:3], instr_i_t0[12], 7'h00 } & _0330_;
assign _0199_ = { instr_i_t0[12], instr_i_t0[8], instr_i_t0[10:9], instr_i_t0[6], instr_i_t0[7], instr_i_t0[2], instr_i_t0[11], instr_i_t0[5:3], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], 4'h0, instr_i_t0[15], 7'h00 } & _0333_;
assign _0202_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[6:2], 8'h00, instr_i_t0[11:7], 7'h00 } & _0298_;
assign _0205_ = _0457_ & _0337_;
assign _0208_ = _0028_ & _0289_;
assign _0217_ = instr_i_t0 & _0344_;
assign _0220_ = { 5'h00, instr_i_t0[5], instr_i_t0[12:10], instr_i_t0[6], 4'h0, instr_i_t0[9:7], 5'h00, instr_i_t0[4:2], 7'h00 } & _0298_;
assign _0223_ = _0466_ & _0348_;
assign _0228_ = _0020_ & _0352_;
assign _0231_ = _0470_ & _0355_;
assign _0234_ = instr_i_t0 & _0358_;
assign _0237_ = _0018_ & _0361_;
assign _0240_ = _0474_ & _0364_;
assign _0250_ = { 7'h00, instr_i_t0[6:2], instr_i_t0[11:7], 3'h0, instr_i_t0[11:7], 7'h00 } & _0368_;
assign _0253_ = { 7'h00, instr_i_t0[6:2], 8'h00, instr_i_t0[11:7], 7'h00 } & _0368_;
assign _0260_ = _0002_ & _0374_;
assign _0267_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[4:3], instr_i_t0[5], instr_i_t0[2], instr_i_t0[6], 24'h000000 } & _0377_;
assign _0287_ = _0148_ | _0149_;
assign _0290_ = _0151_ | _0152_;
assign _0293_ = _0154_ | _0155_;
assign _0296_ = _0157_ | _0158_;
assign _0299_ = _0160_ | _0161_;
assign _0302_ = _0163_ | _0164_;
assign _0305_ = _0166_ | _0167_;
assign _0308_ = _0169_ | _0170_;
assign _0311_ = _0172_ | _0173_;
assign _0314_ = _0175_ | _0176_;
assign _0317_ = _0178_ | _0179_;
assign _0321_ = _0183_ | _0184_;
assign _0324_ = _0186_ | _0187_;
assign _0327_ = _0189_ | _0190_;
assign _0328_ = _0192_ | _0193_;
assign _0331_ = _0195_ | _0196_;
assign _0334_ = _0198_ | _0199_;
assign _0335_ = _0201_ | _0202_;
assign _0338_ = _0204_ | _0205_;
assign _0339_ = _0207_ | _0208_;
assign _0345_ = _0216_ | _0217_;
assign _0346_ = _0219_ | _0220_;
assign _0349_ = _0222_ | _0223_;
assign _0353_ = _0227_ | _0228_;
assign _0356_ = _0230_ | _0231_;
assign _0359_ = _0233_ | _0234_;
assign _0362_ = _0236_ | _0237_;
assign _0365_ = _0239_ | _0240_;
assign _0369_ = _0249_ | _0250_;
assign _0370_ = _0252_ | _0253_;
assign _0375_ = _0259_ | _0260_;
assign _0378_ = _0266_ | _0267_;
assign _0379_ = _0000_ ^ _0003_;
assign _0380_ = _0434_ ^ _0007_;
assign _0381_ = _0436_ ^ _0432_;
assign _0382_ = { 4'h0, instr_i[8:7], instr_i[12], instr_i[6:2], 8'h12, instr_i[11:9], 9'h023 } ^ instr_i;
assign _0383_ = { 7'h00, instr_i[6:2], instr_i[11:7], 3'h1, instr_i[11:7], 7'h13 } ^ { 4'h0, instr_i[3:2], instr_i[12], instr_i[6:4], 10'h012, instr_i[11:7], 7'h03 };
assign _0384_ = _0440_ ^ _0035_;
assign _0385_ = _0442_ ^ _0438_;
assign _0386_ = { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h1d, instr_i[9:7], 7'h33 } ^ instr_i;
assign _0387_ = { 9'h081, instr_i[4:2], 2'h1, instr_i[9:7], 5'h01, instr_i[9:7], 7'h33 } ^ { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h11, instr_i[9:7], 7'h33 };
assign _0388_ = _0446_ ^ { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h19, instr_i[9:7], 7'h33 };
assign _0389_ = _0448_ ^ _0444_;
assign _0390_ = _0450_ ^ _0033_;
assign _0391_ = { 1'h0, instr_i[10], 5'h00, instr_i[6:2], 2'h1, instr_i[9:7], 5'h15, instr_i[9:7], 7'h13 } ^ { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], 2'h1, instr_i[9:7], 5'h1d, instr_i[9:7], 7'h13 };
assign _0392_ = _0452_ ^ _0029_;
assign _0393_ = _0021_ ^ _0025_;
assign _0394_ = _0454_ ^ { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:5], instr_i[2], 7'h01, instr_i[9:7], 2'h0, instr_i[13], instr_i[11:10], instr_i[4:3], instr_i[12], 7'h63 };
assign _0395_ = { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], instr_i[11:7], 3'h0, instr_i[11:7], 7'h13 } ^ { instr_i[12], instr_i[8], instr_i[10:9], instr_i[6], instr_i[7], instr_i[2], instr_i[11], instr_i[5:3], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], 4'h0, _0484_, 7'h6f };
assign _0396_ = _0458_ ^ { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], 8'h00, instr_i[11:7], 7'h13 };
assign _0397_ = _0460_ ^ _0456_;
assign _0398_ = _0023_ ^ _0027_;
assign _0400_ = { 5'h00, instr_i[5], instr_i[12], 2'h1, instr_i[4:2], 2'h1, instr_i[9:7], 3'h2, instr_i[11:10], instr_i[6], 9'h023 } ^ instr_i;
assign _0401_ = { 2'h0, instr_i[10:7], instr_i[12:11], instr_i[5], instr_i[6], 12'h041, instr_i[4:2], 7'h13 } ^ { 5'h00, instr_i[5], instr_i[12:10], instr_i[6], 4'h1, instr_i[9:7], 5'h09, instr_i[4:2], 7'h03 };
assign _0402_ = _0467_ ^ _0465_;
assign _0403_ = _0011_ ^ _0019_;
assign _0404_ = _0471_ ^ _0469_;
assign _0405_ = _0031_ ^ instr_i;
assign _0406_ = _0013_ ^ _0017_;
assign _0407_ = _0475_ ^ _0473_;
assign _0408_ = _0005_ ^ { 7'h00, instr_i[6:2], instr_i[11:7], 3'h0, instr_i[11:7], 7'h33 };
assign _0409_ = { 12'h000, instr_i[11:7], 15'h0067 } ^ { 7'h00, instr_i[6:2], 8'h00, instr_i[11:7], 7'h33 };
assign _0410_ = _0039_ ^ _0001_;
assign _0411_ = { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], instr_i[11:7], 7'h37 } ^ { instr_i[12], instr_i[12], instr_i[12], instr_i[4:3], instr_i[5], instr_i[2], instr_i[6], 24'h010113 };
assign _0150_ = _0490_ & _0379_;
assign _0153_ = _0486_ & _0380_;
assign _0156_ = _0274_ & _0381_;
assign _0159_ = { _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_, _0433_ } & _0382_;
assign _0162_ = { _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_ } & _0383_;
assign _0165_ = { _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_ } & _0384_;
assign _0168_ = { _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_, _0274_ } & _0385_;
assign _0171_ = { _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_, _0034_ } & _0386_;
assign _0174_ = { _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_, _0506_ } & _0387_;
assign _0177_ = { _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_, _0504_ } & _0388_;
assign _0180_ = { _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_, _0276_ } & _0389_;
assign _0182_ = _0512_ & _0000_;
assign _0185_ = _0508_ & _0390_;
assign _0188_ = { _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_, _0512_ } & _0391_;
assign _0191_ = { _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_, _0508_ } & _0392_;
assign _0194_ = { _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_, _0486_ } & _0393_;
assign _0197_ = { _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_, _0514_ } & _0394_;
assign _0200_ = { _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_, _0516_ } & _0395_;
assign _0203_ = { _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_ } & _0396_;
assign _0206_ = { _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_, _0128_ } & _0397_;
assign _0209_ = _0486_ & _0398_;
assign _0211_ = _0132_ & _0399_;
assign _0213_ = _0130_ & _0015_;
assign _0215_ = _0518_ & _0123_;
assign _0218_ = { _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_, _0518_ } & _0400_;
assign _0221_ = { _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_, _0490_ } & _0401_;
assign _0224_ = { _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_, _0278_ } & _0402_;
assign _0226_ = is_compressed_o_t0 & _0037_;
assign _0229_ = _0510_ & _0403_;
assign _0232_ = _0280_ & _0404_;
assign _0235_ = { is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0, is_compressed_o_t0 } & _0405_;
assign _0238_ = { _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_, _0510_ } & _0406_;
assign _0241_ = { _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_, _0280_ } & _0407_;
assign _0248_ = { _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_, _0004_ } & { 12'h001, instr_i[11:7], 15'h0094 };
assign _0251_ = { _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_ } & _0408_;
assign _0254_ = { _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_, _0483_ } & _0409_;
assign _0256_ = _0483_ & _0003_;
assign _0258_ = instr_i_t0[12] & _0009_;
assign _0261_ = { instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12], instr_i_t0[12] } & _0410_;
assign _0268_ = { _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_, _0479_ } & _0411_;
assign _0435_ = _0150_ | _0287_;
assign _0437_ = _0153_ | _0290_;
assign _0038_ = _0156_ | _0293_;
assign _0439_ = _0159_ | _0296_;
assign _0441_ = _0162_ | _0299_;
assign _0443_ = _0165_ | _0302_;
assign _0032_ = _0168_ | _0305_;
assign _0445_ = _0171_ | _0308_;
assign _0447_ = _0174_ | _0311_;
assign _0449_ = _0177_ | _0314_;
assign _0030_ = _0180_ | _0317_;
assign _0451_ = _0182_ | _0181_;
assign _0028_ = _0185_ | _0321_;
assign _0453_ = _0188_ | _0324_;
assign _0026_ = _0191_ | _0327_;
assign _0455_ = _0194_ | _0328_;
assign _0457_ = _0197_ | _0331_;
assign _0459_ = _0200_ | _0334_;
assign _0461_ = _0203_ | _0335_;
assign _0018_ = _0206_ | _0338_;
assign _0462_ = _0209_ | _0339_;
assign _0020_ = _0211_ | _0210_;
assign _0464_ = _0213_ | _0212_;
assign _0012_ = _0215_ | _0214_;
assign _0466_ = _0218_ | _0345_;
assign _0468_ = _0221_ | _0346_;
assign _0014_ = _0224_ | _0349_;
assign _0470_ = _0226_ | _0225_;
assign _0472_ = _0229_ | _0353_;
assign illegal_instr_o_t0 = _0232_ | _0356_;
assign _0474_ = _0235_ | _0359_;
assign _0476_ = _0238_ | _0362_;
assign instr_o_t0 = _0241_ | _0365_;
assign _0006_ = _0248_ | _0247_;
assign _0002_ = _0251_ | _0369_;
assign _0040_ = _0254_ | _0370_;
assign _0010_ = _0256_ | _0255_;
assign _0008_ = _0258_ | _0257_;
assign _0036_ = _0261_ | _0375_;
assign _0022_ = _0268_ | _0378_;
assign _0123_ = ~ _0463_;
assign _0129_ = | { _0496_, _0489_ };
assign _0131_ = | { _0496_, _0493_[3:2], _0493_[0], _0491_, _0489_ };
assign _0124_ = ~ _0496_;
assign _0125_ = ~ _0501_;
assign _0126_ = ~ _0487_;
assign _0135_ = _0497_ & _0086_;
assign _0138_ = _0502_ & _0098_;
assign _0141_ = _0497_ & _0108_;
assign _0144_ = _0488_ & _0111_;
assign _0136_ = _0433_ & _0124_;
assign _0139_ = _0034_ & _0125_;
assign _0142_ = _0518_ & _0124_;
assign _0145_ = is_compressed_o_t0 & _0126_;
assign _0137_ = _0497_ & _0433_;
assign _0140_ = _0502_ & _0034_;
assign _0143_ = _0497_ & _0518_;
assign _0146_ = _0488_ & is_compressed_o_t0;
assign _0281_ = _0135_ | _0136_;
assign _0282_ = _0138_ | _0139_;
assign _0283_ = _0141_ | _0142_;
assign _0284_ = _0144_ | _0145_;
assign _0274_ = _0281_ | _0137_;
assign _0276_ = _0282_ | _0140_;
assign _0278_ = _0283_ | _0143_;
assign _0280_ = _0284_ | _0146_;
assign _0273_ = _0496_ | _0495_;
assign _0275_ = _0501_ | _0500_;
assign _0277_ = _0496_ | _0517_;
assign _0279_ = _0487_ | _0519_;
assign _0127_ = | { _0496_, _0493_[3], _0493_[1], _0485_ };
assign _0432_ = _0495_ ? 1'h1 : 1'h0;
assign _0434_ = _0489_ ? _0003_ : _0000_;
assign _0436_ = _0485_ ? _0007_ : _0434_;
assign _0037_ = _0273_ ? _0432_ : _0436_;
assign _0438_ = _0495_ ? instr_i : { 4'h0, instr_i[8:7], instr_i[12], instr_i[6:2], 8'h12, instr_i[11:9], 9'h023 };
assign _0440_ = _0489_ ? { 4'h0, instr_i[3:2], instr_i[12], instr_i[6:4], 10'h012, instr_i[11:7], 7'h03 } : { 7'h00, instr_i[6:2], instr_i[11:7], 3'h1, instr_i[11:7], 7'h13 };
assign _0442_ = _0485_ ? _0035_ : _0440_;
assign _0031_ = _0273_ ? _0438_ : _0442_;
assign _0444_ = _0500_ ? instr_i : { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h1d, instr_i[9:7], 7'h33 };
assign _0446_ = _0505_ ? { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h11, instr_i[9:7], 7'h33 } : { 9'h081, instr_i[4:2], 2'h1, instr_i[9:7], 5'h01, instr_i[9:7], 7'h33 };
assign _0448_ = _0503_ ? { 9'h001, instr_i[4:2], 2'h1, instr_i[9:7], 5'h19, instr_i[9:7], 7'h33 } : _0446_;
assign _0029_ = _0275_ ? _0444_ : _0448_;
assign _0033_ = _0500_ ? 1'h1 : 1'h0;
assign _0450_ = _0511_ ? 1'h0 : _0000_;
assign _0027_ = _0507_ ? _0033_ : _0450_;
assign _0452_ = _0511_ ? { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], 2'h1, instr_i[9:7], 5'h1d, instr_i[9:7], 7'h13 } : { 1'h0, instr_i[10], 5'h00, instr_i[6:2], 2'h1, instr_i[9:7], 5'h15, instr_i[9:7], 7'h13 };
assign _0025_ = _0507_ ? _0029_ : _0452_;
assign _0454_ = _0485_ ? _0025_ : _0021_;
assign _0456_ = _0513_ ? { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:5], instr_i[2], 7'h01, instr_i[9:7], 2'h0, instr_i[13], instr_i[11:10], instr_i[4:3], instr_i[12], 7'h63 } : _0454_;
assign _0458_ = _0515_ ? { instr_i[12], instr_i[8], instr_i[10:9], instr_i[6], instr_i[7], instr_i[2], instr_i[11], instr_i[5:3], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], 4'h0, _0484_, 7'h6f } : { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], instr_i[11:7], 3'h0, instr_i[11:7], 7'h13 };
assign _0460_ = _0489_ ? { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], 8'h00, instr_i[11:7], 7'h13 } : _0458_;
assign _0017_ = _0127_ ? _0456_ : _0460_;
assign _0399_ = _0485_ ? _0027_ : _0023_;
assign _0019_ = _0131_ ? 1'h0 : _0399_;
assign _0463_ = _0129_ ? 1'h0 : _0015_;
assign _0011_ = _0517_ ? 1'h1 : _0463_;
assign _0465_ = _0517_ ? instr_i : { 5'h00, instr_i[5], instr_i[12], 2'h1, instr_i[4:2], 2'h1, instr_i[9:7], 3'h2, instr_i[11:10], instr_i[6], 9'h023 };
assign _0467_ = _0489_ ? { 5'h00, instr_i[5], instr_i[12:10], instr_i[6], 4'h1, instr_i[9:7], 5'h09, instr_i[4:2], 7'h03 } : { 2'h0, instr_i[10:7], instr_i[12:11], instr_i[5], instr_i[6], 12'h041, instr_i[4:2], 7'h13 };
assign _0013_ = _0277_ ? _0465_ : _0467_;
assign _0469_ = _0519_ ? 1'h0 : _0037_;
assign _0471_ = _0509_ ? _0019_ : _0011_;
assign illegal_instr_o = _0279_ ? _0469_ : _0471_;
assign _0473_ = _0519_ ? instr_i : _0031_;
assign _0475_ = _0509_ ? _0017_ : _0013_;
assign instr_o = _0279_ ? _0473_ : _0475_;
assign _0477_ = ! /* src = "generated/sv2v_out.v:12058.11-12058.39" */ instr_i[12:5];
assign _0478_ = instr_i[11:7] == /* src = "generated/sv2v_out.v:12073.11-12073.33" */ 5'h02;
assign _0480_ = ! /* src = "generated/sv2v_out.v:12075.11-12075.51" */ { instr_i[12], instr_i[6:2] };
assign _0481_ = ! /* src = "generated/sv2v_out.v:12124.16-12124.41" */ instr_i[11:7];
assign _0482_ = | /* src = "generated/sv2v_out.v:12122.16-12122.40" */ instr_i[6:2];
assign is_compressed_o = instr_i[1:0] != /* src = "generated/sv2v_out.v:12137.27-12137.48" */ 2'h3;
assign _0484_ = ~ /* src = "generated/sv2v_out.v:12069.164-12069.176" */ instr_i[15];
assign _0005_ = _0481_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12124.16-12124.41|generated/sv2v_out.v:12124.12-12127.77" */ 32'd1048691 : { 12'h000, instr_i[11:7], 15'h00e7 };
assign _0001_ = _0482_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12122.16-12122.40|generated/sv2v_out.v:12122.12-12127.77" */ { 7'h00, instr_i[6:2], instr_i[11:7], 3'h0, instr_i[11:7], 7'h33 } : _0005_;
assign _0039_ = _0482_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12114.12-12114.36|generated/sv2v_out.v:12114.8-12120.11" */ { 7'h00, instr_i[6:2], 8'h00, instr_i[11:7], 7'h33 } : { 12'h000, instr_i[11:7], 15'h0067 };
assign _0009_ = _0482_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12114.12-12114.36|generated/sv2v_out.v:12114.8-12120.11" */ 1'h0 : _0003_;
assign _0007_ = instr_i[12] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12113.11-12113.30|generated/sv2v_out.v:12113.7-12127.77" */ 1'h0 : _0009_;
assign _0035_ = instr_i[12] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12113.11-12113.30|generated/sv2v_out.v:12113.7-12127.77" */ _0001_ : _0039_;
assign _0003_ = _0481_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12109.11-12109.36|generated/sv2v_out.v:12109.7-12110.31" */ 1'h1 : 1'h0;
assign _0000_ = instr_i[12] ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12104.11-12104.30|generated/sv2v_out.v:12104.7-12105.31" */ 1'h1 : 1'h0;
assign _0495_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12101.5-12131.12" */ _0493_;
assign _0500_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12087.9-12094.16" */ _0498_;
assign _0498_[0] = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12087.9-12094.16" */ 3'h4;
assign _0498_[1] = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12087.9-12094.16" */ 3'h5;
assign _0498_[2] = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12087.9-12094.16" */ 3'h6;
assign _0498_[3] = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12087.9-12094.16" */ 3'h7;
assign _0501_ = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12087.9-12094.16" */ 3'h3;
assign _0503_ = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12087.9-12094.16" */ 3'h2;
assign _0505_ = { instr_i[12], instr_i[6:5] } == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12087.9-12094.16" */ 3'h1;
assign _0507_ = instr_i[11:10] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12079.7-12096.14" */ 2'h3;
assign _0511_ = instr_i[11:10] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12079.7-12096.14" */ 2'h2;
assign _0023_ = _0480_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12075.11-12075.51|generated/sv2v_out.v:12075.7-12076.31" */ 1'h1 : 1'h0;
assign _0021_ = _0478_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12073.11-12073.33|generated/sv2v_out.v:12073.7-12074.126" */ { instr_i[12], instr_i[12], instr_i[12], instr_i[4:3], instr_i[5], instr_i[2], instr_i[6], 24'h010113 } : { instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[12], instr_i[6:2], instr_i[11:7], 7'h37 };
assign _0513_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12067.5-12099.12" */ { _0496_, _0493_[3] };
assign _0515_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12067.5-12099.12" */ { _0493_[2], _0493_[0] };
assign _0015_ = _0477_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:12058.11-12058.39|generated/sv2v_out.v:12058.7-12059.31" */ 1'h1 : 1'h0;
assign _0517_ = | /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ { _0493_, _0485_ };
assign _0493_[0] = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ 3'h1;
assign _0493_[1] = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ 3'h3;
assign _0485_ = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ 3'h4;
assign _0493_[2] = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ 3'h5;
assign _0493_[3] = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ 3'h7;
assign _0496_ = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ 3'h6;
assign _0489_ = instr_i[15:13] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ 3'h2;
assign _0491_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12055.5-12065.12" */ instr_i[15:13];
assign _0509_ = instr_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12053.3-12135.10" */ 2'h1;
assign _0519_ = instr_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12053.3-12135.10" */ 2'h3;
assign _0487_ = instr_i[1:0] == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:12053.3-12135.10" */ 2'h2;
endmodule

module ibex_multdiv_slow(clk_i, rst_ni, mult_en_i, div_en_i, mult_sel_i, div_sel_i, operator_i, signed_mode_i, op_a_i, op_b_i, alu_adder_ext_i, alu_adder_i, equal_to_zero_i, data_ind_timing_i, alu_operand_a_o, alu_operand_b_o, imd_val_q_i, imd_val_d_o, imd_val_we_o, multdiv_ready_id_i, multdiv_result_o
, valid_o, valid_o_t0, data_ind_timing_i_t0, alu_adder_ext_i_t0, alu_adder_i_t0, alu_operand_a_o_t0, alu_operand_b_o_t0, div_en_i_t0, div_sel_i_t0, equal_to_zero_i_t0, imd_val_d_o_t0, imd_val_q_i_t0, imd_val_we_o_t0, mult_en_i_t0, mult_sel_i_t0, multdiv_ready_id_i_t0, multdiv_result_o_t0, op_a_i_t0, op_b_i_t0, operator_i_t0, signed_mode_i_t0
);
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0000_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0001_;
/* src = "generated/sv2v_out.v:19542.2-19575.5" */
wire [32:0] _0002_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19542.2-19575.5" */
wire [32:0] _0003_;
/* src = "generated/sv2v_out.v:19542.2-19575.5" */
wire [32:0] _0004_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19542.2-19575.5" */
wire [32:0] _0005_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [2:0] _0006_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [2:0] _0007_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [4:0] _0008_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [4:0] _0009_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire _0010_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire _0011_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0012_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0013_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0014_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0015_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [31:0] _0016_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [31:0] _0017_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0018_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0019_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire _0020_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire _0021_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [2:0] _0022_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [2:0] _0023_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire _0024_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire _0025_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0026_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0027_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0028_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0029_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0030_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0031_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [2:0] _0032_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [2:0] _0033_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0034_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0035_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0036_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0037_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0038_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0039_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [2:0] _0040_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [2:0] _0041_;
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0042_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19589.2-19701.5" */
wire [32:0] _0043_;
/* src = "generated/sv2v_out.v:19604.55-19604.88" */
wire [31:0] _0044_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19604.55-19604.88" */
wire [31:0] _0045_;
/* src = "generated/sv2v_out.v:19604.28-19604.52" */
wire _0046_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19604.28-19604.52" */
wire _0047_;
/* src = "generated/sv2v_out.v:19610.61-19610.94" */
wire [30:0] _0048_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19610.61-19610.94" */
wire [30:0] _0049_;
/* src = "generated/sv2v_out.v:19718.43-19718.111" */
wire _0050_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19718.43-19718.111" */
wire _0051_;
wire _0052_;
wire _0053_;
wire _0054_;
wire _0055_;
wire _0056_;
wire _0057_;
wire _0058_;
wire _0059_;
wire _0060_;
wire _0061_;
wire _0062_;
wire _0063_;
wire [1:0] _0064_;
wire [1:0] _0065_;
wire [1:0] _0066_;
wire _0067_;
wire [4:0] _0068_;
wire [2:0] _0069_;
wire [1:0] _0070_;
wire _0071_;
wire _0072_;
wire _0073_;
wire _0074_;
wire _0075_;
wire _0076_;
wire _0077_;
wire _0078_;
wire _0079_;
wire _0080_;
wire _0081_;
wire _0082_;
wire [1:0] _0083_;
wire [2:0] _0084_;
wire [2:0] _0085_;
wire [2:0] _0086_;
wire [1:0] _0087_;
wire [1:0] _0088_;
wire [2:0] _0089_;
wire [1:0] _0090_;
wire [3:0] _0091_;
wire [2:0] _0092_;
wire [32:0] _0093_;
wire [32:0] _0094_;
wire _0095_;
wire _0096_;
wire _0097_;
wire _0098_;
wire _0099_;
wire _0100_;
wire _0101_;
wire _0102_;
wire _0103_;
wire _0104_;
wire _0105_;
wire _0106_;
wire _0107_;
wire _0108_;
wire _0109_;
wire _0110_;
wire _0111_;
wire _0112_;
wire [32:0] _0113_;
wire [32:0] _0114_;
wire _0115_;
wire [2:0] _0116_;
wire [2:0] _0117_;
wire [32:0] _0118_;
wire [32:0] _0119_;
wire [2:0] _0120_;
wire [32:0] _0121_;
wire [32:0] _0122_;
wire [32:0] _0123_;
wire [32:0] _0124_;
wire [32:0] _0125_;
wire [32:0] _0126_;
wire [32:0] _0127_;
wire [32:0] _0128_;
wire [2:0] _0129_;
wire [2:0] _0130_;
wire [2:0] _0131_;
wire [2:0] _0132_;
wire _0133_;
wire [32:0] _0134_;
wire _0135_;
wire [31:0] _0136_;
wire [31:0] _0137_;
wire [32:0] _0138_;
wire [32:0] _0139_;
wire _0140_;
wire [31:0] _0141_;
wire [32:0] _0142_;
wire [31:0] _0143_;
wire [32:0] _0144_;
wire [32:0] _0145_;
wire [32:0] _0146_;
wire [31:0] _0147_;
wire [1:0] _0148_;
wire [1:0] _0149_;
wire [4:0] _0150_;
wire [32:0] _0151_;
wire _0152_;
wire _0153_;
wire [32:0] _0154_;
wire _0155_;
wire _0156_;
wire _0157_;
wire _0158_;
wire _0159_;
wire [32:0] _0160_;
wire _0161_;
wire _0162_;
wire _0163_;
wire _0164_;
wire _0165_;
/* cellift = 32'd1 */
wire _0166_;
wire _0167_;
/* cellift = 32'd1 */
wire _0168_;
wire _0169_;
wire _0170_;
wire _0171_;
wire _0172_;
wire _0173_;
wire _0174_;
wire _0175_;
wire _0176_;
wire _0177_;
wire _0178_;
wire _0179_;
wire _0180_;
/* cellift = 32'd1 */
wire _0181_;
wire _0182_;
/* cellift = 32'd1 */
wire _0183_;
wire _0184_;
/* cellift = 32'd1 */
wire _0185_;
wire _0186_;
/* cellift = 32'd1 */
wire _0187_;
wire _0188_;
/* cellift = 32'd1 */
wire _0189_;
wire _0190_;
/* cellift = 32'd1 */
wire _0191_;
wire _0192_;
/* cellift = 32'd1 */
wire _0193_;
wire _0194_;
/* cellift = 32'd1 */
wire _0195_;
wire _0196_;
/* cellift = 32'd1 */
wire _0197_;
wire _0198_;
/* cellift = 32'd1 */
wire _0199_;
wire _0200_;
/* cellift = 32'd1 */
wire _0201_;
wire _0202_;
/* cellift = 32'd1 */
wire _0203_;
wire _0204_;
wire _0205_;
/* cellift = 32'd1 */
wire _0206_;
wire _0207_;
/* cellift = 32'd1 */
wire _0208_;
wire _0209_;
/* cellift = 32'd1 */
wire _0210_;
wire [31:0] _0211_;
wire [31:0] _0212_;
wire [31:0] _0213_;
wire _0214_;
wire _0215_;
wire _0216_;
wire _0217_;
wire _0218_;
wire _0219_;
wire _0220_;
wire _0221_;
wire _0222_;
wire _0223_;
wire _0224_;
wire _0225_;
wire [31:0] _0226_;
wire [31:0] _0227_;
wire [31:0] _0228_;
wire [30:0] _0229_;
wire [30:0] _0230_;
wire [30:0] _0231_;
wire _0232_;
wire _0233_;
wire _0234_;
wire _0235_;
wire _0236_;
wire _0237_;
wire _0238_;
wire _0239_;
wire _0240_;
wire [2:0] _0241_;
wire [2:0] _0242_;
wire [2:0] _0243_;
wire [4:0] _0244_;
wire [4:0] _0245_;
wire [4:0] _0246_;
wire [32:0] _0247_;
wire [32:0] _0248_;
wire [32:0] _0249_;
wire [32:0] _0250_;
wire [32:0] _0251_;
wire [32:0] _0252_;
wire _0253_;
wire _0254_;
wire _0255_;
wire [1:0] _0256_;
wire [1:0] _0257_;
wire [1:0] _0258_;
wire [2:0] _0259_;
wire [1:0] _0260_;
wire [2:0] _0261_;
wire [2:0] _0262_;
wire [1:0] _0263_;
wire [1:0] _0264_;
wire [2:0] _0265_;
wire [1:0] _0266_;
wire [3:0] _0267_;
wire _0268_;
wire _0269_;
wire _0270_;
wire _0271_;
wire _0272_;
wire _0273_;
wire _0274_;
wire _0275_;
wire _0276_;
wire [2:0] _0277_;
wire [32:0] _0278_;
wire [32:0] _0279_;
wire [32:0] _0280_;
wire [32:0] _0281_;
wire [32:0] _0282_;
wire [32:0] _0283_;
wire _0284_;
wire _0285_;
wire [32:0] _0286_;
wire [32:0] _0287_;
wire [32:0] _0288_;
wire [32:0] _0289_;
wire [32:0] _0290_;
wire [32:0] _0291_;
wire [2:0] _0292_;
wire [2:0] _0293_;
wire [2:0] _0294_;
wire [32:0] _0295_;
wire [32:0] _0296_;
wire [32:0] _0297_;
wire [32:0] _0298_;
wire [32:0] _0299_;
wire [32:0] _0300_;
wire [32:0] _0301_;
wire [32:0] _0302_;
wire [32:0] _0303_;
wire [2:0] _0304_;
wire [2:0] _0305_;
wire [2:0] _0306_;
wire [2:0] _0307_;
wire [2:0] _0308_;
wire [32:0] _0309_;
wire [32:0] _0310_;
wire [32:0] _0311_;
wire [32:0] _0312_;
wire [32:0] _0313_;
wire [32:0] _0314_;
wire [32:0] _0315_;
wire [32:0] _0316_;
wire [32:0] _0317_;
wire [32:0] _0318_;
wire [32:0] _0319_;
wire [4:0] _0320_;
wire [4:0] _0321_;
wire [32:0] _0322_;
wire [32:0] _0323_;
wire [32:0] _0324_;
wire [32:0] _0325_;
wire [32:0] _0326_;
wire [32:0] _0327_;
wire [32:0] _0328_;
wire [32:0] _0329_;
wire [32:0] _0330_;
wire [32:0] _0331_;
wire [32:0] _0332_;
wire [32:0] _0333_;
wire [32:0] _0334_;
wire [32:0] _0335_;
wire [32:0] _0336_;
wire [32:0] _0337_;
wire [32:0] _0338_;
wire [32:0] _0339_;
wire [32:0] _0340_;
wire [32:0] _0341_;
wire [32:0] _0342_;
wire [32:0] _0343_;
wire [32:0] _0344_;
wire [32:0] _0345_;
wire [32:0] _0346_;
wire [32:0] _0347_;
wire [2:0] _0348_;
wire [2:0] _0349_;
wire [2:0] _0350_;
wire [2:0] _0351_;
wire [2:0] _0352_;
wire [2:0] _0353_;
wire [2:0] _0354_;
wire [2:0] _0355_;
wire [2:0] _0356_;
wire [2:0] _0357_;
wire [2:0] _0358_;
wire [2:0] _0359_;
wire [2:0] _0360_;
wire _0361_;
wire _0362_;
wire _0363_;
wire _0364_;
wire _0365_;
wire [32:0] _0366_;
wire [32:0] _0367_;
wire [32:0] _0368_;
wire [32:0] _0369_;
wire [32:0] _0370_;
wire [32:0] _0371_;
wire [32:0] _0372_;
wire [32:0] _0373_;
wire [32:0] _0374_;
wire [32:0] _0375_;
wire [32:0] _0376_;
wire [32:0] _0377_;
wire [32:0] _0378_;
wire [32:0] _0379_;
wire [32:0] _0380_;
wire [32:0] _0381_;
wire [32:0] _0382_;
wire [32:0] _0383_;
wire _0384_;
wire _0385_;
wire [32:0] _0386_;
wire [32:0] _0387_;
wire [4:0] _0388_;
wire _0389_;
wire _0390_;
wire _0391_;
wire _0392_;
wire _0393_;
wire _0394_;
wire _0395_;
wire _0396_;
wire _0397_;
wire _0398_;
wire _0399_;
wire _0400_;
wire _0401_;
wire _0402_;
wire _0403_;
wire [32:0] _0404_;
wire [32:0] _0405_;
wire [32:0] _0406_;
wire _0407_;
wire _0408_;
wire _0409_;
wire _0410_;
wire _0411_;
wire _0412_;
wire _0413_;
wire _0414_;
wire _0415_;
wire [2:0] _0416_;
wire [31:0] _0417_;
wire [31:0] _0418_;
wire [31:0] _0419_;
wire _0420_;
wire _0421_;
wire [31:0] _0422_;
wire [31:0] _0423_;
wire [31:0] _0424_;
wire [32:0] _0425_;
wire [32:0] _0426_;
wire [32:0] _0427_;
wire [32:0] _0428_;
wire [32:0] _0429_;
wire [1:0] _0430_;
wire [32:0] _0431_;
wire [32:0] _0432_;
wire [32:0] _0433_;
wire _0434_;
wire _0435_;
wire _0436_;
wire [31:0] _0437_;
wire [31:0] _0438_;
wire [31:0] _0439_;
wire [32:0] _0440_;
wire [32:0] _0441_;
wire [32:0] _0442_;
wire [31:0] _0443_;
wire [31:0] _0444_;
wire [31:0] _0445_;
wire [32:0] _0446_;
wire [32:0] _0447_;
wire [32:0] _0448_;
wire [32:0] _0449_;
wire [32:0] _0450_;
wire [32:0] _0451_;
wire [32:0] _0452_;
wire [32:0] _0453_;
wire [32:0] _0454_;
wire [31:0] _0455_;
wire [31:0] _0456_;
wire [31:0] _0457_;
wire _0458_;
/* cellift = 32'd1 */
wire _0459_;
wire _0460_;
/* cellift = 32'd1 */
wire _0461_;
wire _0462_;
/* cellift = 32'd1 */
wire _0463_;
wire [31:0] _0464_;
wire _0465_;
wire _0466_;
wire _0467_;
wire _0468_;
wire [31:0] _0469_;
wire [30:0] _0470_;
wire _0471_;
wire _0472_;
wire _0473_;
wire [2:0] _0474_;
wire [2:0] _0475_;
wire [2:0] _0476_;
wire [2:0] _0477_;
wire [4:0] _0478_;
wire [4:0] _0479_;
wire [4:0] _0480_;
wire [4:0] _0481_;
wire [32:0] _0482_;
wire [32:0] _0483_;
wire [32:0] _0484_;
wire [32:0] _0485_;
wire [32:0] _0486_;
wire [32:0] _0487_;
wire [32:0] _0488_;
wire [32:0] _0489_;
wire _0490_;
wire _0491_;
wire _0492_;
wire _0493_;
wire [1:0] _0494_;
wire [2:0] _0495_;
wire [4:0] _0496_;
wire [4:0] _0497_;
wire [3:0] _0498_;
wire _0499_;
wire _0500_;
wire _0501_;
wire [32:0] _0502_;
wire [32:0] _0503_;
wire [32:0] _0504_;
wire [32:0] _0505_;
wire [32:0] _0506_;
wire [32:0] _0507_;
wire _0508_;
wire [2:0] _0509_;
wire [2:0] _0510_;
wire [32:0] _0511_;
wire [32:0] _0512_;
wire [2:0] _0513_;
wire [2:0] _0514_;
wire [2:0] _0515_;
wire [32:0] _0516_;
wire [32:0] _0517_;
wire [32:0] _0518_;
wire [32:0] _0519_;
wire [32:0] _0520_;
wire [32:0] _0521_;
wire [32:0] _0522_;
wire [2:0] _0523_;
wire [2:0] _0524_;
wire [32:0] _0525_;
wire [32:0] _0526_;
wire [32:0] _0527_;
wire [32:0] _0528_;
wire [32:0] _0529_;
wire [4:0] _0530_;
wire [32:0] _0531_;
wire [32:0] _0532_;
wire [32:0] _0533_;
wire [32:0] _0534_;
wire [32:0] _0535_;
wire [32:0] _0536_;
wire [32:0] _0537_;
wire [32:0] _0538_;
wire [32:0] _0539_;
wire [32:0] _0540_;
wire [32:0] _0541_;
wire [32:0] _0542_;
wire [32:0] _0543_;
wire [32:0] _0544_;
wire [32:0] _0545_;
wire [32:0] _0546_;
wire [32:0] _0547_;
wire [32:0] _0548_;
wire [32:0] _0549_;
wire [32:0] _0550_;
wire [32:0] _0551_;
wire [32:0] _0552_;
wire [2:0] _0553_;
wire [2:0] _0554_;
wire [2:0] _0555_;
wire [2:0] _0556_;
wire [2:0] _0557_;
wire [2:0] _0558_;
wire [2:0] _0559_;
wire [2:0] _0560_;
wire [2:0] _0561_;
wire [2:0] _0562_;
wire [2:0] _0563_;
wire _0564_;
wire _0565_;
wire _0566_;
wire _0567_;
wire [32:0] _0568_;
wire [32:0] _0569_;
wire [32:0] _0570_;
wire [32:0] _0571_;
wire [32:0] _0572_;
wire [32:0] _0573_;
wire [32:0] _0574_;
wire [32:0] _0575_;
wire _0576_;
wire _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire [32:0] _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire [32:0] _0586_;
wire _0587_;
wire [31:0] _0588_;
wire [31:0] _0589_;
wire [31:0] _0590_;
wire _0591_;
wire [31:0] _0592_;
wire [31:0] _0593_;
wire [31:0] _0594_;
wire [32:0] _0595_;
wire [32:0] _0596_;
wire [32:0] _0597_;
wire [32:0] _0598_;
wire [4:0] _0599_;
wire [32:0] _0600_;
wire _0601_;
wire _0602_;
wire _0603_;
wire [31:0] _0604_;
wire [31:0] _0605_;
wire [31:0] _0606_;
wire [32:0] _0607_;
wire [32:0] _0608_;
wire [32:0] _0609_;
wire [31:0] _0610_;
wire [31:0] _0611_;
wire [31:0] _0612_;
wire [32:0] _0613_;
wire [32:0] _0614_;
wire [32:0] _0615_;
wire [32:0] _0616_;
wire [32:0] _0617_;
wire [32:0] _0618_;
wire [32:0] _0619_;
wire [32:0] _0620_;
wire [32:0] _0621_;
wire [31:0] _0622_;
wire [31:0] _0623_;
wire [31:0] _0624_;
wire [2:0] _0625_;
wire [4:0] _0626_;
wire [32:0] _0627_;
wire [32:0] _0628_;
wire _0629_;
wire [32:0] _0630_;
wire [32:0] _0631_;
wire _0632_;
wire [32:0] _0633_;
wire [32:0] _0634_;
wire [2:0] _0635_;
wire [32:0] _0636_;
wire [32:0] _0637_;
wire [32:0] _0638_;
wire [2:0] _0639_;
wire [2:0] _0640_;
wire [32:0] _0641_;
wire [32:0] _0642_;
wire [32:0] _0643_;
wire [32:0] _0644_;
wire [32:0] _0645_;
wire [32:0] _0646_;
wire [32:0] _0647_;
wire [32:0] _0648_;
wire [32:0] _0649_;
wire [32:0] _0650_;
wire [32:0] _0651_;
wire [2:0] _0652_;
wire [2:0] _0653_;
wire [2:0] _0654_;
wire [2:0] _0655_;
wire _0656_;
wire [32:0] _0657_;
wire [32:0] _0658_;
wire [32:0] _0659_;
wire [32:0] _0660_;
wire [32:0] _0661_;
wire [32:0] _0662_;
wire [31:0] _0663_;
wire [31:0] _0664_;
wire [32:0] _0665_;
wire [4:0] _0666_;
wire [32:0] _0667_;
wire _0668_;
wire [31:0] _0669_;
wire [32:0] _0670_;
wire [31:0] _0671_;
wire [32:0] _0672_;
wire [32:0] _0673_;
wire [31:0] _0674_;
wire _0675_;
wire _0676_;
wire _0677_;
wire _0678_;
wire _0679_;
wire _0680_;
wire _0681_;
wire _0682_;
wire _0683_;
wire _0684_;
wire _0685_;
wire _0686_;
wire _0687_;
wire _0688_;
wire [4:0] _0689_;
wire [4:0] _0690_;
wire [32:0] _0691_;
/* cellift = 32'd1 */
wire [32:0] _0692_;
wire [32:0] _0693_;
/* cellift = 32'd1 */
wire [32:0] _0694_;
wire [32:0] _0695_;
/* cellift = 32'd1 */
wire [32:0] _0696_;
wire [2:0] _0697_;
/* cellift = 32'd1 */
wire [2:0] _0698_;
wire [32:0] _0699_;
/* cellift = 32'd1 */
wire [32:0] _0700_;
wire [32:0] _0701_;
/* cellift = 32'd1 */
wire [32:0] _0702_;
wire [32:0] _0703_;
/* cellift = 32'd1 */
wire [32:0] _0704_;
wire [32:0] _0705_;
/* cellift = 32'd1 */
wire [32:0] _0706_;
wire [32:0] _0707_;
/* cellift = 32'd1 */
wire [32:0] _0708_;
wire [32:0] _0709_;
/* cellift = 32'd1 */
wire [32:0] _0710_;
wire [32:0] _0711_;
/* cellift = 32'd1 */
wire [32:0] _0712_;
wire [32:0] _0713_;
/* cellift = 32'd1 */
wire [32:0] _0714_;
wire [2:0] _0715_;
/* cellift = 32'd1 */
wire [2:0] _0716_;
wire [2:0] _0717_;
/* cellift = 32'd1 */
wire [2:0] _0718_;
wire [2:0] _0719_;
/* cellift = 32'd1 */
wire [2:0] _0720_;
wire [2:0] _0721_;
/* cellift = 32'd1 */
wire [2:0] _0722_;
wire [2:0] _0723_;
/* cellift = 32'd1 */
wire [2:0] _0724_;
wire _0725_;
/* cellift = 32'd1 */
wire _0726_;
wire [32:0] _0727_;
/* cellift = 32'd1 */
wire [32:0] _0728_;
wire [32:0] _0729_;
/* cellift = 32'd1 */
wire [32:0] _0730_;
wire [32:0] _0731_;
/* cellift = 32'd1 */
wire [32:0] _0732_;
wire _0733_;
wire [32:0] _0734_;
/* src = "generated/sv2v_out.v:19546.29-19546.47" */
wire _0735_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19546.29-19546.47" */
wire _0736_;
/* src = "generated/sv2v_out.v:19583.29-19583.67" */
wire _0737_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19583.29-19583.67" */
wire _0738_;
/* src = "generated/sv2v_out.v:19606.45-19606.65" */
wire _0739_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19606.45-19606.65" */
wire _0740_;
/* src = "generated/sv2v_out.v:19645.46-19645.63" */
wire _0741_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19645.46-19645.63" */
wire _0742_;
/* src = "generated/sv2v_out.v:19645.70-19645.93" */
wire _0743_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19645.70-19645.93" */
wire _0744_;
/* src = "generated/sv2v_out.v:19718.20-19718.38" */
wire _0745_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19718.20-19718.38" */
wire _0746_;
/* src = "generated/sv2v_out.v:19718.68-19718.86" */
wire _0747_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19718.68-19718.86" */
wire _0748_;
/* src = "generated/sv2v_out.v:19718.91-19718.109" */
wire _0749_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19718.91-19718.109" */
wire _0750_;
/* src = "generated/sv2v_out.v:19606.22-19606.66" */
wire _0751_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19606.22-19606.66" */
wire _0752_;
/* src = "generated/sv2v_out.v:19616.22-19616.59" */
wire _0753_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19616.22-19616.59" */
wire _0754_;
/* src = "generated/sv2v_out.v:19645.23-19645.64" */
wire _0755_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19645.23-19645.64" */
wire _0756_;
/* src = "generated/sv2v_out.v:19606.22-19606.40" */
wire _0757_;
/* src = "generated/sv2v_out.v:19598.7-19598.30" */
wire _0758_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19598.7-19598.30" */
wire _0759_;
/* src = "generated/sv2v_out.v:19645.22-19645.94" */
wire _0760_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19645.22-19645.94" */
wire _0761_;
/* src = "generated/sv2v_out.v:19551.26-19551.33" */
wire [31:0] _0762_;
/* src = "generated/sv2v_out.v:19555.26-19555.33" */
wire [31:0] _0763_;
/* src = "generated/sv2v_out.v:19563.26-19563.47" */
wire [31:0] _0764_;
/* src = "generated/sv2v_out.v:19567.26-19567.45" */
wire [31:0] _0765_;
/* src = "generated/sv2v_out.v:19583.70-19583.86" */
wire _0766_;
/* src = "generated/sv2v_out.v:19587.47-19587.61" */
wire _0767_;
/* src = "generated/sv2v_out.v:19604.26-19604.53" */
wire _0768_;
/* src = "generated/sv2v_out.v:19586.45-19586.69" */
wire [32:0] _0769_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19586.45-19586.69" */
wire [32:0] _0770_;
/* src = "generated/sv2v_out.v:19702.23-19702.43" */
wire _0771_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19702.23-19702.43" */
wire _0772_;
/* src = "generated/sv2v_out.v:19718.67-19718.110" */
wire _0773_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19718.67-19718.110" */
wire _0774_;
wire _0775_;
/* cellift = 32'd1 */
wire _0776_;
wire _0777_;
/* cellift = 32'd1 */
wire _0778_;
wire _0779_;
/* cellift = 32'd1 */
wire _0780_;
wire _0781_;
/* cellift = 32'd1 */
wire _0782_;
wire _0783_;
/* cellift = 32'd1 */
wire _0784_;
wire _0785_;
/* cellift = 32'd1 */
wire _0786_;
wire _0787_;
/* src = "generated/sv2v_out.v:0.0-0.0" */
wire _0788_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:0.0-0.0" */
wire _0789_;
/* src = "generated/sv2v_out.v:19639.24-19639.47" */
wire [4:0] _0790_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19639.24-19639.47" */
wire [4:0] _0791_;
/* src = "generated/sv2v_out.v:19546.29-19546.78" */
wire [32:0] _0792_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19546.29-19546.78" */
wire [32:0] _0793_;
/* src = "generated/sv2v_out.v:19606.22-19606.80" */
wire [2:0] _0794_;
/* src = "generated/sv2v_out.v:19616.22-19616.73" */
wire [2:0] _0795_;
/* src = "generated/sv2v_out.v:19630.24-19630.53" */
wire [31:0] _0796_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19630.24-19630.53" */
wire [31:0] _0797_;
/* src = "generated/sv2v_out.v:19635.22-19635.67" */
wire [32:0] _0798_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19635.22-19635.67" */
wire [32:0] _0799_;
/* src = "generated/sv2v_out.v:19645.22-19645.108" */
wire [2:0] _0800_;
/* src = "generated/sv2v_out.v:19651.22-19651.59" */
wire [2:0] _0801_;
/* src = "generated/sv2v_out.v:19689.31-19689.85" */
wire [32:0] _0802_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19689.31-19689.85" */
wire [32:0] _0803_;
/* src = "generated/sv2v_out.v:19690.31-19690.85" */
wire [32:0] _0804_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19690.31-19690.85" */
wire [32:0] _0805_;
/* src = "generated/sv2v_out.v:19587.28-19587.43" */
wire _0806_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19587.28-19587.43" */
wire _0807_;
/* src = "generated/sv2v_out.v:19502.13-19502.27" */
wire [32:0] accum_window_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19502.13-19502.27" */
wire [32:0] accum_window_d_t0;
/* src = "generated/sv2v_out.v:19487.20-19487.35" */
input [33:0] alu_adder_ext_i;
wire [33:0] alu_adder_ext_i;
/* cellift = 32'd1 */
input [33:0] alu_adder_ext_i_t0;
wire [33:0] alu_adder_ext_i_t0;
/* src = "generated/sv2v_out.v:19488.20-19488.31" */
input [31:0] alu_adder_i;
wire [31:0] alu_adder_i;
/* cellift = 32'd1 */
input [31:0] alu_adder_i_t0;
wire [31:0] alu_adder_i_t0;
/* src = "generated/sv2v_out.v:19491.20-19491.35" */
output [32:0] alu_operand_a_o;
wire [32:0] alu_operand_a_o;
/* cellift = 32'd1 */
output [32:0] alu_operand_a_o_t0;
wire [32:0] alu_operand_a_o_t0;
/* src = "generated/sv2v_out.v:19492.20-19492.35" */
output [32:0] alu_operand_b_o;
wire [32:0] alu_operand_b_o;
/* cellift = 32'd1 */
output [32:0] alu_operand_b_o_t0;
wire [32:0] alu_operand_b_o_t0;
/* src = "generated/sv2v_out.v:19477.13-19477.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:19490.13-19490.30" */
input data_ind_timing_i;
wire data_ind_timing_i;
/* cellift = 32'd1 */
input data_ind_timing_i_t0;
wire data_ind_timing_i_t0;
/* src = "generated/sv2v_out.v:19529.6-19529.19" */
reg div_by_zero_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19529.6-19529.19" */
reg div_by_zero_q_t0;
/* src = "generated/sv2v_out.v:19526.7-19526.22" */
wire div_change_sign;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19526.7-19526.22" */
wire div_change_sign_t0;
/* src = "generated/sv2v_out.v:19480.13-19480.21" */
input div_en_i;
wire div_en_i;
/* cellift = 32'd1 */
input div_en_i_t0;
wire div_en_i_t0;
/* src = "generated/sv2v_out.v:19482.13-19482.22" */
input div_sel_i;
wire div_sel_i;
/* cellift = 32'd1 */
input div_sel_i_t0;
wire div_sel_i_t0;
/* src = "generated/sv2v_out.v:19489.13-19489.28" */
input equal_to_zero_i;
wire equal_to_zero_i;
/* cellift = 32'd1 */
input equal_to_zero_i_t0;
wire equal_to_zero_i_t0;
/* src = "generated/sv2v_out.v:19494.21-19494.32" */
output [67:0] imd_val_d_o;
wire [67:0] imd_val_d_o;
/* cellift = 32'd1 */
output [67:0] imd_val_d_o_t0;
wire [67:0] imd_val_d_o_t0;
/* src = "generated/sv2v_out.v:19493.20-19493.31" */
input [67:0] imd_val_q_i;
wire [67:0] imd_val_q_i;
/* cellift = 32'd1 */
input [67:0] imd_val_q_i_t0;
wire [67:0] imd_val_q_i_t0;
/* src = "generated/sv2v_out.v:19495.20-19495.32" */
output [1:0] imd_val_we_o;
wire [1:0] imd_val_we_o;
/* cellift = 32'd1 */
output [1:0] imd_val_we_o_t0;
wire [1:0] imd_val_we_o_t0;
/* src = "generated/sv2v_out.v:19525.7-19525.23" */
wire is_greater_equal;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19525.7-19525.23" */
wire is_greater_equal_t0;
/* src = "generated/sv2v_out.v:19499.12-19499.22" */
reg [2:0] md_state_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19499.12-19499.22" */
reg [2:0] md_state_q_t0;
/* src = "generated/sv2v_out.v:19479.13-19479.22" */
input mult_en_i;
wire mult_en_i;
/* cellift = 32'd1 */
input mult_en_i_t0;
wire mult_en_i_t0;
/* src = "generated/sv2v_out.v:19481.13-19481.23" */
input mult_sel_i;
wire mult_sel_i;
/* cellift = 32'd1 */
input mult_sel_i_t0;
wire mult_sel_i_t0;
/* src = "generated/sv2v_out.v:19507.12-19507.27" */
reg [4:0] multdiv_count_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19507.12-19507.27" */
reg [4:0] multdiv_count_q_t0;
/* src = "generated/sv2v_out.v:19531.7-19531.17" */
wire multdiv_en;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19531.7-19531.17" */
wire multdiv_en_t0;
/* src = "generated/sv2v_out.v:19530.6-19530.18" */
wire multdiv_hold;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19530.6-19530.18" */
wire multdiv_hold_t0;
/* src = "generated/sv2v_out.v:19496.13-19496.31" */
input multdiv_ready_id_i;
wire multdiv_ready_id_i;
/* cellift = 32'd1 */
input multdiv_ready_id_i_t0;
wire multdiv_ready_id_i_t0;
/* src = "generated/sv2v_out.v:19497.21-19497.37" */
output [31:0] multdiv_result_o;
wire [31:0] multdiv_result_o;
/* cellift = 32'd1 */
output [31:0] multdiv_result_o_t0;
wire [31:0] multdiv_result_o_t0;
/* src = "generated/sv2v_out.v:19521.14-19521.27" */
wire [32:0] next_quotient;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19521.14-19521.27" */
wire [32:0] next_quotient_t0;
/* src = "generated/sv2v_out.v:19522.14-19522.28" */
wire [31:0] next_remainder;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19522.14-19522.28" */
wire [31:0] next_remainder_t0;
/* src = "generated/sv2v_out.v:19515.14-19515.23" */
wire [32:0] one_shift;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19515.14-19515.23" */
wire [32:0] one_shift_t0;
/* src = "generated/sv2v_out.v:19517.14-19517.29" */
wire [32:0] op_a_bw_last_pp;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19517.14-19517.29" */
wire [32:0] op_a_bw_last_pp_t0;
/* src = "generated/sv2v_out.v:19516.14-19516.24" */
wire [32:0] op_a_bw_pp;
/* src = "generated/sv2v_out.v:19485.20-19485.26" */
input [31:0] op_a_i;
wire [31:0] op_a_i;
/* cellift = 32'd1 */
input [31:0] op_a_i_t0;
wire [31:0] op_a_i_t0;
/* src = "generated/sv2v_out.v:19511.13-19511.25" */
reg [32:0] op_a_shift_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19511.13-19511.25" */
reg [32:0] op_a_shift_q_t0;
/* src = "generated/sv2v_out.v:19486.20-19486.26" */
input [31:0] op_b_i;
wire [31:0] op_b_i;
/* cellift = 32'd1 */
input [31:0] op_b_i_t0;
wire [31:0] op_b_i_t0;
/* src = "generated/sv2v_out.v:19509.13-19509.25" */
reg [32:0] op_b_shift_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19509.13-19509.25" */
reg [32:0] op_b_shift_q_t0;
/* src = "generated/sv2v_out.v:19524.13-19524.27" */
wire [31:0] op_numerator_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19524.13-19524.27" */
wire [31:0] op_numerator_d_t0;
/* src = "generated/sv2v_out.v:19483.19-19483.29" */
input [1:0] operator_i;
wire [1:0] operator_i;
/* cellift = 32'd1 */
input [1:0] operator_i_t0;
wire [1:0] operator_i_t0;
/* src = "generated/sv2v_out.v:19527.7-19527.22" */
wire rem_change_sign;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19527.7-19527.22" */
wire rem_change_sign_t0;
/* src = "generated/sv2v_out.v:19478.13-19478.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:19520.7-19520.13" */
wire sign_b;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:19520.7-19520.13" */
wire sign_b_t0;
/* src = "generated/sv2v_out.v:19484.19-19484.32" */
input [1:0] signed_mode_i;
wire [1:0] signed_mode_i;
/* cellift = 32'd1 */
input [1:0] signed_mode_i_t0;
wire [1:0] signed_mode_i_t0;
/* src = "generated/sv2v_out.v:19498.14-19498.21" */
output valid_o;
wire valid_o;
/* cellift = 32'd1 */
output valid_o_t0;
wire valid_o_t0;
assign op_a_bw_pp[31:0] = op_a_shift_q[31:0] & /* src = "generated/sv2v_out.v:19578.66-19578.90" */ { op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0] };
assign op_a_bw_last_pp[32] = op_a_shift_q[32] & /* src = "generated/sv2v_out.v:19578.28-19578.62" */ op_b_shift_q[0];
assign rem_change_sign = op_a_i[31] & /* src = "generated/sv2v_out.v:19579.18-19579.47" */ signed_mode_i[0];
assign sign_b = op_b_i[31] & /* src = "generated/sv2v_out.v:19580.18-19580.47" */ signed_mode_i[1];
assign div_change_sign = _0806_ & /* src = "generated/sv2v_out.v:19587.27-19587.61" */ _0767_;
assign _0044_ = op_a_i & /* src = "generated/sv2v_out.v:19604.55-19604.88" */ { op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0] };
assign _0048_ = op_a_i[31:1] & /* src = "generated/sv2v_out.v:19610.61-19610.94" */ { op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0] };
assign _0046_ = rem_change_sign & /* src = "generated/sv2v_out.v:19610.34-19610.58" */ op_b_i[0];
assign multdiv_en = _0771_ & /* src = "generated/sv2v_out.v:19702.22-19702.60" */ imd_val_we_o[0];
assign _0050_ = _0735_ & /* src = "generated/sv2v_out.v:19718.43-19718.111" */ _0773_;
assign _0052_ = ~ _0194_;
assign _0053_ = ~ _0196_;
assign _0054_ = ~ _0198_;
assign _0055_ = ~ _0200_;
assign _0056_ = ~ _0202_;
assign _0625_ = _0006_ ^ md_state_q;
assign _0626_ = _0008_ ^ multdiv_count_q;
assign _0627_ = _0014_ ^ op_b_shift_q;
assign _0628_ = _0012_ ^ op_a_shift_q;
assign _0629_ = _0020_ ^ div_by_zero_q;
assign _0474_ = _0007_ | md_state_q_t0;
assign _0478_ = _0009_ | multdiv_count_q_t0;
assign _0482_ = _0015_ | op_b_shift_q_t0;
assign _0486_ = _0013_ | op_a_shift_q_t0;
assign _0490_ = _0021_ | div_by_zero_q_t0;
assign _0475_ = _0625_ | _0474_;
assign _0479_ = _0626_ | _0478_;
assign _0483_ = _0627_ | _0482_;
assign _0487_ = _0628_ | _0486_;
assign _0491_ = _0629_ | _0490_;
assign _0241_ = { _0194_, _0194_, _0194_ } & _0007_;
assign _0244_ = { _0196_, _0196_, _0196_, _0196_, _0196_ } & _0009_;
assign _0247_ = { _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_, _0198_ } & _0015_;
assign _0250_ = { _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_, _0200_ } & _0013_;
assign _0253_ = _0202_ & _0021_;
assign _0242_ = { _0052_, _0052_, _0052_ } & md_state_q_t0;
assign _0245_ = { _0053_, _0053_, _0053_, _0053_, _0053_ } & multdiv_count_q_t0;
assign _0248_ = { _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_, _0054_ } & op_b_shift_q_t0;
assign _0251_ = { _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_, _0055_ } & op_a_shift_q_t0;
assign _0254_ = _0056_ & div_by_zero_q_t0;
assign _0243_ = _0475_ & { _0195_, _0195_, _0195_ };
assign _0246_ = _0479_ & { _0197_, _0197_, _0197_, _0197_, _0197_ };
assign _0249_ = _0483_ & { _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_, _0199_ };
assign _0252_ = _0487_ & { _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_, _0201_ };
assign _0255_ = _0491_ & _0203_;
assign _0476_ = _0241_ | _0242_;
assign _0480_ = _0244_ | _0245_;
assign _0484_ = _0247_ | _0248_;
assign _0488_ = _0250_ | _0251_;
assign _0492_ = _0253_ | _0254_;
assign _0477_ = _0476_ | _0243_;
assign _0481_ = _0480_ | _0246_;
assign _0485_ = _0484_ | _0249_;
assign _0489_ = _0488_ | _0252_;
assign _0493_ = _0492_ | _0255_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME md_state_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) md_state_q_t0 <= 3'h0;
else md_state_q_t0 <= _0477_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME multdiv_count_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) multdiv_count_q_t0 <= 5'h00;
else multdiv_count_q_t0 <= _0481_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME op_b_shift_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) op_b_shift_q_t0 <= 33'h000000000;
else op_b_shift_q_t0 <= _0485_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME op_a_shift_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) op_a_shift_q_t0 <= 33'h000000000;
else op_a_shift_q_t0 <= _0489_;
/* taint_ff = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME div_by_zero_q_t0 */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) div_by_zero_q_t0 <= 1'h0;
else div_by_zero_q_t0 <= _0493_;
assign _0211_ = op_a_shift_q_t0[31:0] & { op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0], op_b_shift_q[0] };
assign _0214_ = op_a_shift_q_t0[32] & op_b_shift_q[0];
assign _0217_ = op_a_i_t0[31] & signed_mode_i[0];
assign _0220_ = op_b_i_t0[31] & signed_mode_i[1];
assign _0223_ = _0807_ & _0767_;
assign _0226_ = op_a_i_t0 & { op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0] };
assign _0229_ = op_a_i_t0[31:1] & { op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0], op_b_i[0] };
assign _0232_ = rem_change_sign_t0 & op_b_i[0];
assign _0235_ = _0772_ & imd_val_we_o[0];
assign _0238_ = _0736_ & _0773_;
assign _0212_ = { op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0] } & op_a_shift_q[31:0];
assign _0215_ = op_b_shift_q_t0[0] & op_a_shift_q[32];
assign _0218_ = signed_mode_i_t0[0] & op_a_i[31];
assign _0221_ = signed_mode_i_t0[1] & op_b_i[31];
assign _0224_ = div_by_zero_q_t0 & _0806_;
assign _0227_ = { op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0] } & op_a_i;
assign _0230_ = { op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0] } & op_a_i[31:1];
assign _0233_ = op_b_i_t0[0] & rem_change_sign;
assign _0236_ = multdiv_hold_t0 & _0771_;
assign _0239_ = _0774_ & _0735_;
assign _0213_ = op_a_shift_q_t0[31:0] & { op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0], op_b_shift_q_t0[0] };
assign _0216_ = op_a_shift_q_t0[32] & op_b_shift_q_t0[0];
assign _0219_ = op_a_i_t0[31] & signed_mode_i_t0[0];
assign _0222_ = op_b_i_t0[31] & signed_mode_i_t0[1];
assign _0225_ = _0807_ & div_by_zero_q_t0;
assign _0228_ = op_a_i_t0 & { op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0] };
assign _0231_ = op_a_i_t0[31:1] & { op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0], op_b_i_t0[0] };
assign _0234_ = rem_change_sign_t0 & op_b_i_t0[0];
assign _0237_ = _0772_ & multdiv_hold_t0;
assign _0240_ = _0736_ & _0774_;
assign _0464_ = _0211_ | _0212_;
assign _0465_ = _0214_ | _0215_;
assign _0466_ = _0217_ | _0218_;
assign _0467_ = _0220_ | _0221_;
assign _0468_ = _0223_ | _0224_;
assign _0469_ = _0226_ | _0227_;
assign _0470_ = _0229_ | _0230_;
assign _0471_ = _0232_ | _0233_;
assign _0472_ = _0235_ | _0236_;
assign _0473_ = _0238_ | _0239_;
assign op_a_bw_last_pp_t0[31:0] = _0464_ | _0213_;
assign op_a_bw_last_pp_t0[32] = _0465_ | _0216_;
assign rem_change_sign_t0 = _0466_ | _0219_;
assign sign_b_t0 = _0467_ | _0222_;
assign div_change_sign_t0 = _0468_ | _0225_;
assign _0045_ = _0469_ | _0228_;
assign _0049_ = _0470_ | _0231_;
assign _0047_ = _0471_ | _0234_;
assign multdiv_en_t0 = _0472_ | _0237_;
assign _0051_ = _0473_ | _0240_;
assign _0057_ = | { _0041_[2], _0782_ };
assign _0058_ = | { _0041_[2], _0784_ };
assign _0059_ = | { _0750_, _0782_ };
assign _0060_ = | { op_b_shift_q_t0[31], imd_val_q_i_t0[65] };
assign _0061_ = | multdiv_count_q_t0;
assign _0576_ = imd_val_q_i_t0[65] | op_b_shift_q_t0[31];
assign _0064_ = ~ { _0782_, _0041_[2] };
assign _0065_ = ~ { _0784_, _0041_[2] };
assign _0066_ = ~ { _0782_, _0750_ };
assign _0067_ = ~ _0576_;
assign _0068_ = ~ multdiv_count_q_t0;
assign _0069_ = ~ md_state_q_t0;
assign _0070_ = ~ operator_i_t0;
assign _0257_ = { _0781_, _0164_ } & _0064_;
assign _0258_ = { _0783_, _0164_ } & _0065_;
assign _0260_ = { _0781_, _0749_ } & _0066_;
assign _0384_ = imd_val_q_i[65] & _0067_;
assign _0388_ = multdiv_count_q & _0068_;
assign _0416_ = md_state_q & _0069_;
assign _0430_ = operator_i & _0070_;
assign _0385_ = op_b_shift_q[31] & _0067_;
assign _0675_ = _0257_ == _0064_;
assign _0676_ = _0258_ == _0065_;
assign _0677_ = _0260_ == _0066_;
assign _0678_ = _0384_ == _0385_;
assign _0679_ = _0388_ == { 4'h0, _0068_[0] };
assign _0680_ = _0416_ == { 1'h0, _0069_[1:0] };
assign _0681_ = _0416_ == { _0069_[2:1], 1'h0 };
assign _0682_ = _0416_ == { _0069_[2], 2'h0 };
assign _0683_ = _0416_ == { _0069_[2], 1'h0, _0069_[0] };
assign _0684_ = _0416_ == { 1'h0, _0069_[1], 1'h0 };
assign _0685_ = _0416_ == { 2'h0, _0069_[0] };
assign _0686_ = _0430_ == { 1'h0, _0070_[0] };
assign _0687_ = _0430_ == { _0070_[1], 1'h0 };
assign _0688_ = _0430_ == _0070_;
assign _0183_ = _0675_ & _0057_;
assign _0185_ = _0676_ & _0058_;
assign _0189_ = _0677_ & _0059_;
assign _0738_ = _0678_ & _0060_;
assign _0744_ = _0679_ & _0061_;
assign _0782_ = _0680_ & _0062_;
assign _0746_ = _0681_ & _0062_;
assign _0736_ = _0682_ & _0062_;
assign _0780_ = _0683_ & _0062_;
assign _0720_[0] = _0684_ & _0062_;
assign _0786_ = _0685_ & _0062_;
assign _0750_ = _0686_ & _0063_;
assign _0778_ = _0687_ & _0063_;
assign _0776_ = _0688_ & _0063_;
/* src = "generated/sv2v_out.v:19703.2-19717.6" */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME md_state_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) md_state_q <= 3'h0;
else if (_0194_) md_state_q <= _0006_;
/* src = "generated/sv2v_out.v:19703.2-19717.6" */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME multdiv_count_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) multdiv_count_q <= 5'h00;
else if (_0196_) multdiv_count_q <= _0008_;
/* src = "generated/sv2v_out.v:19703.2-19717.6" */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME op_b_shift_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) op_b_shift_q <= 33'h000000000;
else if (_0198_) op_b_shift_q <= _0014_;
/* src = "generated/sv2v_out.v:19703.2-19717.6" */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME op_a_shift_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) op_a_shift_q <= 33'h000000000;
else if (_0200_) op_a_shift_q <= _0012_;
/* src = "generated/sv2v_out.v:19703.2-19717.6" */
/* PC_TAINT_INFO MODULE_NAME ibex_multdiv_slow */
/* PC_TAINT_INFO STATE_NAME div_by_zero_q */
always_ff @(posedge clk_i, negedge rst_ni)
if (!rst_ni) div_by_zero_q <= 1'h0;
else if (_0202_) div_by_zero_q <= _0020_;
assign _0389_ = data_ind_timing_i_t0 & _0739_;
assign _0392_ = data_ind_timing_i_t0 & equal_to_zero_i;
assign _0395_ = data_ind_timing_i_t0 & _0741_;
assign _0390_ = _0740_ & _0757_;
assign _0393_ = equal_to_zero_i_t0 & _0757_;
assign _0396_ = _0742_ & _0757_;
assign _0391_ = data_ind_timing_i_t0 & _0740_;
assign _0394_ = data_ind_timing_i_t0 & equal_to_zero_i_t0;
assign _0397_ = data_ind_timing_i_t0 & _0742_;
assign _0577_ = _0389_ | _0390_;
assign _0578_ = _0392_ | _0393_;
assign _0579_ = _0395_ | _0396_;
assign _0752_ = _0577_ | _0391_;
assign _0754_ = _0578_ | _0394_;
assign _0756_ = _0579_ | _0397_;
assign _0071_ = | { _0784_, _0782_ };
assign _0072_ = | { _0720_[0], _0784_, _0782_ };
assign _0073_ = | { _0786_, _0784_, _0782_ };
assign _0074_ = | { _0776_, _0748_, _0750_ };
assign _0075_ = | { _0720_[0], _0784_ };
assign _0076_ = | { _0748_, _0750_ };
assign _0077_ = | { _0778_, _0776_, _0750_ };
assign _0078_ = | { _0778_, _0776_ };
assign _0079_ = | { _0720_[0], _0780_, _0786_, _0784_ };
assign _0080_ = | { _0780_, _0782_, _0736_ };
assign _0081_ = | { sign_b_t0, op_b_i_t0[31:1] };
assign _0082_ = | op_b_shift_q_t0[32:1];
assign _0062_ = | md_state_q_t0;
assign _0063_ = | operator_i_t0;
assign _0083_ = ~ { _0784_, _0782_ };
assign _0084_ = ~ { _0720_[0], _0784_, _0782_ };
assign _0085_ = ~ { _0786_, _0784_, _0782_ };
assign _0086_ = ~ { _0776_, _0750_, _0748_ };
assign _0087_ = ~ { _0720_[0], _0784_ };
assign _0088_ = ~ { _0750_, _0748_ };
assign _0089_ = ~ { _0778_, _0776_, _0750_ };
assign _0090_ = ~ { _0778_, _0776_ };
assign _0091_ = ~ { _0720_[0], _0786_, _0784_, _0780_ };
assign _0092_ = ~ { _0782_, _0780_, _0736_ };
assign _0093_ = ~ { 1'h0, sign_b_t0, op_b_i_t0[31:1] };
assign _0094_ = ~ { 1'h0, op_b_shift_q_t0[32:1] };
assign _0256_ = { _0783_, _0781_ } & _0083_;
assign _0259_ = { _0787_, _0783_, _0781_ } & _0084_;
assign _0261_ = { _0785_, _0783_, _0781_ } & _0085_;
assign _0262_ = { _0775_, _0749_, _0747_ } & _0086_;
assign _0263_ = { _0787_, _0783_ } & _0087_;
assign _0264_ = { _0749_, _0747_ } & _0088_;
assign _0265_ = { _0777_, _0775_, _0749_ } & _0089_;
assign _0266_ = { _0777_, _0775_ } & _0090_;
assign _0267_ = { _0787_, _0785_, _0783_, _0779_ } & _0091_;
assign _0277_ = { _0781_, _0779_, _0735_ } & _0092_;
assign _0386_ = { 1'h0, sign_b, op_b_i[31:1] } & _0093_;
assign _0387_ = { 1'h0, op_b_shift_q[32:1] } & _0094_;
assign _0095_ = ! _0256_;
assign _0096_ = ! _0259_;
assign _0097_ = ! _0261_;
assign _0098_ = ! _0262_;
assign _0099_ = ! _0263_;
assign _0100_ = ! _0264_;
assign _0101_ = ! _0265_;
assign _0102_ = ! _0266_;
assign _0103_ = ! _0267_;
assign _0104_ = ! _0277_;
assign _0105_ = ! _0386_;
assign _0106_ = ! _0387_;
assign _0107_ = ! _0416_;
assign _0108_ = ! _0430_;
assign _0181_ = _0095_ & _0071_;
assign _0187_ = _0096_ & _0072_;
assign _0191_ = _0097_ & _0073_;
assign _0193_ = _0098_ & _0074_;
assign _0208_ = _0099_ & _0075_;
assign _0206_ = _0100_ & _0076_;
assign _0210_ = _0101_ & _0077_;
assign _0041_[2] = _0102_ & _0078_;
assign _0166_ = _0103_ & _0079_;
assign _0168_ = _0104_ & _0080_;
assign _0740_ = _0105_ & _0081_;
assign _0742_ = _0106_ & _0082_;
assign _0784_ = _0107_ & _0062_;
assign _0748_ = _0108_ & _0063_;
assign _0109_ = ~ mult_sel_i;
assign _0110_ = ~ _0755_;
assign _0111_ = ~ div_sel_i;
assign _0112_ = ~ _0743_;
assign _0398_ = mult_sel_i_t0 & _0111_;
assign _0401_ = _0756_ & _0112_;
assign _0399_ = div_sel_i_t0 & _0109_;
assign _0402_ = _0744_ & _0110_;
assign _0400_ = mult_sel_i_t0 & div_sel_i_t0;
assign _0403_ = _0756_ & _0744_;
assign _0580_ = _0398_ | _0399_;
assign _0581_ = _0401_ | _0402_;
assign _0759_ = _0580_ | _0400_;
assign _0761_ = _0581_ | _0403_;
assign _0113_ = ~ { _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_ };
assign _0114_ = ~ { _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_ };
assign _0115_ = ~ _0164_;
assign _0116_ = ~ { _0164_, _0164_, _0164_ };
assign _0117_ = ~ { _0209_, _0209_, _0209_ };
assign _0118_ = ~ { _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_ };
assign _0119_ = ~ { _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_ };
assign _0120_ = ~ { _0749_, _0749_, _0749_ };
assign _0121_ = ~ { _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_ };
assign _0122_ = ~ { _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_ };
assign _0123_ = ~ { _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_ };
assign _0124_ = ~ { _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_ };
assign _0125_ = ~ { _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_ };
assign _0126_ = ~ { _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_ };
assign _0127_ = ~ { _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_ };
assign _0128_ = ~ { _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_ };
assign _0129_ = ~ { _0735_, _0735_, _0735_ };
assign _0130_ = ~ { _0779_, _0779_, _0779_ };
assign _0131_ = ~ { _0460_, _0460_, _0460_ };
assign _0132_ = ~ { _0167_, _0167_, _0167_ };
assign _0133_ = ~ _0745_;
assign _0134_ = ~ { _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_ };
assign _0135_ = ~ _0777_;
assign _0136_ = ~ { _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_ };
assign _0137_ = ~ { _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_ };
assign _0138_ = ~ { _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_ };
assign _0139_ = ~ { _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_, _0165_ };
assign _0140_ = ~ _0737_;
assign _0141_ = ~ { is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal };
assign _0142_ = ~ { is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal };
assign _0143_ = ~ { rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign };
assign _0144_ = ~ { sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b };
assign _0145_ = ~ { div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign };
assign _0146_ = ~ { rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign };
assign _0147_ = ~ { div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i };
assign _0502_ = { _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_ } | _0113_;
assign _0505_ = { _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_ } | _0114_;
assign _0508_ = _0041_[2] | _0115_;
assign _0509_ = { _0041_[2], _0041_[2], _0041_[2] } | _0116_;
assign _0513_ = { _0210_, _0210_, _0210_ } | _0117_;
assign _0516_ = { _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2] } | _0118_;
assign _0519_ = { _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_ } | _0119_;
assign _0523_ = { _0750_, _0750_, _0750_ } | _0120_;
assign _0526_ = { _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_ } | _0121_;
assign _0531_ = { _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_ } | _0122_;
assign _0533_ = { _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_ } | _0123_;
assign _0536_ = { _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0] } | _0124_;
assign _0540_ = { _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_ } | _0125_;
assign _0543_ = { _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_ } | _0126_;
assign _0546_ = { _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_ } | _0127_;
assign _0550_ = { _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_ } | _0128_;
assign _0553_ = { _0736_, _0736_, _0736_ } | _0129_;
assign _0556_ = { _0780_, _0780_, _0780_ } | _0130_;
assign _0558_ = { _0461_, _0461_, _0461_ } | _0131_;
assign _0561_ = { _0168_, _0168_, _0168_ } | _0132_;
assign _0565_ = _0746_ | _0133_;
assign _0570_ = { _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_ } | _0134_;
assign _0588_ = { _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_ } | _0136_;
assign _0592_ = { _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_ } | _0137_;
assign _0595_ = { _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_ } | _0138_;
assign _0598_ = { _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_ } | _0139_;
assign _0601_ = _0738_ | _0140_;
assign _0604_ = { is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0 } | _0141_;
assign _0607_ = { is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0 } | _0142_;
assign _0610_ = { rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0 } | _0143_;
assign _0613_ = { sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0 } | _0144_;
assign _0616_ = { div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0 } | _0145_;
assign _0619_ = { rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0 } | _0146_;
assign _0622_ = { div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0 } | _0147_;
assign _0503_ = { _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_ } | { _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_, _0777_ };
assign _0506_ = { _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_ } | { _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_, _0775_ };
assign _0510_ = { _0041_[2], _0041_[2], _0041_[2] } | { _0164_, _0164_, _0164_ };
assign _0514_ = { _0210_, _0210_, _0210_ } | { _0209_, _0209_, _0209_ };
assign _0517_ = { _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2] } | { _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_, _0164_ };
assign _0520_ = { _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_ } | { _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_, _0749_ };
assign _0527_ = { _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_ } | { _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_, _0458_ };
assign _0530_ = { _0782_, _0782_, _0782_, _0782_, _0782_ } | { _0781_, _0781_, _0781_, _0781_, _0781_ };
assign _0532_ = { _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_ } | { _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_ };
assign _0534_ = { _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_ } | { _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_, _0781_ };
assign _0537_ = { _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0] } | { _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_, _0787_ };
assign _0541_ = { _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_ } | { _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_, _0735_ };
assign _0544_ = { _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_ } | { _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_, _0779_ };
assign _0547_ = { _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_ } | { _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_, _0783_ };
assign _0551_ = { _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_ } | { _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_, _0167_ };
assign _0554_ = { _0736_, _0736_, _0736_ } | { _0735_, _0735_, _0735_ };
assign _0557_ = { _0784_, _0784_, _0784_ } | { _0783_, _0783_, _0783_ };
assign _0559_ = { _0461_, _0461_, _0461_ } | { _0460_, _0460_, _0460_ };
assign _0562_ = { _0168_, _0168_, _0168_ } | { _0167_, _0167_, _0167_ };
assign _0564_ = _0736_ | _0735_;
assign _0566_ = _0746_ | _0745_;
assign _0571_ = { _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_ } | { _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_, _0462_ };
assign _0586_ = { _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_, _0206_ } | { _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_, _0205_ };
assign _0587_ = _0778_ | _0777_;
assign _0589_ = { _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_ } | { _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_, _0785_ };
assign _0591_ = _0759_ | _0758_;
assign _0593_ = { _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_ } | { _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_ };
assign _0596_ = { _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_ } | { _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_, _0758_ };
assign _0602_ = _0738_ | _0737_;
assign _0605_ = { is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0 } | { is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal };
assign _0608_ = { is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0 } | { is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal, is_greater_equal };
assign _0611_ = { rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0 } | { rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign };
assign _0614_ = { sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0 } | { sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b, sign_b };
assign _0617_ = { div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0 } | { div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign, div_change_sign };
assign _0620_ = { rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0 } | { rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign, rem_change_sign };
assign _0623_ = { div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0 } | { div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i, div_en_i };
assign _0278_ = imd_val_q_i_t0[66:34] & _0502_;
assign _0281_ = _0692_ & _0505_;
assign _0284_ = multdiv_ready_id_i_t0 & _0508_;
assign _0286_ = alu_adder_ext_i_t0[32:0] & _0502_;
assign _0289_ = _0694_ & _0505_;
assign _0292_ = { _0761_, _0761_, _0761_ } & _0513_;
assign _0295_ = { op_a_shift_q_t0[31:0], 1'h0 } & _0516_;
assign _0298_ = alu_adder_ext_i_t0[32:0] & _0519_;
assign _0301_ = _0696_ & _0516_;
assign _0304_ = { _0752_, _0752_, _0752_ } & _0523_;
assign _0306_ = _0698_ & _0509_;
assign _0311_ = { _0047_, _0045_ } & _0519_;
assign _0314_ = _0702_ & _0526_;
assign _0317_ = { op_a_i_t0, 1'h0 } & _0519_;
assign _0322_ = _0027_ & _0531_;
assign _0324_ = _0704_ & _0533_;
assign _0327_ = _0029_ & _0536_;
assign _0330_ = _0706_ & _0533_;
assign _0333_ = _0031_ & _0540_;
assign _0336_ = _0708_ & _0543_;
assign _0339_ = imd_val_q_i_t0[66:34] & _0546_;
assign _0342_ = _0712_ & _0536_;
assign _0345_ = _0714_ & _0550_;
assign _0348_ = _0033_ & _0553_;
assign _0351_ = _0716_ & _0556_;
assign _0355_ = _0722_ & _0558_;
assign _0358_ = _0724_ & _0561_;
assign _0363_ = _0726_ & _0565_;
assign _0366_ = { op_b_i_t0, 1'h0 } & _0543_;
assign _0369_ = { op_b_shift_q_t0[31:0], 1'h0 } & _0531_;
assign _0372_ = _0730_ & _0570_;
assign _0375_ = op_a_bw_last_pp_t0 & _0519_;
assign _0378_ = _0732_ & _0516_;
assign _0381_ = imd_val_q_i_t0[66:34] & _0516_;
assign _0417_ = imd_val_q_i_t0[31:0] & _0588_;
assign _0422_ = imd_val_q_i_t0[31:0] & _0592_;
assign _0425_ = imd_val_q_i_t0[66:34] & _0595_;
assign _0428_ = { imd_val_q_i_t0[65:34], 1'h0 } & _0598_;
assign _0431_ = op_a_bw_last_pp_t0 & _0540_;
assign _0434_ = imd_val_q_i_t0[65] & _0601_;
assign _0437_ = imd_val_q_i_t0[65:34] & _0604_;
assign _0440_ = op_a_shift_q_t0 & _0607_;
assign _0443_ = op_a_i_t0 & _0610_;
assign _0446_ = { 1'h0, op_b_i_t0 } & _0613_;
assign _0449_ = imd_val_q_i_t0[66:34] & _0616_;
assign _0452_ = imd_val_q_i_t0[66:34] & _0619_;
assign _0455_ = alu_adder_ext_i_t0[31:0] & _0622_;
assign _0279_ = _0803_ & _0503_;
assign _0282_ = _0805_ & _0506_;
assign _0287_ = next_quotient_t0 & _0503_;
assign _0290_ = { 1'h0, next_remainder_t0 } & _0506_;
assign _0293_ = { _0744_, _0744_, _0744_ } & _0514_;
assign _0296_ = next_quotient_t0 & _0517_;
assign _0299_ = alu_adder_ext_i_t0[33:1] & _0520_;
assign _0302_ = { next_remainder_t0, _0789_ } & _0517_;
assign _0307_ = { _0754_, _0754_, _0754_ } & _0510_;
assign _0309_ = { rem_change_sign_t0, op_a_i_t0 } & _0506_;
assign _0312_ = { 1'h0, _0047_, _0049_ } & _0520_;
assign _0315_ = _0700_ & _0527_;
assign _0318_ = { rem_change_sign_t0, op_a_i_t0 } & _0520_;
assign _0320_ = _0791_ & _0530_;
assign _0325_ = _0035_ & _0534_;
assign _0328_ = _0799_ & _0537_;
assign _0331_ = _0037_ & _0534_;
assign _0334_ = _0039_ & _0541_;
assign _0337_ = _0043_ & _0544_;
assign _0340_ = _0019_ & _0547_;
assign _0343_ = { 32'h00000000, imd_val_q_i_t0[31] } & _0537_;
assign _0346_ = _0710_ & _0551_;
assign _0349_ = { _0041_[2], 1'h0, _0041_[2] } & _0554_;
assign _0353_ = _0023_ & _0557_;
assign _0356_ = { 2'h0, _0720_[0] } & _0559_;
assign _0359_ = _0718_ & _0562_;
assign _0361_ = _0025_ & _0564_;
assign _0364_ = multdiv_ready_id_i_t0 & _0566_;
assign _0367_ = { imd_val_q_i_t0[65:34], 1'h0 } & _0544_;
assign _0370_ = { op_a_i_t0, 1'h0 } & _0532_;
assign _0373_ = _0728_ & _0571_;
assign _0376_ = _0793_ & _0520_;
assign _0379_ = _0005_ & _0517_;
assign _0382_ = _0003_ & _0517_;
assign _0037_ = { 1'h0, op_b_shift_q_t0[32:1] } & _0586_;
assign _0029_ = { 1'h0, sign_b_t0, op_b_i_t0[31:1] } & _0586_;
assign _0021_ = equal_to_zero_i_t0 & _0587_;
assign _0418_ = _0797_ & _0589_;
assign _0420_ = _0011_ & _0591_;
assign _0423_ = _0017_ & _0593_;
assign _0426_ = _0001_ & _0596_;
assign _0432_ = op_a_bw_last_pp_t0 & _0541_;
assign _0435_ = alu_adder_ext_i_t0[32] & _0602_;
assign _0438_ = alu_adder_ext_i_t0[32:1] & _0605_;
assign _0441_ = _0770_ & _0608_;
assign _0444_ = alu_adder_i_t0 & _0611_;
assign _0447_ = { 1'h0, alu_adder_i_t0 } & _0614_;
assign _0450_ = { 1'h0, alu_adder_i_t0 } & _0617_;
assign _0453_ = { 1'h0, alu_adder_i_t0 } & _0620_;
assign _0456_ = imd_val_q_i_t0[65:34] & _0623_;
assign _0504_ = _0278_ | _0279_;
assign _0507_ = _0281_ | _0282_;
assign _0511_ = _0286_ | _0287_;
assign _0512_ = _0289_ | _0290_;
assign _0515_ = _0292_ | _0293_;
assign _0518_ = _0295_ | _0296_;
assign _0521_ = _0298_ | _0299_;
assign _0522_ = _0301_ | _0302_;
assign _0524_ = _0306_ | _0307_;
assign _0525_ = _0311_ | _0312_;
assign _0528_ = _0314_ | _0315_;
assign _0529_ = _0317_ | _0318_;
assign _0535_ = _0324_ | _0325_;
assign _0538_ = _0327_ | _0328_;
assign _0539_ = _0330_ | _0331_;
assign _0542_ = _0333_ | _0334_;
assign _0545_ = _0336_ | _0337_;
assign _0548_ = _0339_ | _0340_;
assign _0549_ = _0342_ | _0343_;
assign _0552_ = _0345_ | _0346_;
assign _0555_ = _0348_ | _0349_;
assign _0560_ = _0355_ | _0356_;
assign _0563_ = _0358_ | _0359_;
assign _0567_ = _0363_ | _0364_;
assign _0568_ = _0366_ | _0367_;
assign _0569_ = _0369_ | _0370_;
assign _0572_ = _0372_ | _0373_;
assign _0573_ = _0375_ | _0376_;
assign _0574_ = _0378_ | _0379_;
assign _0575_ = _0381_ | _0382_;
assign _0590_ = _0417_ | _0418_;
assign _0594_ = _0422_ | _0423_;
assign _0597_ = _0425_ | _0426_;
assign _0600_ = _0431_ | _0432_;
assign _0603_ = _0434_ | _0435_;
assign _0606_ = _0437_ | _0438_;
assign _0609_ = _0440_ | _0441_;
assign _0612_ = _0443_ | _0444_;
assign _0615_ = _0446_ | _0447_;
assign _0618_ = _0449_ | _0450_;
assign _0621_ = _0452_ | _0453_;
assign _0624_ = _0455_ | _0456_;
assign _0630_ = imd_val_q_i[66:34] ^ _0802_;
assign _0631_ = _0691_ ^ _0804_;
assign _0633_ = alu_adder_ext_i[32:0] ^ next_quotient;
assign _0634_ = _0693_ ^ { 1'h0, next_remainder };
assign _0635_ = _0800_ ^ _0801_;
assign _0636_ = { op_a_shift_q[31:0], 1'h0 } ^ next_quotient;
assign _0637_ = alu_adder_ext_i[32:0] ^ alu_adder_ext_i[33:1];
assign _0638_ = _0695_ ^ { next_remainder, _0788_ };
assign _0640_ = _0697_ ^ _0795_;
assign _0641_ = { _0768_, _0044_ } ^ { 1'h1, _0768_, _0048_ };
assign _0642_ = _0701_ ^ _0699_;
assign _0643_ = { op_a_i, 1'h0 } ^ { rem_change_sign, op_a_i };
assign _0644_ = _0703_ ^ _0034_;
assign _0645_ = _0028_ ^ _0798_;
assign _0646_ = _0705_ ^ _0036_;
assign _0647_ = _0030_ ^ _0038_;
assign _0648_ = _0707_ ^ _0042_;
assign _0649_ = imd_val_q_i[66:34] ^ _0018_;
assign _0650_ = _0711_ ^ { 32'h00000000, imd_val_q_i[31] };
assign _0651_ = _0713_ ^ _0709_;
assign _0652_ = _0032_ ^ _0040_;
assign _0654_ = _0721_ ^ _0719_;
assign _0655_ = _0723_ ^ _0717_;
assign _0656_ = _0725_ ^ _0632_;
assign _0657_ = { _0762_, 1'h1 } ^ { _0764_, 1'h1 };
assign _0658_ = { _0765_, 1'h1 } ^ { _0763_, 1'h1 };
assign _0659_ = _0729_ ^ _0727_;
assign _0660_ = op_a_bw_pp ^ _0792_;
assign _0661_ = _0731_ ^ _0004_;
assign _0662_ = imd_val_q_i[66:34] ^ _0002_;
assign _0663_ = imd_val_q_i[31:0] ^ _0796_;
assign _0664_ = imd_val_q_i[31:0] ^ _0016_;
assign _0665_ = imd_val_q_i[66:34] ^ _0000_;
assign _0667_ = op_a_bw_pp ^ op_a_bw_last_pp;
assign _0668_ = imd_val_q_i[65] ^ _0766_;
assign _0669_ = imd_val_q_i[65:34] ^ alu_adder_ext_i[32:1];
assign _0670_ = op_a_shift_q ^ _0769_;
assign _0671_ = op_a_i ^ alu_adder_i;
assign _0672_ = { 1'h0, op_b_i } ^ { 1'h0, alu_adder_i };
assign _0673_ = imd_val_q_i[66:34] ^ { 1'h0, alu_adder_i };
assign _0674_ = alu_adder_ext_i[31:0] ^ imd_val_q_i[65:34];
assign _0280_ = { _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_ } & _0630_;
assign _0283_ = { _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_ } & _0631_;
assign _0285_ = _0041_[2] & _0632_;
assign _0288_ = { _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_, _0778_ } & _0633_;
assign _0291_ = { _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_ } & _0634_;
assign _0294_ = { _0210_, _0210_, _0210_ } & _0635_;
assign _0297_ = { _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2] } & _0636_;
assign _0300_ = { _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_ } & _0637_;
assign _0303_ = { _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2] } & _0638_;
assign _0305_ = { _0750_, _0750_, _0750_ } & { _0639_[2], _0148_ };
assign _0308_ = { _0041_[2], _0041_[2], _0041_[2] } & _0640_;
assign _0310_ = { _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_, _0776_ } & _0151_;
assign _0313_ = { _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_ } & _0641_;
assign _0316_ = { _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_, _0459_ } & _0642_;
assign _0319_ = { _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_ } & _0643_;
assign _0321_ = { _0782_, _0782_, _0782_, _0782_, _0782_ } & _0150_;
assign _0323_ = { _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_ } & _0026_;
assign _0326_ = { _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_ } & _0644_;
assign _0329_ = { _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0] } & _0645_;
assign _0332_ = { _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_, _0782_ } & _0646_;
assign _0335_ = { _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_ } & _0647_;
assign _0338_ = { _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_ } & _0648_;
assign _0341_ = { _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_, _0784_ } & _0649_;
assign _0344_ = { _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0], _0720_[0] } & _0650_;
assign _0347_ = { _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_, _0168_ } & _0651_;
assign _0350_ = { _0736_, _0736_, _0736_ } & _0652_;
assign _0352_ = { _0780_, _0780_, _0780_ } & { _0149_, _0653_[0] };
assign _0354_ = { _0784_, _0784_, _0784_ } & _0022_;
assign _0357_ = { _0461_, _0461_, _0461_ } & _0654_;
assign _0360_ = { _0168_, _0168_, _0168_ } & _0655_;
assign _0362_ = _0736_ & _0024_;
assign _0365_ = _0746_ & _0656_;
assign _0368_ = { _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_, _0780_ } & _0657_;
assign _0371_ = { _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_ } & _0658_;
assign _0374_ = { _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_, _0463_ } & _0659_;
assign _0377_ = { _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_, _0750_ } & _0660_;
assign _0380_ = { _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2] } & _0661_;
assign _0383_ = { _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2], _0041_[2] } & _0662_;
assign _0419_ = { _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_, _0786_ } & _0663_;
assign _0421_ = _0759_ & _0010_;
assign _0424_ = { _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_ } & _0664_;
assign _0427_ = { _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_, _0759_ } & _0665_;
assign _0429_ = { _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_, _0166_ } & { imd_val_q_i[65:34], 1'h0 };
assign _0433_ = { _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_, _0736_ } & _0667_;
assign _0436_ = _0738_ & _0668_;
assign _0439_ = { is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0 } & _0669_;
assign _0442_ = { is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0, is_greater_equal_t0 } & _0670_;
assign _0445_ = { rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0 } & _0671_;
assign _0448_ = { sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0, sign_b_t0 } & _0672_;
assign _0451_ = { div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0, div_change_sign_t0 } & _0673_;
assign _0454_ = { rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0, rem_change_sign_t0 } & _0673_;
assign _0457_ = { div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0, div_en_i_t0 } & _0674_;
assign _0692_ = _0280_ | _0504_;
assign _0043_ = _0283_ | _0507_;
assign _0025_ = _0285_ | _0284_;
assign _0694_ = _0288_ | _0511_;
assign _0039_ = _0291_ | _0512_;
assign _0033_ = _0294_ | _0515_;
assign _0035_ = _0297_ | _0518_;
assign _0696_ = _0300_ | _0521_;
assign _0031_ = _0303_ | _0522_;
assign _0698_ = _0305_ | _0304_;
assign _0023_ = _0308_ | _0524_;
assign _0700_ = _0310_ | _0309_;
assign _0702_ = _0313_ | _0525_;
assign _0019_ = _0316_ | _0528_;
assign _0027_ = _0319_ | _0529_;
assign _0009_ = _0321_ | _0320_;
assign _0704_ = _0323_ | _0322_;
assign _0013_ = _0326_ | _0535_;
assign _0706_ = _0329_ | _0538_;
assign _0015_ = _0332_ | _0539_;
assign _0708_ = _0335_ | _0542_;
assign _0710_ = _0338_ | _0545_;
assign _0712_ = _0341_ | _0548_;
assign _0714_ = _0344_ | _0549_;
assign _0001_ = _0347_ | _0552_;
assign _0716_ = _0350_ | _0555_;
assign _0718_ = _0352_ | _0351_;
assign _0722_ = _0354_ | _0353_;
assign _0724_ = _0357_ | _0560_;
assign _0007_ = _0360_ | _0563_;
assign _0726_ = _0362_ | _0361_;
assign _0011_ = _0365_ | _0567_;
assign _0728_ = _0368_ | _0568_;
assign _0730_ = _0371_ | _0569_;
assign _0005_ = _0374_ | _0572_;
assign _0732_ = _0377_ | _0573_;
assign alu_operand_b_o_t0 = _0380_ | _0574_;
assign alu_operand_a_o_t0 = _0383_ | _0575_;
assign _0017_ = _0419_ | _0590_;
assign multdiv_hold_t0 = _0421_ | _0420_;
assign op_numerator_d_t0 = _0424_ | _0594_;
assign accum_window_d_t0 = _0427_ | _0597_;
assign _0003_ = _0429_ | _0428_;
assign _0793_ = _0433_ | _0600_;
assign is_greater_equal_t0 = _0436_ | _0603_;
assign next_remainder_t0 = _0439_ | _0606_;
assign next_quotient_t0 = _0442_ | _0609_;
assign _0797_ = _0445_ | _0612_;
assign _0799_ = _0448_ | _0615_;
assign _0803_ = _0451_ | _0618_;
assign _0805_ = _0454_ | _0621_;
assign multdiv_result_o_t0 = _0457_ | _0624_;
assign _0180_ = | { _0783_, _0781_ };
assign _0182_ = { _0781_, _0164_ } != 2'h3;
assign _0184_ = { _0783_, _0164_ } != 2'h3;
assign _0186_ = | { _0787_, _0783_, _0781_ };
assign _0188_ = { _0781_, _0749_ } != 2'h3;
assign _0190_ = | { _0785_, _0783_, _0781_ };
assign _0192_ = ~ _0204_;
assign _0194_ = & { _0758_, multdiv_en };
assign _0196_ = & { _0180_, _0758_, multdiv_en };
assign _0198_ = & { _0758_, multdiv_en, _0182_, _0184_, _0186_ };
assign _0200_ = & { _0758_, multdiv_en, _0184_, _0188_, _0190_ };
assign _0202_ = & { _0783_, _0758_, multdiv_en, _0192_ };
assign _0148_ = ~ _0794_[1:0];
assign _0149_ = ~ _0715_[2:1];
assign _0150_ = ~ _0790_;
assign _0151_ = ~ { rem_change_sign, op_a_i };
assign _0204_ = | { _0775_, _0749_, _0747_ };
assign _0207_ = | { _0787_, _0783_ };
assign _0205_ = | { _0749_, _0747_ };
assign _0209_ = | { _0777_, _0775_, _0749_ };
assign _0152_ = ~ _0785_;
assign _0153_ = ~ _0207_;
assign _0154_ = ~ op_a_shift_q;
assign _0155_ = ~ mult_en_i;
assign _0156_ = ~ _0747_;
assign _0157_ = ~ _0775_;
assign _0158_ = ~ _0787_;
assign _0159_ = ~ _0779_;
assign _0160_ = ~ one_shift;
assign _0161_ = ~ div_en_i;
assign _0162_ = ~ _0749_;
assign _0163_ = ~ _0050_;
assign _0268_ = _0778_ & _0157_;
assign _0271_ = _0786_ & _0158_;
assign _0274_ = _0208_ & _0159_;
assign _0404_ = op_a_shift_q_t0 & _0160_;
assign _0407_ = mult_en_i_t0 & _0161_;
assign _0410_ = _0748_ & _0162_;
assign _0413_ = _0746_ & _0163_;
assign _0269_ = _0776_ & _0135_;
assign _0272_ = _0720_[0] & _0152_;
assign _0275_ = _0780_ & _0153_;
assign _0405_ = one_shift_t0 & _0154_;
assign _0408_ = div_en_i_t0 & _0155_;
assign _0411_ = _0750_ & _0156_;
assign _0414_ = _0051_ & _0133_;
assign _0270_ = _0778_ & _0776_;
assign _0273_ = _0786_ & _0720_[0];
assign _0276_ = _0208_ & _0780_;
assign _0406_ = op_a_shift_q_t0 & one_shift_t0;
assign _0409_ = mult_en_i_t0 & div_en_i_t0;
assign _0412_ = _0748_ & _0750_;
assign _0415_ = _0746_ & _0051_;
assign _0499_ = _0268_ | _0269_;
assign _0500_ = _0271_ | _0272_;
assign _0501_ = _0274_ | _0275_;
assign _0582_ = _0404_ | _0405_;
assign _0583_ = _0407_ | _0408_;
assign _0584_ = _0410_ | _0411_;
assign _0585_ = _0413_ | _0414_;
assign _0459_ = _0499_ | _0270_;
assign _0461_ = _0500_ | _0273_;
assign _0463_ = _0501_ | _0276_;
assign _0770_ = _0582_ | _0406_;
assign _0772_ = _0583_ | _0409_;
assign _0774_ = _0584_ | _0412_;
assign valid_o_t0 = _0585_ | _0415_;
assign _0164_ = | { _0777_, _0775_ };
assign _0165_ = | { _0787_, _0785_, _0783_, _0779_ };
assign _0458_ = _0777_ | _0775_;
assign _0460_ = _0785_ | _0787_;
assign _0462_ = _0207_ | _0779_;
assign _0167_ = | { _0781_, _0779_, _0735_ };
assign _0691_ = _0777_ ? _0802_ : imd_val_q_i[66:34];
assign _0042_ = _0775_ ? _0804_ : _0691_;
assign _0024_ = _0164_ ? 1'h0 : _0632_;
assign _0040_ = _0164_ ? 3'h5 : 3'h0;
assign _0693_ = _0777_ ? next_quotient : alu_adder_ext_i[32:0];
assign _0038_ = _0775_ ? { 1'h0, next_remainder } : _0693_;
assign _0032_ = _0209_ ? _0801_ : _0800_;
assign _0034_ = _0164_ ? next_quotient : { op_a_shift_q[31:0], 1'h0 };
assign _0695_ = _0749_ ? alu_adder_ext_i[33:1] : alu_adder_ext_i[32:0];
assign _0030_ = _0164_ ? { next_remainder, _0788_ } : _0695_;
assign _0697_ = _0749_ ? 3'h3 : { _0639_[2], _0794_[1:0] };
assign _0022_ = _0164_ ? _0795_ : _0697_;
assign _0699_ = _0775_ ? { rem_change_sign, op_a_i } : 33'h1ffffffff;
assign _0701_ = _0749_ ? { 1'h1, _0768_, _0048_ } : { _0768_, _0044_ };
assign _0018_ = _0458_ ? _0699_ : _0701_;
assign _0026_ = _0749_ ? { rem_change_sign, op_a_i } : { op_a_i, 1'h0 };
assign _0008_ = _0781_ ? _0790_ : 5'h1f;
assign _0703_ = _0785_ ? 33'h000000000 : _0026_;
assign _0012_ = _0781_ ? _0034_ : _0703_;
assign _0705_ = _0787_ ? _0798_ : _0028_;
assign _0014_ = _0781_ ? _0036_ : _0705_;
assign _0707_ = _0735_ ? _0038_ : _0030_;
assign _0709_ = _0779_ ? _0042_ : _0707_;
assign _0711_ = _0783_ ? _0018_ : imd_val_q_i[66:34];
assign _0713_ = _0787_ ? { 32'h00000000, imd_val_q_i[31] } : _0711_;
assign _0000_ = _0167_ ? _0709_ : _0713_;
assign { _0715_[2:1], _0653_[0] } = _0735_ ? _0040_ : _0032_;
assign _0717_ = _0779_ ? 3'h6 : { _0715_[2:1], _0653_[0] };
assign _0719_ = _0787_ ? 3'h3 : 3'h2;
assign _0721_ = _0783_ ? _0022_ : 3'h0;
assign _0723_ = _0460_ ? _0719_ : _0721_;
assign _0006_ = _0167_ ? _0717_ : _0723_;
assign _0725_ = _0735_ ? _0024_ : 1'h0;
assign _0010_ = _0745_ ? _0632_ : _0725_;
assign _0727_ = _0779_ ? { _0764_, 1'h1 } : { _0762_, 1'h1 };
assign _0729_ = _0785_ ? { _0763_, 1'h1 } : { _0765_, 1'h1 };
assign _0004_ = _0462_ ? _0727_ : _0729_;
assign _0731_ = _0749_ ? _0792_ : op_a_bw_pp;
assign alu_operand_b_o = _0164_ ? _0004_ : _0731_;
assign alu_operand_a_o = _0164_ ? _0002_ : imd_val_q_i[66:34];
assign _0169_ = | { _0759_, multdiv_en_t0 };
assign _0170_ = | { _0759_, _0181_, multdiv_en_t0 };
assign _0171_ = | { _0759_, _0187_, _0185_, _0183_, multdiv_en_t0 };
assign _0172_ = | { _0759_, _0191_, _0189_, _0185_, multdiv_en_t0 };
assign _0173_ = | { _0759_, _0193_, _0784_, multdiv_en_t0 };
assign _0494_ = { _0758_, multdiv_en } | { _0759_, multdiv_en_t0 };
assign _0495_ = { _0180_, _0758_, multdiv_en } | { _0181_, _0759_, multdiv_en_t0 };
assign _0496_ = { _0758_, multdiv_en, _0182_, _0184_, _0186_ } | { _0759_, multdiv_en_t0, _0183_, _0185_, _0187_ };
assign _0497_ = { _0758_, multdiv_en, _0184_, _0188_, _0190_ } | { _0759_, multdiv_en_t0, _0185_, _0189_, _0191_ };
assign _0498_ = { _0783_, _0758_, multdiv_en, _0192_ } | { _0784_, _0759_, multdiv_en_t0, _0193_ };
assign _0174_ = & _0494_;
assign _0175_ = & _0495_;
assign _0176_ = & _0496_;
assign _0177_ = & _0497_;
assign _0178_ = & _0498_;
assign _0195_ = _0169_ & _0174_;
assign _0197_ = _0170_ & _0175_;
assign _0199_ = _0171_ & _0176_;
assign _0201_ = _0172_ & _0177_;
assign _0203_ = _0173_ & _0178_;
assign _0179_ = | _0791_;
wire [31:0] _1661_ = imd_val_q_i_t0[31:0];
assign _0733_ = _1661_[_0790_ +: 1];
assign _0789_ = _0179_ | _0733_;
assign _0734_ = 33'h000000000 << multdiv_count_q;
assign one_shift_t0 = { _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_, _0061_ } | _0734_;
assign _0599_ = multdiv_count_q | multdiv_count_q_t0;
assign _0689_ = _0599_ - 5'h01;
assign _0690_ = _0388_ - 5'h01;
assign _0666_ = _0689_ ^ _0690_;
assign _0791_ = _0666_ | multdiv_count_q_t0;
assign _0807_ = rem_change_sign_t0 | sign_b_t0;
assign _0737_ = imd_val_q_i[65] == /* src = "generated/sv2v_out.v:19583.29-19583.67" */ op_b_shift_q[31];
assign _0739_ = ! /* src = "generated/sv2v_out.v:19606.45-19606.65" */ { 1'h0, sign_b, op_b_i[31:1] };
assign _0741_ = ! /* src = "generated/sv2v_out.v:19645.46-19645.63" */ { 1'h0, op_b_shift_q[32:1] };
assign _0743_ = multdiv_count_q == /* src = "generated/sv2v_out.v:19656.22-19656.45" */ 5'h01;
assign _0751_ = _0757_ && /* src = "generated/sv2v_out.v:19606.22-19606.66" */ _0739_;
assign _0753_ = _0757_ && /* src = "generated/sv2v_out.v:19621.22-19621.59" */ equal_to_zero_i;
assign _0755_ = _0757_ && /* src = "generated/sv2v_out.v:19645.23-19645.64" */ _0741_;
assign _0757_ = ! /* src = "generated/sv2v_out.v:19645.23-19645.41" */ data_ind_timing_i;
assign _0758_ = mult_sel_i || /* src = "generated/sv2v_out.v:19598.7-19598.30" */ div_sel_i;
assign _0760_ = _0755_ || /* src = "generated/sv2v_out.v:19645.22-19645.94" */ _0743_;
assign _0763_ = ~ /* src = "generated/sv2v_out.v:19555.26-19555.33" */ op_a_i;
assign _0762_ = ~ /* src = "generated/sv2v_out.v:19559.26-19559.33" */ op_b_i;
assign _0764_ = ~ /* src = "generated/sv2v_out.v:19563.26-19563.47" */ imd_val_q_i[65:34];
assign _0765_ = ~ /* src = "generated/sv2v_out.v:19572.24-19572.43" */ op_b_shift_q[31:0];
assign op_a_bw_pp[32] = ~ /* src = "generated/sv2v_out.v:19577.23-19577.60" */ op_a_bw_last_pp[32];
assign op_a_bw_last_pp[31:0] = ~ /* src = "generated/sv2v_out.v:19578.64-19578.91" */ op_a_bw_pp[31:0];
assign _0766_ = ~ /* src = "generated/sv2v_out.v:19583.70-19583.86" */ alu_adder_ext_i[32];
assign _0767_ = ~ /* src = "generated/sv2v_out.v:19587.47-19587.61" */ div_by_zero_q;
assign _0768_ = ~ /* src = "generated/sv2v_out.v:19610.32-19610.59" */ _0046_;
assign _0632_ = ~ /* src = "generated/sv2v_out.v:19697.21-19697.40" */ multdiv_ready_id_i;
assign imd_val_we_o[0] = ~ /* src = "generated/sv2v_out.v:19702.47-19702.60" */ multdiv_hold;
assign _0769_ = op_a_shift_q | /* src = "generated/sv2v_out.v:19586.45-19586.69" */ one_shift;
assign _0771_ = mult_en_i | /* src = "generated/sv2v_out.v:19702.23-19702.43" */ div_en_i;
assign _0773_ = _0747_ | /* src = "generated/sv2v_out.v:19718.67-19718.110" */ _0749_;
assign valid_o = _0745_ | /* src = "generated/sv2v_out.v:19718.19-19718.112" */ _0050_;
assign _0036_ = _0205_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19640.6-19660.13" */ { 1'h0, op_b_shift_q[32:1] } : 33'hxxxxxxxxx;
assign _0028_ = _0205_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19601.6-19625.13" */ { 1'h0, sign_b, op_b_i[31:1] } : 33'hxxxxxxxxx;
assign _0020_ = _0777_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19601.6-19625.13" */ equal_to_zero_i : 1'hx;
assign _0781_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19599.4-19700.11" */ 3'h3;
assign _0745_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19599.4-19700.11" */ 3'h6;
assign _0735_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19599.4-19700.11" */ 3'h4;
assign _0016_ = _0785_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19599.4-19700.11" */ _0796_ : imd_val_q_i[31:0];
assign multdiv_hold = _0758_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:19598.7-19598.30|generated/sv2v_out.v:19598.3-19700.11" */ _0010_ : 1'h0;
assign op_numerator_d = _0758_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:19598.7-19598.30|generated/sv2v_out.v:19598.3-19700.11" */ _0016_ : imd_val_q_i[31:0];
assign accum_window_d = _0758_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:19598.7-19598.30|generated/sv2v_out.v:19598.3-19700.11" */ _0000_ : imd_val_q_i[66:34];
assign _0002_ = _0165_ ? /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19548.5-19569.12" */ 33'h000000001 : { imd_val_q_i[65:34], 1'h1 };
assign _0779_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19548.5-19569.12" */ 3'h5;
assign _0787_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19548.5-19569.12" */ 3'h2;
assign _0785_ = md_state_q == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19548.5-19569.12" */ 3'h1;
assign _0783_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19548.5-19569.12" */ md_state_q;
assign _0749_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19544.3-19574.10" */ 2'h1;
assign _0747_ = ! /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19544.3-19574.10" */ operator_i;
assign _0777_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19544.3-19574.10" */ 2'h2;
assign _0775_ = operator_i == /* full_case = 32'd1 */ /* src = "generated/sv2v_out.v:0.0-0.0|generated/sv2v_out.v:19544.3-19574.10" */ 2'h3;
wire [31:0] _1662_ = imd_val_q_i[31:0];
assign _0788_ = _1662_[_0790_ +: 1];
assign one_shift = 33'h000000001 << /* src = "generated/sv2v_out.v:19584.21-19584.77" */ multdiv_count_q;
assign _0790_ = multdiv_count_q - /* src = "generated/sv2v_out.v:19639.24-19639.47" */ 5'h01;
assign _0792_ = _0735_ ? /* src = "generated/sv2v_out.v:19546.29-19546.78" */ op_a_bw_last_pp : op_a_bw_pp;
assign is_greater_equal = _0737_ ? /* src = "generated/sv2v_out.v:19583.29-19583.107" */ _0766_ : imd_val_q_i[65];
assign next_remainder = is_greater_equal ? /* src = "generated/sv2v_out.v:19585.27-19585.86" */ alu_adder_ext_i[32:1] : imd_val_q_i[65:34];
assign next_quotient = is_greater_equal ? /* src = "generated/sv2v_out.v:19586.26-19586.84" */ _0769_ : op_a_shift_q;
assign { _0639_[2], _0794_[1:0] } = _0751_ ? /* src = "generated/sv2v_out.v:19606.22-19606.80" */ 3'h4 : 3'h3;
assign _0795_ = _0753_ ? /* src = "generated/sv2v_out.v:19621.22-19621.73" */ 3'h6 : 3'h1;
assign _0796_ = rem_change_sign ? /* src = "generated/sv2v_out.v:19630.24-19630.53" */ alu_adder_i : op_a_i;
assign _0798_ = sign_b ? /* src = "generated/sv2v_out.v:19635.22-19635.67" */ { 1'h0, alu_adder_i } : { 1'h0, op_b_i };
assign _0800_ = _0760_ ? /* src = "generated/sv2v_out.v:19645.22-19645.108" */ 3'h4 : 3'h3;
assign _0801_ = _0743_ ? /* src = "generated/sv2v_out.v:19656.22-19656.59" */ 3'h4 : 3'h3;
assign _0802_ = div_change_sign ? /* src = "generated/sv2v_out.v:19689.31-19689.85" */ { 1'h0, alu_adder_i } : imd_val_q_i[66:34];
assign _0804_ = rem_change_sign ? /* src = "generated/sv2v_out.v:19690.31-19690.85" */ { 1'h0, alu_adder_i } : imd_val_q_i[66:34];
assign multdiv_result_o = div_en_i ? /* src = "generated/sv2v_out.v:19719.29-19719.80" */ imd_val_q_i[65:34] : alu_adder_ext_i[31:0];
assign _0806_ = rem_change_sign ^ /* src = "generated/sv2v_out.v:19587.28-19587.43" */ sign_b;
assign _0041_[1:0] = { 1'h0, _0041_[2] };
assign _0639_[1:0] = _0148_;
assign _0653_[2:1] = _0149_;
assign _0715_[0] = _0653_[0];
assign _0720_[2:1] = 2'h0;
assign _0794_[2] = _0639_[2];
assign imd_val_d_o = { 1'h0, accum_window_d, 2'h0, op_numerator_d };
assign imd_val_d_o_t0 = { 1'h0, accum_window_d_t0, 2'h0, op_numerator_d_t0 };
assign imd_val_we_o[1] = multdiv_en;
assign imd_val_we_o_t0 = { multdiv_en_t0, multdiv_hold_t0 };
endmodule

module ibex_top(clk_i, rst_ni, test_en_i, ram_cfg_i, hart_id_i, boot_addr_i, instr_req_o, instr_gnt_i, instr_rvalid_i, instr_addr_o, instr_rdata_i, instr_rdata_intg_i, instr_err_i, data_req_o, data_gnt_i, data_rvalid_i, data_we_o, data_be_o, data_addr_o, data_wdata_o, data_wdata_intg_o
, data_rdata_i, data_rdata_intg_i, data_err_i, irq_software_i, irq_timer_i, irq_external_i, irq_fast_i, irq_nm_i, scramble_key_valid_i, scramble_key_i, scramble_nonce_i, scramble_req_o, debug_req_i, crash_dump_o, double_fault_seen_o, fetch_enable_i, alert_minor_o, alert_major_internal_o, alert_major_bus_o, core_sleep_o, scan_rst_ni
, data_we_o_t0, data_req_o_t0, debug_req_i_t0, boot_addr_i_t0, instr_rvalid_i_t0, instr_req_o_t0, instr_rdata_i_t0, instr_gnt_i_t0, instr_err_i_t0, instr_addr_o_t0, test_en_i_t0, irq_nm_i_t0, data_addr_o_t0, data_be_o_t0, data_gnt_i_t0, data_rdata_i_t0, data_rvalid_i_t0, data_wdata_o_t0, double_fault_seen_o_t0, hart_id_i_t0, irq_external_i_t0
, irq_fast_i_t0, irq_software_i_t0, irq_timer_i_t0, alert_major_bus_o_t0, alert_major_internal_o_t0, alert_minor_o_t0, crash_dump_o_t0, data_err_i_t0, fetch_enable_i_t0, core_sleep_o_t0, data_rdata_intg_i_t0, data_wdata_intg_o_t0, instr_rdata_intg_i_t0, ram_cfg_i_t0, scan_rst_ni_t0, scramble_key_i_t0, scramble_key_valid_i_t0, scramble_nonce_i_t0, scramble_req_o_t0);
wire _00_;
wire [3:0] _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
wire _08_;
wire _09_;
wire [3:0] _10_;
wire _11_;
wire _12_;
wire _13_;
wire _14_;
wire _15_;
wire _16_;
wire _17_;
wire _18_;
wire _19_;
wire _20_;
wire _21_;
wire _22_;
wire _23_;
wire _24_;
wire _25_;
wire _26_;
wire _27_;
/* src = "generated/sv2v_out.v:20335.25-20335.60" */
wire _28_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20335.25-20335.60" */
wire _29_;
/* src = "generated/sv2v_out.v:20335.24-20335.75" */
wire _30_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20335.24-20335.75" */
wire _31_;
/* src = "generated/sv2v_out.v:20335.23-20335.90" */
wire _32_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20335.23-20335.90" */
wire _33_;
/* src = "generated/sv2v_out.v:20250.14-20250.31" */
output alert_major_bus_o;
wire alert_major_bus_o;
/* cellift = 32'd1 */
output alert_major_bus_o_t0;
wire alert_major_bus_o_t0;
/* src = "generated/sv2v_out.v:20249.14-20249.36" */
output alert_major_internal_o;
wire alert_major_internal_o;
/* cellift = 32'd1 */
output alert_major_internal_o_t0;
wire alert_major_internal_o_t0;
/* src = "generated/sv2v_out.v:20248.14-20248.27" */
output alert_minor_o;
wire alert_minor_o;
/* cellift = 32'd1 */
output alert_minor_o_t0;
wire alert_minor_o_t0;
/* src = "generated/sv2v_out.v:20216.20-20216.31" */
input [31:0] boot_addr_i;
wire [31:0] boot_addr_i;
/* cellift = 32'd1 */
input [31:0] boot_addr_i_t0;
wire [31:0] boot_addr_i_t0;
/* src = "generated/sv2v_out.v:20278.7-20278.10" */
wire clk;
/* src = "generated/sv2v_out.v:20211.13-20211.18" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:20281.7-20281.15" */
wire clock_en;
/* src = "generated/sv2v_out.v:20308.7-20308.32" */
wire core_alert_major_internal;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20308.7-20308.32" */
wire core_alert_major_internal_t0;
/* src = "generated/sv2v_out.v:20279.13-20279.24" */
wire [3:0] core_busy_d;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20279.13-20279.24" */
wire [3:0] core_busy_d_t0;
/* src = "generated/sv2v_out.v:20280.12-20280.23" */
wire [3:0] core_busy_q;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20280.12-20280.23" */
wire [3:0] core_busy_q_t0;
/* src = "generated/sv2v_out.v:20251.14-20251.26" */
output core_sleep_o;
wire core_sleep_o;
/* cellift = 32'd1 */
output core_sleep_o_t0;
wire core_sleep_o_t0;
/* src = "generated/sv2v_out.v:20245.22-20245.34" */
output [159:0] crash_dump_o;
wire [159:0] crash_dump_o;
/* cellift = 32'd1 */
output [159:0] crash_dump_o_t0;
wire [159:0] crash_dump_o_t0;
/* src = "generated/sv2v_out.v:20229.21-20229.32" */
output [31:0] data_addr_o;
wire [31:0] data_addr_o;
/* cellift = 32'd1 */
output [31:0] data_addr_o_t0;
wire [31:0] data_addr_o_t0;
/* src = "generated/sv2v_out.v:20228.20-20228.29" */
output [3:0] data_be_o;
wire [3:0] data_be_o;
/* cellift = 32'd1 */
output [3:0] data_be_o_t0;
wire [3:0] data_be_o_t0;
/* src = "generated/sv2v_out.v:20234.13-20234.23" */
input data_err_i;
wire data_err_i;
/* cellift = 32'd1 */
input data_err_i_t0;
wire data_err_i_t0;
/* src = "generated/sv2v_out.v:20225.13-20225.23" */
input data_gnt_i;
wire data_gnt_i;
/* cellift = 32'd1 */
input data_gnt_i_t0;
wire data_gnt_i_t0;
/* src = "generated/sv2v_out.v:20232.20-20232.32" */
input [31:0] data_rdata_i;
wire [31:0] data_rdata_i;
/* cellift = 32'd1 */
input [31:0] data_rdata_i_t0;
wire [31:0] data_rdata_i_t0;
/* src = "generated/sv2v_out.v:20233.19-20233.36" */
input [6:0] data_rdata_intg_i;
wire [6:0] data_rdata_intg_i;
/* cellift = 32'd1 */
input [6:0] data_rdata_intg_i_t0;
wire [6:0] data_rdata_intg_i_t0;
/* src = "generated/sv2v_out.v:20224.14-20224.24" */
output data_req_o;
wire data_req_o;
/* cellift = 32'd1 */
output data_req_o_t0;
wire data_req_o_t0;
/* src = "generated/sv2v_out.v:20226.13-20226.26" */
input data_rvalid_i;
wire data_rvalid_i;
/* cellift = 32'd1 */
input data_rvalid_i_t0;
wire data_rvalid_i_t0;
/* src = "generated/sv2v_out.v:20294.28-20294.43" */
wire [38:0] data_wdata_core;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20294.28-20294.43" */
wire [38:0] data_wdata_core_t0;
/* src = "generated/sv2v_out.v:20231.20-20231.37" */
output [6:0] data_wdata_intg_o;
wire [6:0] data_wdata_intg_o;
/* cellift = 32'd1 */
output [6:0] data_wdata_intg_o_t0;
wire [6:0] data_wdata_intg_o_t0;
/* src = "generated/sv2v_out.v:20230.21-20230.33" */
output [31:0] data_wdata_o;
wire [31:0] data_wdata_o;
/* cellift = 32'd1 */
output [31:0] data_wdata_o_t0;
wire [31:0] data_wdata_o_t0;
/* src = "generated/sv2v_out.v:20227.14-20227.23" */
output data_we_o;
wire data_we_o;
/* cellift = 32'd1 */
output data_we_o_t0;
wire data_we_o_t0;
/* src = "generated/sv2v_out.v:20244.13-20244.24" */
input debug_req_i;
wire debug_req_i;
/* cellift = 32'd1 */
input debug_req_i_t0;
wire debug_req_i_t0;
/* src = "generated/sv2v_out.v:20246.14-20246.33" */
output double_fault_seen_o;
wire double_fault_seen_o;
/* cellift = 32'd1 */
output double_fault_seen_o_t0;
wire double_fault_seen_o_t0;
/* src = "generated/sv2v_out.v:20283.7-20283.21" */
wire dummy_instr_id;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20283.7-20283.21" */
wire dummy_instr_id_t0;
/* src = "generated/sv2v_out.v:20284.7-20284.21" */
wire dummy_instr_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20284.7-20284.21" */
wire dummy_instr_wb_t0;
/* src = "generated/sv2v_out.v:20320.13-20320.29" */
wire [3:0] fetch_enable_buf;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20320.13-20320.29" */
wire [3:0] fetch_enable_buf_t0;
/* src = "generated/sv2v_out.v:20247.19-20247.33" */
input [3:0] fetch_enable_i;
wire [3:0] fetch_enable_i;
/* cellift = 32'd1 */
input [3:0] fetch_enable_i_t0;
wire [3:0] fetch_enable_i_t0;
/* src = "generated/sv2v_out.v:20215.20-20215.29" */
input [31:0] hart_id_i;
wire [31:0] hart_id_i;
/* cellift = 32'd1 */
input [31:0] hart_id_i_t0;
wire [31:0] hart_id_i_t0;
/* src = "generated/sv2v_out.v:20304.35-20304.47" */
/* unused_bits = "0 1 2 3 4 5 6 7" */
wire [7:0] ic_data_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20304.35-20304.47" */
/* unused_bits = "0 1 2 3 4 5 6 7" */
wire [7:0] ic_data_addr_t0;
/* src = "generated/sv2v_out.v:20302.13-20302.24" */
/* unused_bits = "0 1" */
wire [1:0] ic_data_req;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20302.13-20302.24" */
/* unused_bits = "0 1" */
wire [1:0] ic_data_req_t0;
/* src = "generated/sv2v_out.v:20305.27-20305.40" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63" */
wire [63:0] ic_data_wdata;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20305.27-20305.40" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63" */
wire [63:0] ic_data_wdata_t0;
/* src = "generated/sv2v_out.v:20303.7-20303.20" */
/* unused_bits = "0" */
wire ic_data_write;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20303.7-20303.20" */
/* unused_bits = "0" */
wire ic_data_write_t0;
/* src = "generated/sv2v_out.v:20307.7-20307.21" */
/* unused_bits = "0" */
wire ic_scr_key_req;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20307.7-20307.21" */
/* unused_bits = "0" */
wire ic_scr_key_req_t0;
/* src = "generated/sv2v_out.v:20299.35-20299.46" */
/* unused_bits = "0 1 2 3 4 5 6 7" */
wire [7:0] ic_tag_addr;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20299.35-20299.46" */
/* unused_bits = "0 1 2 3 4 5 6 7" */
wire [7:0] ic_tag_addr_t0;
/* src = "generated/sv2v_out.v:20297.13-20297.23" */
/* unused_bits = "0 1" */
wire [1:0] ic_tag_req;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20297.13-20297.23" */
/* unused_bits = "0 1" */
wire [1:0] ic_tag_req_t0;
/* src = "generated/sv2v_out.v:20300.26-20300.38" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21" */
wire [21:0] ic_tag_wdata;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20300.26-20300.38" */
/* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21" */
wire [21:0] ic_tag_wdata_t0;
/* src = "generated/sv2v_out.v:20298.7-20298.19" */
/* unused_bits = "0" */
wire ic_tag_write;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20298.7-20298.19" */
/* unused_bits = "0" */
wire ic_tag_write_t0;
/* src = "generated/sv2v_out.v:20220.21-20220.33" */
output [31:0] instr_addr_o;
wire [31:0] instr_addr_o;
/* cellift = 32'd1 */
output [31:0] instr_addr_o_t0;
wire [31:0] instr_addr_o_t0;
/* src = "generated/sv2v_out.v:20223.13-20223.24" */
input instr_err_i;
wire instr_err_i;
/* cellift = 32'd1 */
input instr_err_i_t0;
wire instr_err_i_t0;
/* src = "generated/sv2v_out.v:20218.13-20218.24" */
input instr_gnt_i;
wire instr_gnt_i;
/* cellift = 32'd1 */
input instr_gnt_i_t0;
wire instr_gnt_i_t0;
/* src = "generated/sv2v_out.v:20221.20-20221.33" */
input [31:0] instr_rdata_i;
wire [31:0] instr_rdata_i;
/* cellift = 32'd1 */
input [31:0] instr_rdata_i_t0;
wire [31:0] instr_rdata_i_t0;
/* src = "generated/sv2v_out.v:20222.19-20222.37" */
input [6:0] instr_rdata_intg_i;
wire [6:0] instr_rdata_intg_i;
/* cellift = 32'd1 */
input [6:0] instr_rdata_intg_i_t0;
wire [6:0] instr_rdata_intg_i_t0;
/* src = "generated/sv2v_out.v:20217.14-20217.25" */
output instr_req_o;
wire instr_req_o;
/* cellift = 32'd1 */
output instr_req_o_t0;
wire instr_req_o_t0;
/* src = "generated/sv2v_out.v:20219.13-20219.27" */
input instr_rvalid_i;
wire instr_rvalid_i;
/* cellift = 32'd1 */
input instr_rvalid_i_t0;
wire instr_rvalid_i_t0;
/* src = "generated/sv2v_out.v:20237.13-20237.27" */
input irq_external_i;
wire irq_external_i;
/* cellift = 32'd1 */
input irq_external_i_t0;
wire irq_external_i_t0;
/* src = "generated/sv2v_out.v:20238.20-20238.30" */
input [14:0] irq_fast_i;
wire [14:0] irq_fast_i;
/* cellift = 32'd1 */
input [14:0] irq_fast_i_t0;
wire [14:0] irq_fast_i_t0;
/* src = "generated/sv2v_out.v:20239.13-20239.21" */
input irq_nm_i;
wire irq_nm_i;
/* cellift = 32'd1 */
input irq_nm_i_t0;
wire irq_nm_i_t0;
/* src = "generated/sv2v_out.v:20282.7-20282.18" */
wire irq_pending;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20282.7-20282.18" */
wire irq_pending_t0;
/* src = "generated/sv2v_out.v:20235.13-20235.27" */
input irq_software_i;
wire irq_software_i;
/* cellift = 32'd1 */
input irq_software_i_t0;
wire irq_software_i_t0;
/* src = "generated/sv2v_out.v:20236.13-20236.24" */
input irq_timer_i;
wire irq_timer_i;
/* cellift = 32'd1 */
input irq_timer_i_t0;
wire irq_timer_i_t0;
/* src = "generated/sv2v_out.v:20214.19-20214.28" */
input [9:0] ram_cfg_i;
wire [9:0] ram_cfg_i;
/* cellift = 32'd1 */
input [9:0] ram_cfg_i_t0;
wire [9:0] ram_cfg_i_t0;
/* src = "generated/sv2v_out.v:20465.7-20465.30" */
wire rf_alert_major_internal;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20465.7-20465.30" */
wire rf_alert_major_internal_t0;
/* src = "generated/sv2v_out.v:20285.13-20285.23" */
wire [4:0] rf_raddr_a;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20285.13-20285.23" */
wire [4:0] rf_raddr_a_t0;
/* src = "generated/sv2v_out.v:20286.13-20286.23" */
wire [4:0] rf_raddr_b;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20286.13-20286.23" */
wire [4:0] rf_raddr_b_t0;
/* src = "generated/sv2v_out.v:20290.32-20290.46" */
wire [38:0] rf_rdata_a_ecc;
/* src = "generated/sv2v_out.v:20291.32-20291.50" */
wire [38:0] rf_rdata_a_ecc_buf;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20291.32-20291.50" */
wire [38:0] rf_rdata_a_ecc_buf_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20290.32-20290.46" */
wire [38:0] rf_rdata_a_ecc_t0;
/* src = "generated/sv2v_out.v:20292.32-20292.46" */
wire [38:0] rf_rdata_b_ecc;
/* src = "generated/sv2v_out.v:20293.32-20293.50" */
wire [38:0] rf_rdata_b_ecc_buf;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20293.32-20293.50" */
wire [38:0] rf_rdata_b_ecc_buf_t0;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20292.32-20292.46" */
wire [38:0] rf_rdata_b_ecc_t0;
/* src = "generated/sv2v_out.v:20287.13-20287.24" */
wire [4:0] rf_waddr_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20287.13-20287.24" */
wire [4:0] rf_waddr_wb_t0;
/* src = "generated/sv2v_out.v:20289.32-20289.47" */
wire [38:0] rf_wdata_wb_ecc;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20289.32-20289.47" */
wire [38:0] rf_wdata_wb_ecc_t0;
/* src = "generated/sv2v_out.v:20288.7-20288.15" */
wire rf_we_wb;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:20288.7-20288.15" */
wire rf_we_wb_t0;
/* src = "generated/sv2v_out.v:20212.13-20212.19" */
input rst_ni;
wire rst_ni;
/* src = "generated/sv2v_out.v:20252.13-20252.24" */
input scan_rst_ni;
wire scan_rst_ni;
/* cellift = 32'd1 */
input scan_rst_ni_t0;
wire scan_rst_ni_t0;
/* src = "generated/sv2v_out.v:20241.21-20241.35" */
input [127:0] scramble_key_i;
wire [127:0] scramble_key_i;
/* cellift = 32'd1 */
input [127:0] scramble_key_i_t0;
wire [127:0] scramble_key_i_t0;
/* src = "generated/sv2v_out.v:20240.13-20240.33" */
input scramble_key_valid_i;
wire scramble_key_valid_i;
/* cellift = 32'd1 */
input scramble_key_valid_i_t0;
wire scramble_key_valid_i_t0;
/* src = "generated/sv2v_out.v:20242.20-20242.36" */
input [63:0] scramble_nonce_i;
wire [63:0] scramble_nonce_i;
/* cellift = 32'd1 */
input [63:0] scramble_nonce_i_t0;
wire [63:0] scramble_nonce_i_t0;
/* src = "generated/sv2v_out.v:20243.14-20243.28" */
output scramble_req_o;
wire scramble_req_o;
/* cellift = 32'd1 */
output scramble_req_o_t0;
wire scramble_req_o_t0;
/* src = "generated/sv2v_out.v:20213.13-20213.22" */
input test_en_i;
wire test_en_i;
/* cellift = 32'd1 */
input test_en_i_t0;
wire test_en_i_t0;
assign _00_ = | core_busy_q_t0;
assign _01_ = ~ core_busy_q_t0;
assign _10_ = core_busy_q & _01_;
assign _27_ = _10_ == { _01_[3], 1'h0, _01_[1], 1'h0 };
assign _29_ = _27_ & _00_;
assign _02_ = ~ _28_;
assign _03_ = ~ _30_;
assign _04_ = ~ _32_;
assign _05_ = ~ core_alert_major_internal;
assign _06_ = ~ debug_req_i;
assign _07_ = ~ irq_pending;
assign _08_ = ~ irq_nm_i;
assign _09_ = ~ rf_alert_major_internal;
assign _11_ = _29_ & _06_;
assign _14_ = _31_ & _07_;
assign _17_ = _33_ & _08_;
assign _20_ = core_alert_major_internal_t0 & _09_;
assign _12_ = debug_req_i_t0 & _02_;
assign _15_ = irq_pending_t0 & _03_;
assign _18_ = irq_nm_i_t0 & _04_;
assign _21_ = rf_alert_major_internal_t0 & _05_;
assign _13_ = _29_ & debug_req_i_t0;
assign _16_ = _31_ & irq_pending_t0;
assign _19_ = _33_ & irq_nm_i_t0;
assign _22_ = core_alert_major_internal_t0 & rf_alert_major_internal_t0;
assign _23_ = _11_ | _12_;
assign _24_ = _14_ | _15_;
assign _25_ = _17_ | _18_;
assign _26_ = _20_ | _21_;
assign _31_ = _23_ | _13_;
assign _33_ = _24_ | _16_;
assign core_sleep_o_t0 = _25_ | _19_;
assign alert_major_internal_o_t0 = _26_ | _22_;
assign _28_ = core_busy_q != /* src = "generated/sv2v_out.v:20335.25-20335.60" */ 4'ha;
assign core_sleep_o = ~ /* src = "generated/sv2v_out.v:20348.24-20348.33" */ clock_en;
assign _30_ = _28_ | /* src = "generated/sv2v_out.v:20335.24-20335.75" */ debug_req_i;
assign _32_ = _30_ | /* src = "generated/sv2v_out.v:20335.23-20335.90" */ irq_pending;
assign clock_en = _32_ | /* src = "generated/sv2v_out.v:20335.22-20335.102" */ irq_nm_i;
assign alert_major_internal_o = core_alert_major_internal | /* src = "generated/sv2v_out.v:20877.34-20877.119" */ rf_alert_major_internal;
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20349.20-20354.3" */
prim_clock_gating core_clock_gate_i (
.clk_i(clk_i),
.clk_o(clk),
.en_i(clock_en),
.en_i_t0(core_sleep_o_t0),
.test_en_i(test_en_i),
.test_en_i_t0(test_en_i_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20329.6-20334.5" */
\$paramod$46c6ade532ce01738802967926171b52e9aa3bc1\prim_flop  \g_clock_en_secure.u_prim_core_busy_flop  (
.clk_i(clk_i),
.d_i(core_busy_d),
.d_i_t0(core_busy_d_t0),
.q_o(core_busy_q),
.q_o_t0(core_busy_q_t0),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20688.26-20691.5" */
\$paramod\prim_buf\Width=s32'00000000000000000000000000000111  \gen_mem_wdata_ecc.u_prim_buf_data_wdata_intg  (
.in_i(data_wdata_core[38:32]),
.in_i_t0(data_wdata_core_t0[38:32]),
.out_o(data_wdata_intg_o),
.out_o_t0(data_wdata_intg_o_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20479.6-20493.5" */
\$paramod$a575b78552d69534d7f9dc1a7d63a5588d1a8b59\ibex_register_file_ff  \gen_regfile_ff.register_file_i  (
.clk_i(clk),
.dummy_instr_id_i(dummy_instr_id),
.dummy_instr_id_i_t0(dummy_instr_id_t0),
.dummy_instr_wb_i(dummy_instr_wb),
.dummy_instr_wb_i_t0(dummy_instr_wb_t0),
.err_o(rf_alert_major_internal),
.err_o_t0(rf_alert_major_internal_t0),
.raddr_a_i(rf_raddr_a),
.raddr_a_i_t0(rf_raddr_a_t0),
.raddr_b_i(rf_raddr_b),
.raddr_b_i_t0(rf_raddr_b_t0),
.rdata_a_o(rf_rdata_a_ecc),
.rdata_a_o_t0(rf_rdata_a_ecc_t0),
.rdata_b_o(rf_rdata_b_ecc),
.rdata_b_o_t0(rf_rdata_b_ecc_t0),
.rst_ni(rst_ni),
.test_en_i(test_en_i),
.test_en_i_t0(test_en_i_t0),
.waddr_a_i(rf_waddr_wb),
.waddr_a_i_t0(rf_waddr_wb_t0),
.wdata_a_i(rf_wdata_wb_ecc),
.wdata_a_i_t0(rf_wdata_wb_ecc_t0),
.we_a_i(rf_we_wb),
.we_a_i_t0(rf_we_wb_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20355.24-20358.3" */
\$paramod\prim_buf\Width=s32'00000000000000000000000000000100  u_fetch_enable_buf (
.in_i(fetch_enable_i),
.in_i_t0(fetch_enable_i_t0),
.out_o(fetch_enable_buf),
.out_o_t0(fetch_enable_buf_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20409.4-20464.3" */
\$paramod$5c0dc9f9e0551018f7d8916b4fcabdef94a17390\ibex_core  u_ibex_core (
.alert_major_bus_o(alert_major_bus_o),
.alert_major_bus_o_t0(alert_major_bus_o_t0),
.alert_major_internal_o(core_alert_major_internal),
.alert_major_internal_o_t0(core_alert_major_internal_t0),
.alert_minor_o(alert_minor_o),
.alert_minor_o_t0(alert_minor_o_t0),
.boot_addr_i(boot_addr_i),
.boot_addr_i_t0(boot_addr_i_t0),
.clk_i(clk),
.core_busy_o(core_busy_d),
.core_busy_o_t0(core_busy_d_t0),
.crash_dump_o(crash_dump_o),
.crash_dump_o_t0(crash_dump_o_t0),
.data_addr_o(data_addr_o),
.data_addr_o_t0(data_addr_o_t0),
.data_be_o(data_be_o),
.data_be_o_t0(data_be_o_t0),
.data_err_i(data_err_i),
.data_err_i_t0(data_err_i_t0),
.data_gnt_i(data_gnt_i),
.data_gnt_i_t0(data_gnt_i_t0),
.data_rdata_i({ data_rdata_intg_i, data_rdata_i }),
.data_rdata_i_t0({ data_rdata_intg_i_t0, data_rdata_i_t0 }),
.data_req_o(data_req_o),
.data_req_o_t0(data_req_o_t0),
.data_rvalid_i(data_rvalid_i),
.data_rvalid_i_t0(data_rvalid_i_t0),
.data_wdata_o(data_wdata_core),
.data_wdata_o_t0(data_wdata_core_t0),
.data_we_o(data_we_o),
.data_we_o_t0(data_we_o_t0),
.debug_req_i(debug_req_i),
.debug_req_i_t0(debug_req_i_t0),
.double_fault_seen_o(double_fault_seen_o),
.double_fault_seen_o_t0(double_fault_seen_o_t0),
.dummy_instr_id_o(dummy_instr_id),
.dummy_instr_id_o_t0(dummy_instr_id_t0),
.dummy_instr_wb_o(dummy_instr_wb),
.dummy_instr_wb_o_t0(dummy_instr_wb_t0),
.fetch_enable_i(fetch_enable_buf),
.fetch_enable_i_t0(fetch_enable_buf_t0),
.hart_id_i(hart_id_i),
.hart_id_i_t0(hart_id_i_t0),
.ic_data_addr_o(ic_data_addr),
.ic_data_addr_o_t0(ic_data_addr_t0),
.ic_data_rdata_i(128'h00000000000000000000000000000000),
.ic_data_rdata_i_t0(128'h00000000000000000000000000000000),
.ic_data_req_o(ic_data_req),
.ic_data_req_o_t0(ic_data_req_t0),
.ic_data_wdata_o(ic_data_wdata),
.ic_data_wdata_o_t0(ic_data_wdata_t0),
.ic_data_write_o(ic_data_write),
.ic_data_write_o_t0(ic_data_write_t0),
.ic_scr_key_req_o(ic_scr_key_req),
.ic_scr_key_req_o_t0(ic_scr_key_req_t0),
.ic_scr_key_valid_i(1'h1),
.ic_scr_key_valid_i_t0(1'h0),
.ic_tag_addr_o(ic_tag_addr),
.ic_tag_addr_o_t0(ic_tag_addr_t0),
.ic_tag_rdata_i(44'h00000000000),
.ic_tag_rdata_i_t0(44'h00000000000),
.ic_tag_req_o(ic_tag_req),
.ic_tag_req_o_t0(ic_tag_req_t0),
.ic_tag_wdata_o(ic_tag_wdata),
.ic_tag_wdata_o_t0(ic_tag_wdata_t0),
.ic_tag_write_o(ic_tag_write),
.ic_tag_write_o_t0(ic_tag_write_t0),
.instr_addr_o(instr_addr_o),
.instr_addr_o_t0(instr_addr_o_t0),
.instr_err_i(instr_err_i),
.instr_err_i_t0(instr_err_i_t0),
.instr_gnt_i(instr_gnt_i),
.instr_gnt_i_t0(instr_gnt_i_t0),
.instr_rdata_i({ instr_rdata_intg_i, instr_rdata_i }),
.instr_rdata_i_t0({ instr_rdata_intg_i_t0, instr_rdata_i_t0 }),
.instr_req_o(instr_req_o),
.instr_req_o_t0(instr_req_o_t0),
.instr_rvalid_i(instr_rvalid_i),
.instr_rvalid_i_t0(instr_rvalid_i_t0),
.irq_external_i(irq_external_i),
.irq_external_i_t0(irq_external_i_t0),
.irq_fast_i(irq_fast_i),
.irq_fast_i_t0(irq_fast_i_t0),
.irq_nm_i(irq_nm_i),
.irq_nm_i_t0(irq_nm_i_t0),
.irq_pending_o(irq_pending),
.irq_pending_o_t0(irq_pending_t0),
.irq_software_i(irq_software_i),
.irq_software_i_t0(irq_software_i_t0),
.irq_timer_i(irq_timer_i),
.irq_timer_i_t0(irq_timer_i_t0),
.rf_raddr_a_o(rf_raddr_a),
.rf_raddr_a_o_t0(rf_raddr_a_t0),
.rf_raddr_b_o(rf_raddr_b),
.rf_raddr_b_o_t0(rf_raddr_b_t0),
.rf_rdata_a_ecc_i(rf_rdata_a_ecc_buf),
.rf_rdata_a_ecc_i_t0(rf_rdata_a_ecc_buf_t0),
.rf_rdata_b_ecc_i(rf_rdata_b_ecc_buf),
.rf_rdata_b_ecc_i_t0(rf_rdata_b_ecc_buf_t0),
.rf_waddr_wb_o(rf_waddr_wb),
.rf_waddr_wb_o_t0(rf_waddr_wb_t0),
.rf_wdata_wb_ecc_o(rf_wdata_wb_ecc),
.rf_wdata_wb_ecc_o_t0(rf_wdata_wb_ecc_t0),
.rf_we_wb_o(rf_we_wb),
.rf_we_wb_o_t0(rf_we_wb_t0),
.rst_ni(rst_ni)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20359.39-20362.3" */
\$paramod\prim_buf\Width=32'00000000000000000000000000100111  u_rf_rdata_a_ecc_buf (
.in_i(rf_rdata_a_ecc),
.in_i_t0(rf_rdata_a_ecc_t0),
.out_o(rf_rdata_a_ecc_buf),
.out_o_t0(rf_rdata_a_ecc_buf_t0)
);
/* module_not_derived = 32'd1 */
/* src = "generated/sv2v_out.v:20363.39-20366.3" */
\$paramod\prim_buf\Width=32'00000000000000000000000000100111  u_rf_rdata_b_ecc_buf (
.in_i(rf_rdata_b_ecc),
.in_i_t0(rf_rdata_b_ecc_t0),
.out_o(rf_rdata_b_ecc_buf),
.out_o_t0(rf_rdata_b_ecc_buf_t0)
);
assign data_wdata_o = data_wdata_core[31:0];
assign data_wdata_o_t0 = data_wdata_core_t0[31:0];
assign scramble_req_o = 1'h0;
assign scramble_req_o_t0 = 1'h0;
endmodule

module prim_clock_gating(clk_i, en_i, test_en_i, clk_o, clk_o_t0, en_i_t0, test_en_i_t0);
/* src = "generated/sv2v_out.v:23060.2-23062.32" */
wire _00_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:23060.2-23062.32" */
wire _01_;
wire _02_;
wire _03_;
wire _04_;
wire _05_;
wire _06_;
wire _07_;
/* src = "generated/sv2v_out.v:23055.8-23055.13" */
input clk_i;
wire clk_i;
/* src = "generated/sv2v_out.v:23058.14-23058.19" */
output clk_o;
wire clk_o;
/* cellift = 32'd1 */
output clk_o_t0;
wire clk_o_t0;
/* src = "generated/sv2v_out.v:23056.8-23056.12" */
input en_i;
wire en_i;
/* cellift = 32'd1 */
input en_i_t0;
wire en_i_t0;
/* src = "generated/sv2v_out.v:23059.6-23059.14" */
reg en_latch;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:23059.6-23059.14" */
reg en_latch_t0;
/* src = "generated/sv2v_out.v:23057.8-23057.17" */
input test_en_i;
wire test_en_i;
/* cellift = 32'd1 */
input test_en_i_t0;
wire test_en_i_t0;
assign clk_o = en_latch & /* src = "generated/sv2v_out.v:23063.17-23063.33" */ clk_i;
assign clk_o_t0 = en_latch_t0 & clk_i;
/* taint_latch = 32'd1 */
/* PC_TAINT_INFO MODULE_NAME prim_clock_gating */
/* PC_TAINT_INFO STATE_NAME en_latch_t0 */
always_latch
if (!clk_i) en_latch_t0 = _01_;
assign _02_ = ~ en_i;
assign _03_ = ~ test_en_i;
assign _04_ = en_i_t0 & _03_;
assign _05_ = test_en_i_t0 & _02_;
assign _06_ = en_i_t0 & test_en_i_t0;
assign _07_ = _04_ | _05_;
assign _01_ = _07_ | _06_;
/* src = "generated/sv2v_out.v:23060.2-23062.32" */
/* PC_TAINT_INFO MODULE_NAME prim_clock_gating */
/* PC_TAINT_INFO STATE_NAME en_latch */
always_latch
if (!clk_i) en_latch = _00_;
assign _00_ = en_i | /* src = "generated/sv2v_out.v:23062.15-23062.31" */ test_en_i;
endmodule

module prim_secded_inv_39_32_dec(data_i, data_o, syndrome_o, err_o, syndrome_o_t0, err_o_t0, data_o_t0, data_i_t0);
/* src = "generated/sv2v_out.v:29273.21-29273.63" */
wire [38:0] _000_;
/* src = "generated/sv2v_out.v:29275.21-29275.63" */
wire [38:0] _001_;
/* src = "generated/sv2v_out.v:29277.21-29277.63" */
wire [38:0] _002_;
wire [6:0] _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire [6:0] _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
/* src = "generated/sv2v_out.v:29279.16-29279.35" */
wire _042_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29279.16-29279.35" */
wire _043_;
/* src = "generated/sv2v_out.v:29280.16-29280.35" */
wire _044_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29280.16-29280.35" */
wire _045_;
/* src = "generated/sv2v_out.v:29281.16-29281.35" */
wire _046_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29281.16-29281.35" */
wire _047_;
/* src = "generated/sv2v_out.v:29282.16-29282.35" */
wire _048_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29282.16-29282.35" */
wire _049_;
/* src = "generated/sv2v_out.v:29283.16-29283.35" */
wire _050_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29283.16-29283.35" */
wire _051_;
/* src = "generated/sv2v_out.v:29284.16-29284.35" */
wire _052_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29284.16-29284.35" */
wire _053_;
/* src = "generated/sv2v_out.v:29285.16-29285.35" */
wire _054_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29285.16-29285.35" */
wire _055_;
/* src = "generated/sv2v_out.v:29286.16-29286.35" */
wire _056_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29286.16-29286.35" */
wire _057_;
/* src = "generated/sv2v_out.v:29287.16-29287.35" */
wire _058_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29287.16-29287.35" */
wire _059_;
/* src = "generated/sv2v_out.v:29288.16-29288.35" */
wire _060_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29288.16-29288.35" */
wire _061_;
/* src = "generated/sv2v_out.v:29289.17-29289.36" */
wire _062_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29289.17-29289.36" */
wire _063_;
/* src = "generated/sv2v_out.v:29290.17-29290.36" */
wire _064_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29290.17-29290.36" */
wire _065_;
/* src = "generated/sv2v_out.v:29291.17-29291.36" */
wire _066_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29291.17-29291.36" */
wire _067_;
/* src = "generated/sv2v_out.v:29292.17-29292.36" */
wire _068_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29292.17-29292.36" */
wire _069_;
/* src = "generated/sv2v_out.v:29293.17-29293.36" */
wire _070_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29293.17-29293.36" */
wire _071_;
/* src = "generated/sv2v_out.v:29294.17-29294.36" */
wire _072_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29294.17-29294.36" */
wire _073_;
/* src = "generated/sv2v_out.v:29295.17-29295.36" */
wire _074_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29295.17-29295.36" */
wire _075_;
/* src = "generated/sv2v_out.v:29296.17-29296.36" */
wire _076_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29296.17-29296.36" */
wire _077_;
/* src = "generated/sv2v_out.v:29297.17-29297.36" */
wire _078_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29297.17-29297.36" */
wire _079_;
/* src = "generated/sv2v_out.v:29298.17-29298.36" */
wire _080_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29298.17-29298.36" */
wire _081_;
/* src = "generated/sv2v_out.v:29299.17-29299.36" */
wire _082_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29299.17-29299.36" */
wire _083_;
/* src = "generated/sv2v_out.v:29300.17-29300.36" */
wire _084_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29300.17-29300.36" */
wire _085_;
/* src = "generated/sv2v_out.v:29301.17-29301.36" */
wire _086_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29301.17-29301.36" */
wire _087_;
/* src = "generated/sv2v_out.v:29302.17-29302.36" */
wire _088_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29302.17-29302.36" */
wire _089_;
/* src = "generated/sv2v_out.v:29303.17-29303.36" */
wire _090_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29303.17-29303.36" */
wire _091_;
/* src = "generated/sv2v_out.v:29304.17-29304.36" */
wire _092_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29304.17-29304.36" */
wire _093_;
/* src = "generated/sv2v_out.v:29305.17-29305.36" */
wire _094_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29305.17-29305.36" */
wire _095_;
/* src = "generated/sv2v_out.v:29306.17-29306.36" */
wire _096_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29306.17-29306.36" */
wire _097_;
/* src = "generated/sv2v_out.v:29307.17-29307.36" */
wire _098_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29307.17-29307.36" */
wire _099_;
/* src = "generated/sv2v_out.v:29308.17-29308.36" */
wire _100_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29308.17-29308.36" */
wire _101_;
/* src = "generated/sv2v_out.v:29309.17-29309.36" */
wire _102_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29309.17-29309.36" */
wire _103_;
/* src = "generated/sv2v_out.v:29310.17-29310.36" */
wire _104_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29310.17-29310.36" */
wire _105_;
/* src = "generated/sv2v_out.v:29312.14-29312.23" */
wire _106_;
/* src = "generated/sv2v_out.v:29312.26-29312.37" */
wire _107_;
/* cellift = 32'd1 */
/* src = "generated/sv2v_out.v:29312.26-29312.37" */
wire _108_;
/* src = "generated/sv2v_out.v:29267.15-29267.21" */
input [38:0] data_i;
wire [38:0] data_i;
/* cellift = 32'd1 */
input [38:0] data_i_t0;
wire [38:0] data_i_t0;
/* src = "generated/sv2v_out.v:29268.20-29268.26" */
output [31:0] data_o;
wire [31:0] data_o;
/* cellift = 32'd1 */
output [31:0] data_o_t0;
wire [31:0] data_o_t0;
/* src = "generated/sv2v_out.v:29270.19-29270.24" */
output [1:0] err_o;
wire [1:0] err_o;
/* cellift = 32'd1 */
output [1:0] err_o_t0;
wire [1:0] err_o_t0;
/* src = "generated/sv2v_out.v:29269.19-29269.29" */
output [6:0] syndrome_o;
wire [6:0] syndrome_o;
/* cellift = 32'd1 */
output [6:0] syndrome_o_t0;
wire [6:0] syndrome_o_t0;
assign err_o[1] = _106_ & /* src = "generated/sv2v_out.v:29312.14-29312.37" */ _107_;
assign _005_ = err_o_t0[0] & _107_;
assign _006_ = _108_ & _106_;
assign _007_ = err_o_t0[0] & _108_;
assign _009_ = _005_ | _006_;
assign err_o_t0[1] = _009_ | _007_;
assign err_o_t0[0] = | data_i_t0;
assign _003_ = ~ syndrome_o_t0;
assign _008_ = syndrome_o & _003_;
assign _010_ = _008_ == { 2'h0, _003_[4:3], 2'h0, _003_[0] };
assign _011_ = _008_ == { _003_[6], 1'h0, _003_[4], 1'h0, _003_[2], 2'h0 };
assign _012_ = _008_ == { _003_[6:5], 4'h0, _003_[0] };
assign _013_ = _008_ == { 1'h0, _003_[5:4], 1'h0, _003_[2], 2'h0 };
assign _014_ = _008_ == { 2'h0, _003_[4:3], 1'h0, _003_[1], 1'h0 };
assign _015_ = _008_ == { 2'h0, _003_[4], 1'h0, _003_[2], 1'h0, _003_[0] };
assign _016_ = _008_ == { 1'h0, _003_[5], 1'h0, _003_[3], 1'h0, _003_[1], 1'h0 };
assign _017_ = _008_ == { _003_[6], 2'h0, _003_[3:2], 2'h0 };
assign _018_ = _008_ == { _003_[6], 3'h0, _003_[2], 1'h0, _003_[0] };
assign _019_ = _008_ == { 1'h0, _003_[5:3], 3'h0 };
assign _020_ = _008_ == { _003_[6], 2'h0, _003_[3], 2'h0, _003_[0] };
assign _021_ = _008_ == { 3'h0, _003_[3:2], 1'h0, _003_[0] };
assign _022_ = _008_ == { _003_[6], 1'h0, _003_[4], 3'h0, _003_[0] };
assign _023_ = _008_ == { 1'h0, _003_[5:4], 3'h0, _003_[0] };
assign _024_ = _008_ == { _003_[6:5], 1'h0, _003_[3], 3'h0 };
assign _025_ = _008_ == { 4'h0, _003_[2:0] };
assign _026_ = _008_ == { 2'h0, _003_[4:2], 2'h0 };
assign _027_ = _008_ == { 3'h0, _003_[3], 1'h0, _003_[1:0] };
assign _028_ = _008_ == { 1'h0, _003_[5], 2'h0, _003_[2], 1'h0, _003_[0] };
assign _029_ = _008_ == { 1'h0, _003_[5], 2'h0, _003_[2:1], 1'h0 };
assign _030_ = _008_ == { _003_[6], 3'h0, _003_[2:1], 1'h0 };
assign _031_ = _008_ == { 3'h0, _003_[3:1], 1'h0 };
assign _032_ = _008_ == { _003_[6:4], 4'h0 };
assign _033_ = _008_ == { 1'h0, _003_[5:4], 2'h0, _003_[1], 1'h0 };
assign _034_ = _008_ == { 1'h0, _003_[5], 1'h0, _003_[3:2], 2'h0 };
assign _035_ = _008_ == { 2'h0, _003_[4], 2'h0, _003_[1:0] };
assign _036_ = _008_ == { 1'h0, _003_[5], 3'h0, _003_[1:0] };
assign _037_ = _008_ == { _003_[6:5], 3'h0, _003_[1], 1'h0 };
assign _038_ = _008_ == { _003_[6], 2'h0, _003_[3], 1'h0, _003_[1], 1'h0 };
assign _039_ = _008_ == { 1'h0, _003_[5], 1'h0, _003_[3], 2'h0, _003_[0] };
assign _040_ = _008_ == { 2'h0, _003_[4], 1'h0, _003_[2:1], 1'h0 };
assign _041_ = _008_ == { _003_[6], 1'h0, _003_[4], 2'h0, _003_[1], 1'h0 };
assign _043_ = _010_ & err_o_t0[0];
assign _045_ = _011_ & err_o_t0[0];
assign _047_ = _012_ & err_o_t0[0];
assign _049_ = _013_ & err_o_t0[0];
assign _051_ = _014_ & err_o_t0[0];
assign _053_ = _015_ & err_o_t0[0];
assign _055_ = _016_ & err_o_t0[0];
assign _057_ = _017_ & err_o_t0[0];
assign _059_ = _018_ & err_o_t0[0];
assign _061_ = _019_ & err_o_t0[0];
assign _063_ = _020_ & err_o_t0[0];
assign _065_ = _021_ & err_o_t0[0];
assign _067_ = _022_ & err_o_t0[0];
assign _069_ = _023_ & err_o_t0[0];
assign _071_ = _024_ & err_o_t0[0];
assign _073_ = _025_ & err_o_t0[0];
assign _075_ = _026_ & err_o_t0[0];
assign _077_ = _027_ & err_o_t0[0];
assign _079_ = _028_ & err_o_t0[0];
assign _081_ = _029_ & err_o_t0[0];
assign _083_ = _030_ & err_o_t0[0];
assign _085_ = _031_ & err_o_t0[0];
assign _087_ = _032_ & err_o_t0[0];
assign _089_ = _033_ & err_o_t0[0];
assign _091_ = _034_ & err_o_t0[0];
assign _093_ = _035_ & err_o_t0[0];
assign _095_ = _036_ & err_o_t0[0];
assign _097_ = _037_ & err_o_t0[0];
assign _099_ = _038_ & err_o_t0[0];
assign _101_ = _039_ & err_o_t0[0];
assign _103_ = _040_ & err_o_t0[0];
assign _105_ = _041_ & err_o_t0[0];
assign _004_ = ! _008_;
assign _108_ = _004_ & err_o_t0[0];
assign { _002_[37], _001_[35], _000_[33] } = ~ { data_i[37], data_i[35], data_i[33] };
assign syndrome_o_t0[0] = | { data_i_t0[32], data_i_t0[29], data_i_t0[26:25], data_i_t0[18:17], data_i_t0[15], data_i_t0[13:10], data_i_t0[8], data_i_t0[5], data_i_t0[2], data_i_t0[0] };
assign syndrome_o_t0[1] = | { data_i_t0[33], data_i_t0[31:30], data_i_t0[28:25], data_i_t0[23], data_i_t0[21:19], data_i_t0[17], data_i_t0[15], data_i_t0[6], data_i_t0[4] };
assign syndrome_o_t0[2] = | { data_i_t0[34], data_i_t0[30], data_i_t0[24], data_i_t0[21:18], data_i_t0[16:15], data_i_t0[11], data_i_t0[8:7], data_i_t0[5], data_i_t0[3], data_i_t0[1] };
assign syndrome_o_t0[3] = | { data_i_t0[35], data_i_t0[29:28], data_i_t0[24], data_i_t0[21], data_i_t0[17:16], data_i_t0[14], data_i_t0[11:9], data_i_t0[7:6], data_i_t0[4], data_i_t0[0] };
assign syndrome_o_t0[4] = | { data_i_t0[36], data_i_t0[31:30], data_i_t0[25], data_i_t0[23:22], data_i_t0[16], data_i_t0[13:12], data_i_t0[9], data_i_t0[5:3], data_i_t0[1:0] };
assign syndrome_o_t0[5] = | { data_i_t0[37], data_i_t0[29], data_i_t0[27:26], data_i_t0[24:22], data_i_t0[19:18], data_i_t0[14:13], data_i_t0[9], data_i_t0[6], data_i_t0[3:2] };
assign syndrome_o_t0[6] = | { data_i_t0[38], data_i_t0[31], data_i_t0[28:27], data_i_t0[22], data_i_t0[20], data_i_t0[14], data_i_t0[12], data_i_t0[10], data_i_t0[8:7], data_i_t0[2:1] };
assign data_o_t0[0] = _043_ | data_i_t0[0];
assign data_o_t0[1] = _045_ | data_i_t0[1];
assign data_o_t0[2] = _047_ | data_i_t0[2];
assign data_o_t0[3] = _049_ | data_i_t0[3];
assign data_o_t0[4] = _051_ | data_i_t0[4];
assign data_o_t0[5] = _053_ | data_i_t0[5];
assign data_o_t0[6] = _055_ | data_i_t0[6];
assign data_o_t0[7] = _057_ | data_i_t0[7];
assign data_o_t0[8] = _059_ | data_i_t0[8];
assign data_o_t0[9] = _061_ | data_i_t0[9];
assign data_o_t0[10] = _063_ | data_i_t0[10];
assign data_o_t0[11] = _065_ | data_i_t0[11];
assign data_o_t0[12] = _067_ | data_i_t0[12];
assign data_o_t0[13] = _069_ | data_i_t0[13];
assign data_o_t0[14] = _071_ | data_i_t0[14];
assign data_o_t0[15] = _073_ | data_i_t0[15];
assign data_o_t0[16] = _075_ | data_i_t0[16];
assign data_o_t0[17] = _077_ | data_i_t0[17];
assign data_o_t0[18] = _079_ | data_i_t0[18];
assign data_o_t0[19] = _081_ | data_i_t0[19];
assign data_o_t0[20] = _083_ | data_i_t0[20];
assign data_o_t0[21] = _085_ | data_i_t0[21];
assign data_o_t0[22] = _087_ | data_i_t0[22];
assign data_o_t0[23] = _089_ | data_i_t0[23];
assign data_o_t0[24] = _091_ | data_i_t0[24];
assign data_o_t0[25] = _093_ | data_i_t0[25];
assign data_o_t0[26] = _095_ | data_i_t0[26];
assign data_o_t0[27] = _097_ | data_i_t0[27];
assign data_o_t0[28] = _099_ | data_i_t0[28];
assign data_o_t0[29] = _101_ | data_i_t0[29];
assign data_o_t0[30] = _103_ | data_i_t0[30];
assign data_o_t0[31] = _105_ | data_i_t0[31];
assign _042_ = syndrome_o == /* src = "generated/sv2v_out.v:29279.16-29279.35" */ 7'h19;
assign _044_ = syndrome_o == /* src = "generated/sv2v_out.v:29280.16-29280.35" */ 7'h54;
assign _046_ = syndrome_o == /* src = "generated/sv2v_out.v:29281.16-29281.35" */ 7'h61;
assign _048_ = syndrome_o == /* src = "generated/sv2v_out.v:29282.16-29282.35" */ 7'h34;
assign _050_ = syndrome_o == /* src = "generated/sv2v_out.v:29283.16-29283.35" */ 7'h1a;
assign _052_ = syndrome_o == /* src = "generated/sv2v_out.v:29284.16-29284.35" */ 7'h15;
assign _054_ = syndrome_o == /* src = "generated/sv2v_out.v:29285.16-29285.35" */ 7'h2a;
assign _056_ = syndrome_o == /* src = "generated/sv2v_out.v:29286.16-29286.35" */ 7'h4c;
assign _058_ = syndrome_o == /* src = "generated/sv2v_out.v:29287.16-29287.35" */ 7'h45;
assign _060_ = syndrome_o == /* src = "generated/sv2v_out.v:29288.16-29288.35" */ 7'h38;
assign _062_ = syndrome_o == /* src = "generated/sv2v_out.v:29289.17-29289.36" */ 7'h49;
assign _064_ = syndrome_o == /* src = "generated/sv2v_out.v:29290.17-29290.36" */ 7'h0d;
assign _066_ = syndrome_o == /* src = "generated/sv2v_out.v:29291.17-29291.36" */ 7'h51;
assign _068_ = syndrome_o == /* src = "generated/sv2v_out.v:29292.17-29292.36" */ 7'h31;
assign _070_ = syndrome_o == /* src = "generated/sv2v_out.v:29293.17-29293.36" */ 7'h68;
assign _072_ = syndrome_o == /* src = "generated/sv2v_out.v:29294.17-29294.36" */ 7'h07;
assign _074_ = syndrome_o == /* src = "generated/sv2v_out.v:29295.17-29295.36" */ 7'h1c;
assign _076_ = syndrome_o == /* src = "generated/sv2v_out.v:29296.17-29296.36" */ 7'h0b;
assign _078_ = syndrome_o == /* src = "generated/sv2v_out.v:29297.17-29297.36" */ 7'h25;
assign _080_ = syndrome_o == /* src = "generated/sv2v_out.v:29298.17-29298.36" */ 7'h26;
assign _082_ = syndrome_o == /* src = "generated/sv2v_out.v:29299.17-29299.36" */ 7'h46;
assign _084_ = syndrome_o == /* src = "generated/sv2v_out.v:29300.17-29300.36" */ 7'h0e;
assign _086_ = syndrome_o == /* src = "generated/sv2v_out.v:29301.17-29301.36" */ 7'h70;
assign _088_ = syndrome_o == /* src = "generated/sv2v_out.v:29302.17-29302.36" */ 7'h32;
assign _090_ = syndrome_o == /* src = "generated/sv2v_out.v:29303.17-29303.36" */ 7'h2c;
assign _092_ = syndrome_o == /* src = "generated/sv2v_out.v:29304.17-29304.36" */ 7'h13;
assign _094_ = syndrome_o == /* src = "generated/sv2v_out.v:29305.17-29305.36" */ 7'h23;
assign _096_ = syndrome_o == /* src = "generated/sv2v_out.v:29306.17-29306.36" */ 7'h62;
assign _098_ = syndrome_o == /* src = "generated/sv2v_out.v:29307.17-29307.36" */ 7'h4a;
assign _100_ = syndrome_o == /* src = "generated/sv2v_out.v:29308.17-29308.36" */ 7'h29;
assign _102_ = syndrome_o == /* src = "generated/sv2v_out.v:29309.17-29309.36" */ 7'h16;
assign _104_ = syndrome_o == /* src = "generated/sv2v_out.v:29310.17-29310.36" */ 7'h52;
assign _106_ = ~ /* src = "generated/sv2v_out.v:29312.14-29312.23" */ err_o[0];
assign _107_ = | /* src = "generated/sv2v_out.v:29312.26-29312.37" */ syndrome_o;
assign syndrome_o[0] = ^ /* src = "generated/sv2v_out.v:29272.19-29272.64" */ { 6'h00, data_i[32], 2'h0, data_i[29], 2'h0, data_i[26:25], 6'h00, data_i[18:17], 1'h0, data_i[15], 1'h0, data_i[13:10], 1'h0, data_i[8], 2'h0, data_i[5], 2'h0, data_i[2], 1'h0, data_i[0] };
assign syndrome_o[1] = ^ /* src = "generated/sv2v_out.v:29273.19-29273.64" */ { 5'h00, _000_[33], 1'h0, data_i[31:30], 1'h0, data_i[28:25], 1'h0, data_i[23], 1'h0, data_i[21:19], 1'h0, data_i[17], 1'h0, data_i[15], 8'h00, data_i[6], 1'h0, data_i[4], 4'h0 };
assign syndrome_o[2] = ^ /* src = "generated/sv2v_out.v:29274.19-29274.64" */ { 4'h0, data_i[34], 3'h0, data_i[30], 5'h00, data_i[24], 2'h0, data_i[21:18], 1'h0, data_i[16:15], 3'h0, data_i[11], 2'h0, data_i[8:7], 1'h0, data_i[5], 1'h0, data_i[3], 1'h0, data_i[1], 1'h0 };
assign syndrome_o[3] = ^ /* src = "generated/sv2v_out.v:29275.19-29275.64" */ { 3'h0, _001_[35], 5'h00, data_i[29:28], 3'h0, data_i[24], 2'h0, data_i[21], 3'h0, data_i[17:16], 1'h0, data_i[14], 2'h0, data_i[11:9], 1'h0, data_i[7:6], 1'h0, data_i[4], 3'h0, data_i[0] };
assign syndrome_o[4] = ^ /* src = "generated/sv2v_out.v:29276.19-29276.64" */ { 2'h0, data_i[36], 4'h0, data_i[31:30], 4'h0, data_i[25], 1'h0, data_i[23:22], 5'h00, data_i[16], 2'h0, data_i[13:12], 2'h0, data_i[9], 3'h0, data_i[5:3], 1'h0, data_i[1:0] };
assign syndrome_o[5] = ^ /* src = "generated/sv2v_out.v:29277.19-29277.64" */ { 1'h0, _002_[37], 7'h00, data_i[29], 1'h0, data_i[27:26], 1'h0, data_i[24:22], 2'h0, data_i[19:18], 3'h0, data_i[14:13], 3'h0, data_i[9], 2'h0, data_i[6], 2'h0, data_i[3:2], 2'h0 };
assign syndrome_o[6] = ^ /* src = "generated/sv2v_out.v:29278.19-29278.64" */ { data_i[38], 6'h00, data_i[31], 2'h0, data_i[28:27], 4'h0, data_i[22], 1'h0, data_i[20], 5'h00, data_i[14], 1'h0, data_i[12], 1'h0, data_i[10], 1'h0, data_i[8:7], 4'h0, data_i[2:1], 1'h0 };
assign err_o[0] = ^ /* src = "generated/sv2v_out.v:29311.14-29311.25" */ syndrome_o;
assign data_o[0] = _042_ ^ /* src = "generated/sv2v_out.v:29279.15-29279.48" */ data_i[0];
assign data_o[1] = _044_ ^ /* src = "generated/sv2v_out.v:29280.15-29280.48" */ data_i[1];
assign data_o[2] = _046_ ^ /* src = "generated/sv2v_out.v:29281.15-29281.48" */ data_i[2];
assign data_o[3] = _048_ ^ /* src = "generated/sv2v_out.v:29282.15-29282.48" */ data_i[3];
assign data_o[4] = _050_ ^ /* src = "generated/sv2v_out.v:29283.15-29283.48" */ data_i[4];
assign data_o[5] = _052_ ^ /* src = "generated/sv2v_out.v:29284.15-29284.48" */ data_i[5];
assign data_o[6] = _054_ ^ /* src = "generated/sv2v_out.v:29285.15-29285.48" */ data_i[6];
assign data_o[7] = _056_ ^ /* src = "generated/sv2v_out.v:29286.15-29286.48" */ data_i[7];
assign data_o[8] = _058_ ^ /* src = "generated/sv2v_out.v:29287.15-29287.48" */ data_i[8];
assign data_o[9] = _060_ ^ /* src = "generated/sv2v_out.v:29288.15-29288.48" */ data_i[9];
assign data_o[10] = _062_ ^ /* src = "generated/sv2v_out.v:29289.16-29289.50" */ data_i[10];
assign data_o[11] = _064_ ^ /* src = "generated/sv2v_out.v:29290.16-29290.50" */ data_i[11];
assign data_o[12] = _066_ ^ /* src = "generated/sv2v_out.v:29291.16-29291.50" */ data_i[12];
assign data_o[13] = _068_ ^ /* src = "generated/sv2v_out.v:29292.16-29292.50" */ data_i[13];
assign data_o[14] = _070_ ^ /* src = "generated/sv2v_out.v:29293.16-29293.50" */ data_i[14];
assign data_o[15] = _072_ ^ /* src = "generated/sv2v_out.v:29294.16-29294.50" */ data_i[15];
assign data_o[16] = _074_ ^ /* src = "generated/sv2v_out.v:29295.16-29295.50" */ data_i[16];
assign data_o[17] = _076_ ^ /* src = "generated/sv2v_out.v:29296.16-29296.50" */ data_i[17];
assign data_o[18] = _078_ ^ /* src = "generated/sv2v_out.v:29297.16-29297.50" */ data_i[18];
assign data_o[19] = _080_ ^ /* src = "generated/sv2v_out.v:29298.16-29298.50" */ data_i[19];
assign data_o[20] = _082_ ^ /* src = "generated/sv2v_out.v:29299.16-29299.50" */ data_i[20];
assign data_o[21] = _084_ ^ /* src = "generated/sv2v_out.v:29300.16-29300.50" */ data_i[21];
assign data_o[22] = _086_ ^ /* src = "generated/sv2v_out.v:29301.16-29301.50" */ data_i[22];
assign data_o[23] = _088_ ^ /* src = "generated/sv2v_out.v:29302.16-29302.50" */ data_i[23];
assign data_o[24] = _090_ ^ /* src = "generated/sv2v_out.v:29303.16-29303.50" */ data_i[24];
assign data_o[25] = _092_ ^ /* src = "generated/sv2v_out.v:29304.16-29304.50" */ data_i[25];
assign data_o[26] = _094_ ^ /* src = "generated/sv2v_out.v:29305.16-29305.50" */ data_i[26];
assign data_o[27] = _096_ ^ /* src = "generated/sv2v_out.v:29306.16-29306.50" */ data_i[27];
assign data_o[28] = _098_ ^ /* src = "generated/sv2v_out.v:29307.16-29307.50" */ data_i[28];
assign data_o[29] = _100_ ^ /* src = "generated/sv2v_out.v:29308.16-29308.50" */ data_i[29];
assign data_o[30] = _102_ ^ /* src = "generated/sv2v_out.v:29309.16-29309.50" */ data_i[30];
assign data_o[31] = _104_ ^ /* src = "generated/sv2v_out.v:29310.16-29310.50" */ data_i[31];
assign { _000_[38:34], _000_[32:0] } = { 6'h00, data_i[31:30], 1'h0, data_i[28:25], 1'h0, data_i[23], 1'h0, data_i[21:19], 1'h0, data_i[17], 1'h0, data_i[15], 8'h00, data_i[6], 1'h0, data_i[4], 4'h0 };
assign { _001_[38:36], _001_[34:0] } = { 8'h00, data_i[29:28], 3'h0, data_i[24], 2'h0, data_i[21], 3'h0, data_i[17:16], 1'h0, data_i[14], 2'h0, data_i[11:9], 1'h0, data_i[7:6], 1'h0, data_i[4], 3'h0, data_i[0] };
assign { _002_[38], _002_[36:0] } = { 8'h00, data_i[29], 1'h0, data_i[27:26], 1'h0, data_i[24:22], 2'h0, data_i[19:18], 3'h0, data_i[14:13], 3'h0, data_i[9], 2'h0, data_i[6], 2'h0, data_i[3:2], 2'h0 };
endmodule

module prim_secded_inv_39_32_enc(data_i, data_o, data_o_t0, data_i_t0);
/* src = "generated/sv2v_out.v:29328.16-29328.42" */
wire _00_;
/* src = "generated/sv2v_out.v:29330.16-29330.42" */
wire _01_;
/* src = "generated/sv2v_out.v:29332.16-29332.42" */
wire _02_;
/* src = "generated/sv2v_out.v:29319.15-29319.21" */
input [31:0] data_i;
wire [31:0] data_i;
/* cellift = 32'd1 */
input [31:0] data_i_t0;
wire [31:0] data_i_t0;
/* src = "generated/sv2v_out.v:29320.20-29320.26" */
output [38:0] data_o;
wire [38:0] data_o;
/* cellift = 32'd1 */
output [38:0] data_o_t0;
wire [38:0] data_o_t0;
assign { data_o[37], data_o[35], data_o[33] } = ~ { _02_, _01_, _00_ };
assign data_o_t0[32] = | { data_i_t0[29], data_i_t0[26:25], data_i_t0[18:17], data_i_t0[15], data_i_t0[13:10], data_i_t0[8], data_i_t0[5], data_i_t0[2], data_i_t0[0] };
assign data_o_t0[33] = | { data_i_t0[31:30], data_i_t0[28:25], data_i_t0[23], data_i_t0[21:19], data_i_t0[17], data_i_t0[15], data_i_t0[6], data_i_t0[4] };
assign data_o_t0[34] = | { data_i_t0[30], data_i_t0[24], data_i_t0[21:18], data_i_t0[16:15], data_i_t0[11], data_i_t0[8:7], data_i_t0[5], data_i_t0[3], data_i_t0[1] };
assign data_o_t0[35] = | { data_i_t0[29:28], data_i_t0[24], data_i_t0[21], data_i_t0[17:16], data_i_t0[14], data_i_t0[11:9], data_i_t0[7:6], data_i_t0[4], data_i_t0[0] };
assign data_o_t0[36] = | { data_i_t0[31:30], data_i_t0[25], data_i_t0[23:22], data_i_t0[16], data_i_t0[13:12], data_i_t0[9], data_i_t0[5:3], data_i_t0[1:0] };
assign data_o_t0[37] = | { data_i_t0[29], data_i_t0[27:26], data_i_t0[24:22], data_i_t0[19:18], data_i_t0[14:13], data_i_t0[9], data_i_t0[6], data_i_t0[3:2] };
assign data_o_t0[38] = | { data_i_t0[31], data_i_t0[28:27], data_i_t0[22], data_i_t0[20], data_i_t0[14], data_i_t0[12], data_i_t0[10], data_i_t0[8:7], data_i_t0[2:1] };
assign data_o[32] = ^ /* src = "generated/sv2v_out.v:29327.16-29327.42" */ { 9'h000, data_i[29], 2'h0, data_i[26:25], 6'h00, data_i[18:17], 1'h0, data_i[15], 1'h0, data_i[13:10], 1'h0, data_i[8], 2'h0, data_i[5], 2'h0, data_i[2], 1'h0, data_i[0] };
assign _00_ = ^ /* src = "generated/sv2v_out.v:29328.16-29328.42" */ { 7'h00, data_i[31:30], 1'h0, data_i[28:25], 1'h0, data_i[23], 1'h0, data_i[21:19], 1'h0, data_i[17], 1'h0, data_i[15], 8'h00, data_i[6], 1'h0, data_i[4], 4'h0 };
assign data_o[34] = ^ /* src = "generated/sv2v_out.v:29329.16-29329.42" */ { 8'h00, data_i[30], 5'h00, data_i[24], 2'h0, data_i[21:18], 1'h0, data_i[16:15], 3'h0, data_i[11], 2'h0, data_i[8:7], 1'h0, data_i[5], 1'h0, data_i[3], 1'h0, data_i[1], 1'h0 };
assign _01_ = ^ /* src = "generated/sv2v_out.v:29330.16-29330.42" */ { 9'h000, data_i[29:28], 3'h0, data_i[24], 2'h0, data_i[21], 3'h0, data_i[17:16], 1'h0, data_i[14], 2'h0, data_i[11:9], 1'h0, data_i[7:6], 1'h0, data_i[4], 3'h0, data_i[0] };
assign data_o[36] = ^ /* src = "generated/sv2v_out.v:29331.16-29331.42" */ { 7'h00, data_i[31:30], 4'h0, data_i[25], 1'h0, data_i[23:22], 5'h00, data_i[16], 2'h0, data_i[13:12], 2'h0, data_i[9], 3'h0, data_i[5:3], 1'h0, data_i[1:0] };
assign _02_ = ^ /* src = "generated/sv2v_out.v:29332.16-29332.42" */ { 9'h000, data_i[29], 1'h0, data_i[27:26], 1'h0, data_i[24:22], 2'h0, data_i[19:18], 3'h0, data_i[14:13], 3'h0, data_i[9], 2'h0, data_i[6], 2'h0, data_i[3:2], 2'h0 };
assign data_o[38] = ^ /* src = "generated/sv2v_out.v:29333.16-29333.42" */ { 7'h00, data_i[31], 2'h0, data_i[28:27], 4'h0, data_i[22], 1'h0, data_i[20], 5'h00, data_i[14], 1'h0, data_i[12], 1'h0, data_i[10], 1'h0, data_i[8:7], 4'h0, data_i[2:1], 1'h0 };
assign data_o[31:0] = data_i;
assign data_o_t0[31:0] = data_i_t0;
endmodule